

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6387, n6388, n6389, n6390, n6392, n6394, n6395, n6396, n6398, n6399,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6415, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173;

  AND2_X1 U7135 ( .A1(n13901), .A2(n13902), .ZN(n14125) );
  NOR2_X1 U7136 ( .A1(n14370), .A2(n14369), .ZN(n14371) );
  INV_X1 U7137 ( .A(n14130), .ZN(n13926) );
  NAND3_X1 U7138 ( .A1(n6931), .A2(n14022), .A3(n6930), .ZN(n13963) );
  NAND2_X1 U7140 ( .A1(n11885), .A2(n11884), .ZN(n13969) );
  CLKBUF_X1 U7141 ( .A(n12488), .Z(n6403) );
  AND2_X1 U7142 ( .A1(n10712), .A2(n10723), .ZN(n10849) );
  NOR2_X1 U7143 ( .A1(n10496), .A2(n10495), .ZN(n10524) );
  NAND2_X1 U7144 ( .A1(n11025), .A2(n11023), .ZN(n7165) );
  AND2_X1 U7145 ( .A1(n9658), .A2(n8734), .ZN(n10680) );
  INV_X2 U7146 ( .A(n9450), .ZN(n9078) );
  NAND2_X1 U7147 ( .A1(n10691), .A2(n10771), .ZN(n9116) );
  INV_X1 U7149 ( .A(n9167), .ZN(n9177) );
  CLKBUF_X2 U7150 ( .A(n8175), .Z(n6411) );
  CLKBUF_X2 U7151 ( .A(n7596), .Z(n6410) );
  INV_X2 U7152 ( .A(n11471), .ZN(n9436) );
  INV_X2 U7154 ( .A(n11849), .ZN(n11085) );
  INV_X1 U7155 ( .A(n12167), .ZN(n11548) );
  NAND2_X1 U7156 ( .A1(n7541), .A2(n7540), .ZN(n13564) );
  NAND2_X1 U7157 ( .A1(n6942), .A2(n6941), .ZN(n7541) );
  INV_X4 U7158 ( .A(n6396), .ZN(n9812) );
  INV_X4 U7159 ( .A(n6395), .ZN(n9828) );
  NAND2_X2 U7160 ( .A1(n9791), .A2(n14238), .ZN(n11835) );
  OR2_X1 U7161 ( .A1(n9679), .A2(n9668), .ZN(n9681) );
  NAND4_X1 U7162 ( .A1(n12625), .A2(n9465), .A3(n9713), .A4(n6927), .ZN(n9696)
         );
  INV_X2 U7163 ( .A(n13420), .ZN(n13394) );
  INV_X1 U7164 ( .A(n12037), .ZN(n12033) );
  INV_X1 U7165 ( .A(n12173), .ZN(n12128) );
  AOI21_X1 U7166 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10525), .A(n10524), .ZN(
        n10651) );
  NOR2_X1 U7167 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8198) );
  NOR2_X1 U7168 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7819) );
  INV_X1 U7169 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9849) );
  INV_X2 U7170 ( .A(n6401), .ZN(n8764) );
  OR2_X1 U7171 ( .A1(n15082), .A2(n15069), .ZN(n8987) );
  AND2_X1 U7172 ( .A1(n8420), .A2(n8419), .ZN(n8447) );
  INV_X1 U7173 ( .A(n7589), .ZN(n7854) );
  INV_X2 U7174 ( .A(n6410), .ZN(n7855) );
  CLKBUF_X2 U7175 ( .A(n11746), .Z(n11863) );
  NAND2_X1 U7176 ( .A1(n6591), .A2(n11138), .ZN(n14590) );
  INV_X1 U7177 ( .A(n8609), .ZN(n8523) );
  CLKBUF_X3 U7179 ( .A(n6411), .Z(n8587) );
  OAI21_X1 U7180 ( .B1(n8477), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8478) );
  BUF_X1 U7181 ( .A(n11832), .Z(n6395) );
  INV_X2 U7182 ( .A(n11928), .ZN(n9756) );
  INV_X1 U7183 ( .A(n11709), .ZN(n9682) );
  NAND2_X1 U7184 ( .A1(n9683), .A2(n11709), .ZN(n9745) );
  NOR2_X1 U7185 ( .A1(n13901), .A2(n13859), .ZN(n13860) );
  XNOR2_X1 U7186 ( .A(n7512), .B(n7510), .ZN(n7909) );
  XNOR2_X1 U7187 ( .A(n10312), .B(n10311), .ZN(n10313) );
  OAI22_X1 U7188 ( .A1(n10313), .A2(n14866), .B1(n10312), .B2(n10311), .ZN(
        n10339) );
  XNOR2_X1 U7189 ( .A(n7109), .B(n12474), .ZN(n14369) );
  NOR2_X1 U7190 ( .A1(n14371), .A2(n12436), .ZN(n14387) );
  NAND2_X1 U7191 ( .A1(n7897), .A2(n7896), .ZN(n13299) );
  INV_X1 U7192 ( .A(n10885), .ZN(n14623) );
  AND4_X1 U7193 ( .A1(n9790), .A2(n9789), .A3(n9788), .A4(n9787), .ZN(n12011)
         );
  NAND2_X1 U7194 ( .A1(n14017), .A2(n6479), .ZN(n14001) );
  NAND2_X1 U7195 ( .A1(n11519), .A2(n11518), .ZN(n14481) );
  AOI21_X1 U7196 ( .B1(n14122), .B2(n14625), .A(n6453), .ZN(n6702) );
  XNOR2_X1 U7197 ( .A(n6880), .B(n9349), .ZN(n14226) );
  INV_X1 U7198 ( .A(n6621), .ZN(n8875) );
  NAND2_X1 U7199 ( .A1(n11835), .A2(n14251), .ZN(n14007) );
  XNOR2_X1 U7200 ( .A(n8875), .B(n6966), .ZN(n14291) );
  CLKBUF_X3 U7201 ( .A(n7626), .Z(n6390) );
  XOR2_X1 U7202 ( .A(n13856), .B(n12181), .Z(n6387) );
  AND2_X1 U7203 ( .A1(n7003), .A2(n6468), .ZN(n6388) );
  XNOR2_X2 U7204 ( .A(n8108), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8366) );
  XNOR2_X2 U7205 ( .A(n7539), .B(n7538), .ZN(n8033) );
  NAND2_X2 U7206 ( .A1(n11457), .A2(n6492), .ZN(n11497) );
  NOR2_X2 U7207 ( .A1(n14044), .A2(n6648), .ZN(n14018) );
  AOI21_X2 U7208 ( .B1(n7009), .B2(n7007), .A(n6537), .ZN(n7008) );
  NAND2_X2 U7209 ( .A1(n6879), .A2(n7444), .ZN(n7633) );
  XNOR2_X2 U7211 ( .A(n8149), .B(n12969), .ZN(n8152) );
  AOI21_X1 U7212 ( .B1(n12358), .B2(n12743), .A(n8788), .ZN(n8789) );
  NOR2_X2 U7213 ( .A1(n13254), .A2(n6498), .ZN(n13240) );
  NAND2_X2 U7214 ( .A1(n7742), .A2(n7413), .ZN(n7471) );
  NAND2_X2 U7215 ( .A1(n8107), .A2(n6710), .ZN(n8108) );
  INV_X2 U7216 ( .A(n9683), .ZN(n14233) );
  XNOR2_X2 U7217 ( .A(n9678), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9683) );
  INV_X4 U7218 ( .A(n9167), .ZN(n9369) );
  INV_X8 U7219 ( .A(n9190), .ZN(n9167) );
  INV_X2 U7220 ( .A(n10471), .ZN(n10559) );
  XNOR2_X1 U7221 ( .A(n13733), .B(n14589), .ZN(n14582) );
  NAND4_X2 U7222 ( .A1(n9750), .A2(n9749), .A3(n9748), .A4(n9747), .ZN(n13733)
         );
  XNOR2_X2 U7223 ( .A(n9571), .B(n9572), .ZN(n11603) );
  NAND2_X2 U7224 ( .A1(n11557), .A2(n9570), .ZN(n9571) );
  BUF_X1 U7225 ( .A(n7626), .Z(n6389) );
  AND2_X2 U7226 ( .A1(n6925), .A2(n6388), .ZN(n8652) );
  AND2_X2 U7227 ( .A1(n6926), .A2(n7002), .ZN(n6925) );
  NAND2_X1 U7228 ( .A1(n12547), .A2(n8568), .ZN(n12532) );
  NAND2_X2 U7229 ( .A1(n7909), .A2(SI_23_), .ZN(n7911) );
  AOI211_X2 U7230 ( .C1(n6950), .C2(n13189), .A(n13394), .B(n13188), .ZN(
        n13433) );
  XNOR2_X2 U7231 ( .A(n15060), .B(n8229), .ZN(n15043) );
  OAI21_X2 U7232 ( .B1(n7728), .B2(n7727), .A(n7466), .ZN(n7742) );
  NAND2_X2 U7233 ( .A1(n7462), .A2(n7461), .ZN(n7728) );
  XNOR2_X2 U7234 ( .A(n7458), .B(SI_9_), .ZN(n7690) );
  OAI21_X2 U7235 ( .B1(n10950), .B2(n10949), .A(n10948), .ZN(n13690) );
  AOI21_X2 U7236 ( .B1(n10802), .B2(n10801), .A(n6818), .ZN(n10950) );
  XNOR2_X2 U7237 ( .A(n13752), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n8847) );
  INV_X4 U7238 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n13752) );
  OAI22_X2 U7239 ( .A1(n14874), .A2(n14873), .B1(n10490), .B2(n6844), .ZN(
        n10518) );
  AOI21_X2 U7240 ( .B1(n10489), .B2(n10488), .A(n6641), .ZN(n14874) );
  OAI222_X1 U7242 ( .A1(P3_U3151), .A2(n10311), .B1(n14275), .B2(n9821), .C1(
        n14277), .C2(n9820), .ZN(P3_U3294) );
  XNOR2_X2 U7243 ( .A(n9681), .B(n9680), .ZN(n11709) );
  NAND2_X2 U7244 ( .A1(n8973), .A2(n12900), .ZN(n15088) );
  AND2_X2 U7246 ( .A1(n8981), .A2(n8985), .ZN(n15087) );
  AOI21_X2 U7247 ( .B1(n7086), .B2(n8223), .A(n7084), .ZN(n7083) );
  XNOR2_X2 U7248 ( .A(n7433), .B(SI_2_), .ZN(n7593) );
  XNOR2_X2 U7249 ( .A(n7439), .B(SI_3_), .ZN(n7614) );
  NAND2_X2 U7250 ( .A1(n6582), .A2(n7437), .ZN(n7439) );
  NAND2_X2 U7251 ( .A1(n15012), .A2(n8299), .ZN(n11317) );
  NAND2_X2 U7252 ( .A1(n7165), .A2(n7164), .ZN(n15012) );
  AOI21_X2 U7253 ( .B1(n10898), .B2(n10899), .A(n8741), .ZN(n10928) );
  XNOR2_X2 U7254 ( .A(n13126), .B(n6760), .ZN(n10594) );
  XNOR2_X2 U7255 ( .A(n7427), .B(SI_1_), .ZN(n7586) );
  NAND2_X2 U7256 ( .A1(n6580), .A2(n6699), .ZN(n7427) );
  BUF_X4 U7257 ( .A(n6675), .Z(n6413) );
  AND2_X2 U7258 ( .A1(n8987), .A2(n8989), .ZN(n15059) );
  CLKBUF_X1 U7259 ( .A(n14238), .Z(n6394) );
  NAND4_X2 U7260 ( .A1(n8174), .A2(n8173), .A3(n8172), .A4(n8171), .ZN(n15083)
         );
  NAND2_X1 U7261 ( .A1(n15063), .A2(n8216), .ZN(n15040) );
  XNOR2_X2 U7262 ( .A(n6819), .B(n7385), .ZN(n10802) );
  OAI21_X2 U7263 ( .B1(n14091), .B2(n13868), .A(n13869), .ZN(n14076) );
  NAND2_X2 U7264 ( .A1(n6590), .A2(n13866), .ZN(n14091) );
  XNOR2_X1 U7265 ( .A(n8735), .B(n15082), .ZN(n10679) );
  XNOR2_X2 U7266 ( .A(n8822), .B(n10480), .ZN(n8856) );
  AND3_X2 U7267 ( .A1(n6955), .A2(n6954), .A3(n6546), .ZN(n8822) );
  NAND2_X2 U7268 ( .A1(n12513), .A2(n9092), .ZN(n12505) );
  BUF_X2 U7269 ( .A(n11832), .Z(n6396) );
  INV_X1 U7270 ( .A(n7476), .ZN(n11832) );
  NOR2_X4 U7271 ( .A1(n14523), .A2(n6786), .ZN(n14526) );
  AND2_X1 U7272 ( .A1(n10290), .A2(n9828), .ZN(n8175) );
  CLKBUF_X1 U7273 ( .A(n13008), .Z(n6398) );
  OAI211_X1 U7276 ( .C1(n7589), .C2(n13154), .A(n7617), .B(n7616), .ZN(n13008)
         );
  OAI22_X2 U7277 ( .A1(n8289), .A2(n8099), .B1(P1_DATAO_REG_8__SCAN_IN), .B2(
        n9860), .ZN(n8308) );
  OAI21_X2 U7278 ( .B1(n8273), .B2(n8272), .A(n8098), .ZN(n8289) );
  AND2_X4 U7279 ( .A1(n11929), .A2(n11966), .ZN(n11928) );
  OAI22_X2 U7280 ( .A1(n7476), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n7432), .ZN(n7433) );
  AND2_X2 U7281 ( .A1(n9760), .A2(n9775), .ZN(n9494) );
  OAI22_X2 U7282 ( .A1(n10473), .A2(n10474), .B1(n10316), .B2(n7120), .ZN(
        n10489) );
  AOI22_X2 U7283 ( .A1(n10339), .A2(n10340), .B1(n10351), .B2(n10315), .ZN(
        n10473) );
  BUF_X4 U7284 ( .A(n12296), .Z(n6401) );
  BUF_X4 U7285 ( .A(n12296), .Z(n6402) );
  NAND2_X2 U7286 ( .A1(n8726), .A2(n9116), .ZN(n12296) );
  XNOR2_X1 U7287 ( .A(n8478), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12488) );
  OAI22_X2 U7288 ( .A1(n8197), .A2(n8088), .B1(P2_DATAO_REG_2__SCAN_IN), .B2(
        n9825), .ZN(n8211) );
  XNOR2_X2 U7289 ( .A(n7544), .B(n13552), .ZN(n12247) );
  NAND2_X2 U7290 ( .A1(n13551), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7544) );
  XNOR2_X2 U7291 ( .A(n8151), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8153) );
  OR2_X2 U7292 ( .A1(n8150), .A2(n8416), .ZN(n8151) );
  NOR2_X2 U7293 ( .A1(n8859), .A2(n8860), .ZN(n8863) );
  XNOR2_X2 U7294 ( .A(n6783), .B(n8879), .ZN(n14292) );
  NAND2_X2 U7295 ( .A1(n8877), .A2(n8878), .ZN(n6783) );
  OR2_X1 U7296 ( .A1(n13180), .A2(n13183), .ZN(n9385) );
  INV_X1 U7297 ( .A(n9388), .ZN(n13517) );
  INV_X2 U7298 ( .A(n12511), .ZN(n12518) );
  NAND2_X1 U7299 ( .A1(n7567), .A2(n7566), .ZN(n13267) );
  NOR2_X2 U7300 ( .A1(n13335), .A2(n13319), .ZN(n13318) );
  INV_X1 U7301 ( .A(n14170), .ZN(n14028) );
  NAND2_X1 U7302 ( .A1(n10006), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13096) );
  INV_X1 U7303 ( .A(n10623), .ZN(n6760) );
  XNOR2_X1 U7304 ( .A(n10681), .B(n6401), .ZN(n8735) );
  CLKBUF_X2 U7305 ( .A(n13026), .Z(n6712) );
  NAND4_X1 U7306 ( .A1(n8239), .A2(n8238), .A3(n8237), .A4(n8236), .ZN(n11052)
         );
  NAND2_X1 U7307 ( .A1(n8104), .A2(n7091), .ZN(n8342) );
  CLKBUF_X2 U7308 ( .A(n7599), .Z(n8036) );
  BUF_X1 U7309 ( .A(n10290), .Z(n6675) );
  NAND2_X1 U7310 ( .A1(n7589), .A2(n9812), .ZN(n7596) );
  NAND2_X2 U7311 ( .A1(n11059), .A2(n9428), .ZN(n9500) );
  INV_X2 U7312 ( .A(n14559), .ZN(n12226) );
  BUF_X2 U7313 ( .A(n7578), .Z(n8038) );
  NOR2_X1 U7314 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8124) );
  AND3_X1 U7315 ( .A1(n7187), .A2(n12221), .A3(n7185), .ZN(n7184) );
  AND2_X1 U7316 ( .A1(n6531), .A2(n7060), .ZN(n8723) );
  OAI21_X1 U7317 ( .B1(n9384), .B2(n9383), .A(n6674), .ZN(n6714) );
  AND2_X1 U7318 ( .A1(n12491), .A2(n15136), .ZN(n7422) );
  NOR2_X1 U7319 ( .A1(n12515), .A2(n12514), .ZN(n12523) );
  AOI21_X1 U7320 ( .B1(n7200), .B2(n12180), .A(n7199), .ZN(n7198) );
  OAI21_X1 U7321 ( .B1(n7072), .B2(n9117), .A(n7071), .ZN(n7068) );
  AND3_X1 U7322 ( .A1(n13189), .A2(n8716), .A3(n13420), .ZN(n13436) );
  AND2_X1 U7323 ( .A1(n7171), .A2(n7170), .ZN(n12833) );
  OAI21_X1 U7324 ( .B1(n13517), .B2(n9177), .A(n9361), .ZN(n9382) );
  AOI21_X1 U7325 ( .B1(n13934), .B2(n14625), .A(n13933), .ZN(n14137) );
  NAND2_X1 U7326 ( .A1(n6581), .A2(n9350), .ZN(n13180) );
  OR2_X1 U7327 ( .A1(n7031), .A2(n7027), .ZN(n7026) );
  NAND2_X1 U7328 ( .A1(n12162), .A2(n12161), .ZN(n13859) );
  CLKBUF_X1 U7329 ( .A(n12546), .Z(n6409) );
  AOI21_X1 U7330 ( .B1(n6768), .B2(n7330), .A(n7327), .ZN(n13237) );
  NOR2_X1 U7331 ( .A1(n13240), .A2(n13239), .ZN(n13238) );
  AOI21_X1 U7332 ( .B1(n6766), .B2(n6764), .A(n6505), .ZN(n6763) );
  INV_X1 U7333 ( .A(n7256), .ZN(n7255) );
  AND2_X1 U7334 ( .A1(n9357), .A2(n9356), .ZN(n12245) );
  OR2_X1 U7335 ( .A1(n13958), .A2(n13961), .ZN(n7361) );
  NAND2_X1 U7336 ( .A1(n12182), .A2(n13878), .ZN(n13961) );
  NOR2_X1 U7337 ( .A1(n13931), .A2(n6622), .ZN(n7258) );
  INV_X1 U7338 ( .A(n13939), .ZN(n6701) );
  NAND2_X1 U7339 ( .A1(n6881), .A2(n9346), .ZN(n9357) );
  NAND2_X1 U7340 ( .A1(n12150), .A2(n12149), .ZN(n14126) );
  NAND2_X1 U7341 ( .A1(n7962), .A2(n7961), .ZN(n13199) );
  OAI211_X1 U7342 ( .C1(n7042), .C2(n13308), .A(n7043), .B(n7040), .ZN(n13255)
         );
  AND2_X1 U7343 ( .A1(n13974), .A2(n13973), .ZN(n13976) );
  NAND2_X1 U7344 ( .A1(n6605), .A2(n6604), .ZN(n12305) );
  XNOR2_X1 U7345 ( .A(n13267), .B(n13242), .ZN(n13256) );
  OR2_X1 U7346 ( .A1(n12830), .A2(n12265), .ZN(n9100) );
  CLKBUF_X1 U7347 ( .A(n12830), .Z(n6688) );
  NAND2_X1 U7348 ( .A1(n7929), .A2(n7928), .ZN(n13246) );
  NOR2_X1 U7349 ( .A1(n13983), .A2(n6932), .ZN(n6931) );
  NAND2_X1 U7350 ( .A1(n13657), .A2(n13656), .ZN(n13655) );
  NAND2_X1 U7351 ( .A1(n11711), .A2(n11710), .ZN(n14135) );
  AOI21_X1 U7352 ( .B1(n12978), .B2(n6411), .A(n8586), .ZN(n12494) );
  XNOR2_X1 U7353 ( .A(n9341), .B(n9340), .ZN(n12147) );
  AND2_X1 U7354 ( .A1(n6918), .A2(n6543), .ZN(n12755) );
  XNOR2_X1 U7355 ( .A(n8691), .B(n8690), .ZN(n14235) );
  NAND2_X1 U7356 ( .A1(n7543), .A2(n7542), .ZN(n13229) );
  AND2_X1 U7357 ( .A1(n6958), .A2(n14828), .ZN(n6618) );
  NAND2_X1 U7358 ( .A1(n8943), .A2(n8942), .ZN(n14411) );
  NAND2_X1 U7359 ( .A1(n7399), .A2(n6491), .ZN(n13603) );
  XNOR2_X1 U7360 ( .A(n8931), .B(n7101), .ZN(n12978) );
  NAND2_X1 U7361 ( .A1(n6596), .A2(n6882), .ZN(n9341) );
  NOR2_X1 U7362 ( .A1(n14159), .A2(n6934), .ZN(n6933) );
  NAND2_X1 U7363 ( .A1(n13318), .A2(n13532), .ZN(n13301) );
  NAND2_X1 U7364 ( .A1(n13680), .A2(n13679), .ZN(n7399) );
  NAND2_X2 U7365 ( .A1(n11853), .A2(n11852), .ZN(n14159) );
  XNOR2_X1 U7366 ( .A(n7940), .B(n7523), .ZN(n13565) );
  OAI21_X1 U7367 ( .B1(n7940), .B2(n6564), .A(n7939), .ZN(n7957) );
  AND2_X1 U7368 ( .A1(n7925), .A2(n7367), .ZN(n13572) );
  INV_X1 U7369 ( .A(n9096), .ZN(n12512) );
  NAND2_X1 U7370 ( .A1(n7364), .A2(n7565), .ZN(n7925) );
  NAND2_X1 U7371 ( .A1(n6703), .A2(n7522), .ZN(n7940) );
  NAND2_X1 U7372 ( .A1(n13637), .A2(n11752), .ZN(n13680) );
  OR2_X1 U7373 ( .A1(n11850), .A2(n6647), .ZN(n11853) );
  AND2_X1 U7374 ( .A1(n12838), .A2(n12550), .ZN(n9096) );
  OAI21_X1 U7375 ( .B1(n7911), .B2(n7519), .A(n7518), .ZN(n6703) );
  AND2_X1 U7376 ( .A1(n8574), .A2(n8573), .ZN(n12838) );
  AOI21_X1 U7377 ( .B1(n7517), .B2(n7564), .A(n7516), .ZN(n7518) );
  XNOR2_X1 U7378 ( .A(n11834), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14251) );
  NAND2_X1 U7379 ( .A1(n8560), .A2(n8559), .ZN(n12845) );
  AND2_X1 U7380 ( .A1(n7512), .A2(n7511), .ZN(n7517) );
  NAND2_X1 U7381 ( .A1(n8629), .A2(n9044), .ZN(n12823) );
  NOR2_X1 U7382 ( .A1(n13357), .A2(n13337), .ZN(n6953) );
  NOR2_X1 U7383 ( .A1(n14065), .A2(n6480), .ZN(n14051) );
  NAND2_X1 U7384 ( .A1(n11815), .A2(n11814), .ZN(n14170) );
  NAND2_X1 U7385 ( .A1(n7504), .A2(SI_22_), .ZN(n7509) );
  NAND2_X1 U7386 ( .A1(n6588), .A2(n6984), .ZN(n13865) );
  NAND2_X1 U7387 ( .A1(n7162), .A2(n6488), .ZN(n12764) );
  AND2_X1 U7388 ( .A1(n6471), .A2(n6794), .ZN(n14516) );
  NAND2_X1 U7389 ( .A1(n7882), .A2(n7503), .ZN(n7504) );
  NAND2_X1 U7390 ( .A1(n7880), .A2(n7879), .ZN(n7882) );
  NAND2_X1 U7391 ( .A1(n11537), .A2(n11536), .ZN(n14113) );
  CLKBUF_X1 U7392 ( .A(n11715), .Z(n6609) );
  NAND2_X1 U7393 ( .A1(n7363), .A2(n7498), .ZN(n6878) );
  NAND2_X1 U7394 ( .A1(n6625), .A2(SI_20_), .ZN(n7499) );
  NAND2_X1 U7395 ( .A1(n7497), .A2(n10770), .ZN(n7363) );
  CLKBUF_X1 U7396 ( .A(n11651), .Z(n6671) );
  OR2_X1 U7397 ( .A1(n8503), .A2(n8502), .ZN(n7075) );
  AND2_X1 U7398 ( .A1(n14970), .A2(n12463), .ZN(n14994) );
  NAND2_X1 U7399 ( .A1(n7772), .A2(n7771), .ZN(n11490) );
  AND2_X1 U7400 ( .A1(n6679), .A2(n6680), .ZN(n14511) );
  NAND2_X1 U7401 ( .A1(n7493), .A2(SI_18_), .ZN(n7372) );
  NAND2_X1 U7402 ( .A1(n7371), .A2(n7370), .ZN(n7369) );
  XNOR2_X1 U7403 ( .A(n7787), .B(n7786), .ZN(n11520) );
  NAND2_X1 U7404 ( .A1(n7492), .A2(n10637), .ZN(n7371) );
  AND2_X1 U7405 ( .A1(n14955), .A2(n12459), .ZN(n14972) );
  OR2_X1 U7406 ( .A1(n14954), .A2(n14953), .ZN(n14955) );
  OAI21_X1 U7407 ( .B1(n7784), .B2(n7783), .A(n7782), .ZN(n7787) );
  NAND2_X1 U7408 ( .A1(n6896), .A2(n6897), .ZN(n7764) );
  OR2_X1 U7409 ( .A1(n7471), .A2(n6900), .ZN(n6896) );
  NAND2_X1 U7410 ( .A1(n6651), .A2(n6649), .ZN(n8414) );
  NAND2_X1 U7411 ( .A1(n11084), .A2(n11083), .ZN(n14666) );
  NAND2_X2 U7412 ( .A1(n13907), .A2(n14555), .ZN(n14562) );
  OR2_X1 U7413 ( .A1(n10527), .A2(n10526), .ZN(n6840) );
  INV_X2 U7414 ( .A(n15109), .ZN(n15005) );
  NAND2_X2 U7415 ( .A1(n7654), .A2(n7653), .ZN(n10698) );
  NAND2_X1 U7416 ( .A1(n7666), .A2(n7665), .ZN(n10766) );
  NAND2_X1 U7417 ( .A1(n7453), .A2(n7452), .ZN(n7678) );
  AND2_X1 U7418 ( .A1(n8495), .A2(n8494), .ZN(n8507) );
  NOR2_X1 U7419 ( .A1(n8865), .A2(n8864), .ZN(n8867) );
  NAND2_X1 U7420 ( .A1(n10870), .A2(n10869), .ZN(n12183) );
  AND2_X1 U7421 ( .A1(n10778), .A2(n10777), .ZN(n14634) );
  INV_X2 U7422 ( .A(n11929), .ZN(n9737) );
  NAND2_X1 U7423 ( .A1(n8342), .A2(n6554), .ZN(n8107) );
  OAI211_X1 U7424 ( .C1(n7589), .C2(n13136), .A(n7598), .B(n7597), .ZN(n10266)
         );
  NOR2_X1 U7425 ( .A1(n8828), .A2(n8829), .ZN(n8869) );
  NAND4_X2 U7426 ( .A1(n10786), .A2(n10785), .A3(n10784), .A4(n10783), .ZN(
        n13730) );
  NAND2_X1 U7427 ( .A1(n9501), .A2(n9500), .ZN(n13026) );
  NAND3_X1 U7428 ( .A1(n9727), .A2(n9726), .A3(n6589), .ZN(n11139) );
  NAND4_X1 U7429 ( .A1(n8208), .A2(n8207), .A3(n8206), .A4(n8205), .ZN(n15082)
         );
  INV_X2 U7430 ( .A(n8234), .ZN(n8547) );
  NAND4_X1 U7431 ( .A1(n7611), .A2(n7610), .A3(n7609), .A4(n7608), .ZN(n13128)
         );
  NAND2_X1 U7432 ( .A1(n6979), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6928) );
  NAND2_X2 U7433 ( .A1(n9494), .A2(n9765), .ZN(n9701) );
  OAI21_X1 U7434 ( .B1(n8308), .B2(n8101), .A(n8100), .ZN(n8325) );
  CLKBUF_X1 U7435 ( .A(n11849), .Z(n6647) );
  AND2_X1 U7436 ( .A1(n9493), .A2(n6445), .ZN(n9765) );
  AOI21_X1 U7437 ( .B1(n7457), .B2(n7344), .A(n6518), .ZN(n7343) );
  NAND2_X1 U7438 ( .A1(n7589), .A2(n11832), .ZN(n7595) );
  NAND2_X1 U7439 ( .A1(n8155), .A2(n8153), .ZN(n8234) );
  INV_X1 U7440 ( .A(n12488), .ZN(n10691) );
  NAND2_X1 U7441 ( .A1(n10285), .A2(n8604), .ZN(n10290) );
  INV_X2 U7442 ( .A(n7576), .ZN(n9351) );
  NAND2_X1 U7443 ( .A1(n11835), .A2(n9812), .ZN(n11849) );
  NAND2_X1 U7444 ( .A1(n11976), .A2(n11982), .ZN(n11966) );
  NAND2_X2 U7445 ( .A1(n8033), .A2(n13564), .ZN(n7589) );
  XNOR2_X1 U7446 ( .A(n9481), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9760) );
  NOR2_X1 U7447 ( .A1(n9777), .A2(n11982), .ZN(n11985) );
  NAND2_X1 U7448 ( .A1(n14233), .A2(n11709), .ZN(n11178) );
  XNOR2_X1 U7449 ( .A(n8140), .B(n8139), .ZN(n8604) );
  AOI21_X1 U7450 ( .B1(n7448), .B2(n7348), .A(n6519), .ZN(n7347) );
  NAND2_X1 U7451 ( .A1(n6614), .A2(n6612), .ZN(n10285) );
  NAND2_X1 U7452 ( .A1(n9495), .A2(n9675), .ZN(n11976) );
  NAND2_X4 U7453 ( .A1(n12247), .A2(n7552), .ZN(n7577) );
  NOR2_X1 U7454 ( .A1(n8823), .A2(n8824), .ZN(n8826) );
  OR2_X1 U7455 ( .A1(n7976), .A2(n12614), .ZN(n7979) );
  XNOR2_X1 U7456 ( .A(n7853), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U7457 ( .A1(n8062), .A2(n7303), .ZN(n11471) );
  NAND2_X1 U7458 ( .A1(n8138), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8140) );
  MUX2_X1 U7459 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8648), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8650) );
  NAND2_X1 U7460 ( .A1(n9692), .A2(n9693), .ZN(n14238) );
  NAND2_X2 U7461 ( .A1(n6396), .A2(P1_U3086), .ZN(n14245) );
  NAND2_X1 U7462 ( .A1(n8447), .A2(n8446), .ZN(n8477) );
  OR2_X1 U7463 ( .A1(n8649), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n6442) );
  XNOR2_X1 U7464 ( .A(n7547), .B(P2_IR_REG_29__SCAN_IN), .ZN(n7552) );
  OR2_X1 U7466 ( .A1(n7545), .A2(n7980), .ZN(n7547) );
  NOR2_X1 U7467 ( .A1(n10687), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n9702) );
  AND4_X1 U7468 ( .A1(n7743), .A2(n7339), .A3(n7532), .A4(n6545), .ZN(n7545)
         );
  AND2_X1 U7469 ( .A1(n10582), .A2(n9474), .ZN(n10385) );
  AND2_X1 U7470 ( .A1(n6926), .A2(n6924), .ZN(n6923) );
  AND2_X1 U7471 ( .A1(n8369), .A2(n8415), .ZN(n8420) );
  AND2_X1 U7472 ( .A1(n7002), .A2(n8148), .ZN(n6924) );
  OR2_X1 U7473 ( .A1(n7431), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6580) );
  AND2_X1 U7474 ( .A1(n7340), .A2(n7536), .ZN(n7339) );
  NOR2_X1 U7475 ( .A1(n7006), .A2(n7005), .ZN(n8369) );
  NAND2_X1 U7476 ( .A1(n6876), .A2(n6875), .ZN(n7431) );
  AND2_X1 U7477 ( .A1(n7174), .A2(n8212), .ZN(n7003) );
  AND2_X1 U7478 ( .A1(n8133), .A2(n8127), .ZN(n7002) );
  AND2_X1 U7479 ( .A1(n8128), .A2(n8132), .ZN(n6926) );
  NAND4_X1 U7480 ( .A1(n9704), .A2(n9476), .A3(n9475), .A4(n9477), .ZN(n9486)
         );
  AND4_X1 U7481 ( .A1(n8131), .A2(n8130), .A3(n8129), .A4(n8400), .ZN(n8132)
         );
  AND2_X1 U7482 ( .A1(n8126), .A2(n8125), .ZN(n8127) );
  AND4_X2 U7483 ( .A1(n8124), .A2(n8225), .A3(n8123), .A4(n12632), .ZN(n8128)
         );
  AND2_X2 U7484 ( .A1(n8198), .A2(n6847), .ZN(n8212) );
  NAND2_X1 U7485 ( .A1(n7537), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6941) );
  AND2_X1 U7486 ( .A1(n7176), .A2(n7175), .ZN(n7174) );
  AND2_X1 U7487 ( .A1(n8086), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U7488 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n6711), .ZN(n6710) );
  INV_X4 U7489 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7490 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n7818) );
  NOR2_X1 U7491 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8130) );
  INV_X1 U7492 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9839) );
  INV_X1 U7493 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n12614) );
  NOR2_X1 U7494 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8131) );
  INV_X1 U7495 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7627) );
  INV_X1 U7496 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9704) );
  INV_X1 U7497 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n12654) );
  INV_X1 U7498 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9856) );
  INV_X1 U7499 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7591) );
  NOR2_X1 U7500 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7590) );
  INV_X1 U7501 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8225) );
  INV_X2 U7502 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n12625) );
  INV_X4 U7503 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U7504 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7505 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n12632) );
  INV_X1 U7506 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7981) );
  INV_X1 U7507 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7176) );
  INV_X1 U7508 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8063) );
  INV_X1 U7509 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7423) );
  INV_X1 U7510 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7424) );
  INV_X1 U7511 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8647) );
  INV_X1 U7512 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8400) );
  INV_X1 U7513 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8123) );
  NOR2_X1 U7514 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8125) );
  NOR2_X1 U7515 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8126) );
  OR2_X1 U7516 ( .A1(n11923), .A2(n10895), .ZN(n10783) );
  OR2_X1 U7517 ( .A1(n7909), .A2(SI_23_), .ZN(n7910) );
  NAND2_X2 U7518 ( .A1(n13670), .A2(n11848), .ZN(n13580) );
  OAI21_X2 U7519 ( .B1(n11651), .B2(n6522), .A(n6821), .ZN(n11667) );
  NAND2_X1 U7520 ( .A1(n10871), .A2(n12001), .ZN(n11149) );
  NOR2_X2 U7521 ( .A1(n13940), .A2(n6700), .ZN(n13921) );
  XNOR2_X2 U7522 ( .A(n6666), .B(n13899), .ZN(n14127) );
  NAND2_X2 U7523 ( .A1(n8974), .A2(n8972), .ZN(n8973) );
  NAND2_X1 U7524 ( .A1(n15026), .A2(n15027), .ZN(n15025) );
  OAI21_X2 U7525 ( .B1(n11317), .B2(n7143), .A(n7140), .ZN(n11504) );
  NAND2_X2 U7526 ( .A1(n11504), .A2(n8349), .ZN(n8351) );
  AND2_X2 U7527 ( .A1(n13232), .A2(n13215), .ZN(n13216) );
  AND2_X2 U7528 ( .A1(n13951), .A2(n13939), .ZN(n13935) );
  XNOR2_X2 U7529 ( .A(n8161), .B(n7096), .ZN(n12984) );
  NAND2_X2 U7530 ( .A1(n8121), .A2(n6708), .ZN(n8161) );
  NAND2_X1 U7531 ( .A1(n8632), .A2(n6407), .ZN(n6404) );
  AND2_X2 U7532 ( .A1(n6404), .A2(n6405), .ZN(n12744) );
  OR2_X1 U7533 ( .A1(n6406), .A2(n6543), .ZN(n6405) );
  INV_X1 U7534 ( .A(n9071), .ZN(n6406) );
  AND2_X1 U7535 ( .A1(n8631), .A2(n9071), .ZN(n6407) );
  CLKBUF_X1 U7536 ( .A(n11044), .Z(n6408) );
  NAND2_X1 U7537 ( .A1(n8621), .A2(n8996), .ZN(n11044) );
  NAND2_X1 U7538 ( .A1(n8620), .A2(n8619), .ZN(n15024) );
  INV_X1 U7539 ( .A(n7595), .ZN(n7626) );
  AND2_X1 U7540 ( .A1(n9653), .A2(n6906), .ZN(n9122) );
  INV_X4 U7541 ( .A(n12033), .ZN(n12173) );
  NOR2_X2 U7542 ( .A1(n14576), .A2(n14651), .ZN(n14574) );
  AOI21_X2 U7543 ( .B1(n12733), .B2(n12732), .A(n8637), .ZN(n12575) );
  OAI21_X2 U7544 ( .B1(n12744), .B2(n8964), .A(n8636), .ZN(n12733) );
  OAI21_X2 U7545 ( .B1(n12783), .B2(n8474), .A(n9057), .ZN(n12772) );
  NAND2_X2 U7546 ( .A1(n8630), .A2(n8967), .ZN(n12783) );
  AND2_X1 U7547 ( .A1(n8155), .A2(n8153), .ZN(n6412) );
  XNOR2_X1 U7549 ( .A(n9689), .B(n9688), .ZN(n9791) );
  NOR2_X2 U7550 ( .A1(n10671), .A2(n10698), .ZN(n10712) );
  BUF_X4 U7551 ( .A(n8240), .Z(n8572) );
  INV_X2 U7552 ( .A(n7432), .ZN(n7476) );
  INV_X1 U7553 ( .A(n7431), .ZN(n7432) );
  NOR2_X2 U7554 ( .A1(n10365), .A2(n6399), .ZN(n10452) );
  OR2_X1 U7555 ( .A1(n10260), .A2(n10266), .ZN(n10365) );
  NAND2_X1 U7556 ( .A1(n8325), .A2(n8324), .ZN(n8104) );
  INV_X1 U7557 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8597) );
  INV_X1 U7558 ( .A(n12998), .ZN(n7300) );
  INV_X1 U7559 ( .A(n9613), .ZN(n7301) );
  AND2_X1 U7560 ( .A1(n7197), .A2(n7205), .ZN(n7196) );
  NAND2_X1 U7561 ( .A1(n12178), .A2(n12179), .ZN(n7205) );
  NAND2_X1 U7562 ( .A1(n7198), .A2(n7201), .ZN(n7197) );
  NAND2_X1 U7563 ( .A1(n9683), .A2(n9682), .ZN(n9721) );
  AND2_X1 U7564 ( .A1(n7244), .A2(n9476), .ZN(n7243) );
  OR2_X1 U7565 ( .A1(n12493), .A2(n8234), .ZN(n8949) );
  AND2_X1 U7566 ( .A1(n8676), .A2(n8603), .ZN(n15052) );
  OR2_X1 U7567 ( .A1(n11007), .A2(n9117), .ZN(n15076) );
  NAND2_X1 U7568 ( .A1(n8161), .A2(n8160), .ZN(n7104) );
  AND2_X1 U7569 ( .A1(n7092), .A2(n8103), .ZN(n7091) );
  INV_X1 U7570 ( .A(n8339), .ZN(n7092) );
  AOI21_X1 U7571 ( .B1(n7083), .B2(n7085), .A(n7081), .ZN(n7080) );
  NAND2_X1 U7572 ( .A1(n6450), .A2(n6745), .ZN(n6743) );
  NAND2_X1 U7573 ( .A1(n7133), .A2(n7132), .ZN(n6740) );
  NOR2_X1 U7574 ( .A1(n6449), .A2(n7134), .ZN(n7133) );
  NOR2_X1 U7575 ( .A1(n7183), .A2(n6500), .ZN(n7178) );
  MUX2_X1 U7576 ( .A(n14159), .B(n13876), .S(n12037), .Z(n12111) );
  OAI21_X1 U7577 ( .B1(n9316), .B2(n7137), .A(n7136), .ZN(n9321) );
  AND2_X1 U7578 ( .A1(n9314), .A2(n9315), .ZN(n7137) );
  OR2_X1 U7579 ( .A1(n9315), .A2(n9314), .ZN(n7136) );
  NAND2_X1 U7580 ( .A1(n12127), .A2(n12124), .ZN(n7231) );
  OR2_X1 U7581 ( .A1(n12409), .A2(n15010), .ZN(n9015) );
  INV_X1 U7582 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7175) );
  AOI21_X1 U7583 ( .B1(n6889), .B2(n6887), .A(n6886), .ZN(n6885) );
  INV_X1 U7584 ( .A(n8690), .ZN(n6886) );
  INV_X1 U7585 ( .A(n6891), .ZN(n6887) );
  INV_X1 U7586 ( .A(n10655), .ZN(n6838) );
  AND2_X1 U7587 ( .A1(n9132), .A2(n7149), .ZN(n7148) );
  OR2_X1 U7588 ( .A1(n7151), .A2(n7150), .ZN(n7149) );
  OR2_X1 U7589 ( .A1(n11027), .A2(n10929), .ZN(n9002) );
  INV_X1 U7590 ( .A(SI_14_), .ZN(n8386) );
  NOR2_X1 U7591 ( .A1(n7087), .A2(n8241), .ZN(n7086) );
  INV_X1 U7592 ( .A(n8092), .ZN(n7087) );
  NAND2_X1 U7593 ( .A1(n9831), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8094) );
  AOI21_X1 U7594 ( .B1(n13466), .B2(n7922), .A(n7045), .ZN(n7044) );
  AOI21_X1 U7595 ( .B1(n7337), .B2(n9406), .A(n6558), .ZN(n7336) );
  OAI21_X1 U7596 ( .B1(n6448), .B2(n7038), .A(n8011), .ZN(n7037) );
  NOR2_X1 U7597 ( .A1(n13206), .A2(n7322), .ZN(n6766) );
  OR2_X1 U7598 ( .A1(n7696), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U7599 ( .A1(n11256), .A2(n7403), .ZN(n7406) );
  NOR2_X1 U7600 ( .A1(n11258), .A2(n7404), .ZN(n7403) );
  INV_X1 U7601 ( .A(n11255), .ZN(n7404) );
  INV_X1 U7602 ( .A(n11985), .ZN(n9673) );
  INV_X1 U7603 ( .A(n13946), .ZN(n6622) );
  NAND2_X1 U7604 ( .A1(n14153), .A2(n6983), .ZN(n6982) );
  INV_X1 U7605 ( .A(n13893), .ZN(n6983) );
  INV_X1 U7606 ( .A(n14021), .ZN(n7264) );
  INV_X1 U7607 ( .A(n14090), .ZN(n6870) );
  AND2_X1 U7608 ( .A1(n12078), .A2(n12200), .ZN(n6869) );
  OR2_X1 U7609 ( .A1(n14481), .A2(n11723), .ZN(n12073) );
  INV_X1 U7610 ( .A(n11068), .ZN(n6854) );
  INV_X1 U7611 ( .A(n10888), .ZN(n6855) );
  AOI21_X1 U7612 ( .B1(n12197), .B2(n6861), .A(n6514), .ZN(n6860) );
  INV_X1 U7613 ( .A(n11299), .ZN(n6861) );
  NAND2_X1 U7614 ( .A1(n6526), .A2(n10385), .ZN(n9495) );
  INV_X1 U7615 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9478) );
  INV_X1 U7616 ( .A(n7355), .ZN(n7354) );
  XNOR2_X1 U7617 ( .A(n8826), .B(n8825), .ZN(n8846) );
  AOI21_X1 U7618 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n8898), .A(n8897), .ZN(
        n8903) );
  NAND2_X1 U7619 ( .A1(n8142), .A2(n8141), .ZN(n12830) );
  INV_X1 U7620 ( .A(n12308), .ZN(n6604) );
  INV_X1 U7621 ( .A(n8605), .ZN(n8946) );
  INV_X1 U7622 ( .A(n8509), .ZN(n8605) );
  NAND2_X1 U7623 ( .A1(n6827), .A2(n6464), .ZN(n7118) );
  AOI21_X1 U7624 ( .B1(n7142), .B2(n7141), .A(n6467), .ZN(n7140) );
  INV_X1 U7625 ( .A(n8314), .ZN(n7141) );
  AND2_X1 U7626 ( .A1(n9002), .A2(n9001), .ZN(n11048) );
  NAND2_X1 U7627 ( .A1(n10290), .A2(n11832), .ZN(n8240) );
  AND2_X1 U7628 ( .A1(n8657), .A2(n6999), .ZN(n10109) );
  XNOR2_X1 U7629 ( .A(n8673), .B(P3_IR_REG_23__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U7630 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n6709), .ZN(n6708) );
  INV_X1 U7631 ( .A(n8598), .ZN(n8596) );
  NAND2_X1 U7632 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n7077), .ZN(n7076) );
  NAND2_X1 U7633 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n6707), .ZN(n6706) );
  AND2_X1 U7634 ( .A1(n9945), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8101) );
  AND2_X1 U7635 ( .A1(n8096), .A2(n8095), .ZN(n8256) );
  NOR2_X1 U7636 ( .A1(n10607), .A2(n7293), .ZN(n7292) );
  INV_X1 U7637 ( .A(n9522), .ZN(n7293) );
  AND2_X1 U7638 ( .A1(n11559), .A2(n6472), .ZN(n7283) );
  OAI21_X1 U7639 ( .B1(n9612), .B2(n6461), .A(n7295), .ZN(n7298) );
  NAND2_X1 U7640 ( .A1(n9613), .A2(n12998), .ZN(n7299) );
  NOR2_X1 U7641 ( .A1(n10374), .A2(n7271), .ZN(n7270) );
  INV_X1 U7642 ( .A(n7274), .ZN(n7271) );
  INV_X1 U7643 ( .A(n7314), .ZN(n9507) );
  INV_X1 U7644 ( .A(n13106), .ZN(n13223) );
  NAND2_X1 U7645 ( .A1(n11405), .A2(n11059), .ZN(n9627) );
  OR2_X1 U7646 ( .A1(n12247), .A2(n7552), .ZN(n7578) );
  NAND2_X1 U7647 ( .A1(n7548), .A2(n7552), .ZN(n7599) );
  INV_X1 U7648 ( .A(n13228), .ZN(n7325) );
  INV_X1 U7649 ( .A(n13256), .ZN(n13259) );
  NAND2_X1 U7650 ( .A1(n13275), .A2(n13274), .ZN(n13273) );
  NAND2_X1 U7651 ( .A1(n6748), .A2(n6747), .ZN(n7318) );
  AOI21_X1 U7652 ( .B1(n6750), .B2(n6752), .A(n13307), .ZN(n6747) );
  NAND2_X1 U7653 ( .A1(n8034), .A2(n9864), .ZN(n13404) );
  INV_X1 U7654 ( .A(n13352), .ZN(n13405) );
  NAND2_X1 U7655 ( .A1(n7123), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7853) );
  INV_X1 U7656 ( .A(n6824), .ZN(n6822) );
  OR2_X1 U7657 ( .A1(n11872), .A2(n13650), .ZN(n11887) );
  AOI21_X1 U7658 ( .B1(n7375), .B2(n7377), .A(n6474), .ZN(n7373) );
  AND2_X1 U7659 ( .A1(n11984), .A2(n7193), .ZN(n7192) );
  NAND2_X1 U7660 ( .A1(n7196), .A2(n7194), .ZN(n7193) );
  AND2_X1 U7661 ( .A1(n11785), .A2(n11784), .ZN(n13682) );
  CLKBUF_X3 U7662 ( .A(n9721), .Z(n9744) );
  XNOR2_X1 U7663 ( .A(n13926), .B(n13904), .ZN(n13920) );
  NOR2_X1 U7664 ( .A1(n11976), .A2(n14559), .ZN(n11971) );
  INV_X1 U7665 ( .A(n14575), .ZN(n14591) );
  NAND2_X1 U7666 ( .A1(n11745), .A2(n11744), .ZN(n14192) );
  INV_X1 U7667 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U7668 ( .A1(n7372), .A2(n7369), .ZN(n7852) );
  NAND2_X1 U7669 ( .A1(n7471), .A2(n7470), .ZN(n7754) );
  OAI21_X1 U7670 ( .B1(n14516), .B2(n6791), .A(n6469), .ZN(n8892) );
  INV_X1 U7671 ( .A(n6792), .ZN(n6791) );
  NAND2_X1 U7672 ( .A1(n6600), .A2(n6494), .ZN(n8918) );
  NAND2_X1 U7673 ( .A1(n8915), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n6600) );
  INV_X1 U7674 ( .A(n12581), .ZN(n12743) );
  AOI21_X1 U7675 ( .B1(n12503), .B2(n15081), .A(n12502), .ZN(n7170) );
  NAND2_X1 U7676 ( .A1(n7173), .A2(n7172), .ZN(n7171) );
  OR2_X1 U7677 ( .A1(n9184), .A2(n9185), .ZN(n6724) );
  NAND2_X1 U7678 ( .A1(n12036), .A2(n7218), .ZN(n7217) );
  INV_X1 U7679 ( .A(n12035), .ZN(n7218) );
  OR2_X1 U7680 ( .A1(n9205), .A2(n9206), .ZN(n6732) );
  NAND2_X1 U7681 ( .A1(n12049), .A2(n12047), .ZN(n7215) );
  INV_X1 U7682 ( .A(n9233), .ZN(n6745) );
  NAND2_X1 U7683 ( .A1(n7237), .A2(n12058), .ZN(n7236) );
  NAND2_X1 U7684 ( .A1(n12070), .A2(n7240), .ZN(n7239) );
  INV_X1 U7685 ( .A(n12069), .ZN(n7240) );
  NAND2_X1 U7686 ( .A1(n6734), .A2(n6738), .ZN(n9237) );
  AOI21_X1 U7687 ( .B1(n6738), .B2(n6737), .A(n6736), .ZN(n6735) );
  INV_X1 U7688 ( .A(n9236), .ZN(n6736) );
  INV_X1 U7689 ( .A(n6741), .ZN(n6737) );
  NAND2_X1 U7690 ( .A1(n6454), .A2(n6424), .ZN(n9298) );
  OAI21_X1 U7691 ( .B1(n7129), .B2(n7127), .A(n7128), .ZN(n7126) );
  NOR2_X1 U7692 ( .A1(n12101), .A2(n12100), .ZN(n7225) );
  NAND2_X1 U7693 ( .A1(n12098), .A2(n7226), .ZN(n7224) );
  AOI21_X1 U7694 ( .B1(n12101), .B2(n12100), .A(n7227), .ZN(n7226) );
  INV_X1 U7695 ( .A(n12097), .ZN(n7227) );
  OR2_X1 U7696 ( .A1(n12108), .A2(n12109), .ZN(n7210) );
  AND2_X1 U7697 ( .A1(n12109), .A2(n12108), .ZN(n7211) );
  OAI21_X1 U7698 ( .B1(n12110), .B2(n7211), .A(n7210), .ZN(n12112) );
  NAND2_X1 U7699 ( .A1(n7209), .A2(n12111), .ZN(n7208) );
  NAND2_X1 U7700 ( .A1(n7210), .A2(n7211), .ZN(n7209) );
  NOR2_X1 U7701 ( .A1(n9326), .A2(n9327), .ZN(n6729) );
  AOI22_X1 U7702 ( .A1(n13437), .A2(n9369), .B1(n9167), .B2(n13104), .ZN(n9372) );
  AOI21_X1 U7703 ( .B1(n7232), .B2(n7231), .A(n7229), .ZN(n7228) );
  NOR2_X1 U7704 ( .A1(n12127), .A2(n12124), .ZN(n7232) );
  AND2_X1 U7705 ( .A1(n6897), .A2(n6529), .ZN(n6895) );
  AOI21_X1 U7706 ( .B1(n6443), .B2(n6899), .A(n6898), .ZN(n6897) );
  INV_X1 U7707 ( .A(n7475), .ZN(n6898) );
  INV_X1 U7708 ( .A(n7470), .ZN(n6899) );
  INV_X1 U7709 ( .A(n6443), .ZN(n6900) );
  NOR2_X1 U7710 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7107) );
  NAND2_X1 U7711 ( .A1(n7999), .A2(n10594), .ZN(n6758) );
  INV_X1 U7712 ( .A(n7999), .ZN(n7025) );
  INV_X1 U7713 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7534) );
  NOR2_X1 U7714 ( .A1(n11985), .A2(n11971), .ZN(n9738) );
  INV_X1 U7715 ( .A(n6889), .ZN(n6888) );
  NAND2_X1 U7716 ( .A1(n7500), .A2(SI_21_), .ZN(n7503) );
  NOR2_X1 U7717 ( .A1(n7356), .A2(n7352), .ZN(n7351) );
  INV_X1 U7718 ( .A(n7482), .ZN(n7352) );
  INV_X1 U7719 ( .A(n12324), .ZN(n7014) );
  NAND2_X1 U7720 ( .A1(n8938), .A2(n7093), .ZN(n9113) );
  AND2_X1 U7721 ( .A1(n12396), .A2(n8937), .ZN(n7093) );
  AND2_X1 U7722 ( .A1(n7107), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10317) );
  NOR2_X1 U7723 ( .A1(n10498), .A2(n10331), .ZN(n6643) );
  INV_X1 U7724 ( .A(n14896), .ZN(n12446) );
  NOR2_X1 U7725 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6613) );
  OR2_X1 U7726 ( .A1(n12338), .A2(n12742), .ZN(n9071) );
  OR2_X1 U7727 ( .A1(n12364), .A2(n12792), .ZN(n9057) );
  INV_X1 U7728 ( .A(n12822), .ZN(n6911) );
  INV_X1 U7729 ( .A(n9054), .ZN(n6913) );
  OR2_X1 U7730 ( .A1(n12964), .A2(n12405), .ZN(n9041) );
  NAND2_X1 U7731 ( .A1(n15083), .A2(n12908), .ZN(n8972) );
  INV_X1 U7732 ( .A(n9653), .ZN(n6908) );
  AND2_X1 U7733 ( .A1(n9037), .A2(n9035), .ZN(n11677) );
  NAND2_X1 U7734 ( .A1(n11317), .A2(n8314), .ZN(n7144) );
  AND2_X1 U7735 ( .A1(n7144), .A2(n6456), .ZN(n11476) );
  NOR2_X1 U7736 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7166) );
  OAI21_X1 U7737 ( .B1(n8211), .B2(n8209), .A(n8090), .ZN(n8224) );
  INV_X1 U7738 ( .A(n13035), .ZN(n7282) );
  AOI21_X1 U7739 ( .B1(n13017), .B2(n13013), .A(n13014), .ZN(n13064) );
  INV_X1 U7740 ( .A(n7032), .ZN(n7031) );
  OAI21_X1 U7741 ( .B1(n7033), .B2(n9390), .A(n13206), .ZN(n7032) );
  INV_X1 U7742 ( .A(n7035), .ZN(n7027) );
  AOI21_X1 U7743 ( .B1(n7335), .B2(n7334), .A(n7760), .ZN(n7332) );
  NOR2_X1 U7744 ( .A1(n11360), .A2(n13119), .ZN(n7335) );
  NAND2_X1 U7745 ( .A1(n11360), .A2(n13119), .ZN(n7334) );
  NAND2_X1 U7746 ( .A1(n7984), .A2(n11405), .ZN(n9501) );
  OAI22_X1 U7747 ( .A1(n10706), .A2(n8000), .B1(n10752), .B2(n10766), .ZN(
        n10844) );
  INV_X1 U7748 ( .A(n10594), .ZN(n6759) );
  NAND2_X1 U7749 ( .A1(n7540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7539) );
  INV_X1 U7750 ( .A(n7822), .ZN(n7824) );
  NAND2_X1 U7751 ( .A1(n7743), .A2(n7755), .ZN(n7766) );
  INV_X1 U7752 ( .A(n11918), .ZN(n7397) );
  CLKBUF_X1 U7753 ( .A(n9738), .Z(n11652) );
  INV_X1 U7754 ( .A(n7198), .ZN(n7194) );
  INV_X1 U7755 ( .A(n11080), .ZN(n6972) );
  NAND2_X1 U7756 ( .A1(n6859), .A2(n6857), .ZN(n14096) );
  AND2_X1 U7757 ( .A1(n14112), .A2(n6858), .ZN(n6857) );
  NAND2_X1 U7758 ( .A1(n11534), .A2(n6860), .ZN(n6858) );
  INV_X1 U7759 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9477) );
  INV_X1 U7760 ( .A(n7836), .ZN(n7370) );
  OR2_X1 U7761 ( .A1(n10183), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U7762 ( .A1(n8832), .A2(n8833), .ZN(n8874) );
  AOI21_X1 U7763 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n8835), .A(n8834), .ZN(
        n8845) );
  NOR2_X1 U7764 ( .A1(n8874), .A2(n8873), .ZN(n8834) );
  AOI21_X1 U7765 ( .B1(n8763), .B2(n6994), .A(n6993), .ZN(n6992) );
  INV_X1 U7766 ( .A(n12346), .ZN(n6993) );
  INV_X1 U7767 ( .A(n8761), .ZN(n6994) );
  INV_X1 U7768 ( .A(n8763), .ZN(n6995) );
  NAND2_X1 U7769 ( .A1(n6402), .A2(n8974), .ZN(n8727) );
  NAND2_X1 U7770 ( .A1(n15086), .A2(n6603), .ZN(n6602) );
  INV_X1 U7771 ( .A(n6401), .ZN(n6603) );
  NAND2_X1 U7772 ( .A1(n8725), .A2(n9446), .ZN(n8726) );
  NAND2_X1 U7773 ( .A1(n6996), .A2(n8724), .ZN(n8725) );
  NOR2_X1 U7774 ( .A1(n12332), .A2(n7017), .ZN(n7016) );
  INV_X1 U7775 ( .A(n8775), .ZN(n7017) );
  NAND2_X1 U7776 ( .A1(n7007), .A2(n8737), .ZN(n7010) );
  AND2_X1 U7777 ( .A1(n8949), .A2(n8948), .ZN(n14394) );
  NAND2_X1 U7778 ( .A1(n7119), .A2(n7122), .ZN(n7121) );
  NAND2_X1 U7779 ( .A1(n10329), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7122) );
  NOR2_X1 U7780 ( .A1(n6425), .A2(n10499), .ZN(n10493) );
  NAND2_X1 U7781 ( .A1(n6843), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6842) );
  NAND2_X1 U7782 ( .A1(n6425), .A2(n10499), .ZN(n6843) );
  NAND2_X1 U7783 ( .A1(n6840), .A2(n6426), .ZN(n6839) );
  INV_X1 U7784 ( .A(n12427), .ZN(n6837) );
  NOR2_X1 U7785 ( .A1(n14906), .A2(n7112), .ZN(n12431) );
  AND2_X1 U7786 ( .A1(n14914), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7112) );
  NAND2_X1 U7787 ( .A1(n7116), .A2(n6566), .ZN(n6828) );
  OR2_X1 U7788 ( .A1(n7116), .A2(n12461), .ZN(n6829) );
  NAND2_X1 U7789 ( .A1(n14949), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7115) );
  NAND2_X1 U7790 ( .A1(n7118), .A2(n7117), .ZN(n7116) );
  INV_X1 U7791 ( .A(n14942), .ZN(n7117) );
  OR2_X1 U7792 ( .A1(n14979), .A2(n14978), .ZN(n7106) );
  NAND2_X1 U7793 ( .A1(n7106), .A2(n12466), .ZN(n12434) );
  OR2_X1 U7794 ( .A1(n14325), .A2(n14326), .ZN(n6835) );
  NAND2_X1 U7795 ( .A1(n6834), .A2(n6833), .ZN(n7111) );
  INV_X1 U7796 ( .A(n14342), .ZN(n6833) );
  NAND2_X1 U7797 ( .A1(n7111), .A2(n7110), .ZN(n7109) );
  NAND2_X1 U7798 ( .A1(n14349), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7110) );
  AOI22_X1 U7799 ( .A1(n12532), .A2(n8584), .B1(n12550), .B2(n12380), .ZN(
        n12519) );
  AOI21_X1 U7800 ( .B1(n7148), .B2(n7150), .A(n6482), .ZN(n7146) );
  NAND2_X1 U7801 ( .A1(n12789), .A2(n12790), .ZN(n7162) );
  AND2_X1 U7802 ( .A1(n9057), .A2(n9063), .ZN(n12782) );
  INV_X1 U7803 ( .A(n12793), .ZN(n12790) );
  INV_X1 U7804 ( .A(n12401), .ZN(n12808) );
  AND2_X1 U7805 ( .A1(n9048), .A2(n9052), .ZN(n12822) );
  NAND2_X1 U7806 ( .A1(n12823), .A2(n12822), .ZN(n12821) );
  AOI21_X1 U7807 ( .B1(n7155), .B2(n7154), .A(n6508), .ZN(n7153) );
  INV_X1 U7808 ( .A(n7158), .ZN(n7154) );
  OR2_X1 U7809 ( .A1(n11461), .A2(n11499), .ZN(n11508) );
  AND2_X1 U7810 ( .A1(n9011), .A2(n8279), .ZN(n7164) );
  NAND2_X1 U7811 ( .A1(n15025), .A2(n7163), .ZN(n11051) );
  AND2_X1 U7812 ( .A1(n8263), .A2(n8248), .ZN(n7163) );
  AND2_X1 U7813 ( .A1(n10286), .A2(n14410), .ZN(n10631) );
  AND2_X1 U7814 ( .A1(n8808), .A2(n9078), .ZN(n15081) );
  INV_X1 U7815 ( .A(n9122), .ZN(n12905) );
  NAND2_X1 U7816 ( .A1(n6908), .A2(n6906), .ZN(n12900) );
  NAND2_X1 U7817 ( .A1(n8406), .A2(n8405), .ZN(n12384) );
  INV_X1 U7818 ( .A(n14914), .ZN(n12451) );
  AND2_X1 U7819 ( .A1(n9497), .A2(n12967), .ZN(n10286) );
  AND2_X1 U7820 ( .A1(n9442), .A2(n9440), .ZN(n8811) );
  INV_X1 U7821 ( .A(n12967), .ZN(n10108) );
  NAND2_X1 U7822 ( .A1(n6999), .A2(n6998), .ZN(n6997) );
  NOR2_X1 U7823 ( .A1(n12990), .A2(P3_D_REG_0__SCAN_IN), .ZN(n6998) );
  INV_X1 U7824 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U7825 ( .A1(n8598), .A2(n7000), .ZN(n8649) );
  AND2_X1 U7826 ( .A1(n6549), .A2(n8597), .ZN(n7000) );
  INV_X1 U7827 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7001) );
  XNOR2_X1 U7828 ( .A(n8119), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U7829 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n8085), .ZN(n6607) );
  NAND2_X1 U7830 ( .A1(n8518), .A2(n8516), .ZN(n6608) );
  NAND2_X1 U7831 ( .A1(n8598), .A2(n8597), .ZN(n8646) );
  INV_X1 U7832 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8129) );
  INV_X1 U7833 ( .A(n7006), .ZN(n7004) );
  NAND2_X1 U7834 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n6632), .ZN(n6631) );
  INV_X1 U7835 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U7836 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n6650), .ZN(n6649) );
  INV_X1 U7837 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8102) );
  XNOR2_X1 U7838 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8324) );
  OR2_X1 U7839 ( .A1(n8310), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8343) );
  AND2_X1 U7840 ( .A1(n9860), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8099) );
  INV_X1 U7841 ( .A(n8094), .ZN(n7084) );
  INV_X1 U7842 ( .A(n7086), .ZN(n7085) );
  INV_X1 U7843 ( .A(n6576), .ZN(n7090) );
  INV_X1 U7844 ( .A(n8223), .ZN(n7089) );
  CLKBUF_X1 U7845 ( .A(n8224), .Z(n6576) );
  INV_X1 U7846 ( .A(n9560), .ZN(n7285) );
  INV_X1 U7847 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8118) );
  INV_X1 U7848 ( .A(n7313), .ZN(n7311) );
  INV_X1 U7849 ( .A(n13091), .ZN(n7308) );
  NOR2_X1 U7850 ( .A1(n7288), .A2(n7291), .ZN(n7287) );
  INV_X1 U7851 ( .A(n10761), .ZN(n7291) );
  INV_X1 U7852 ( .A(n9527), .ZN(n7290) );
  NAND2_X1 U7853 ( .A1(n6691), .A2(n6690), .ZN(n10747) );
  INV_X1 U7854 ( .A(n10749), .ZN(n6690) );
  INV_X1 U7855 ( .A(n10750), .ZN(n6691) );
  NAND2_X1 U7856 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  INV_X1 U7857 ( .A(n9642), .ZN(n7297) );
  NAND2_X1 U7859 ( .A1(n6644), .A2(n13063), .ZN(n13062) );
  NAND2_X1 U7860 ( .A1(n11341), .A2(n11342), .ZN(n11340) );
  XNOR2_X1 U7861 ( .A(n13026), .B(n10266), .ZN(n7314) );
  XNOR2_X1 U7862 ( .A(n13026), .B(n10238), .ZN(n9503) );
  INV_X1 U7863 ( .A(n13517), .ZN(n6950) );
  AND2_X1 U7864 ( .A1(n8694), .A2(n8693), .ZN(n9364) );
  INV_X1 U7865 ( .A(n6766), .ZN(n6765) );
  INV_X1 U7866 ( .A(n7324), .ZN(n6764) );
  OAI22_X1 U7867 ( .A1(n13237), .A2(n7936), .B1(n13526), .B2(n13258), .ZN(
        n13228) );
  NOR2_X2 U7868 ( .A1(n13244), .A2(n13229), .ZN(n13232) );
  NAND2_X1 U7869 ( .A1(n13572), .A2(n7626), .ZN(n7567) );
  INV_X1 U7870 ( .A(n7923), .ZN(n7331) );
  NAND2_X1 U7871 ( .A1(n7044), .A2(n7041), .ZN(n7040) );
  AOI21_X1 U7872 ( .B1(n7044), .B2(n6422), .A(n6524), .ZN(n7043) );
  NOR2_X2 U7873 ( .A1(n13301), .A2(n13466), .ZN(n13279) );
  AND2_X1 U7874 ( .A1(n7046), .A2(n6458), .ZN(n13294) );
  NOR2_X1 U7875 ( .A1(n13293), .A2(n7317), .ZN(n7316) );
  INV_X1 U7876 ( .A(n7892), .ZN(n7317) );
  INV_X1 U7877 ( .A(n6754), .ZN(n6753) );
  OAI21_X1 U7878 ( .B1(n9410), .B2(n6755), .A(n6495), .ZN(n6754) );
  OAI21_X1 U7879 ( .B1(n13385), .B2(n7049), .A(n7047), .ZN(n13330) );
  INV_X1 U7880 ( .A(n7051), .ZN(n7049) );
  AOI21_X1 U7881 ( .B1(n7051), .B2(n7048), .A(n6503), .ZN(n7047) );
  NOR2_X1 U7882 ( .A1(n7053), .A2(n8023), .ZN(n7051) );
  OAI21_X1 U7883 ( .B1(n11491), .B2(n6523), .A(n6779), .ZN(n13390) );
  AND2_X1 U7884 ( .A1(n7336), .A2(n6541), .ZN(n6779) );
  OAI21_X1 U7885 ( .B1(n11483), .B2(n7058), .A(n7057), .ZN(n13402) );
  AOI21_X1 U7886 ( .B1(n7059), .B2(n9405), .A(n6504), .ZN(n7057) );
  INV_X1 U7887 ( .A(n7059), .ZN(n7058) );
  NAND2_X1 U7888 ( .A1(n11482), .A2(n8015), .ZN(n11588) );
  AND2_X1 U7889 ( .A1(n9406), .A2(n8015), .ZN(n7059) );
  AND2_X1 U7890 ( .A1(n14434), .A2(n7781), .ZN(n11593) );
  NAND2_X1 U7891 ( .A1(n11593), .A2(n7799), .ZN(n11592) );
  NAND2_X1 U7892 ( .A1(n11483), .A2(n6780), .ZN(n11482) );
  OAI21_X1 U7893 ( .B1(n8008), .B2(n7038), .A(n7036), .ZN(n8013) );
  INV_X1 U7894 ( .A(n7037), .ZN(n7036) );
  NAND2_X1 U7895 ( .A1(n6945), .A2(n6944), .ZN(n11239) );
  NAND2_X1 U7896 ( .A1(n10842), .A2(n7689), .ZN(n10828) );
  NAND2_X1 U7897 ( .A1(n10703), .A2(n7326), .ZN(n10842) );
  AND2_X1 U7898 ( .A1(n9400), .A2(n7676), .ZN(n7326) );
  NAND2_X1 U7899 ( .A1(n6746), .A2(n7320), .ZN(n10704) );
  AOI21_X1 U7900 ( .B1(n7321), .B2(n10665), .A(n6502), .ZN(n7320) );
  NAND2_X1 U7901 ( .A1(n10593), .A2(n7319), .ZN(n6746) );
  INV_X1 U7902 ( .A(n9398), .ZN(n10705) );
  NAND2_X1 U7903 ( .A1(n10704), .A2(n10705), .ZN(n10703) );
  INV_X1 U7904 ( .A(n9396), .ZN(n10665) );
  NAND2_X1 U7905 ( .A1(n10593), .A2(n10594), .ZN(n10592) );
  INV_X1 U7906 ( .A(n10238), .ZN(n7587) );
  NAND2_X1 U7907 ( .A1(n7589), .A2(n7020), .ZN(n7021) );
  AND2_X1 U7908 ( .A1(n9812), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7020) );
  INV_X1 U7909 ( .A(n8713), .ZN(n7064) );
  AND2_X1 U7910 ( .A1(n6767), .A2(n7323), .ZN(n13211) );
  NAND2_X1 U7911 ( .A1(n6767), .A2(n6766), .ZN(n13441) );
  OAI21_X1 U7912 ( .B1(n6663), .B2(n13405), .A(n6660), .ZN(n13448) );
  AND2_X1 U7913 ( .A1(n6662), .A2(n6661), .ZN(n6660) );
  OR2_X1 U7914 ( .A1(n13258), .A2(n13404), .ZN(n6661) );
  NAND2_X1 U7915 ( .A1(n7884), .A2(n7883), .ZN(n13319) );
  NAND2_X1 U7916 ( .A1(n7870), .A2(n7869), .ZN(n13337) );
  AND2_X1 U7917 ( .A1(n10254), .A2(n13355), .ZN(n14428) );
  NOR2_X1 U7918 ( .A1(n7977), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U7919 ( .A1(n7824), .A2(n7823), .ZN(n7840) );
  AND2_X1 U7920 ( .A1(n7697), .A2(n7729), .ZN(n9984) );
  AND2_X1 U7921 ( .A1(n11728), .A2(n6808), .ZN(n6807) );
  NAND2_X1 U7922 ( .A1(n13662), .A2(n6809), .ZN(n6808) );
  INV_X1 U7923 ( .A(n11714), .ZN(n6809) );
  INV_X1 U7924 ( .A(n13662), .ZN(n6810) );
  INV_X1 U7925 ( .A(n7410), .ZN(n7384) );
  INV_X1 U7926 ( .A(n7396), .ZN(n7395) );
  OAI21_X1 U7927 ( .B1(n13699), .B2(n7397), .A(n12231), .ZN(n7396) );
  NAND2_X1 U7928 ( .A1(n13655), .A2(n6493), .ZN(n13609) );
  NAND2_X1 U7929 ( .A1(n13627), .A2(n11741), .ZN(n13638) );
  NAND2_X1 U7930 ( .A1(n7401), .A2(n9733), .ZN(n10269) );
  NAND2_X1 U7931 ( .A1(n11139), .A2(n11928), .ZN(n7401) );
  AOI21_X1 U7932 ( .B1(n6622), .B2(n7357), .A(n6512), .ZN(n7360) );
  INV_X1 U7933 ( .A(n13878), .ZN(n7357) );
  NAND2_X1 U7934 ( .A1(n13978), .A2(n6980), .ZN(n7359) );
  NOR2_X1 U7935 ( .A1(n6447), .A2(n6981), .ZN(n6980) );
  INV_X1 U7936 ( .A(n6982), .ZN(n6981) );
  AND2_X1 U7937 ( .A1(n7359), .A2(n7358), .ZN(n13940) );
  AND2_X1 U7938 ( .A1(n7360), .A2(n13931), .ZN(n7358) );
  NAND2_X1 U7939 ( .A1(n13960), .A2(n6484), .ZN(n13947) );
  AND2_X1 U7940 ( .A1(n11905), .A2(n11888), .ZN(n13965) );
  XNOR2_X1 U7941 ( .A(n13983), .B(n13893), .ZN(n13973) );
  AOI21_X1 U7942 ( .B1(n13890), .B2(n14001), .A(n6490), .ZN(n13996) );
  NAND2_X1 U7943 ( .A1(n7264), .A2(n6455), .ZN(n7261) );
  NOR2_X1 U7944 ( .A1(n7262), .A2(n6874), .ZN(n6872) );
  NAND2_X1 U7945 ( .A1(n7264), .A2(n7263), .ZN(n7262) );
  INV_X1 U7946 ( .A(n14041), .ZN(n7263) );
  AOI21_X1 U7947 ( .B1(n14048), .B2(n13873), .A(n13872), .ZN(n14042) );
  NAND2_X1 U7948 ( .A1(n14049), .A2(n6873), .ZN(n14033) );
  NOR2_X1 U7949 ( .A1(n14033), .A2(n14041), .ZN(n14032) );
  NOR2_X1 U7950 ( .A1(n14084), .A2(n14192), .ZN(n6937) );
  OAI21_X1 U7951 ( .B1(n11685), .B2(n6867), .A(n6864), .ZN(n7259) );
  AOI21_X1 U7952 ( .B1(n6866), .B2(n6865), .A(n6465), .ZN(n6864) );
  INV_X1 U7953 ( .A(n6869), .ZN(n6865) );
  AND2_X1 U7954 ( .A1(n7259), .A2(n13885), .ZN(n14065) );
  NAND2_X1 U7955 ( .A1(n11685), .A2(n6869), .ZN(n6868) );
  AND2_X1 U7956 ( .A1(n13867), .A2(n13869), .ZN(n14090) );
  NAND2_X1 U7957 ( .A1(n11699), .A2(n13881), .ZN(n14084) );
  AND4_X1 U7958 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n14099) );
  INV_X1 U7959 ( .A(n14112), .ZN(n11538) );
  AND2_X1 U7960 ( .A1(n12073), .A2(n12072), .ZN(n14112) );
  NAND2_X1 U7961 ( .A1(n11283), .A2(n11282), .ZN(n11535) );
  NAND2_X1 U7962 ( .A1(n14300), .A2(n14299), .ZN(n14298) );
  NAND2_X1 U7963 ( .A1(n11206), .A2(n11183), .ZN(n11208) );
  AND2_X1 U7964 ( .A1(n12191), .A2(n11099), .ZN(n7260) );
  NAND2_X1 U7965 ( .A1(n6973), .A2(n6974), .ZN(n14567) );
  OR2_X1 U7966 ( .A1(n14641), .A2(n10874), .ZN(n10875) );
  AOI21_X1 U7967 ( .B1(n10891), .B2(n6855), .A(n6854), .ZN(n6850) );
  NAND2_X1 U7968 ( .A1(n6852), .A2(n6851), .ZN(n14564) );
  NAND2_X1 U7969 ( .A1(n10889), .A2(n6853), .ZN(n6852) );
  NOR2_X1 U7970 ( .A1(n6855), .A2(n6854), .ZN(n6853) );
  NAND2_X1 U7971 ( .A1(n10889), .A2(n10888), .ZN(n10890) );
  INV_X1 U7972 ( .A(n14634), .ZN(n7265) );
  XNOR2_X1 U7973 ( .A(n13731), .B(n10885), .ZN(n12003) );
  NAND2_X1 U7974 ( .A1(n10862), .A2(n11977), .ZN(n14575) );
  NAND2_X1 U7975 ( .A1(n11139), .A2(n10411), .ZN(n11134) );
  NAND2_X1 U7976 ( .A1(n14126), .A2(n14652), .ZN(n6939) );
  INV_X1 U7977 ( .A(n14131), .ZN(n6594) );
  AND2_X1 U7978 ( .A1(n10862), .A2(n9781), .ZN(n14652) );
  AND2_X1 U7979 ( .A1(n14568), .A2(n14656), .ZN(n14644) );
  INV_X1 U7980 ( .A(n14625), .ZN(n14635) );
  NAND2_X1 U7981 ( .A1(n9357), .A2(n9347), .ZN(n6880) );
  NAND2_X1 U7982 ( .A1(n14228), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9678) );
  AND2_X1 U7983 ( .A1(n8692), .A2(n7960), .ZN(n8690) );
  NOR2_X1 U7984 ( .A1(n7956), .A2(n6892), .ZN(n6891) );
  INV_X1 U7985 ( .A(n7939), .ZN(n6892) );
  AOI21_X1 U7986 ( .B1(n6891), .B2(n6564), .A(n6890), .ZN(n6889) );
  INV_X1 U7987 ( .A(n7955), .ZN(n6890) );
  XNOR2_X1 U7988 ( .A(n7927), .B(n7926), .ZN(n13568) );
  NAND2_X1 U7989 ( .A1(n7925), .A2(n7924), .ZN(n7927) );
  XNOR2_X1 U7990 ( .A(n9496), .B(P1_IR_REG_23__SCAN_IN), .ZN(n9937) );
  MUX2_X1 U7991 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9674), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n9675) );
  INV_X1 U7992 ( .A(n7865), .ZN(n7498) );
  NAND2_X1 U7993 ( .A1(n7363), .A2(n7499), .ZN(n7866) );
  OR2_X1 U7994 ( .A1(n6473), .A2(n9669), .ZN(n9670) );
  AND2_X1 U7995 ( .A1(n9668), .A2(n9475), .ZN(n9669) );
  INV_X1 U7996 ( .A(n7369), .ZN(n7368) );
  INV_X1 U7997 ( .A(n7353), .ZN(n7816) );
  AOI21_X1 U7998 ( .B1(n7801), .B2(n7415), .A(n7356), .ZN(n7353) );
  NOR2_X1 U7999 ( .A1(n9940), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n10104) );
  NAND2_X1 U8000 ( .A1(n7345), .A2(n7456), .ZN(n7691) );
  NAND2_X1 U8001 ( .A1(n7678), .A2(n7454), .ZN(n7345) );
  XNOR2_X1 U8002 ( .A(n7678), .B(n7677), .ZN(n11081) );
  INV_X1 U8003 ( .A(n6967), .ZN(n8827) );
  AOI21_X1 U8004 ( .B1(n8880), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n8837), .ZN(
        n8885) );
  AOI21_X1 U8005 ( .B1(n6599), .B2(n6598), .A(n6597), .ZN(n8842) );
  AND2_X1 U8006 ( .A1(n8839), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n6597) );
  INV_X1 U8007 ( .A(n8888), .ZN(n6598) );
  INV_X1 U8008 ( .A(n8889), .ZN(n6599) );
  INV_X1 U8009 ( .A(n6964), .ZN(n8890) );
  NAND2_X1 U8010 ( .A1(n8911), .A2(n14811), .ZN(n8912) );
  AOI22_X1 U8011 ( .A1(n12295), .A2(n12294), .B1(n12536), .B2(n12293), .ZN(
        n12298) );
  NAND2_X1 U8012 ( .A1(n8505), .A2(n8504), .ZN(n12746) );
  NAND2_X1 U8013 ( .A1(n8452), .A2(n8451), .ZN(n12795) );
  AND3_X1 U8014 ( .A1(n8512), .A2(n8511), .A3(n8510), .ZN(n12754) );
  NAND2_X1 U8015 ( .A1(n8520), .A2(n8519), .ZN(n12734) );
  AND3_X1 U8016 ( .A1(n8486), .A2(n8485), .A3(n8484), .ZN(n12781) );
  AND3_X1 U8017 ( .A1(n8262), .A2(n8261), .A3(n8260), .ZN(n10929) );
  INV_X1 U8018 ( .A(n12395), .ZN(n14859) );
  INV_X1 U8019 ( .A(n14861), .ZN(n12382) );
  AND2_X1 U8020 ( .A1(n9144), .A2(n8724), .ZN(n7071) );
  NAND2_X1 U8021 ( .A1(n8528), .A2(n8527), .ZN(n12581) );
  AND2_X1 U8022 ( .A1(n14984), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U8023 ( .A1(n14867), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14866) );
  INV_X1 U8024 ( .A(n10329), .ZN(n10351) );
  NOR2_X1 U8025 ( .A1(n14376), .A2(n12440), .ZN(n6642) );
  AND2_X1 U8026 ( .A1(n10300), .A2(n10293), .ZN(n14385) );
  XNOR2_X1 U8027 ( .A(n6626), .B(n6569), .ZN(n12490) );
  NAND2_X1 U8028 ( .A1(n14377), .A2(n6627), .ZN(n6626) );
  OR2_X1 U8029 ( .A1(n14376), .A2(n12875), .ZN(n6627) );
  NOR2_X1 U8030 ( .A1(n8614), .A2(n8613), .ZN(n8615) );
  AND2_X1 U8031 ( .A1(n8348), .A2(n8347), .ZN(n14413) );
  NAND2_X1 U8032 ( .A1(n15159), .A2(n14410), .ZN(n12899) );
  NAND2_X1 U8033 ( .A1(n12832), .A2(n12833), .ZN(n12911) );
  AND2_X1 U8034 ( .A1(n12994), .A2(n12990), .ZN(n8659) );
  NAND2_X1 U8035 ( .A1(n7097), .A2(n6568), .ZN(n8931) );
  NAND2_X1 U8036 ( .A1(n7104), .A2(n6437), .ZN(n7097) );
  NAND2_X1 U8037 ( .A1(n7857), .A2(n7856), .ZN(n13360) );
  INV_X1 U8038 ( .A(n9510), .ZN(n7273) );
  INV_X1 U8039 ( .A(n9511), .ZN(n7275) );
  INV_X1 U8040 ( .A(n9512), .ZN(n7276) );
  INV_X1 U8041 ( .A(n13108), .ZN(n13258) );
  NAND2_X1 U8042 ( .A1(n9623), .A2(n9622), .ZN(n13088) );
  NAND4_X1 U8043 ( .A1(n7604), .A2(n7603), .A3(n7602), .A4(n7601), .ZN(n9166)
         );
  NAND2_X1 U8044 ( .A1(n7875), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7579) );
  CLKBUF_X1 U8045 ( .A(n9157), .Z(n13131) );
  OR2_X1 U8046 ( .A1(n7743), .A2(n7980), .ZN(n7744) );
  INV_X1 U8047 ( .A(n7063), .ZN(n7062) );
  OAI21_X1 U8048 ( .B1(n7064), .B2(n13352), .A(n13427), .ZN(n7063) );
  INV_X1 U8049 ( .A(n7030), .ZN(n13207) );
  AOI21_X1 U8050 ( .B1(n13238), .B2(n9390), .A(n7033), .ZN(n7030) );
  AND2_X1 U8051 ( .A1(n13273), .A2(n7330), .ZN(n13459) );
  NAND2_X1 U8052 ( .A1(n13273), .A2(n7923), .ZN(n13260) );
  INV_X1 U8053 ( .A(n13229), .ZN(n13522) );
  INV_X1 U8054 ( .A(n9423), .ZN(n11405) );
  NAND2_X1 U8055 ( .A1(n7399), .A2(n11771), .ZN(n13602) );
  NAND2_X1 U8056 ( .A1(n6822), .A2(n7378), .ZN(n6821) );
  INV_X1 U8057 ( .A(n7378), .ZN(n6823) );
  NAND2_X1 U8058 ( .A1(n13603), .A2(n11793), .ZN(n13657) );
  OR2_X1 U8059 ( .A1(n12177), .A2(n7190), .ZN(n7189) );
  NAND2_X1 U8060 ( .A1(n11862), .A2(n11861), .ZN(n13876) );
  NAND2_X1 U8061 ( .A1(n11825), .A2(n11824), .ZN(n13874) );
  OR2_X1 U8062 ( .A1(n12167), .A2(n10016), .ZN(n9711) );
  OR2_X1 U8063 ( .A1(n11178), .A2(n9707), .ZN(n9708) );
  INV_X1 U8064 ( .A(n13859), .ZN(n14121) );
  NAND2_X1 U8065 ( .A1(n13926), .A2(n13897), .ZN(n6667) );
  NAND2_X1 U8066 ( .A1(n11289), .A2(n11288), .ZN(n12068) );
  NAND2_X1 U8067 ( .A1(n6578), .A2(n6577), .ZN(n9692) );
  NAND2_X1 U8068 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9676), .ZN(n6577) );
  NAND2_X1 U8069 ( .A1(n6784), .A2(n8853), .ZN(n14260) );
  AOI21_X1 U8070 ( .B1(n8821), .B2(n6957), .A(n8820), .ZN(n8848) );
  NOR2_X1 U8071 ( .A1(n14260), .A2(n14259), .ZN(n14258) );
  NAND2_X1 U8072 ( .A1(n6620), .A2(n6619), .ZN(n6795) );
  INV_X1 U8073 ( .A(n14510), .ZN(n6619) );
  INV_X1 U8074 ( .A(n14511), .ZN(n6620) );
  INV_X1 U8075 ( .A(n8900), .ZN(n6789) );
  AND2_X1 U8076 ( .A1(n8901), .A2(n8900), .ZN(n14523) );
  OR2_X1 U8077 ( .A1(n8912), .A2(n8916), .ZN(n6960) );
  XNOR2_X1 U8078 ( .A(n8922), .B(n12642), .ZN(n7414) );
  INV_X1 U8079 ( .A(n10870), .ZN(n11994) );
  OR2_X1 U8080 ( .A1(n9174), .A2(n9173), .ZN(n9181) );
  OR2_X1 U8081 ( .A1(n9165), .A2(n9164), .ZN(n9172) );
  NAND2_X1 U8082 ( .A1(n7139), .A2(n7138), .ZN(n9197) );
  OR2_X1 U8083 ( .A1(n9188), .A2(n9189), .ZN(n7138) );
  NOR2_X1 U8084 ( .A1(n6429), .A2(n6520), .ZN(n6723) );
  NAND2_X1 U8085 ( .A1(n7220), .A2(n12035), .ZN(n7219) );
  NAND2_X1 U8086 ( .A1(n12048), .A2(n7214), .ZN(n7213) );
  INV_X1 U8087 ( .A(n12047), .ZN(n7214) );
  NAND2_X1 U8088 ( .A1(n6731), .A2(n6730), .ZN(n9216) );
  AOI21_X1 U8089 ( .B1(n6417), .B2(n6733), .A(n6431), .ZN(n6730) );
  AND2_X1 U8090 ( .A1(n9205), .A2(n9206), .ZN(n6733) );
  NAND2_X1 U8091 ( .A1(n12059), .A2(n7235), .ZN(n7234) );
  INV_X1 U8092 ( .A(n12058), .ZN(n7235) );
  INV_X1 U8093 ( .A(n9229), .ZN(n7134) );
  NAND2_X1 U8094 ( .A1(n6449), .A2(n7134), .ZN(n7132) );
  NOR2_X1 U8095 ( .A1(n6450), .A2(n6745), .ZN(n6744) );
  NOR2_X1 U8096 ( .A1(n6744), .A2(n6742), .ZN(n6741) );
  INV_X1 U8097 ( .A(n7132), .ZN(n6742) );
  NAND2_X1 U8098 ( .A1(n7242), .A2(n12069), .ZN(n7241) );
  NOR2_X1 U8099 ( .A1(n9282), .A2(n7131), .ZN(n7130) );
  AND2_X1 U8100 ( .A1(n9288), .A2(n9287), .ZN(n7131) );
  OR2_X1 U8101 ( .A1(n9237), .A2(n9236), .ZN(n9258) );
  NAND2_X1 U8102 ( .A1(n6525), .A2(n7182), .ZN(n7179) );
  INV_X1 U8103 ( .A(n12080), .ZN(n7180) );
  INV_X1 U8104 ( .A(n12083), .ZN(n7183) );
  NOR2_X1 U8105 ( .A1(n9287), .A2(n9288), .ZN(n7129) );
  INV_X1 U8106 ( .A(n9292), .ZN(n7127) );
  INV_X1 U8107 ( .A(n9291), .ZN(n7128) );
  INV_X1 U8108 ( .A(n7225), .ZN(n7221) );
  NOR2_X1 U8109 ( .A1(n7225), .A2(n7223), .ZN(n7222) );
  NAND2_X1 U8110 ( .A1(n6721), .A2(n6434), .ZN(n6718) );
  OR2_X1 U8111 ( .A1(n12112), .A2(n12111), .ZN(n12115) );
  AND2_X1 U8112 ( .A1(n6637), .A2(n6636), .ZN(n6635) );
  NAND2_X1 U8113 ( .A1(n9101), .A2(n9078), .ZN(n6637) );
  NAND2_X1 U8114 ( .A1(n9102), .A2(n9450), .ZN(n6636) );
  AND2_X1 U8115 ( .A1(n11968), .A2(n11967), .ZN(n12171) );
  NAND2_X1 U8116 ( .A1(n12171), .A2(n11969), .ZN(n12163) );
  OR2_X1 U8117 ( .A1(n8433), .A2(n12804), .ZN(n8435) );
  NAND2_X1 U8118 ( .A1(n9327), .A2(n9326), .ZN(n6728) );
  NAND2_X1 U8119 ( .A1(n9372), .A2(n9373), .ZN(n6665) );
  NOR2_X1 U8120 ( .A1(n9371), .A2(n9370), .ZN(n7135) );
  NAND2_X1 U8121 ( .A1(n9385), .A2(n6704), .ZN(n6674) );
  INV_X1 U8122 ( .A(n11234), .ZN(n7039) );
  AND2_X1 U8123 ( .A1(n7229), .A2(n7231), .ZN(n6616) );
  NOR2_X1 U8124 ( .A1(n7203), .A2(n7202), .ZN(n7201) );
  INV_X1 U8125 ( .A(n12176), .ZN(n7202) );
  INV_X1 U8126 ( .A(n12175), .ZN(n7203) );
  NOR2_X1 U8127 ( .A1(n9486), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n7408) );
  OAI21_X1 U8128 ( .B1(n7415), .B2(n7356), .A(n7489), .ZN(n7355) );
  AOI21_X1 U8129 ( .B1(n6895), .B2(n6900), .A(n6521), .ZN(n6893) );
  NAND2_X1 U8130 ( .A1(n7484), .A2(n8423), .ZN(n7487) );
  NAND2_X1 U8131 ( .A1(n7472), .A2(n14276), .ZN(n7475) );
  INV_X1 U8132 ( .A(n7456), .ZN(n7344) );
  NAND2_X1 U8133 ( .A1(n9828), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n6668) );
  NOR2_X1 U8134 ( .A1(n7647), .A2(n7632), .ZN(n7346) );
  INV_X1 U8135 ( .A(n7447), .ZN(n7348) );
  AND2_X1 U8136 ( .A1(n7107), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10327) );
  OR2_X1 U8137 ( .A1(n12413), .A2(n6628), .ZN(n12415) );
  NOR2_X1 U8138 ( .A1(n12414), .A2(n15155), .ZN(n6628) );
  OAI21_X1 U8139 ( .B1(n12451), .B2(n12417), .A(n14909), .ZN(n12418) );
  OAI21_X1 U8140 ( .B1(n12433), .B2(n12420), .A(n14944), .ZN(n12421) );
  NOR2_X1 U8141 ( .A1(n12501), .A2(n12504), .ZN(n12500) );
  AND2_X1 U8142 ( .A1(n8957), .A2(n8641), .ZN(n9134) );
  INV_X1 U8143 ( .A(n8529), .ZN(n7150) );
  NOR2_X1 U8144 ( .A1(n8530), .A2(n7152), .ZN(n7151) );
  INV_X1 U8145 ( .A(n8514), .ZN(n7152) );
  OR2_X1 U8146 ( .A1(n8521), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U8147 ( .A1(n8507), .A2(n8506), .ZN(n8521) );
  INV_X1 U8148 ( .A(n11576), .ZN(n7160) );
  NOR2_X1 U8149 ( .A1(n8365), .A2(n7159), .ZN(n7158) );
  INV_X1 U8150 ( .A(n8350), .ZN(n7159) );
  NAND2_X1 U8151 ( .A1(n12352), .A2(n11684), .ZN(n7161) );
  NAND2_X1 U8152 ( .A1(n8351), .A2(n7158), .ZN(n7157) );
  NOR2_X1 U8153 ( .A1(n11475), .A2(n9024), .ZN(n6920) );
  NAND2_X1 U8154 ( .A1(n8730), .A2(n8974), .ZN(n15075) );
  INV_X1 U8155 ( .A(SI_15_), .ZN(n8403) );
  INV_X1 U8156 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U8157 ( .A1(n7101), .A2(n6568), .ZN(n7100) );
  NOR2_X1 U8158 ( .A1(n7100), .A2(n7096), .ZN(n7095) );
  NOR2_X2 U8159 ( .A1(n8117), .A2(n7105), .ZN(n8119) );
  AND2_X1 U8160 ( .A1(n8118), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7105) );
  INV_X1 U8161 ( .A(n8256), .ZN(n7081) );
  NOR2_X1 U8162 ( .A1(n8258), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8275) );
  OR2_X1 U8163 ( .A1(n8244), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8258) );
  NOR2_X1 U8164 ( .A1(n7808), .A2(n7807), .ZN(n7806) );
  AOI21_X1 U8165 ( .B1(n7280), .B2(n7279), .A(n7278), .ZN(n7277) );
  INV_X1 U8166 ( .A(n9607), .ZN(n7278) );
  INV_X1 U8167 ( .A(n13063), .ZN(n7279) );
  AND2_X1 U8168 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7619) );
  NOR2_X1 U8169 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7525) );
  INV_X1 U8170 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7524) );
  NAND2_X1 U8171 ( .A1(n13229), .A2(n13107), .ZN(n7324) );
  AND2_X1 U8172 ( .A1(n13246), .A2(n13258), .ZN(n8029) );
  INV_X1 U8173 ( .A(n8028), .ZN(n7041) );
  NAND2_X1 U8174 ( .A1(n13290), .A2(n7908), .ZN(n6768) );
  INV_X1 U8175 ( .A(n7055), .ZN(n7048) );
  NOR2_X1 U8176 ( .A1(n7860), .A2(n7859), .ZN(n7858) );
  NOR2_X1 U8177 ( .A1(n8021), .A2(n7056), .ZN(n7055) );
  INV_X1 U8178 ( .A(n8019), .ZN(n7056) );
  OAI21_X1 U8179 ( .B1(n8021), .B2(n7054), .A(n8022), .ZN(n7053) );
  NAND2_X1 U8180 ( .A1(n8020), .A2(n8019), .ZN(n7054) );
  INV_X1 U8181 ( .A(n8010), .ZN(n7038) );
  AND2_X1 U8182 ( .A1(n7714), .A2(n7550), .ZN(n7736) );
  NAND2_X1 U8183 ( .A1(n7722), .A2(n11351), .ZN(n6775) );
  OR2_X1 U8184 ( .A1(n6776), .A2(n11337), .ZN(n6772) );
  INV_X1 U8185 ( .A(n6777), .ZN(n6776) );
  OAI21_X1 U8186 ( .B1(n10935), .B2(n6778), .A(n13120), .ZN(n6777) );
  OR2_X1 U8187 ( .A1(n10935), .A2(n6775), .ZN(n6771) );
  NAND2_X1 U8188 ( .A1(n8008), .A2(n6448), .ZN(n11231) );
  NOR2_X1 U8189 ( .A1(n7716), .A2(n7715), .ZN(n7714) );
  AND2_X1 U8190 ( .A1(n10665), .A2(n10594), .ZN(n7319) );
  INV_X1 U8191 ( .A(n7646), .ZN(n7321) );
  NOR2_X1 U8192 ( .A1(n13238), .A2(n8029), .ZN(n13222) );
  OR2_X1 U8193 ( .A1(n13223), .A2(n13408), .ZN(n6662) );
  AOI21_X1 U8194 ( .B1(n6421), .B2(n7025), .A(n6509), .ZN(n7023) );
  NOR2_X1 U8195 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n7536) );
  INV_X1 U8196 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7124) );
  INV_X1 U8197 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U8198 ( .A1(n7743), .A2(n7820), .ZN(n7822) );
  OR2_X1 U8199 ( .A1(n7679), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7692) );
  OR2_X1 U8200 ( .A1(n7634), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7649) );
  INV_X1 U8201 ( .A(n7376), .ZN(n7375) );
  OAI21_X1 U8202 ( .B1(n13579), .B2(n7377), .A(n13648), .ZN(n7376) );
  INV_X1 U8203 ( .A(n11869), .ZN(n7377) );
  NOR2_X1 U8204 ( .A1(n12175), .A2(n12176), .ZN(n7199) );
  NAND2_X1 U8205 ( .A1(n6387), .A2(n12220), .ZN(n7204) );
  OR2_X1 U8206 ( .A1(n11923), .A2(n11129), .ZN(n9787) );
  INV_X1 U8207 ( .A(n6933), .ZN(n6932) );
  NAND2_X1 U8208 ( .A1(n7517), .A2(n7565), .ZN(n6901) );
  INV_X1 U8209 ( .A(n10873), .ZN(n6978) );
  AND2_X1 U8210 ( .A1(n14559), .A2(n11976), .ZN(n11970) );
  INV_X1 U8211 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9466) );
  AOI21_X1 U8212 ( .B1(n6885), .B2(n6888), .A(n6883), .ZN(n6882) );
  NAND2_X1 U8213 ( .A1(n7940), .A2(n6885), .ZN(n6596) );
  INV_X1 U8214 ( .A(n8692), .ZN(n6883) );
  XNOR2_X1 U8215 ( .A(n9342), .B(SI_29_), .ZN(n9340) );
  NAND2_X1 U8216 ( .A1(n7911), .A2(n6902), .ZN(n7364) );
  INV_X1 U8217 ( .A(n7517), .ZN(n6902) );
  NAND2_X1 U8218 ( .A1(n7911), .A2(n7365), .ZN(n7367) );
  NOR2_X1 U8219 ( .A1(n7517), .A2(n7565), .ZN(n7365) );
  MUX2_X1 U8220 ( .A(n8118), .B(n11851), .S(n9812), .Z(n7510) );
  NAND2_X1 U8221 ( .A1(n7895), .A2(n7509), .ZN(n7512) );
  AND2_X1 U8222 ( .A1(n7408), .A2(n6816), .ZN(n7407) );
  AND2_X1 U8223 ( .A1(n7408), .A2(n9474), .ZN(n6814) );
  NAND2_X1 U8224 ( .A1(n6878), .A2(n7499), .ZN(n7880) );
  AND2_X1 U8225 ( .A1(n7503), .A2(n7502), .ZN(n7879) );
  INV_X1 U8226 ( .A(n7487), .ZN(n7356) );
  INV_X1 U8227 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9474) );
  AND2_X1 U8228 ( .A1(n9474), .A2(n12612), .ZN(n7244) );
  OR2_X1 U8229 ( .A1(n7764), .A2(n8386), .ZN(n7765) );
  NAND4_X1 U8230 ( .A1(n7423), .A2(n7362), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6875) );
  INV_X1 U8231 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7362) );
  OAI21_X1 U8232 ( .B1(n8846), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6511), .ZN(
        n6967) );
  XNOR2_X1 U8233 ( .A(n6967), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n8861) );
  AOI21_X1 U8234 ( .B1(n6678), .B2(n6677), .A(n6676), .ZN(n8831) );
  AND2_X1 U8235 ( .A1(n13800), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6676) );
  INV_X1 U8236 ( .A(n8868), .ZN(n6677) );
  INV_X1 U8237 ( .A(n8869), .ZN(n6678) );
  AND2_X1 U8238 ( .A1(n6682), .A2(n6681), .ZN(n8836) );
  NAND2_X1 U8239 ( .A1(n10039), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n6681) );
  AOI21_X1 U8240 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n13820), .A(n8838), .ZN(
        n8889) );
  NOR2_X1 U8241 ( .A1(n8885), .A2(n8884), .ZN(n8838) );
  NOR2_X1 U8242 ( .A1(n8407), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8427) );
  AND2_X1 U8243 ( .A1(n8427), .A2(n12326), .ZN(n8454) );
  INV_X1 U8244 ( .A(n10793), .ZN(n7007) );
  INV_X1 U8245 ( .A(SI_17_), .ZN(n8449) );
  INV_X1 U8246 ( .A(n14361), .ZN(n12474) );
  NAND2_X1 U8247 ( .A1(n6908), .A2(n10588), .ZN(n9120) );
  NAND2_X1 U8248 ( .A1(n11497), .A2(n6481), .ZN(n11614) );
  INV_X1 U8249 ( .A(n8758), .ZN(n7018) );
  INV_X1 U8250 ( .A(n7016), .ZN(n7015) );
  AOI21_X1 U8251 ( .B1(n7016), .B2(n7014), .A(n6556), .ZN(n7013) );
  OR2_X1 U8252 ( .A1(n8468), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8482) );
  AOI21_X1 U8253 ( .B1(n10308), .B2(n10301), .A(n10317), .ZN(n10302) );
  INV_X1 U8254 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n10480) );
  AOI21_X1 U8255 ( .B1(n10475), .B2(n6440), .A(n10332), .ZN(n10491) );
  AND2_X1 U8256 ( .A1(n6841), .A2(n6842), .ZN(n10496) );
  OR2_X1 U8257 ( .A1(n14888), .A2(n12429), .ZN(n7114) );
  OR2_X1 U8258 ( .A1(n14925), .A2(n14926), .ZN(n6827) );
  NAND2_X1 U8259 ( .A1(n14967), .A2(n6831), .ZN(n6830) );
  INV_X1 U8260 ( .A(n7115), .ZN(n6831) );
  NAND2_X1 U8261 ( .A1(n8137), .A2(n6606), .ZN(n6614) );
  NOR2_X1 U8262 ( .A1(n8150), .A2(n6613), .ZN(n6612) );
  NOR2_X1 U8263 ( .A1(n6615), .A2(n8416), .ZN(n6606) );
  NAND2_X1 U8264 ( .A1(n6835), .A2(n6489), .ZN(n6834) );
  AOI21_X1 U8265 ( .B1(n6688), .B2(n12516), .A(n12500), .ZN(n8595) );
  INV_X1 U8266 ( .A(n12500), .ZN(n7173) );
  AOI21_X1 U8267 ( .B1(n12555), .B2(n8547), .A(n8567), .ZN(n12535) );
  INV_X1 U8268 ( .A(n9134), .ZN(n12548) );
  OR2_X1 U8269 ( .A1(n8535), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U8270 ( .A1(n9085), .A2(n8638), .ZN(n12561) );
  INV_X1 U8271 ( .A(n9132), .ZN(n12578) );
  NAND2_X1 U8272 ( .A1(n7147), .A2(n8529), .ZN(n12579) );
  NAND2_X1 U8273 ( .A1(n8515), .A2(n7151), .ZN(n7147) );
  AND2_X1 U8274 ( .A1(n8488), .A2(n9062), .ZN(n12771) );
  AOI21_X1 U8275 ( .B1(n12810), .B2(n6914), .A(n6913), .ZN(n6912) );
  INV_X1 U8276 ( .A(n9052), .ZN(n6914) );
  AND2_X1 U8277 ( .A1(n8966), .A2(n8967), .ZN(n12793) );
  AND2_X1 U8278 ( .A1(n9045), .A2(n9044), .ZN(n11628) );
  OR2_X1 U8279 ( .A1(n8390), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8407) );
  AND2_X1 U8280 ( .A1(n9041), .A2(n9040), .ZN(n11576) );
  NAND2_X1 U8281 ( .A1(n7157), .A2(n7161), .ZN(n11571) );
  NAND2_X1 U8282 ( .A1(n7157), .A2(n7155), .ZN(n11573) );
  INV_X1 U8283 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n12350) );
  NAND2_X1 U8284 ( .A1(n8300), .A2(n14891), .ZN(n8316) );
  OR2_X1 U8285 ( .A1(n8316), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8332) );
  INV_X1 U8286 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8280) );
  AND2_X1 U8287 ( .A1(n8281), .A2(n8280), .ZN(n8300) );
  AND3_X1 U8288 ( .A1(n8298), .A2(n8297), .A3(n8296), .ZN(n15010) );
  AND2_X1 U8289 ( .A1(n9008), .A2(n9007), .ZN(n11026) );
  NOR2_X1 U8290 ( .A1(n8265), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U8291 ( .A1(n15025), .A2(n8248), .ZN(n11049) );
  NAND2_X1 U8292 ( .A1(n12908), .A2(n6694), .ZN(n15086) );
  NAND2_X1 U8293 ( .A1(n15084), .A2(n6908), .ZN(n12902) );
  NAND2_X1 U8294 ( .A1(n8493), .A2(n8492), .ZN(n12338) );
  NAND2_X1 U8295 ( .A1(n8467), .A2(n8466), .ZN(n12364) );
  NAND2_X1 U8296 ( .A1(n8426), .A2(n8425), .ZN(n12322) );
  NAND2_X1 U8297 ( .A1(n8351), .A2(n8350), .ZN(n11678) );
  NAND2_X1 U8298 ( .A1(n7144), .A2(n7142), .ZN(n11474) );
  NAND2_X1 U8299 ( .A1(n7094), .A2(n7098), .ZN(n8941) );
  INV_X1 U8300 ( .A(n7099), .ZN(n7098) );
  OAI22_X1 U8301 ( .A1(n6437), .A2(n7100), .B1(n11944), .B2(
        P2_DATAO_REG_29__SCAN_IN), .ZN(n7099) );
  NAND2_X1 U8302 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7103), .ZN(n7102) );
  NAND2_X1 U8303 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n6685), .ZN(n6684) );
  NAND2_X1 U8304 ( .A1(n11326), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U8305 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n12228), .ZN(n8115) );
  NAND2_X1 U8306 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n12704), .ZN(n8111) );
  NAND2_X1 U8307 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n6630), .ZN(n6629) );
  INV_X1 U8308 ( .A(n8128), .ZN(n7005) );
  AND2_X1 U8309 ( .A1(n8291), .A2(n8290), .ZN(n8294) );
  AND2_X1 U8310 ( .A1(n8275), .A2(n8274), .ZN(n8291) );
  INV_X1 U8311 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8274) );
  OR2_X1 U8312 ( .A1(n11951), .A2(n11952), .ZN(n7313) );
  INV_X1 U8313 ( .A(n7899), .ZN(n7917) );
  NAND2_X1 U8314 ( .A1(n11603), .A2(n11602), .ZN(n7306) );
  NAND2_X1 U8315 ( .A1(n7917), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U8316 ( .A1(n13053), .A2(n13054), .ZN(n13052) );
  AND2_X1 U8317 ( .A1(n9436), .A2(n9428), .ZN(n9864) );
  CLKBUF_X1 U8318 ( .A(n7862), .Z(n7887) );
  OR2_X1 U8319 ( .A1(n7577), .A2(n9871), .ZN(n7581) );
  OR2_X1 U8320 ( .A1(n7599), .A2(n10246), .ZN(n7571) );
  OR2_X1 U8321 ( .A1(n7578), .A2(n7568), .ZN(n7570) );
  NOR2_X1 U8322 ( .A1(n6950), .A2(n6949), .ZN(n6947) );
  NAND2_X1 U8323 ( .A1(n7029), .A2(n7035), .ZN(n7028) );
  INV_X1 U8324 ( .A(n7033), .ZN(n7029) );
  AND2_X1 U8325 ( .A1(n9390), .A2(n9389), .ZN(n13227) );
  INV_X1 U8326 ( .A(n6768), .ZN(n13275) );
  AND2_X1 U8327 ( .A1(n6751), .A2(n7878), .ZN(n6750) );
  NAND2_X1 U8328 ( .A1(n6462), .A2(n6753), .ZN(n6752) );
  INV_X1 U8329 ( .A(n13331), .ZN(n8025) );
  OR2_X1 U8330 ( .A1(n7845), .A2(n7844), .ZN(n7860) );
  NAND2_X1 U8331 ( .A1(n7052), .A2(n7050), .ZN(n13347) );
  INV_X1 U8332 ( .A(n7053), .ZN(n7050) );
  NAND2_X1 U8333 ( .A1(n13385), .A2(n7055), .ZN(n7052) );
  INV_X1 U8334 ( .A(n13359), .ZN(n13374) );
  INV_X1 U8335 ( .A(n6952), .ZN(n13395) );
  OR2_X1 U8336 ( .A1(n7793), .A2(n11604), .ZN(n7808) );
  OR2_X1 U8337 ( .A1(n7775), .A2(n7774), .ZN(n7793) );
  NAND2_X1 U8338 ( .A1(n7333), .A2(n7332), .ZN(n7759) );
  OAI21_X1 U8339 ( .B1(n10934), .B2(n6773), .A(n6770), .ZN(n11348) );
  AOI21_X1 U8340 ( .B1(n7722), .B2(n11333), .A(n6774), .ZN(n6773) );
  AND2_X1 U8341 ( .A1(n6772), .A2(n6771), .ZN(n6770) );
  INV_X1 U8342 ( .A(n6775), .ZN(n6774) );
  NAND2_X1 U8343 ( .A1(n11231), .A2(n8010), .ZN(n11350) );
  NAND2_X1 U8344 ( .A1(n8008), .A2(n8007), .ZN(n11233) );
  NAND2_X1 U8345 ( .A1(n6946), .A2(n6760), .ZN(n10671) );
  INV_X1 U8346 ( .A(n10601), .ZN(n6946) );
  XNOR2_X1 U8347 ( .A(n13127), .B(n10559), .ZN(n10446) );
  NAND2_X1 U8348 ( .A1(n10452), .A2(n10559), .ZN(n10601) );
  XNOR2_X1 U8349 ( .A(n13128), .B(n10563), .ZN(n10366) );
  XNOR2_X1 U8350 ( .A(n7605), .B(n9166), .ZN(n10263) );
  NAND2_X1 U8351 ( .A1(n13131), .A2(n10243), .ZN(n10231) );
  CLKBUF_X1 U8352 ( .A(n9501), .Z(n13355) );
  INV_X1 U8353 ( .A(n9364), .ZN(n13437) );
  OR2_X1 U8354 ( .A1(n8714), .A2(n7985), .ZN(n13201) );
  NOR2_X1 U8355 ( .A1(n13294), .A2(n6422), .ZN(n13283) );
  NAND2_X1 U8356 ( .A1(n10242), .A2(n9627), .ZN(n14849) );
  NAND2_X1 U8357 ( .A1(n7024), .A2(n7999), .ZN(n10666) );
  NAND2_X1 U8358 ( .A1(n10595), .A2(n6759), .ZN(n7024) );
  INV_X1 U8359 ( .A(n14849), .ZN(n13506) );
  NAND4_X1 U8360 ( .A1(n7743), .A2(n7339), .A3(n7532), .A4(n7537), .ZN(n7540)
         );
  INV_X1 U8361 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8051) );
  INV_X1 U8362 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7767) );
  INV_X1 U8363 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7817) );
  INV_X1 U8364 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10967) );
  NAND2_X1 U8365 ( .A1(n6671), .A2(n11650), .ZN(n13589) );
  OAI22_X1 U8366 ( .A1(n12006), .A2(n9728), .B1(n9737), .B2(n14623), .ZN(n9706) );
  AOI21_X1 U8367 ( .B1(n7395), .B2(n7397), .A(n6475), .ZN(n7393) );
  OR2_X1 U8368 ( .A1(n10968), .A2(n10967), .ZN(n10981) );
  OAI22_X1 U8369 ( .A1(n9737), .A2(n6591), .B1(n9728), .B2(n10881), .ZN(n6820)
         );
  NAND2_X1 U8370 ( .A1(n11659), .A2(n11660), .ZN(n7378) );
  INV_X1 U8371 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12613) );
  OR2_X1 U8372 ( .A1(n11546), .A2(n12613), .ZN(n11692) );
  AND2_X1 U8373 ( .A1(n11736), .A2(n7382), .ZN(n7381) );
  INV_X1 U8374 ( .A(n13629), .ZN(n7382) );
  AND2_X1 U8375 ( .A1(n6819), .A2(n10800), .ZN(n6818) );
  NAND2_X1 U8376 ( .A1(n11854), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11872) );
  INV_X1 U8377 ( .A(n11856), .ZN(n11854) );
  INV_X1 U8378 ( .A(n10800), .ZN(n7385) );
  OR2_X1 U8379 ( .A1(n10981), .A2(n10980), .ZN(n11090) );
  NOR2_X1 U8380 ( .A1(n11090), .A2(n11435), .ZN(n11106) );
  NAND2_X1 U8381 ( .A1(n11425), .A2(n11426), .ZN(n7405) );
  INV_X1 U8382 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U8383 ( .A1(n11797), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11818) );
  INV_X1 U8384 ( .A(n11798), .ZN(n11797) );
  NAND2_X1 U8385 ( .A1(n13609), .A2(n11831), .ZN(n13671) );
  INV_X1 U8386 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11174) );
  OR2_X1 U8387 ( .A1(n11175), .A2(n11174), .ZN(n11187) );
  NAND2_X1 U8388 ( .A1(n7406), .A2(n7402), .ZN(n11651) );
  AND2_X1 U8389 ( .A1(n11432), .A2(n7405), .ZN(n7402) );
  NAND2_X1 U8390 ( .A1(n11690), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11757) );
  INV_X1 U8391 ( .A(n11692), .ZN(n11690) );
  OR2_X1 U8392 ( .A1(n11757), .A2(n11756), .ZN(n11778) );
  OR2_X1 U8393 ( .A1(n11303), .A2(n11302), .ZN(n11525) );
  NAND2_X1 U8394 ( .A1(n11523), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11546) );
  INV_X1 U8395 ( .A(n11525), .ZN(n11523) );
  AOI21_X1 U8396 ( .B1(n6807), .B2(n6810), .A(n6506), .ZN(n6805) );
  NAND2_X1 U8397 ( .A1(n7196), .A2(n7191), .ZN(n7190) );
  INV_X1 U8398 ( .A(n7204), .ZN(n7191) );
  INV_X1 U8399 ( .A(n7196), .ZN(n7195) );
  NAND2_X1 U8400 ( .A1(n7196), .A2(n7186), .ZN(n7185) );
  NOR2_X1 U8401 ( .A1(n7204), .A2(n7198), .ZN(n7186) );
  AND2_X1 U8402 ( .A1(n11843), .A2(n11842), .ZN(n13875) );
  INV_X1 U8403 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n13800) );
  AND2_X2 U8404 ( .A1(n7268), .A2(n9473), .ZN(n10582) );
  NAND2_X1 U8405 ( .A1(n9793), .A2(n9792), .ZN(n13903) );
  INV_X1 U8406 ( .A(n7258), .ZN(n7252) );
  NOR2_X1 U8407 ( .A1(n7249), .A2(n13899), .ZN(n7248) );
  OAI22_X1 U8408 ( .A1(n13931), .A2(n7257), .B1(n13896), .B2(n13939), .ZN(
        n7256) );
  NOR2_X1 U8409 ( .A1(n6701), .A2(n13896), .ZN(n6700) );
  NOR2_X2 U8410 ( .A1(n13963), .A2(n14142), .ZN(n13951) );
  NAND2_X1 U8411 ( .A1(n13962), .A2(n13961), .ZN(n13960) );
  NAND2_X1 U8412 ( .A1(n13978), .A2(n6982), .ZN(n13958) );
  NAND2_X1 U8413 ( .A1(n14022), .A2(n6931), .ZN(n13981) );
  AOI22_X1 U8414 ( .A1(n13989), .A2(n13997), .B1(n13892), .B2(n14159), .ZN(
        n13974) );
  XNOR2_X1 U8415 ( .A(n14159), .B(n13876), .ZN(n13997) );
  NAND2_X1 U8416 ( .A1(n14022), .A2(n14007), .ZN(n14002) );
  AND2_X1 U8417 ( .A1(n14175), .A2(n13888), .ZN(n6648) );
  INV_X1 U8418 ( .A(n6935), .ZN(n14052) );
  INV_X1 U8419 ( .A(n13873), .ZN(n14050) );
  AOI21_X1 U8420 ( .B1(n6985), .B2(n14112), .A(n6507), .ZN(n6984) );
  NAND2_X1 U8421 ( .A1(n14113), .A2(n6985), .ZN(n6588) );
  NOR2_X2 U8422 ( .A1(n14107), .A2(n11704), .ZN(n11699) );
  NOR2_X1 U8423 ( .A1(n11187), .A2(n11671), .ZN(n11291) );
  NAND2_X1 U8424 ( .A1(n11291), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11303) );
  AND4_X1 U8425 ( .A1(n11308), .A2(n11307), .A3(n11306), .A4(n11305), .ZN(
        n11723) );
  AOI21_X1 U8426 ( .B1(n6971), .B2(n6972), .A(n6501), .ZN(n6969) );
  NAND2_X1 U8427 ( .A1(n14552), .A2(n11102), .ZN(n11103) );
  NOR2_X1 U8428 ( .A1(n12193), .A2(n6863), .ZN(n6862) );
  INV_X1 U8429 ( .A(n11102), .ZN(n6863) );
  OR2_X1 U8430 ( .A1(n11125), .A2(n14641), .ZN(n14576) );
  NAND2_X1 U8431 ( .A1(n6579), .A2(n14634), .ZN(n11125) );
  INV_X1 U8432 ( .A(n11157), .ZN(n6579) );
  NOR2_X1 U8433 ( .A1(n11979), .A2(n9792), .ZN(n13691) );
  NAND2_X1 U8434 ( .A1(n6856), .A2(n6860), .ZN(n14097) );
  OR2_X1 U8435 ( .A1(n14298), .A2(n11534), .ZN(n6856) );
  INV_X1 U8436 ( .A(n14240), .ZN(n9775) );
  XNOR2_X1 U8437 ( .A(n7957), .B(n7956), .ZN(n13562) );
  AND2_X1 U8438 ( .A1(n6812), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n6811) );
  OR2_X1 U8439 ( .A1(n6814), .A2(n9668), .ZN(n6812) );
  NAND2_X1 U8440 ( .A1(n10582), .A2(n7244), .ZN(n9667) );
  OR2_X1 U8441 ( .A1(n9855), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9858) );
  OR2_X1 U8442 ( .A1(n9858), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U8443 ( .A1(n7349), .A2(n7447), .ZN(n7648) );
  NAND2_X1 U8444 ( .A1(n7633), .A2(n7445), .ZN(n7349) );
  CLKBUF_X1 U8445 ( .A(n9696), .Z(n9697) );
  NOR2_X1 U8446 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9751) );
  INV_X1 U8447 ( .A(n6957), .ZN(n8849) );
  INV_X1 U8448 ( .A(n8850), .ZN(n8821) );
  XNOR2_X1 U8449 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n6957) );
  AND2_X1 U8450 ( .A1(n8819), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U8451 ( .A1(n6672), .A2(n8870), .ZN(n8872) );
  NAND2_X1 U8452 ( .A1(n6965), .A2(n6795), .ZN(n6964) );
  NAND2_X1 U8453 ( .A1(n8886), .A2(n8887), .ZN(n6965) );
  OAI22_X1 U8454 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n8841), .B1(n8842), .B2(
        n8840), .ZN(n8895) );
  OR2_X1 U8455 ( .A1(n14515), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6793) );
  AOI21_X1 U8456 ( .B1(n6992), .B2(n6995), .A(n6990), .ZN(n6989) );
  INV_X1 U8457 ( .A(n12347), .ZN(n6990) );
  NAND2_X1 U8458 ( .A1(n11457), .A2(n8755), .ZN(n11496) );
  NAND2_X1 U8459 ( .A1(n10680), .A2(n10679), .ZN(n10678) );
  AND2_X1 U8460 ( .A1(n8732), .A2(n8728), .ZN(n6987) );
  AND3_X1 U8461 ( .A1(n8499), .A2(n8498), .A3(n8497), .ZN(n12742) );
  NAND2_X1 U8462 ( .A1(n12259), .A2(n7421), .ZN(n12314) );
  NAND2_X1 U8463 ( .A1(n12325), .A2(n12324), .ZN(n12323) );
  INV_X1 U8464 ( .A(n12402), .ZN(n12820) );
  NAND2_X1 U8465 ( .A1(n12323), .A2(n8775), .ZN(n12331) );
  NAND2_X1 U8466 ( .A1(n10678), .A2(n8737), .ZN(n10792) );
  NAND2_X1 U8467 ( .A1(n6991), .A2(n8763), .ZN(n12348) );
  NAND2_X1 U8468 ( .A1(n11636), .A2(n8761), .ZN(n6991) );
  AOI21_X1 U8469 ( .B1(n12525), .B2(n8547), .A(n8169), .ZN(n12536) );
  INV_X1 U8470 ( .A(n12838), .ZN(n12380) );
  INV_X1 U8471 ( .A(n12404), .ZN(n12819) );
  NAND2_X1 U8472 ( .A1(n8797), .A2(n10631), .ZN(n12395) );
  AND2_X1 U8473 ( .A1(n8795), .A2(n10286), .ZN(n14861) );
  NAND2_X1 U8474 ( .A1(n8806), .A2(n8805), .ZN(n12392) );
  INV_X1 U8475 ( .A(n14407), .ZN(n8956) );
  NAND2_X1 U8476 ( .A1(n8583), .A2(n8582), .ZN(n12550) );
  INV_X1 U8477 ( .A(n9084), .ZN(n12582) );
  INV_X1 U8478 ( .A(n12742), .ZN(n12767) );
  NAND2_X1 U8479 ( .A1(n8605), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U8480 ( .A1(n6419), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8206) );
  OR2_X1 U8481 ( .A1(n8509), .A2(n8170), .ZN(n8171) );
  NAND2_X1 U8482 ( .A1(n6419), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8172) );
  AND4_X2 U8483 ( .A1(n8185), .A2(n8184), .A3(n8182), .A4(n8183), .ZN(n9653)
         );
  OR2_X1 U8484 ( .A1(n8509), .A2(n10585), .ZN(n8182) );
  NAND2_X1 U8485 ( .A1(n10476), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10475) );
  AND2_X1 U8486 ( .A1(n10487), .A2(n10498), .ZN(n6641) );
  NAND2_X1 U8487 ( .A1(n6843), .A2(n6841), .ZN(n14879) );
  NOR2_X1 U8488 ( .A1(n6842), .A2(n10493), .ZN(n14878) );
  XNOR2_X1 U8489 ( .A(n10639), .B(n10652), .ZN(n10521) );
  NAND2_X1 U8490 ( .A1(n10521), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n10640) );
  INV_X1 U8491 ( .A(n6839), .ZN(n10656) );
  NOR2_X1 U8492 ( .A1(n10642), .A2(n10643), .ZN(n12413) );
  AND2_X1 U8493 ( .A1(n7114), .A2(n7113), .ZN(n14906) );
  INV_X1 U8494 ( .A(n14907), .ZN(n7113) );
  INV_X1 U8495 ( .A(n7114), .ZN(n14908) );
  INV_X1 U8496 ( .A(n6827), .ZN(n14924) );
  INV_X1 U8497 ( .A(n7116), .ZN(n14941) );
  INV_X1 U8498 ( .A(n7118), .ZN(n14943) );
  AND2_X1 U8499 ( .A1(n6832), .A2(n6653), .ZN(n14979) );
  NAND2_X1 U8500 ( .A1(n6418), .A2(n14967), .ZN(n6653) );
  XNOR2_X1 U8501 ( .A(n12434), .B(n14331), .ZN(n14325) );
  INV_X1 U8502 ( .A(n6835), .ZN(n14324) );
  NAND2_X1 U8503 ( .A1(P3_U3897), .A2(n10285), .ZN(n14952) );
  INV_X1 U8504 ( .A(n7111), .ZN(n14341) );
  INV_X1 U8505 ( .A(n6834), .ZN(n14343) );
  INV_X1 U8506 ( .A(n7109), .ZN(n12435) );
  NAND2_X1 U8507 ( .A1(n8938), .A2(n8937), .ZN(n14407) );
  AOI21_X1 U8508 ( .B1(n11569), .B2(n8587), .A(n8543), .ZN(n12572) );
  NAND2_X1 U8509 ( .A1(n8515), .A2(n8514), .ZN(n12729) );
  NAND2_X1 U8510 ( .A1(n6918), .A2(n8634), .ZN(n12756) );
  NAND2_X1 U8511 ( .A1(n7162), .A2(n8460), .ZN(n12779) );
  NAND2_X1 U8512 ( .A1(n12811), .A2(n12810), .ZN(n12809) );
  NAND2_X1 U8513 ( .A1(n12821), .A2(n9052), .ZN(n12811) );
  INV_X1 U8514 ( .A(n12498), .ZN(n15020) );
  NAND2_X1 U8515 ( .A1(n7165), .A2(n8279), .ZN(n15014) );
  AND2_X1 U8516 ( .A1(n15109), .A2(n15097), .ZN(n12586) );
  INV_X1 U8517 ( .A(n15078), .ZN(n15103) );
  INV_X1 U8518 ( .A(n12524), .ZN(n12915) );
  AND2_X1 U8519 ( .A1(n8534), .A2(n8533), .ZN(n12924) );
  NAND2_X1 U8520 ( .A1(n8481), .A2(n8480), .ZN(n12940) );
  INV_X1 U8521 ( .A(n12364), .ZN(n12944) );
  INV_X1 U8522 ( .A(n12322), .ZN(n12952) );
  INV_X1 U8523 ( .A(n12384), .ZN(n12956) );
  NAND2_X1 U8524 ( .A1(n8374), .A2(n8373), .ZN(n12964) );
  NAND2_X1 U8525 ( .A1(n8330), .A2(n8329), .ZN(n11499) );
  AND2_X1 U8526 ( .A1(n6997), .A2(n6460), .ZN(n12968) );
  AND2_X1 U8527 ( .A1(n8674), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12967) );
  INV_X1 U8528 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8148) );
  XNOR2_X1 U8529 ( .A(n8585), .B(n8122), .ZN(n12980) );
  NAND2_X1 U8530 ( .A1(n8654), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U8531 ( .A1(n8653), .A2(n8654), .ZN(n12994) );
  XOR2_X1 U8532 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8542), .Z(n11569) );
  XNOR2_X1 U8533 ( .A(n8599), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U8534 ( .A1(n7004), .A2(n6430), .ZN(n8601) );
  INV_X1 U8535 ( .A(n12471), .ZN(n14349) );
  INV_X1 U8536 ( .A(n12469), .ZN(n14331) );
  INV_X1 U8537 ( .A(SI_13_), .ZN(n14276) );
  XNOR2_X1 U8538 ( .A(n8354), .B(n7176), .ZN(n14949) );
  NAND2_X1 U8539 ( .A1(n8104), .A2(n8103), .ZN(n8340) );
  XNOR2_X1 U8540 ( .A(n8327), .B(n8326), .ZN(n14914) );
  INV_X1 U8541 ( .A(n14277), .ZN(n14288) );
  INV_X1 U8542 ( .A(n10520), .ZN(n10525) );
  NAND2_X1 U8543 ( .A1(n7083), .A2(n7079), .ZN(n8257) );
  NAND2_X1 U8544 ( .A1(n6576), .A2(n7086), .ZN(n7079) );
  NAND2_X1 U8545 ( .A1(n8092), .A2(n7088), .ZN(n8243) );
  NAND2_X1 U8546 ( .A1(n7089), .A2(n7090), .ZN(n7088) );
  NAND3_X1 U8547 ( .A1(n6848), .A2(n6846), .A3(n6845), .ZN(n10329) );
  OAI211_X1 U8548 ( .C1(P3_IR_REG_0__SCAN_IN), .C2(P3_IR_REG_1__SCAN_IN), .A(
        P3_IR_REG_2__SCAN_IN), .B(P3_IR_REG_31__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U8549 ( .A1(n6847), .A2(n8416), .ZN(n6846) );
  NAND2_X1 U8550 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8177) );
  NAND2_X1 U8551 ( .A1(n9812), .A2(P3_U3151), .ZN(n14277) );
  NAND2_X1 U8552 ( .A1(n7294), .A2(n9527), .ZN(n10762) );
  NAND2_X1 U8553 ( .A1(n10570), .A2(n7292), .ZN(n7294) );
  NAND2_X1 U8554 ( .A1(n13444), .A2(n13086), .ZN(n11961) );
  AND2_X1 U8555 ( .A1(n7284), .A2(n6472), .ZN(n11558) );
  XNOR2_X1 U8556 ( .A(n7302), .B(n9613), .ZN(n12997) );
  NAND2_X1 U8557 ( .A1(n13070), .A2(n9612), .ZN(n7302) );
  NAND2_X2 U8558 ( .A1(n7914), .A2(n7913), .ZN(n13466) );
  INV_X1 U8559 ( .A(n13122), .ZN(n10937) );
  NAND2_X1 U8560 ( .A1(n10190), .A2(n9510), .ZN(n13003) );
  AOI21_X1 U8561 ( .B1(n7309), .B2(n7308), .A(n13024), .ZN(n7307) );
  AOI21_X1 U8562 ( .B1(n7290), .B2(n10761), .A(n6476), .ZN(n7289) );
  NAND2_X1 U8563 ( .A1(n7682), .A2(n7681), .ZN(n10853) );
  NAND2_X1 U8564 ( .A1(n13062), .A2(n9601), .ZN(n13036) );
  NAND2_X1 U8565 ( .A1(n13062), .A2(n7280), .ZN(n13037) );
  INV_X1 U8566 ( .A(n13107), .ZN(n13243) );
  INV_X1 U8567 ( .A(n13109), .ZN(n13242) );
  NAND2_X1 U8568 ( .A1(n7306), .A2(n9574), .ZN(n13046) );
  INV_X1 U8569 ( .A(n7298), .ZN(n9641) );
  NAND2_X1 U8570 ( .A1(n11340), .A2(n9560), .ZN(n11364) );
  NAND2_X1 U8571 ( .A1(n7315), .A2(n7314), .ZN(n9509) );
  INV_X1 U8572 ( .A(n9508), .ZN(n7315) );
  NAND2_X1 U8573 ( .A1(n10570), .A2(n9522), .ZN(n10608) );
  OR2_X1 U8574 ( .A1(n9422), .A2(n9428), .ZN(n6673) );
  NAND2_X1 U8575 ( .A1(n7062), .A2(n7064), .ZN(n7061) );
  XNOR2_X1 U8576 ( .A(n8696), .B(n8695), .ZN(n13440) );
  OAI21_X1 U8577 ( .B1(n7325), .B2(n6765), .A(n6763), .ZN(n7973) );
  INV_X1 U8578 ( .A(n13422), .ZN(n13269) );
  NAND2_X1 U8579 ( .A1(n7318), .A2(n7892), .ZN(n13291) );
  AND2_X1 U8580 ( .A1(n14835), .A2(n8700), .ZN(n13339) );
  NAND2_X1 U8581 ( .A1(n6749), .A2(n6753), .ZN(n13327) );
  NAND2_X1 U8582 ( .A1(n13372), .A2(n6420), .ZN(n6749) );
  NAND2_X1 U8583 ( .A1(n6756), .A2(n7850), .ZN(n13346) );
  NAND2_X1 U8584 ( .A1(n6757), .A2(n9410), .ZN(n6756) );
  INV_X1 U8585 ( .A(n13372), .ZN(n6757) );
  OAI21_X1 U8586 ( .B1(n13385), .B2(n8020), .A(n8019), .ZN(n13368) );
  NAND2_X1 U8587 ( .A1(n7827), .A2(n7826), .ZN(n13500) );
  NAND2_X1 U8588 ( .A1(n11592), .A2(n7337), .ZN(n13409) );
  AND2_X1 U8589 ( .A1(n11592), .A2(n7800), .ZN(n13410) );
  NAND2_X1 U8590 ( .A1(n7805), .A2(n7804), .ZN(n13505) );
  NAND2_X1 U8591 ( .A1(n11482), .A2(n7059), .ZN(n11590) );
  NAND2_X1 U8592 ( .A1(n7791), .A2(n7790), .ZN(n11610) );
  NAND2_X1 U8593 ( .A1(n6781), .A2(n9405), .ZN(n14434) );
  INV_X1 U8594 ( .A(n11491), .ZN(n6781) );
  INV_X1 U8595 ( .A(n13425), .ZN(n13373) );
  NAND2_X1 U8596 ( .A1(n7758), .A2(n7757), .ZN(n11420) );
  NAND2_X1 U8597 ( .A1(n7746), .A2(n7745), .ZN(n11360) );
  NAND2_X1 U8598 ( .A1(n6769), .A2(n7722), .ZN(n11230) );
  NAND2_X1 U8599 ( .A1(n10934), .A2(n10935), .ZN(n6769) );
  NAND2_X1 U8600 ( .A1(n13356), .A2(n8717), .ZN(n13376) );
  NAND2_X1 U8601 ( .A1(n10703), .A2(n7676), .ZN(n10840) );
  NAND2_X1 U8602 ( .A1(n10664), .A2(n10665), .ZN(n10663) );
  NAND2_X1 U8603 ( .A1(n10592), .A2(n7646), .ZN(n10664) );
  NOR2_X1 U8604 ( .A1(n10234), .A2(n6570), .ZN(n10237) );
  INV_X2 U8605 ( .A(n13339), .ZN(n13412) );
  AND2_X1 U8606 ( .A1(n9423), .A2(n11059), .ZN(n10245) );
  INV_X1 U8607 ( .A(n6692), .ZN(n6940) );
  OAI21_X1 U8608 ( .B1(n7595), .B2(n9845), .A(n7021), .ZN(n6692) );
  INV_X1 U8609 ( .A(n13246), .ZN(n13526) );
  OR3_X1 U8610 ( .A1(n13464), .A2(n13463), .A3(n13462), .ZN(n13527) );
  INV_X1 U8611 ( .A(n13319), .ZN(n13536) );
  INV_X1 U8612 ( .A(n13337), .ZN(n13540) );
  INV_X1 U8613 ( .A(n13360), .ZN(n13544) );
  NAND2_X1 U8614 ( .A1(n7699), .A2(n7698), .ZN(n11003) );
  INV_X1 U8615 ( .A(n10238), .ZN(n10554) );
  INV_X1 U8616 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13552) );
  INV_X1 U8617 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11944) );
  INV_X1 U8618 ( .A(n7552), .ZN(n11946) );
  AND2_X1 U8619 ( .A1(n8048), .A2(n8049), .ZN(n13571) );
  INV_X1 U8620 ( .A(n7304), .ZN(n7303) );
  OAI22_X1 U8621 ( .A1(n7982), .A2(n7305), .B1(P2_IR_REG_31__SCAN_IN), .B2(
        P2_IR_REG_22__SCAN_IN), .ZN(n7304) );
  NAND2_X1 U8622 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n7305) );
  INV_X1 U8623 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11326) );
  INV_X1 U8624 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10251) );
  INV_X1 U8625 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10102) );
  INV_X1 U8626 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9945) );
  INV_X1 U8627 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9838) );
  INV_X1 U8628 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U8629 ( .A1(n13688), .A2(n10961), .ZN(n10978) );
  NAND2_X1 U8630 ( .A1(n6804), .A2(n6807), .ZN(n14460) );
  OR2_X1 U8631 ( .A1(n6609), .A2(n6810), .ZN(n6804) );
  NAND2_X1 U8632 ( .A1(n10389), .A2(n7410), .ZN(n9779) );
  OAI22_X1 U8633 ( .A1(n7391), .A2(n7390), .B1(n7398), .B2(n7393), .ZN(n7389)
         );
  NOR2_X1 U8634 ( .A1(n7395), .A2(n7398), .ZN(n7391) );
  INV_X1 U8635 ( .A(n7393), .ZN(n7390) );
  AND2_X1 U8636 ( .A1(n7395), .A2(n7398), .ZN(n7388) );
  NAND2_X1 U8637 ( .A1(n7393), .A2(n12236), .ZN(n7392) );
  NAND2_X1 U8638 ( .A1(n11256), .A2(n11255), .ZN(n11257) );
  NAND2_X1 U8639 ( .A1(n9740), .A2(n7400), .ZN(n10357) );
  NAND2_X1 U8640 ( .A1(n10268), .A2(n10269), .ZN(n7400) );
  NAND2_X1 U8641 ( .A1(n13655), .A2(n11811), .ZN(n13611) );
  INV_X1 U8642 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11671) );
  CLKBUF_X1 U8643 ( .A(n13618), .Z(n13619) );
  NAND2_X1 U8644 ( .A1(n11689), .A2(n11688), .ZN(n14197) );
  INV_X1 U8645 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10824) );
  NAND2_X1 U8646 ( .A1(n13580), .A2(n13579), .ZN(n7374) );
  AND2_X1 U8647 ( .A1(n7406), .A2(n7405), .ZN(n11433) );
  NAND2_X1 U8648 ( .A1(n13663), .A2(n13662), .ZN(n14459) );
  NAND2_X1 U8649 ( .A1(n6609), .A2(n11714), .ZN(n13663) );
  NAND2_X1 U8650 ( .A1(n11173), .A2(n11172), .ZN(n14474) );
  NOR2_X1 U8651 ( .A1(n7380), .A2(n6466), .ZN(n6824) );
  OR2_X1 U8652 ( .A1(n14467), .A2(n14468), .ZN(n7380) );
  INV_X1 U8653 ( .A(n11650), .ZN(n6825) );
  INV_X1 U8654 ( .A(n13590), .ZN(n6826) );
  NAND2_X1 U8655 ( .A1(n9786), .A2(n14555), .ZN(n14475) );
  OR3_X1 U8656 ( .A1(n9778), .A2(n9793), .A3(n14652), .ZN(n13705) );
  CLKBUF_X1 U8657 ( .A(n13707), .Z(n13708) );
  INV_X1 U8658 ( .A(n14479), .ZN(n13714) );
  INV_X1 U8659 ( .A(n12225), .ZN(n6586) );
  NAND2_X1 U8660 ( .A1(n11894), .A2(n11893), .ZN(n13894) );
  NAND2_X1 U8661 ( .A1(n11878), .A2(n11877), .ZN(n13893) );
  INV_X1 U8662 ( .A(n13875), .ZN(n13891) );
  INV_X1 U8663 ( .A(n12011), .ZN(n7266) );
  NAND4_X1 U8664 ( .A1(n9687), .A2(n9686), .A3(n9685), .A4(n9684), .ZN(n13731)
         );
  AND2_X1 U8665 ( .A1(n9724), .A2(n9725), .ZN(n6589) );
  OR2_X1 U8666 ( .A1(n9744), .A2(n10863), .ZN(n9727) );
  NAND2_X1 U8667 ( .A1(n11965), .A2(n11964), .ZN(n13856) );
  NAND2_X1 U8668 ( .A1(n13861), .A2(n6658), .ZN(n14120) );
  AND2_X1 U8669 ( .A1(n6659), .A2(n14591), .ZN(n6658) );
  OR2_X1 U8670 ( .A1(n6640), .A2(n14121), .ZN(n6659) );
  NAND2_X1 U8671 ( .A1(n7359), .A2(n7360), .ZN(n13941) );
  NAND2_X1 U8672 ( .A1(n13568), .A2(n11085), .ZN(n11885) );
  AND2_X1 U8673 ( .A1(n6871), .A2(n6433), .ZN(n14009) );
  NAND2_X1 U8674 ( .A1(n6871), .A2(n7261), .ZN(n14020) );
  NAND2_X1 U8675 ( .A1(n11776), .A2(n11775), .ZN(n14060) );
  INV_X1 U8676 ( .A(n6937), .ZN(n14071) );
  INV_X1 U8677 ( .A(n7259), .ZN(n14066) );
  NAND2_X1 U8678 ( .A1(n6868), .A2(n6444), .ZN(n14080) );
  NAND2_X1 U8679 ( .A1(n11685), .A2(n12078), .ZN(n13883) );
  INV_X1 U8680 ( .A(n11704), .ZN(n14202) );
  NAND2_X1 U8681 ( .A1(n14483), .A2(n6985), .ZN(n11705) );
  NAND2_X1 U8682 ( .A1(n11539), .A2(n11538), .ZN(n14483) );
  INV_X1 U8683 ( .A(n14113), .ZN(n11539) );
  NAND2_X1 U8684 ( .A1(n14298), .A2(n11299), .ZN(n11300) );
  NAND2_X1 U8685 ( .A1(n11280), .A2(n11279), .ZN(n14304) );
  NAND2_X1 U8686 ( .A1(n11089), .A2(n11088), .ZN(n12046) );
  NOR2_X1 U8687 ( .A1(n12232), .A2(n10408), .ZN(n14561) );
  NAND2_X1 U8688 ( .A1(n11100), .A2(n11099), .ZN(n14550) );
  NAND2_X1 U8689 ( .A1(n6970), .A2(n11080), .ZN(n14546) );
  NAND2_X1 U8690 ( .A1(n11079), .A2(n11078), .ZN(n6970) );
  OAI21_X1 U8691 ( .B1(n10889), .B2(n12188), .A(n6850), .ZN(n14565) );
  OR2_X1 U8692 ( .A1(n9946), .A2(n10399), .ZN(n14555) );
  NAND2_X1 U8693 ( .A1(n6975), .A2(n10873), .ZN(n11060) );
  NAND2_X1 U8694 ( .A1(n11124), .A2(n12186), .ZN(n6975) );
  NAND2_X1 U8695 ( .A1(n10890), .A2(n10891), .ZN(n11069) );
  AND2_X1 U8696 ( .A1(n14562), .A2(n14625), .ZN(n14063) );
  OAI211_X2 U8697 ( .C1(n6647), .C2(n9829), .A(n9754), .B(n9753), .ZN(n14589)
         );
  INV_X1 U8698 ( .A(n14585), .ZN(n14088) );
  INV_X1 U8699 ( .A(n11966), .ZN(n10862) );
  AND2_X1 U8700 ( .A1(n14562), .A2(n12226), .ZN(n14595) );
  AND2_X1 U8701 ( .A1(n14562), .A2(n14557), .ZN(n14585) );
  AND2_X2 U8702 ( .A1(n10417), .A2(n10416), .ZN(n14709) );
  NAND2_X1 U8703 ( .A1(n14120), .A2(n6656), .ZN(n14209) );
  INV_X1 U8704 ( .A(n6657), .ZN(n6656) );
  OAI21_X1 U8705 ( .B1(n14121), .B2(n14686), .A(n14119), .ZN(n6657) );
  NAND2_X1 U8706 ( .A1(n6939), .A2(n6486), .ZN(n6938) );
  INV_X1 U8707 ( .A(n6593), .ZN(n6592) );
  NAND2_X1 U8708 ( .A1(n14132), .A2(n14683), .ZN(n6595) );
  AND2_X2 U8709 ( .A1(n10417), .A2(n10860), .ZN(n14693) );
  AND2_X1 U8710 ( .A1(n6427), .A2(n9680), .ZN(n7267) );
  INV_X1 U8711 ( .A(n9690), .ZN(n9677) );
  AND4_X1 U8712 ( .A1(n9488), .A2(n6986), .A3(n7268), .A4(n6427), .ZN(n9679)
         );
  INV_X1 U8713 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14236) );
  NAND2_X1 U8714 ( .A1(n6884), .A2(n6889), .ZN(n8691) );
  NAND2_X1 U8715 ( .A1(n7940), .A2(n6891), .ZN(n6884) );
  OR2_X1 U8716 ( .A1(n11833), .A2(n11832), .ZN(n11834) );
  NAND2_X1 U8717 ( .A1(n9672), .A2(n6441), .ZN(n11982) );
  NAND2_X1 U8718 ( .A1(n6817), .A2(n6815), .ZN(n9672) );
  NAND2_X1 U8719 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6816), .ZN(n6815) );
  NAND2_X1 U8720 ( .A1(n6813), .A2(n6811), .ZN(n6817) );
  NAND2_X1 U8721 ( .A1(n6877), .A2(n7499), .ZN(n7868) );
  INV_X1 U8722 ( .A(n6878), .ZN(n6877) );
  NAND2_X1 U8723 ( .A1(n7372), .A2(n7368), .ZN(n7839) );
  NAND2_X1 U8724 ( .A1(n7372), .A2(n7371), .ZN(n7837) );
  INV_X1 U8725 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11285) );
  INV_X1 U8726 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10107) );
  INV_X1 U8727 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9943) );
  INV_X1 U8728 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9860) );
  INV_X1 U8729 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9852) );
  INV_X1 U8730 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9844) );
  INV_X1 U8731 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9834) );
  INV_X1 U8732 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9848) );
  AOI21_X1 U8733 ( .B1(n8855), .B2(n8854), .A(n14258), .ZN(n15168) );
  INV_X1 U8734 ( .A(n8876), .ZN(n6966) );
  XNOR2_X1 U8735 ( .A(n6964), .B(n6963), .ZN(n14513) );
  INV_X1 U8736 ( .A(n8891), .ZN(n6963) );
  AND2_X1 U8737 ( .A1(n6787), .A2(n6788), .ZN(n6786) );
  INV_X1 U8738 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8739 ( .A1(n14320), .A2(n8917), .ZN(n6958) );
  OAI21_X1 U8740 ( .B1(n9653), .B2(n12399), .A(n6907), .ZN(P3_U3491) );
  NAND2_X1 U8741 ( .A1(n12399), .A2(P3_DATAO_REG_0__SCAN_IN), .ZN(n6907) );
  AOI21_X1 U8742 ( .B1(n14865), .B2(P3_IR_REG_0__SCAN_IN), .A(n7108), .ZN(
        n14871) );
  OAI21_X1 U8743 ( .B1(n14867), .B2(P3_IR_REG_0__SCAN_IN), .A(n14866), .ZN(
        n14868) );
  OR2_X1 U8744 ( .A1(n12490), .A2(n14877), .ZN(n6573) );
  AOI211_X1 U8745 ( .C1(n6403), .C2(n14865), .A(n12487), .B(n12486), .ZN(
        n12489) );
  OAI21_X1 U8746 ( .B1(n9458), .B2(n9457), .A(n9462), .ZN(P3_U3488) );
  NAND2_X1 U8747 ( .A1(n12911), .A2(n15159), .ZN(n7169) );
  INV_X1 U8748 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n7168) );
  NAND2_X1 U8749 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_STATE_REG_SCAN_IN), .ZN(
        n9802) );
  NAND2_X1 U8750 ( .A1(n7272), .A2(n7274), .ZN(n10375) );
  AND3_X1 U8751 ( .A1(n13220), .A2(n13219), .A3(n13218), .ZN(n13221) );
  AOI21_X1 U8752 ( .B1(n13199), .B2(n11336), .A(n8927), .ZN(n8928) );
  NOR2_X1 U8753 ( .A1(n8081), .A2(n8083), .ZN(n8084) );
  NOR2_X1 U8754 ( .A1(n8925), .A2(n13548), .ZN(n8081) );
  AOI21_X1 U8755 ( .B1(n13229), .B2(n11002), .A(n6697), .ZN(n6696) );
  NOR2_X1 U8756 ( .A1(n6800), .A2(n6799), .ZN(n6798) );
  INV_X1 U8757 ( .A(n11943), .ZN(n6799) );
  OR2_X1 U8758 ( .A1(n12224), .A2(n12223), .ZN(n6584) );
  INV_X1 U8759 ( .A(n6795), .ZN(n14509) );
  NOR2_X1 U8760 ( .A1(n14516), .A2(n14515), .ZN(n14514) );
  INV_X1 U8761 ( .A(n6787), .ZN(n14522) );
  OAI21_X1 U8762 ( .B1(n6451), .B2(n8916), .A(n6617), .ZN(n6790) );
  AND2_X1 U8763 ( .A1(n6510), .A2(n6732), .ZN(n6417) );
  NAND2_X1 U8764 ( .A1(n7116), .A2(n7115), .ZN(n6418) );
  INV_X1 U8765 ( .A(n9405), .ZN(n6780) );
  INV_X1 U8766 ( .A(n8604), .ZN(n12480) );
  AND2_X1 U8767 ( .A1(n7850), .A2(n6459), .ZN(n6420) );
  AND2_X1 U8768 ( .A1(n6758), .A2(n9396), .ZN(n6421) );
  AND2_X1 U8769 ( .A1(n13532), .A2(n13313), .ZN(n6422) );
  AND2_X1 U8770 ( .A1(n14022), .A2(n6933), .ZN(n6423) );
  OR2_X1 U8771 ( .A1(n9293), .A2(n9292), .ZN(n6424) );
  INV_X1 U8772 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8139) );
  INV_X1 U8773 ( .A(n9410), .ZN(n13371) );
  NOR2_X1 U8774 ( .A1(n10491), .A2(n6643), .ZN(n6425) );
  NAND2_X1 U8775 ( .A1(n13308), .A2(n8028), .ZN(n7046) );
  INV_X1 U8776 ( .A(n10014), .ZN(n10243) );
  XNOR2_X1 U8777 ( .A(n13466), .B(n7922), .ZN(n13274) );
  INV_X1 U8778 ( .A(n13274), .ZN(n7329) );
  OR2_X1 U8779 ( .A1(n10652), .A2(n10651), .ZN(n6426) );
  AND2_X1 U8780 ( .A1(n9676), .A2(n9688), .ZN(n6427) );
  INV_X1 U8781 ( .A(n12104), .ZN(n7223) );
  XNOR2_X1 U8782 ( .A(n8656), .B(n8655), .ZN(n12990) );
  AND2_X1 U8783 ( .A1(n12141), .A2(n12140), .ZN(n14130) );
  AND2_X1 U8784 ( .A1(n14130), .A2(n13897), .ZN(n6428) );
  AND2_X1 U8785 ( .A1(n9184), .A2(n9185), .ZN(n6429) );
  AND2_X1 U8786 ( .A1(n8132), .A2(n8128), .ZN(n6430) );
  AND2_X1 U8787 ( .A1(n9211), .A2(n6477), .ZN(n6431) );
  NAND2_X1 U8788 ( .A1(n12080), .A2(n12082), .ZN(n7182) );
  OR2_X1 U8789 ( .A1(n9298), .A2(n9297), .ZN(n6432) );
  INV_X1 U8790 ( .A(n13466), .ZN(n13281) );
  NAND2_X1 U8791 ( .A1(n14515), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6792) );
  AND2_X1 U8792 ( .A1(n7261), .A2(n13889), .ZN(n6433) );
  AND2_X1 U8793 ( .A1(n9301), .A2(n9300), .ZN(n6434) );
  AND2_X1 U8794 ( .A1(n6901), .A2(n11085), .ZN(n6435) );
  NAND2_X1 U8795 ( .A1(n7713), .A2(n7712), .ZN(n10945) );
  INV_X1 U8796 ( .A(n10945), .ZN(n6944) );
  NAND2_X1 U8797 ( .A1(n6921), .A2(n6920), .ZN(n6436) );
  INV_X1 U8798 ( .A(n8932), .ZN(n7101) );
  AND2_X1 U8799 ( .A1(n6572), .A2(n7102), .ZN(n6437) );
  XNOR2_X1 U8800 ( .A(n8602), .B(n8133), .ZN(n10771) );
  NAND2_X2 U8801 ( .A1(n10242), .A2(n11059), .ZN(n9498) );
  INV_X1 U8802 ( .A(n8588), .ZN(n8609) );
  OR2_X1 U8803 ( .A1(n14547), .A2(n14666), .ZN(n6438) );
  NAND2_X2 U8804 ( .A1(n9701), .A2(n11985), .ZN(n9728) );
  AND3_X1 U8805 ( .A1(n9708), .A2(n9709), .A3(n9710), .ZN(n6439) );
  INV_X1 U8806 ( .A(n9777), .ZN(n11977) );
  NAND2_X1 U8807 ( .A1(n7121), .A2(n7120), .ZN(n6440) );
  NAND2_X1 U8808 ( .A1(n10385), .A2(n7407), .ZN(n6441) );
  AND2_X1 U8809 ( .A1(n7475), .A2(n7474), .ZN(n6443) );
  OR2_X1 U8810 ( .A1(n13881), .A2(n13880), .ZN(n6444) );
  NAND2_X1 U8811 ( .A1(n10582), .A2(n9488), .ZN(n6445) );
  NAND2_X1 U8812 ( .A1(n13319), .A2(n13334), .ZN(n6446) );
  INV_X1 U8813 ( .A(n7338), .ZN(n7337) );
  NAND2_X1 U8814 ( .A1(n13411), .A2(n7800), .ZN(n7338) );
  OR2_X1 U8815 ( .A1(n13946), .A2(n13961), .ZN(n6447) );
  AND2_X1 U8816 ( .A1(n12199), .A2(n11540), .ZN(n6985) );
  AND2_X1 U8817 ( .A1(n7039), .A2(n8007), .ZN(n6448) );
  INV_X2 U8818 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8416) );
  AND2_X1 U8819 ( .A1(n9228), .A2(n9227), .ZN(n6449) );
  AND2_X1 U8820 ( .A1(n9232), .A2(n9231), .ZN(n6450) );
  AND2_X1 U8821 ( .A1(n8913), .A2(n8912), .ZN(n6451) );
  AND4_X1 U8822 ( .A1(n7525), .A2(n7524), .A3(n7650), .A4(n7627), .ZN(n6452)
         );
  AND2_X1 U8824 ( .A1(n7125), .A2(n7126), .ZN(n6454) );
  INV_X1 U8825 ( .A(n13180), .ZN(n13513) );
  NAND2_X1 U8826 ( .A1(n7374), .A2(n11869), .ZN(n13647) );
  INV_X1 U8827 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9476) );
  AND2_X1 U8828 ( .A1(n14040), .A2(n13888), .ZN(n6455) );
  OR2_X1 U8829 ( .A1(n12408), .A2(n8315), .ZN(n6456) );
  OR2_X1 U8830 ( .A1(n7589), .A2(n9929), .ZN(n6457) );
  INV_X1 U8831 ( .A(n9738), .ZN(n11721) );
  INV_X1 U8832 ( .A(n10499), .ZN(n6844) );
  AND2_X1 U8833 ( .A1(n13293), .A2(n6446), .ZN(n6458) );
  OR2_X1 U8834 ( .A1(n13360), .A2(n13112), .ZN(n6459) );
  NAND2_X1 U8835 ( .A1(n11567), .A2(n12990), .ZN(n6460) );
  AND2_X1 U8836 ( .A1(n7301), .A2(n7300), .ZN(n6461) );
  NAND2_X1 U8837 ( .A1(n13337), .A2(n13310), .ZN(n6462) );
  OR2_X1 U8838 ( .A1(n13440), .A2(n13425), .ZN(n6463) );
  INV_X1 U8839 ( .A(n10588), .ZN(n6906) );
  OR2_X1 U8840 ( .A1(n12455), .A2(n12431), .ZN(n6464) );
  AND2_X1 U8841 ( .A1(n14089), .A2(n13884), .ZN(n6465) );
  AND2_X1 U8842 ( .A1(n13590), .A2(n6825), .ZN(n6466) );
  AND2_X1 U8843 ( .A1(n11461), .A2(n15002), .ZN(n6467) );
  AND4_X1 U8844 ( .A1(n8136), .A2(n8647), .A3(n8135), .A4(n8134), .ZN(n6468)
         );
  INV_X1 U8845 ( .A(n13969), .ZN(n6930) );
  INV_X1 U8846 ( .A(n7577), .ZN(n7862) );
  AND2_X1 U8847 ( .A1(n14519), .A2(n6793), .ZN(n6469) );
  INV_X1 U8848 ( .A(n8916), .ZN(n8917) );
  NAND2_X1 U8849 ( .A1(n12247), .A2(n11946), .ZN(n7576) );
  AND2_X1 U8850 ( .A1(n14142), .A2(n13895), .ZN(n6470) );
  OR2_X1 U8851 ( .A1(n8890), .A2(n8891), .ZN(n6471) );
  NAND2_X1 U8852 ( .A1(n9564), .A2(n9563), .ZN(n6472) );
  AND2_X1 U8853 ( .A1(n10582), .A2(n6814), .ZN(n6473) );
  NAND2_X1 U8854 ( .A1(n7732), .A2(n7731), .ZN(n11337) );
  NAND2_X1 U8855 ( .A1(n11755), .A2(n11754), .ZN(n14187) );
  INV_X1 U8856 ( .A(n14187), .ZN(n6936) );
  INV_X1 U8857 ( .A(n12236), .ZN(n7398) );
  AND2_X1 U8858 ( .A1(n11883), .A2(n11882), .ZN(n6474) );
  AND2_X1 U8859 ( .A1(n12230), .A2(n12229), .ZN(n6475) );
  INV_X1 U8860 ( .A(n13983), .ZN(n14153) );
  NAND2_X1 U8861 ( .A1(n11871), .A2(n11870), .ZN(n13983) );
  NAND2_X1 U8862 ( .A1(n9751), .A2(n12625), .ZN(n9694) );
  AND2_X1 U8863 ( .A1(n9530), .A2(n9529), .ZN(n6476) );
  AND2_X1 U8864 ( .A1(n9209), .A2(n9208), .ZN(n6477) );
  OR2_X1 U8865 ( .A1(n14130), .A2(n13897), .ZN(n6478) );
  OR2_X1 U8866 ( .A1(n14170), .A2(n13874), .ZN(n6479) );
  AND2_X1 U8867 ( .A1(n6936), .A2(n13886), .ZN(n6480) );
  NAND2_X1 U8868 ( .A1(n8357), .A2(n8356), .ZN(n11684) );
  AND2_X1 U8869 ( .A1(n8757), .A2(n7018), .ZN(n6481) );
  NAND2_X1 U8870 ( .A1(n11927), .A2(n11926), .ZN(n13896) );
  INV_X1 U8871 ( .A(n13720), .ZN(n13895) );
  NAND2_X1 U8872 ( .A1(n11912), .A2(n11911), .ZN(n13720) );
  INV_X1 U8873 ( .A(n12131), .ZN(n7229) );
  AND2_X1 U8874 ( .A1(n12282), .A2(n12564), .ZN(n6482) );
  AND2_X1 U8875 ( .A1(n6426), .A2(n12427), .ZN(n6483) );
  OR2_X1 U8876 ( .A1(n6930), .A2(n13894), .ZN(n6484) );
  AND2_X1 U8877 ( .A1(n11471), .A2(n9428), .ZN(n6485) );
  AND2_X1 U8878 ( .A1(n14124), .A2(n14123), .ZN(n6486) );
  AND2_X1 U8879 ( .A1(n6433), .A2(n14010), .ZN(n6487) );
  AND2_X1 U8880 ( .A1(n8474), .A2(n8460), .ZN(n6488) );
  NAND2_X1 U8881 ( .A1(n14331), .A2(n12434), .ZN(n6489) );
  AND2_X1 U8882 ( .A1(n14007), .A2(n13875), .ZN(n6490) );
  AND2_X1 U8883 ( .A1(n11790), .A2(n11771), .ZN(n6491) );
  AND2_X1 U8884 ( .A1(n7019), .A2(n8755), .ZN(n6492) );
  AND2_X1 U8885 ( .A1(n11827), .A2(n11811), .ZN(n6493) );
  OR2_X1 U8886 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n8914), .ZN(n6494) );
  OR2_X1 U8887 ( .A1(n13544), .A2(n13333), .ZN(n6495) );
  OR2_X1 U8888 ( .A1(n11835), .A2(n13738), .ZN(n6496) );
  AND2_X1 U8889 ( .A1(n7166), .A2(n6615), .ZN(n6497) );
  AND2_X1 U8890 ( .A1(n13267), .A2(n13242), .ZN(n6498) );
  OR2_X1 U8891 ( .A1(n9181), .A2(n9180), .ZN(n6499) );
  INV_X1 U8892 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9676) );
  INV_X1 U8893 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7538) );
  INV_X1 U8894 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9688) );
  AND2_X1 U8895 ( .A1(n12082), .A2(n7181), .ZN(n6500) );
  NOR2_X1 U8896 ( .A1(n14666), .A2(n13727), .ZN(n6501) );
  NOR2_X1 U8897 ( .A1(n10698), .A2(n13125), .ZN(n6502) );
  NOR2_X1 U8898 ( .A1(n13360), .A2(n13333), .ZN(n6503) );
  NOR2_X1 U8899 ( .A1(n11610), .A2(n13403), .ZN(n6504) );
  NOR2_X1 U8900 ( .A1(n13215), .A2(n13223), .ZN(n6505) );
  NOR2_X1 U8901 ( .A1(n11731), .A2(n11730), .ZN(n6506) );
  NOR2_X1 U8902 ( .A1(n11704), .A2(n13721), .ZN(n6507) );
  NOR2_X1 U8903 ( .A1(n12964), .A2(n12273), .ZN(n6508) );
  INV_X1 U8904 ( .A(n7722), .ZN(n6778) );
  AND2_X1 U8905 ( .A1(n10698), .A2(n9194), .ZN(n6509) );
  OR2_X1 U8906 ( .A1(n9211), .A2(n6477), .ZN(n6510) );
  OR2_X1 U8907 ( .A1(n8826), .A2(n8825), .ZN(n6511) );
  AND3_X1 U8908 ( .A1(n6925), .A2(n6497), .A3(n6388), .ZN(n8150) );
  AND2_X1 U8909 ( .A1(n14142), .A2(n13720), .ZN(n6512) );
  AND2_X1 U8910 ( .A1(n9574), .A2(n9580), .ZN(n6513) );
  NOR2_X1 U8911 ( .A1(n12068), .A2(n11717), .ZN(n6514) );
  NAND2_X1 U8912 ( .A1(n7255), .A2(n6478), .ZN(n7253) );
  INV_X1 U8913 ( .A(n7253), .ZN(n7249) );
  INV_X1 U8914 ( .A(n6874), .ZN(n6873) );
  NOR2_X1 U8915 ( .A1(n14181), .A2(n13887), .ZN(n6874) );
  OR2_X1 U8916 ( .A1(n9216), .A2(n9215), .ZN(n6515) );
  NAND2_X2 U8917 ( .A1(n9711), .A2(n6439), .ZN(n13734) );
  INV_X1 U8918 ( .A(n13734), .ZN(n10881) );
  NAND2_X1 U8919 ( .A1(n11796), .A2(n11795), .ZN(n14175) );
  NAND2_X1 U8920 ( .A1(n7224), .A2(n7221), .ZN(n6516) );
  XOR2_X1 U8921 ( .A(n7414), .B(n7418), .Z(n6517) );
  INV_X1 U8922 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8655) );
  AND2_X1 U8923 ( .A1(n7458), .A2(SI_9_), .ZN(n6518) );
  AND2_X1 U8924 ( .A1(n7449), .A2(SI_6_), .ZN(n6519) );
  INV_X1 U8925 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n12612) );
  INV_X1 U8926 ( .A(n6949), .ZN(n6948) );
  NAND2_X1 U8927 ( .A1(n9364), .A2(n8925), .ZN(n6949) );
  AND2_X1 U8928 ( .A1(n9188), .A2(n9189), .ZN(n6520) );
  INV_X1 U8929 ( .A(n12908), .ZN(n6695) );
  INV_X1 U8930 ( .A(n7143), .ZN(n7142) );
  NAND2_X1 U8931 ( .A1(n11475), .A2(n6456), .ZN(n7143) );
  INV_X1 U8932 ( .A(n7281), .ZN(n7280) );
  NAND2_X1 U8933 ( .A1(n7282), .A2(n9601), .ZN(n7281) );
  INV_X1 U8934 ( .A(n6867), .ZN(n6866) );
  NAND2_X1 U8935 ( .A1(n6870), .A2(n6444), .ZN(n6867) );
  INV_X1 U8936 ( .A(n7156), .ZN(n7155) );
  NAND2_X1 U8937 ( .A1(n7160), .A2(n7161), .ZN(n7156) );
  OR2_X1 U8938 ( .A1(n7785), .A2(n7481), .ZN(n6521) );
  INV_X1 U8939 ( .A(n12059), .ZN(n7237) );
  OR2_X1 U8940 ( .A1(n6826), .A2(n6823), .ZN(n6522) );
  OR2_X1 U8941 ( .A1(n7338), .A2(n6780), .ZN(n6523) );
  INV_X1 U8942 ( .A(n12178), .ZN(n7200) );
  NOR2_X1 U8943 ( .A1(n13466), .A2(n7922), .ZN(n6524) );
  INV_X1 U8944 ( .A(n12070), .ZN(n7242) );
  OR2_X1 U8945 ( .A1(n7180), .A2(n12084), .ZN(n6525) );
  AND2_X1 U8946 ( .A1(n7407), .A2(n9478), .ZN(n6526) );
  INV_X1 U8947 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7537) );
  INV_X1 U8948 ( .A(n12036), .ZN(n7220) );
  INV_X1 U8949 ( .A(n12191), .ZN(n14549) );
  AND2_X1 U8950 ( .A1(n8342), .A2(n8106), .ZN(n6527) );
  OR2_X1 U8951 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n8872), .ZN(n6528) );
  OR2_X1 U8952 ( .A1(n7783), .A2(SI_14_), .ZN(n6529) );
  OR2_X1 U8953 ( .A1(n14411), .A2(n10746), .ZN(n9140) );
  INV_X1 U8954 ( .A(n9140), .ZN(n6687) );
  AND2_X1 U8955 ( .A1(n7361), .A2(n13878), .ZN(n6530) );
  AND2_X1 U8956 ( .A1(n8722), .A2(n7061), .ZN(n6531) );
  NOR2_X1 U8957 ( .A1(n14641), .A2(n13730), .ZN(n6532) );
  AND2_X1 U8958 ( .A1(n9058), .A2(n9054), .ZN(n12810) );
  INV_X1 U8959 ( .A(n12810), .ZN(n12804) );
  INV_X1 U8960 ( .A(n7677), .ZN(n7454) );
  XNOR2_X1 U8961 ( .A(n7455), .B(SI_8_), .ZN(n7677) );
  AND2_X1 U8962 ( .A1(n13267), .A2(n13109), .ZN(n6533) );
  NOR2_X1 U8963 ( .A1(n11363), .A2(n7285), .ZN(n6534) );
  NOR2_X1 U8964 ( .A1(n14032), .A2(n6455), .ZN(n6535) );
  AND2_X1 U8965 ( .A1(n7130), .A2(n7128), .ZN(n6536) );
  AND2_X1 U8966 ( .A1(n8739), .A2(n15029), .ZN(n6537) );
  AND2_X1 U8967 ( .A1(n14153), .A2(n13893), .ZN(n6538) );
  AND2_X1 U8968 ( .A1(n7046), .A2(n6446), .ZN(n6539) );
  AND2_X1 U8969 ( .A1(n8625), .A2(n6920), .ZN(n6540) );
  OR2_X1 U8970 ( .A1(n7338), .A2(n7781), .ZN(n6541) );
  INV_X1 U8971 ( .A(n9011), .ZN(n15018) );
  INV_X1 U8972 ( .A(n6739), .ZN(n6738) );
  OAI21_X1 U8973 ( .B1(n6744), .B2(n6740), .A(n6743), .ZN(n6739) );
  NAND2_X1 U8974 ( .A1(n10774), .A2(n10773), .ZN(n6542) );
  AND2_X1 U8975 ( .A1(n8635), .A2(n8634), .ZN(n6543) );
  AND2_X1 U8976 ( .A1(n9337), .A2(n9336), .ZN(n6544) );
  AND2_X1 U8977 ( .A1(n7537), .A2(n7538), .ZN(n6545) );
  NAND2_X1 U8978 ( .A1(n13752), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6546) );
  OR2_X1 U8979 ( .A1(n6721), .A2(n6434), .ZN(n6547) );
  AND2_X1 U8980 ( .A1(n7823), .A2(n7124), .ZN(n6548) );
  AND2_X1 U8981 ( .A1(n8647), .A2(n7001), .ZN(n6549) );
  INV_X1 U8982 ( .A(n7323), .ZN(n7322) );
  NAND2_X1 U8983 ( .A1(n13522), .A2(n13243), .ZN(n7323) );
  INV_X1 U8984 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n12631) );
  INV_X1 U8985 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9680) );
  AND2_X1 U8986 ( .A1(n6460), .A2(n11024), .ZN(n6550) );
  INV_X1 U8987 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n6615) );
  INV_X1 U8988 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6816) );
  INV_X1 U8989 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n6847) );
  OR2_X1 U8990 ( .A1(n6838), .A2(n6837), .ZN(n6551) );
  OR2_X1 U8991 ( .A1(n7253), .A2(n13898), .ZN(n6552) );
  INV_X1 U8992 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n8190) );
  INV_X1 U8993 ( .A(n7310), .ZN(n7309) );
  OR2_X1 U8994 ( .A1(n11955), .A2(n7311), .ZN(n7310) );
  NAND2_X1 U8995 ( .A1(n9371), .A2(n9370), .ZN(n6553) );
  INV_X1 U8996 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9827) );
  INV_X1 U8997 ( .A(n10330), .ZN(n7120) );
  INV_X1 U8998 ( .A(n14007), .ZN(n6934) );
  AND2_X1 U8999 ( .A1(n13589), .A2(n13590), .ZN(n13587) );
  INV_X1 U9000 ( .A(n13119), .ZN(n11225) );
  INV_X1 U9001 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6632) );
  INV_X1 U9002 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U9003 ( .A1(n13708), .A2(n11736), .ZN(n13626) );
  NAND2_X1 U9004 ( .A1(n11300), .A2(n12197), .ZN(n11515) );
  AND2_X1 U9005 ( .A1(n8352), .A2(n8106), .ZN(n6554) );
  OR2_X1 U9006 ( .A1(n12915), .A2(n12965), .ZN(n6555) );
  AND2_X1 U9007 ( .A1(n11939), .A2(n11938), .ZN(n13904) );
  INV_X1 U9008 ( .A(n13904), .ZN(n13897) );
  AND2_X1 U9009 ( .A1(n8776), .A2(n12808), .ZN(n6556) );
  AND2_X1 U9010 ( .A1(n14483), .A2(n11540), .ZN(n6557) );
  AND2_X1 U9011 ( .A1(n13505), .A2(n13115), .ZN(n6558) );
  AND2_X1 U9012 ( .A1(n12323), .A2(n7016), .ZN(n6559) );
  INV_X1 U9013 ( .A(n6420), .ZN(n6755) );
  OAI21_X1 U9014 ( .B1(n6671), .B2(n6826), .A(n6824), .ZN(n7379) );
  OR2_X1 U9015 ( .A1(n8646), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n6560) );
  NOR2_X1 U9016 ( .A1(n14306), .A2(n14304), .ZN(n6929) );
  INV_X1 U9017 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n12681) );
  INV_X1 U9018 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10443) );
  INV_X1 U9019 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10189) );
  INV_X1 U9020 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6711) );
  INV_X1 U9021 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6630) );
  OR2_X1 U9022 ( .A1(n12915), .A2(n12899), .ZN(n6561) );
  AND2_X1 U9023 ( .A1(n6868), .A2(n6866), .ZN(n6562) );
  AND2_X1 U9024 ( .A1(n11961), .A2(n11960), .ZN(n6563) );
  INV_X1 U9025 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7103) );
  INV_X1 U9026 ( .A(n13384), .ZN(n13356) );
  INV_X1 U9027 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U9028 ( .A1(n7843), .A2(n7842), .ZN(n13375) );
  INV_X1 U9029 ( .A(n13375), .ZN(n6951) );
  NAND2_X1 U9030 ( .A1(n14854), .A2(n13506), .ZN(n13548) );
  NOR2_X1 U9031 ( .A1(n7977), .A2(n7535), .ZN(n8047) );
  NOR2_X2 U9032 ( .A1(n10850), .A2(n11003), .ZN(n6945) );
  NOR2_X1 U9033 ( .A1(n7938), .A2(SI_26_), .ZN(n6564) );
  INV_X1 U9034 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7077) );
  INV_X1 U9035 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6707) );
  AND2_X1 U9036 ( .A1(n6921), .A2(n9022), .ZN(n6565) );
  AND2_X1 U9037 ( .A1(n12461), .A2(n7115), .ZN(n6566) );
  INV_X1 U9038 ( .A(n7565), .ZN(n7366) );
  AND2_X1 U9039 ( .A1(n6839), .A2(n6838), .ZN(n6567) );
  INV_X1 U9040 ( .A(SI_20_), .ZN(n10770) );
  INV_X1 U9041 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12660) );
  INV_X1 U9042 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11470) );
  INV_X1 U9043 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10589) );
  INV_X1 U9044 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10701) );
  AND2_X1 U9045 ( .A1(n10245), .A2(n11471), .ZN(n9151) );
  OR2_X1 U9046 ( .A1(n9497), .A2(n10108), .ZN(n12399) );
  INV_X1 U9047 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U9048 ( .A1(n7637), .A2(n7636), .ZN(n10623) );
  INV_X1 U9049 ( .A(n7010), .ZN(n7012) );
  OR2_X1 U9050 ( .A1(n14236), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6568) );
  XOR2_X1 U9051 ( .A(n6403), .B(P3_REG1_REG_19__SCAN_IN), .Z(n6569) );
  AND2_X1 U9052 ( .A1(n7986), .A2(n10235), .ZN(n6570) );
  INV_X1 U9053 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14246) );
  INV_X1 U9054 ( .A(n14967), .ZN(n12461) );
  AOI22_X1 U9055 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13563), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n7103), .ZN(n8160) );
  INV_X1 U9056 ( .A(n8160), .ZN(n7096) );
  AND2_X1 U9057 ( .A1(n10678), .A2(n7012), .ZN(n6571) );
  OR2_X1 U9058 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13560), .ZN(n6572) );
  INV_X1 U9059 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13563) );
  INV_X1 U9060 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13566) );
  NAND2_X1 U9061 ( .A1(n6403), .A2(n10771), .ZN(n15101) );
  INV_X1 U9062 ( .A(n14376), .ZN(n12477) );
  INV_X1 U9063 ( .A(n9117), .ZN(n11024) );
  INV_X1 U9064 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6961) );
  INV_X1 U9065 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6785) );
  INV_X1 U9066 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8819) );
  INV_X1 U9067 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6669) );
  NOR2_X1 U9068 ( .A1(n14457), .A2(n13521), .ZN(n6697) );
  OR2_X2 U9069 ( .A1(n9701), .A2(n10081), .ZN(n13732) );
  OR2_X1 U9070 ( .A1(n9937), .A2(P1_U3086), .ZN(n10081) );
  NAND2_X1 U9071 ( .A1(n14972), .A2(n14971), .ZN(n14970) );
  NAND2_X1 U9072 ( .A1(n14936), .A2(n14935), .ZN(n14934) );
  NAND2_X1 U9073 ( .A1(n14919), .A2(n14918), .ZN(n14917) );
  NAND2_X1 U9074 ( .A1(n14992), .A2(n12467), .ZN(n12468) );
  INV_X4 U9075 ( .A(n12480), .ZN(n12449) );
  NOR2_X1 U9076 ( .A1(n14366), .A2(n14365), .ZN(n14364) );
  AOI21_X1 U9077 ( .B1(n12470), .B2(n12469), .A(n14334), .ZN(n14357) );
  XNOR2_X1 U9078 ( .A(n12478), .B(n12477), .ZN(n14382) );
  NAND3_X1 U9079 ( .A1(n6652), .A2(n12489), .A3(n6573), .ZN(P3_U3201) );
  NAND2_X1 U9080 ( .A1(n12448), .A2(n14893), .ZN(n14919) );
  NAND2_X1 U9081 ( .A1(n6574), .A2(n6792), .ZN(n14520) );
  NAND3_X1 U9082 ( .A1(n6794), .A2(n6471), .A3(n6793), .ZN(n6574) );
  NOR2_X1 U9083 ( .A1(n14295), .A2(n14294), .ZN(n14293) );
  NAND2_X1 U9084 ( .A1(n14511), .A2(n14510), .ZN(n8886) );
  OAI21_X1 U9085 ( .B1(n15166), .B2(n15165), .A(n6528), .ZN(n6621) );
  OAI22_X1 U9086 ( .A1(n14292), .A2(P2_ADDR_REG_9__SCAN_IN), .B1(n8879), .B2(
        n6783), .ZN(n6782) );
  NAND3_X1 U9087 ( .A1(n6575), .A2(n6635), .A3(n6686), .ZN(n6683) );
  NAND3_X1 U9088 ( .A1(n6654), .A2(n6639), .A3(n12504), .ZN(n6575) );
  NAND2_X1 U9089 ( .A1(n8163), .A2(n8162), .ZN(n12524) );
  NAND2_X1 U9090 ( .A1(n8399), .A2(n8397), .ZN(n6651) );
  NAND2_X1 U9091 ( .A1(n6705), .A2(n6684), .ZN(n8571) );
  OAI22_X1 U9092 ( .A1(n12518), .A2(n9099), .B1(n9450), .B2(n9098), .ZN(n6655)
         );
  NAND2_X1 U9093 ( .A1(n8463), .A2(n8461), .ZN(n8114) );
  NAND2_X1 U9094 ( .A1(n8632), .A2(n8631), .ZN(n6918) );
  NAND2_X1 U9095 ( .A1(n11577), .A2(n11576), .ZN(n11579) );
  AOI21_X1 U9096 ( .B1(n12546), .B2(n9134), .A(n8959), .ZN(n12531) );
  NAND2_X1 U9097 ( .A1(n9691), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n6578) );
  NOR2_X4 U9099 ( .A1(n14023), .A2(n14170), .ZN(n14022) );
  NOR2_X2 U9101 ( .A1(n9696), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U9102 ( .A1(n12531), .A2(n12533), .ZN(n12530) );
  NAND2_X1 U9103 ( .A1(n11509), .A2(n9030), .ZN(n11676) );
  NAND2_X1 U9104 ( .A1(n6915), .A2(n8640), .ZN(n12546) );
  OAI22_X1 U9105 ( .A1(n8953), .A2(n12396), .B1(n8952), .B2(n9137), .ZN(n8954)
         );
  NAND2_X1 U9106 ( .A1(n8113), .A2(n6631), .ZN(n8463) );
  NAND2_X1 U9107 ( .A1(n7078), .A2(n7076), .ZN(n8503) );
  NAND2_X1 U9108 ( .A1(n8112), .A2(n8111), .ZN(n8443) );
  NAND2_X1 U9109 ( .A1(n8116), .A2(n8115), .ZN(n8491) );
  NAND2_X1 U9110 ( .A1(n8110), .A2(n6629), .ZN(n8399) );
  NOR2_X1 U9111 ( .A1(n9103), .A2(n6687), .ZN(n6686) );
  NAND2_X1 U9112 ( .A1(n8593), .A2(n12301), .ZN(n8950) );
  NAND2_X1 U9113 ( .A1(n13707), .A2(n7381), .ZN(n13627) );
  NAND2_X1 U9114 ( .A1(n11667), .A2(n11666), .ZN(n11715) );
  NAND2_X1 U9115 ( .A1(n7593), .A2(n7594), .ZN(n7436) );
  NAND2_X1 U9116 ( .A1(n7491), .A2(n7490), .ZN(n7492) );
  NAND2_X1 U9117 ( .A1(n7341), .A2(n7343), .ZN(n7710) );
  NAND2_X1 U9118 ( .A1(n14226), .A2(n6389), .ZN(n6581) );
  NAND3_X1 U9119 ( .A1(n7507), .A2(n7509), .A3(n7508), .ZN(n7895) );
  NAND2_X1 U9120 ( .A1(n7506), .A2(n7505), .ZN(n7507) );
  NAND2_X1 U9121 ( .A1(n6623), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U9122 ( .A1(n7660), .A2(n7450), .ZN(n7453) );
  NAND2_X1 U9123 ( .A1(n7436), .A2(n7435), .ZN(n7615) );
  NAND2_X1 U9124 ( .A1(n7441), .A2(n7440), .ZN(n7625) );
  OAI211_X1 U9125 ( .C1(n13947), .C2(n6552), .A(n7245), .B(n7247), .ZN(n14122)
         );
  NAND2_X1 U9126 ( .A1(n6583), .A2(n6586), .ZN(n6585) );
  NAND3_X1 U9127 ( .A1(n7189), .A2(n7184), .A3(n7188), .ZN(n6583) );
  OAI21_X1 U9128 ( .B1(n7208), .B2(n7210), .A(n12113), .ZN(n7207) );
  NOR2_X1 U9129 ( .A1(n13899), .A2(n7250), .ZN(n7246) );
  OAI21_X1 U9130 ( .B1(n12110), .B2(n7208), .A(n7206), .ZN(n12114) );
  AOI22_X1 U9131 ( .A1(n12139), .A2(n12138), .B1(n12137), .B2(n12136), .ZN(
        n12144) );
  NAND2_X1 U9132 ( .A1(n6624), .A2(n7347), .ZN(n7660) );
  INV_X1 U9133 ( .A(n7492), .ZN(n7493) );
  OR2_X1 U9134 ( .A1(n13440), .A2(n14428), .ZN(n6689) );
  AOI21_X1 U9135 ( .B1(n6763), .B2(n6765), .A(n9415), .ZN(n6762) );
  NOR4_X1 U9136 ( .A1(n13920), .A2(n13931), .A3(n6622), .A4(n12204), .ZN(
        n12207) );
  NAND2_X1 U9137 ( .A1(n6585), .A2(n6584), .ZN(P1_U3242) );
  XNOR2_X1 U9138 ( .A(n6670), .B(n12226), .ZN(n12217) );
  NAND2_X1 U9139 ( .A1(n6587), .A2(n9439), .ZN(P2_U3328) );
  OAI21_X1 U9140 ( .B1(n6693), .B2(n9435), .A(n9434), .ZN(n6587) );
  INV_X1 U9141 ( .A(n7251), .ZN(n7250) );
  NAND2_X1 U9142 ( .A1(n12114), .A2(n12115), .ZN(n12118) );
  NAND2_X1 U9143 ( .A1(n7633), .A2(n7346), .ZN(n6624) );
  NOR2_X1 U9144 ( .A1(n13976), .A2(n6538), .ZN(n13962) );
  NAND2_X1 U9145 ( .A1(n6595), .A2(n6592), .ZN(n14211) );
  INV_X1 U9146 ( .A(n7207), .ZN(n7206) );
  OAI21_X1 U9147 ( .B1(n12144), .B2(n12143), .A(n12142), .ZN(n12146) );
  NAND2_X1 U9148 ( .A1(n7255), .A2(n7254), .ZN(n13918) );
  OAI21_X1 U9149 ( .B1(n14133), .B2(n14635), .A(n6594), .ZN(n6593) );
  NAND2_X1 U9150 ( .A1(n14018), .A2(n14021), .ZN(n14017) );
  AOI21_X1 U9151 ( .B1(n12189), .B2(n11080), .A(n12191), .ZN(n6971) );
  NAND3_X2 U9152 ( .A1(n9714), .A2(n6928), .A3(n6496), .ZN(n11992) );
  NAND2_X1 U9153 ( .A1(n13865), .A2(n13882), .ZN(n6590) );
  OAI21_X2 U9154 ( .B1(n14076), .B2(n13871), .A(n13870), .ZN(n14048) );
  NAND2_X1 U9155 ( .A1(n13980), .A2(n13979), .ZN(n13978) );
  INV_X1 U9156 ( .A(n6977), .ZN(n6976) );
  AOI22_X1 U9157 ( .A1(n13996), .A2(n13877), .B1(n13876), .B2(n14159), .ZN(
        n13980) );
  OAI21_X2 U9158 ( .B1(n12183), .B2(n11135), .A(n10870), .ZN(n14588) );
  NAND2_X1 U9159 ( .A1(n6968), .A2(n6969), .ZN(n11161) );
  NAND2_X1 U9160 ( .A1(n11170), .A2(n11169), .ZN(n11274) );
  NAND2_X1 U9161 ( .A1(n10881), .A2(n6591), .ZN(n10870) );
  NAND2_X1 U9162 ( .A1(n7192), .A2(n7195), .ZN(n7187) );
  NAND3_X1 U9163 ( .A1(n6689), .A2(n13439), .A3(n13438), .ZN(n13518) );
  INV_X1 U9164 ( .A(n7328), .ZN(n7327) );
  NAND3_X1 U9165 ( .A1(n7369), .A2(n7372), .A3(n6903), .ZN(n6610) );
  NAND2_X1 U9166 ( .A1(n11221), .A2(n9554), .ZN(n11341) );
  NAND2_X1 U9167 ( .A1(n13090), .A2(n7309), .ZN(n11963) );
  INV_X1 U9168 ( .A(n7292), .ZN(n7288) );
  INV_X1 U9169 ( .A(n6713), .ZN(n6717) );
  OAI22_X1 U9170 ( .A1(n7250), .A2(n7248), .B1(n13899), .B2(n7251), .ZN(n7247)
         );
  INV_X1 U9171 ( .A(n6470), .ZN(n7257) );
  AOI21_X1 U9172 ( .B1(n7330), .B2(n7329), .A(n6533), .ZN(n7328) );
  OR2_X1 U9173 ( .A1(n8845), .A2(n8844), .ZN(n6682) );
  NOR2_X1 U9174 ( .A1(n8896), .A2(n8895), .ZN(n8897) );
  AOI22_X1 U9175 ( .A1(n14545), .A2(P3_ADDR_REG_15__SCAN_IN), .B1(n8904), .B2(
        n8903), .ZN(n8908) );
  NAND2_X1 U9176 ( .A1(n8972), .A2(n9122), .ZN(n8730) );
  OAI22_X1 U9177 ( .A1(n8954), .A2(n9119), .B1(n8956), .B2(n8955), .ZN(n6611)
         );
  NAND2_X1 U9178 ( .A1(n12914), .A2(n6555), .ZN(P3_U3454) );
  NAND2_X1 U9179 ( .A1(n12837), .A2(n6561), .ZN(P3_U3486) );
  NAND2_X1 U9180 ( .A1(n9652), .A2(n6601), .ZN(n8985) );
  INV_X1 U9181 ( .A(n15077), .ZN(n6601) );
  NAND2_X1 U9182 ( .A1(n8623), .A2(n9008), .ZN(n15019) );
  NAND2_X2 U9183 ( .A1(n8760), .A2(n11613), .ZN(n11636) );
  NAND2_X1 U9184 ( .A1(n8727), .A2(n6602), .ZN(n8732) );
  NAND2_X1 U9185 ( .A1(n11037), .A2(n11036), .ZN(n11035) );
  NAND2_X1 U9186 ( .A1(n12271), .A2(n12270), .ZN(n12269) );
  NAND2_X1 U9187 ( .A1(n12287), .A2(n12286), .ZN(n12285) );
  INV_X1 U9188 ( .A(n12307), .ZN(n6605) );
  OAI21_X1 U9189 ( .B1(n12325), .B2(n7015), .A(n7013), .ZN(n12366) );
  INV_X1 U9190 ( .A(n8737), .ZN(n7011) );
  NAND2_X2 U9191 ( .A1(n6608), .A2(n6607), .ZN(n8531) );
  INV_X1 U9192 ( .A(n10354), .ZN(n9742) );
  NAND2_X1 U9193 ( .A1(n9743), .A2(n9720), .ZN(n10354) );
  NOR2_X2 U9194 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9468) );
  NAND2_X1 U9195 ( .A1(n7386), .A2(n6542), .ZN(n6819) );
  NAND3_X1 U9196 ( .A1(n6905), .A2(n6904), .A3(n6674), .ZN(n6715) );
  NAND2_X1 U9197 ( .A1(n6610), .A2(n7496), .ZN(n7497) );
  NAND2_X1 U9198 ( .A1(n6717), .A2(n6715), .ZN(n6716) );
  NAND3_X1 U9199 ( .A1(n6986), .A2(n7268), .A3(n9488), .ZN(n9690) );
  NOR2_X2 U9200 ( .A1(n9487), .A2(n9486), .ZN(n9488) );
  XNOR2_X1 U9201 ( .A(n6611), .B(n6403), .ZN(n9146) );
  NOR2_X2 U9202 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9484) );
  NAND2_X1 U9203 ( .A1(n10872), .A2(n12007), .ZN(n11124) );
  NAND2_X1 U9204 ( .A1(n11063), .A2(n11062), .ZN(n11079) );
  AOI211_X2 U9205 ( .C1(n13450), .C2(n14440), .A(n13449), .B(n13448), .ZN(
        n13520) );
  XNOR2_X1 U9206 ( .A(n13222), .B(n13227), .ZN(n6663) );
  NAND3_X1 U9207 ( .A1(n8894), .A2(n6789), .A3(n8893), .ZN(n6787) );
  XNOR2_X1 U9208 ( .A(n8846), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n8858) );
  NOR2_X1 U9209 ( .A1(n15162), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n8865) );
  XNOR2_X1 U9210 ( .A(n8863), .B(n8862), .ZN(n15162) );
  OAI21_X1 U9211 ( .B1(n12125), .B2(n7232), .A(n6616), .ZN(n12132) );
  NAND3_X1 U9212 ( .A1(n6960), .A2(n6959), .A3(n6618), .ZN(n6617) );
  NAND2_X1 U9213 ( .A1(n7507), .A2(n7509), .ZN(n11833) );
  INV_X1 U9214 ( .A(n14513), .ZN(n6962) );
  NOR2_X1 U9215 ( .A1(n14526), .A2(n14527), .ZN(n14525) );
  NOR2_X1 U9216 ( .A1(n14519), .A2(n14520), .ZN(n14518) );
  NOR2_X1 U9217 ( .A1(n7690), .A2(n7677), .ZN(n7342) );
  INV_X1 U9218 ( .A(n9427), .ZN(n9431) );
  NAND2_X1 U9219 ( .A1(n6646), .A2(n6716), .ZN(n9427) );
  XNOR2_X2 U9220 ( .A(n14142), .B(n13720), .ZN(n13946) );
  INV_X1 U9221 ( .A(n7476), .ZN(n6623) );
  INV_X1 U9222 ( .A(n7497), .ZN(n6625) );
  NOR2_X1 U9223 ( .A1(n9368), .A2(n7135), .ZN(n6904) );
  AOI22_X2 U9224 ( .A1(n9385), .A2(n6633), .B1(n6664), .B2(n6665), .ZN(n9379)
         );
  AOI21_X1 U9225 ( .B1(n13180), .B2(n9369), .A(n6634), .ZN(n6633) );
  AND2_X1 U9226 ( .A1(n13183), .A2(n9167), .ZN(n6634) );
  NAND2_X1 U9227 ( .A1(n7476), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7437) );
  AND2_X2 U9228 ( .A1(n6925), .A2(n7003), .ZN(n8598) );
  NAND2_X1 U9229 ( .A1(n6550), .A2(n6997), .ZN(n6996) );
  NOR2_X1 U9230 ( .A1(n7011), .A2(n10679), .ZN(n7009) );
  NAND2_X1 U9231 ( .A1(n6638), .A2(n8109), .ZN(n8384) );
  NOR2_X1 U9232 ( .A1(n12563), .A2(n6917), .ZN(n6916) );
  NAND2_X1 U9233 ( .A1(n8366), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U9234 ( .A1(n7065), .A2(n8087), .ZN(n8197) );
  NAND2_X1 U9235 ( .A1(n12577), .A2(n6916), .ZN(n6915) );
  NOR2_X2 U9236 ( .A1(n14322), .A2(n14321), .ZN(n14320) );
  XNOR2_X1 U9237 ( .A(n8852), .B(n6785), .ZN(n15172) );
  NAND2_X1 U9238 ( .A1(n15172), .A2(n15173), .ZN(n6784) );
  NAND2_X1 U9239 ( .A1(n7070), .A2(n7073), .ZN(n9118) );
  NAND2_X1 U9240 ( .A1(n7066), .A2(n15101), .ZN(n7070) );
  OR2_X1 U9241 ( .A1(n9097), .A2(n9078), .ZN(n6639) );
  NAND2_X1 U9242 ( .A1(n8414), .A2(n8412), .ZN(n8112) );
  NAND2_X1 U9243 ( .A1(n12575), .A2(n12578), .ZN(n12577) );
  NAND2_X1 U9244 ( .A1(n6935), .A2(n14040), .ZN(n14023) );
  NOR2_X2 U9245 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9467) );
  NAND2_X1 U9246 ( .A1(n6937), .A2(n6936), .ZN(n14069) );
  INV_X1 U9247 ( .A(n6640), .ZN(n13901) );
  NOR2_X2 U9248 ( .A1(n13900), .A2(n14126), .ZN(n6640) );
  NAND2_X1 U9249 ( .A1(n6419), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8185) );
  INV_X1 U9250 ( .A(n12160), .ZN(n6979) );
  NAND2_X1 U9251 ( .A1(n8176), .A2(n8187), .ZN(n7065) );
  NAND2_X1 U9252 ( .A1(n14895), .A2(n14892), .ZN(n12448) );
  NAND2_X1 U9253 ( .A1(n12444), .A2(n12445), .ZN(n14895) );
  XNOR2_X1 U9254 ( .A(n10651), .B(n10652), .ZN(n10527) );
  NOR2_X1 U9255 ( .A1(n14388), .A2(n6642), .ZN(n12438) );
  XNOR2_X1 U9256 ( .A(n12431), .B(n12455), .ZN(n14925) );
  NOR2_X1 U9257 ( .A1(n14890), .A2(n14889), .ZN(n14888) );
  NAND2_X1 U9258 ( .A1(n8056), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6943) );
  AND2_X1 U9259 ( .A1(n9509), .A2(n9510), .ZN(n10192) );
  NAND2_X1 U9260 ( .A1(n6645), .A2(n6563), .ZN(P2_U3186) );
  NAND2_X1 U9261 ( .A1(n11962), .A2(n11963), .ZN(n6645) );
  NOR2_X2 U9262 ( .A1(n11949), .A2(n11948), .ZN(n13092) );
  NOR2_X2 U9263 ( .A1(n9625), .A2(n9624), .ZN(n11949) );
  NAND2_X1 U9264 ( .A1(n12367), .A2(n8779), .ZN(n12287) );
  NAND2_X1 U9265 ( .A1(n11265), .A2(n8752), .ZN(n11459) );
  NAND2_X1 U9266 ( .A1(n12339), .A2(n8784), .ZN(n12307) );
  NAND2_X1 U9268 ( .A1(n13418), .A2(n13417), .ZN(n13421) );
  NAND2_X1 U9269 ( .A1(n6952), .A2(n6951), .ZN(n13359) );
  NAND2_X1 U9270 ( .A1(n11357), .A2(n14444), .ZN(n11416) );
  INV_X1 U9271 ( .A(n6953), .ZN(n13335) );
  NOR2_X2 U9272 ( .A1(n13181), .A2(n13394), .ZN(n13429) );
  NAND2_X1 U9273 ( .A1(n6717), .A2(n6544), .ZN(n6646) );
  NAND2_X1 U9274 ( .A1(n13919), .A2(n6667), .ZN(n6666) );
  INV_X1 U9275 ( .A(n9379), .ZN(n6905) );
  INV_X1 U9276 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8091) );
  NAND2_X1 U9277 ( .A1(n8571), .A2(n8569), .ZN(n8121) );
  OR2_X2 U9278 ( .A1(n12524), .A2(n12536), .ZN(n9094) );
  NAND2_X1 U9279 ( .A1(n12439), .A2(n14385), .ZN(n6652) );
  NAND2_X1 U9280 ( .A1(n6836), .A2(n6551), .ZN(n12428) );
  INV_X1 U9281 ( .A(n6655), .ZN(n6654) );
  INV_X1 U9282 ( .A(n7083), .ZN(n7082) );
  NAND2_X1 U9283 ( .A1(n11543), .A2(n11542), .ZN(n14107) );
  NOR2_X2 U9284 ( .A1(n6438), .A2(n12046), .ZN(n11211) );
  INV_X1 U9285 ( .A(n6929), .ZN(n14307) );
  NAND2_X4 U9286 ( .A1(n11835), .A2(n6396), .ZN(n12160) );
  NAND2_X1 U9287 ( .A1(n7910), .A2(n7911), .ZN(n11850) );
  NAND2_X1 U9288 ( .A1(n9382), .A2(n9381), .ZN(n6664) );
  NOR2_X2 U9289 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n9483) );
  INV_X1 U9290 ( .A(n7044), .ZN(n7042) );
  NOR2_X1 U9291 ( .A1(n6458), .A2(n6422), .ZN(n7045) );
  OAI21_X1 U9292 ( .B1(n9828), .B2(n6669), .A(n6668), .ZN(n7451) );
  NAND4_X1 U9293 ( .A1(n12207), .A2(n6387), .A3(n12206), .A4(n13898), .ZN(
        n6670) );
  NAND2_X1 U9294 ( .A1(n13638), .A2(n13639), .ZN(n13637) );
  XNOR2_X1 U9295 ( .A(n6820), .B(n11721), .ZN(n9717) );
  NAND2_X1 U9296 ( .A1(n7383), .A2(n10389), .ZN(n7386) );
  NAND2_X1 U9297 ( .A1(n14282), .A2(n14281), .ZN(n6672) );
  INV_X1 U9298 ( .A(n6782), .ZN(n14295) );
  AOI21_X1 U9299 ( .B1(n9431), .B2(n10245), .A(n6673), .ZN(n9435) );
  NAND2_X1 U9300 ( .A1(n13710), .A2(n13709), .ZN(n13707) );
  NAND2_X1 U9301 ( .A1(n6806), .A2(n6805), .ZN(n11733) );
  NAND2_X1 U9302 ( .A1(n6797), .A2(n7373), .ZN(n13618) );
  NOR2_X1 U9303 ( .A1(n12804), .A2(n6911), .ZN(n6910) );
  NAND2_X1 U9304 ( .A1(n6962), .A2(n6961), .ZN(n6794) );
  NOR2_X1 U9305 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8861), .ZN(n8828) );
  INV_X1 U9306 ( .A(n14518), .ZN(n8894) );
  NAND2_X1 U9307 ( .A1(n8882), .A2(n8883), .ZN(n6679) );
  INV_X1 U9308 ( .A(n14293), .ZN(n6680) );
  NOR2_X1 U9309 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8871), .ZN(n8832) );
  INV_X1 U9310 ( .A(n14320), .ZN(n8913) );
  NAND2_X1 U9311 ( .A1(n6683), .A2(n9106), .ZN(n9108) );
  NAND2_X1 U9312 ( .A1(n8476), .A2(n8475), .ZN(n8116) );
  NAND2_X1 U9313 ( .A1(n8114), .A2(n6706), .ZN(n8476) );
  NAND2_X1 U9314 ( .A1(n9118), .A2(n9117), .ZN(n9145) );
  OAI21_X1 U9315 ( .B1(n8224), .B2(n7082), .A(n7080), .ZN(n8097) );
  AOI21_X1 U9316 ( .B1(n6976), .B2(n6978), .A(n6532), .ZN(n6974) );
  OAI21_X1 U9317 ( .B1(n12186), .B2(n6978), .A(n12188), .ZN(n6977) );
  NAND2_X1 U9318 ( .A1(n11161), .A2(n12193), .ZN(n11163) );
  NAND2_X1 U9319 ( .A1(n10372), .A2(n9516), .ZN(n10571) );
  NAND2_X1 U9320 ( .A1(n10571), .A2(n10572), .ZN(n10570) );
  NAND2_X1 U9321 ( .A1(n6943), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6942) );
  OAI21_X2 U9322 ( .B1(n13064), .B2(n7281), .A(n7277), .ZN(n9611) );
  INV_X1 U9323 ( .A(n7296), .ZN(n7295) );
  NAND2_X1 U9324 ( .A1(n9432), .A2(n9433), .ZN(n6693) );
  NAND2_X1 U9325 ( .A1(n9359), .A2(n9358), .ZN(n9388) );
  XNOR2_X2 U9326 ( .A(n14135), .B(n13879), .ZN(n13931) );
  INV_X1 U9327 ( .A(n7851), .ZN(n6903) );
  NAND2_X2 U9328 ( .A1(n6695), .A2(n6694), .ZN(n8974) );
  INV_X2 U9329 ( .A(n15083), .ZN(n6694) );
  NAND2_X1 U9330 ( .A1(n6921), .A2(n6540), .ZN(n11509) );
  NAND2_X1 U9331 ( .A1(n6698), .A2(n6696), .ZN(P2_U3493) );
  OR2_X1 U9332 ( .A1(n13520), .A2(n14450), .ZN(n6698) );
  NAND2_X1 U9333 ( .A1(n6909), .A2(n6912), .ZN(n12794) );
  NAND2_X1 U9334 ( .A1(n6922), .A2(n9018), .ZN(n6921) );
  OAI21_X1 U9335 ( .B1(n9146), .B2(n9145), .A(n7067), .ZN(n6919) );
  NAND2_X1 U9336 ( .A1(n7431), .A2(n9846), .ZN(n6699) );
  OAI21_X1 U9337 ( .B1(n14127), .B2(n14644), .A(n6702), .ZN(n14210) );
  OAI21_X1 U9338 ( .B1(n6715), .B2(n6553), .A(n6714), .ZN(n6713) );
  NAND2_X1 U9339 ( .A1(n6894), .A2(n6893), .ZN(n7483) );
  AOI21_X1 U9340 ( .B1(n13180), .B2(n9167), .A(n9386), .ZN(n6704) );
  NAND2_X1 U9341 ( .A1(n8558), .A2(n8556), .ZN(n6705) );
  NAND2_X1 U9342 ( .A1(n8384), .A2(n8382), .ZN(n8110) );
  NAND2_X1 U9343 ( .A1(n8443), .A2(n8441), .ZN(n8113) );
  AND2_X2 U9344 ( .A1(n7075), .A2(n7074), .ZN(n8518) );
  NAND2_X1 U9345 ( .A1(n8491), .A2(n8489), .ZN(n7078) );
  NAND2_X1 U9346 ( .A1(n6919), .A2(n9150), .ZN(P3_U3296) );
  NAND2_X1 U9347 ( .A1(n7272), .A2(n7270), .ZN(n10372) );
  NAND2_X1 U9348 ( .A1(n7284), .A2(n7283), .ZN(n11557) );
  NAND2_X1 U9349 ( .A1(n7286), .A2(n7289), .ZN(n10750) );
  NOR2_X1 U9350 ( .A1(n13004), .A2(n7273), .ZN(n7269) );
  NAND2_X1 U9351 ( .A1(n6719), .A2(n6718), .ZN(n9306) );
  NAND3_X1 U9352 ( .A1(n6720), .A2(n6432), .A3(n6547), .ZN(n6719) );
  INV_X1 U9353 ( .A(n9299), .ZN(n6720) );
  INV_X1 U9354 ( .A(n9302), .ZN(n6721) );
  NAND3_X1 U9355 ( .A1(n9182), .A2(n6724), .A3(n6499), .ZN(n6722) );
  NAND2_X1 U9356 ( .A1(n6722), .A2(n6723), .ZN(n7139) );
  NAND2_X1 U9357 ( .A1(n6725), .A2(n6728), .ZN(n9333) );
  NAND2_X1 U9358 ( .A1(n6727), .A2(n6726), .ZN(n6725) );
  INV_X1 U9359 ( .A(n9323), .ZN(n6726) );
  NOR2_X1 U9360 ( .A1(n9322), .A2(n6729), .ZN(n6727) );
  MUX2_X1 U9361 ( .A(n9931), .B(n13577), .S(n7589), .Z(n10014) );
  NAND2_X1 U9362 ( .A1(n9207), .A2(n6417), .ZN(n6731) );
  NAND2_X1 U9363 ( .A1(n9230), .A2(n6741), .ZN(n6734) );
  OAI21_X1 U9364 ( .B1(n9230), .B2(n6739), .A(n6735), .ZN(n9240) );
  NAND2_X1 U9365 ( .A1(n13372), .A2(n6750), .ZN(n6748) );
  OAI21_X1 U9366 ( .B1(n13372), .B2(n6752), .A(n6750), .ZN(n13317) );
  NAND3_X1 U9367 ( .A1(n6462), .A2(n6753), .A3(n6755), .ZN(n6751) );
  NAND4_X1 U9368 ( .A1(n9397), .A2(n9398), .A3(n9396), .A4(n6759), .ZN(n9399)
         );
  NAND2_X1 U9369 ( .A1(n7325), .A2(n6763), .ZN(n6761) );
  NAND2_X1 U9370 ( .A1(n6761), .A2(n6762), .ZN(n8689) );
  NAND2_X1 U9371 ( .A1(n7325), .A2(n7324), .ZN(n6767) );
  NAND3_X1 U9372 ( .A1(n7743), .A2(n7532), .A3(n7339), .ZN(n8056) );
  NAND2_X1 U9373 ( .A1(n8893), .A2(n8894), .ZN(n8901) );
  XNOR2_X1 U9374 ( .A(n6790), .B(n6517), .ZN(SUB_1596_U4) );
  NAND3_X1 U9375 ( .A1(n8912), .A2(n8913), .A3(n8916), .ZN(n6959) );
  XNOR2_X1 U9376 ( .A(n8872), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15166) );
  NAND2_X2 U9377 ( .A1(n6796), .A2(n11900), .ZN(n13698) );
  NAND2_X1 U9378 ( .A1(n13618), .A2(n13620), .ZN(n6796) );
  NAND2_X1 U9379 ( .A1(n13580), .A2(n7375), .ZN(n6797) );
  NAND2_X1 U9380 ( .A1(n6801), .A2(n6798), .ZN(P1_U3214) );
  NOR2_X1 U9381 ( .A1(n13939), .A2(n13718), .ZN(n6800) );
  NAND2_X1 U9382 ( .A1(n6802), .A2(n14470), .ZN(n6801) );
  XNOR2_X1 U9383 ( .A(n6803), .B(n12231), .ZN(n6802) );
  NAND2_X1 U9384 ( .A1(n7394), .A2(n11918), .ZN(n6803) );
  NAND2_X1 U9385 ( .A1(n11715), .A2(n6807), .ZN(n6806) );
  OR2_X1 U9386 ( .A1(n10582), .A2(n9668), .ZN(n6813) );
  INV_X1 U9387 ( .A(n9717), .ZN(n9718) );
  NAND3_X1 U9388 ( .A1(n6829), .A2(n6830), .A3(n6828), .ZN(n14961) );
  NAND4_X1 U9389 ( .A1(n6829), .A2(n6830), .A3(n6828), .A4(
        P3_REG2_REG_13__SCAN_IN), .ZN(n6832) );
  INV_X1 U9390 ( .A(n6832), .ZN(n14960) );
  NAND2_X1 U9391 ( .A1(n6840), .A2(n6483), .ZN(n6836) );
  INV_X1 U9392 ( .A(n6840), .ZN(n10653) );
  INV_X1 U9393 ( .A(n10493), .ZN(n6841) );
  NAND3_X1 U9394 ( .A1(n6847), .A2(n8178), .A3(n8190), .ZN(n6845) );
  OAI21_X1 U9395 ( .B1(n10891), .B2(n6854), .A(n14566), .ZN(n6849) );
  INV_X1 U9396 ( .A(n6849), .ZN(n6851) );
  NAND2_X1 U9397 ( .A1(n14298), .A2(n6860), .ZN(n6859) );
  NAND2_X1 U9398 ( .A1(n14552), .A2(n6862), .ZN(n11206) );
  NAND2_X1 U9399 ( .A1(n14049), .A2(n6872), .ZN(n6871) );
  NAND2_X1 U9400 ( .A1(n6871), .A2(n6487), .ZN(n14008) );
  NAND4_X1 U9401 ( .A1(n7424), .A2(n13851), .A3(n14257), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U9402 ( .A1(n7625), .A2(n7442), .ZN(n6879) );
  INV_X1 U9403 ( .A(n9355), .ZN(n6881) );
  NAND2_X1 U9404 ( .A1(n7471), .A2(n6895), .ZN(n6894) );
  NAND2_X1 U9405 ( .A1(n12823), .A2(n6910), .ZN(n6909) );
  NAND2_X1 U9406 ( .A1(n12577), .A2(n8962), .ZN(n12562) );
  INV_X1 U9407 ( .A(n6915), .ZN(n8639) );
  INV_X1 U9408 ( .A(n8962), .ZN(n6917) );
  INV_X1 U9409 ( .A(n11315), .ZN(n6922) );
  NAND3_X1 U9410 ( .A1(n6497), .A2(n6923), .A3(n6388), .ZN(n12974) );
  INV_X2 U9411 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6927) );
  NOR2_X2 U9412 ( .A1(n14307), .A2(n12068), .ZN(n11543) );
  NOR2_X2 U9413 ( .A1(n14069), .A2(n14060), .ZN(n6935) );
  NAND2_X2 U9414 ( .A1(n6457), .A2(n6940), .ZN(n10238) );
  NOR2_X2 U9415 ( .A1(n11337), .A2(n11239), .ZN(n11357) );
  NAND2_X1 U9416 ( .A1(n13216), .A2(n6948), .ZN(n13189) );
  NAND2_X1 U9417 ( .A1(n13216), .A2(n6947), .ZN(n13187) );
  AND2_X1 U9418 ( .A1(n13216), .A2(n8925), .ZN(n8714) );
  NOR2_X2 U9419 ( .A1(n13421), .A2(n13500), .ZN(n6952) );
  NOR2_X2 U9420 ( .A1(n11595), .A2(n11610), .ZN(n13418) );
  NAND2_X1 U9421 ( .A1(n6956), .A2(n8820), .ZN(n6954) );
  INV_X1 U9422 ( .A(n8847), .ZN(n6956) );
  NAND3_X1 U9423 ( .A1(n6956), .A2(n6957), .A3(n8821), .ZN(n6955) );
  NAND3_X1 U9424 ( .A1(n6959), .A2(n6960), .A3(n6958), .ZN(n14254) );
  INV_X2 U9425 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U9426 ( .A1(n11079), .A2(n6971), .ZN(n6968) );
  NAND2_X1 U9427 ( .A1(n11124), .A2(n6976), .ZN(n6973) );
  NAND2_X1 U9428 ( .A1(n9693), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9689) );
  NAND4_X1 U9429 ( .A1(n9488), .A2(n6986), .A3(n9676), .A4(n7268), .ZN(n9693)
         );
  NAND3_X1 U9430 ( .A1(n8732), .A2(n8728), .A3(n8731), .ZN(n9649) );
  OAI211_X1 U9431 ( .C1(n6987), .C2(n12900), .A(n9649), .B(n9648), .ZN(n9650)
         );
  NAND2_X1 U9432 ( .A1(n11636), .A2(n6992), .ZN(n6988) );
  NAND2_X1 U9433 ( .A1(n6988), .A2(n6989), .ZN(n12271) );
  NAND2_X1 U9434 ( .A1(n8658), .A2(n12994), .ZN(n6999) );
  NAND2_X1 U9435 ( .A1(n8649), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8648) );
  NAND3_X1 U9436 ( .A1(n7174), .A2(n8212), .A3(n8127), .ZN(n7006) );
  OAI21_X2 U9437 ( .B1(n10680), .B2(n7010), .A(n7008), .ZN(n10898) );
  NAND2_X1 U9438 ( .A1(n11497), .A2(n8757), .ZN(n8759) );
  INV_X1 U9439 ( .A(n11495), .ZN(n7019) );
  INV_X1 U9440 ( .A(n7986), .ZN(n9394) );
  OAI21_X1 U9441 ( .B1(n7986), .B2(n10231), .A(n10230), .ZN(n10534) );
  NAND2_X1 U9442 ( .A1(n10595), .A2(n6421), .ZN(n7022) );
  NAND2_X1 U9443 ( .A1(n7022), .A2(n7023), .ZN(n10706) );
  OAI21_X1 U9444 ( .B1(n13238), .B2(n7028), .A(n7026), .ZN(n8032) );
  OAI21_X2 U9445 ( .B1(n8030), .B2(n7034), .A(n9389), .ZN(n7033) );
  INV_X1 U9446 ( .A(n8029), .ZN(n7034) );
  NAND2_X1 U9447 ( .A1(n8032), .A2(n9415), .ZN(n8705) );
  NAND2_X1 U9448 ( .A1(n13444), .A2(n13223), .ZN(n7035) );
  NAND2_X1 U9449 ( .A1(n8707), .A2(n7062), .ZN(n7060) );
  AOI21_X1 U9450 ( .B1(n8707), .B2(n13352), .A(n7064), .ZN(n13439) );
  AND3_X4 U9451 ( .A1(n6452), .A2(n7612), .A3(n7528), .ZN(n7743) );
  NAND2_X1 U9452 ( .A1(n9115), .A2(n9116), .ZN(n7073) );
  INV_X1 U9453 ( .A(n9115), .ZN(n7066) );
  XNOR2_X1 U9454 ( .A(n9143), .B(n6403), .ZN(n7072) );
  NAND2_X1 U9455 ( .A1(n7069), .A2(n7068), .ZN(n7067) );
  NAND3_X1 U9456 ( .A1(n7070), .A2(n9144), .A3(n7073), .ZN(n7069) );
  NAND2_X1 U9457 ( .A1(n8951), .A2(n9113), .ZN(n9119) );
  NAND2_X1 U9458 ( .A1(n8161), .A2(n7095), .ZN(n7094) );
  NAND2_X1 U9459 ( .A1(n7104), .A2(n7102), .ZN(n8585) );
  AOI21_X2 U9460 ( .B1(n8542), .B2(n13574), .A(n8120), .ZN(n8558) );
  INV_X1 U9461 ( .A(n7106), .ZN(n14977) );
  XNOR2_X1 U9462 ( .A(n7121), .B(n10330), .ZN(n10476) );
  INV_X1 U9463 ( .A(n10341), .ZN(n7119) );
  NAND2_X1 U9464 ( .A1(n7824), .A2(n6548), .ZN(n7123) );
  NAND2_X1 U9465 ( .A1(n9283), .A2(n6536), .ZN(n7125) );
  AOI21_X1 U9466 ( .B1(n9283), .B2(n7130), .A(n7129), .ZN(n9293) );
  NOR2_X1 U9467 ( .A1(n9321), .A2(n9320), .ZN(n9322) );
  NAND2_X2 U9468 ( .A1(n10245), .A2(n6485), .ZN(n9190) );
  NAND2_X1 U9469 ( .A1(n6419), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U9470 ( .A1(n8515), .A2(n7148), .ZN(n7145) );
  NAND2_X1 U9471 ( .A1(n7145), .A2(n7146), .ZN(n12560) );
  OAI21_X2 U9472 ( .B1(n8351), .B2(n7156), .A(n7153), .ZN(n11625) );
  NAND2_X1 U9473 ( .A1(n8652), .A2(n7166), .ZN(n8137) );
  NAND2_X1 U9474 ( .A1(n8652), .A2(n8655), .ZN(n8138) );
  NAND2_X1 U9475 ( .A1(n7169), .A2(n7167), .ZN(P3_U3487) );
  OR2_X1 U9476 ( .A1(n15159), .A2(n7168), .ZN(n7167) );
  AOI21_X1 U9477 ( .B1(n12501), .B2(n12504), .A(n15052), .ZN(n7172) );
  NAND4_X1 U9478 ( .A1(n8128), .A2(n8127), .A3(n8212), .A4(n7176), .ZN(n8367)
         );
  NAND3_X1 U9479 ( .A1(n8128), .A2(n8127), .A3(n8212), .ZN(n8353) );
  NAND2_X1 U9480 ( .A1(n7177), .A2(n7178), .ZN(n12094) );
  NAND2_X1 U9481 ( .A1(n12081), .A2(n7179), .ZN(n7177) );
  INV_X1 U9482 ( .A(n12084), .ZN(n7181) );
  NAND2_X1 U9483 ( .A1(n12177), .A2(n7192), .ZN(n7188) );
  NAND2_X1 U9484 ( .A1(n7212), .A2(n7215), .ZN(n12052) );
  NAND3_X1 U9485 ( .A1(n12045), .A2(n7213), .A3(n12044), .ZN(n7212) );
  NAND2_X1 U9486 ( .A1(n7216), .A2(n7219), .ZN(n12040) );
  NAND3_X1 U9487 ( .A1(n12032), .A2(n7217), .A3(n12031), .ZN(n7216) );
  NAND2_X1 U9488 ( .A1(n7224), .A2(n7222), .ZN(n12103) );
  NAND2_X1 U9489 ( .A1(n7230), .A2(n7228), .ZN(n12130) );
  NAND2_X1 U9490 ( .A1(n12125), .A2(n7231), .ZN(n7230) );
  NAND2_X1 U9491 ( .A1(n7233), .A2(n7236), .ZN(n12062) );
  NAND3_X1 U9492 ( .A1(n12057), .A2(n7234), .A3(n12056), .ZN(n7233) );
  NAND2_X1 U9493 ( .A1(n7238), .A2(n7241), .ZN(n12071) );
  NAND3_X1 U9494 ( .A1(n12067), .A2(n7239), .A3(n12066), .ZN(n7238) );
  NAND2_X1 U9495 ( .A1(n10582), .A2(n7243), .ZN(n10687) );
  XNOR2_X2 U9496 ( .A(n9705), .B(P1_IR_REG_19__SCAN_IN), .ZN(n14559) );
  NAND2_X1 U9497 ( .A1(n13947), .A2(n7246), .ZN(n7245) );
  NAND2_X1 U9498 ( .A1(n13947), .A2(n7258), .ZN(n7254) );
  AOI21_X1 U9499 ( .B1(n13947), .B2(n13946), .A(n6470), .ZN(n13932) );
  AOI21_X2 U9500 ( .B1(n7249), .B2(n7252), .A(n6428), .ZN(n7251) );
  NAND2_X1 U9501 ( .A1(n11100), .A2(n7260), .ZN(n14552) );
  XNOR2_X2 U9502 ( .A(n12011), .B(n7265), .ZN(n12186) );
  MUX2_X1 U9503 ( .A(n7266), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13732), .Z(
        P1_U3564) );
  MUX2_X1 U9504 ( .A(n7266), .B(n7265), .S(n12173), .Z(n12012) );
  NAND2_X1 U9505 ( .A1(n9677), .A2(n7267), .ZN(n14228) );
  NOR2_X2 U9506 ( .A1(n9472), .A2(n9471), .ZN(n7268) );
  NAND2_X1 U9507 ( .A1(n10190), .A2(n7269), .ZN(n7272) );
  NAND2_X1 U9508 ( .A1(n7276), .A2(n7275), .ZN(n7274) );
  NAND2_X1 U9509 ( .A1(n11340), .A2(n6534), .ZN(n7284) );
  NAND2_X1 U9510 ( .A1(n10570), .A2(n7287), .ZN(n7286) );
  OAI21_X1 U9511 ( .B1(n13070), .B2(n6461), .A(n7299), .ZN(n7296) );
  AND2_X2 U9512 ( .A1(n7298), .A2(n7297), .ZN(n9640) );
  NAND2_X1 U9513 ( .A1(n6513), .A2(n7306), .ZN(n13044) );
  OAI21_X1 U9514 ( .B1(n13092), .B2(n7310), .A(n7307), .ZN(n7312) );
  NAND2_X1 U9515 ( .A1(n13092), .A2(n13091), .ZN(n13090) );
  NAND2_X1 U9516 ( .A1(n13090), .A2(n7313), .ZN(n11956) );
  INV_X1 U9517 ( .A(n7312), .ZN(n13029) );
  INV_X2 U9518 ( .A(n13026), .ZN(n9588) );
  NAND2_X1 U9519 ( .A1(n7318), .A2(n7316), .ZN(n13290) );
  NOR2_X2 U9520 ( .A1(n13259), .A2(n7331), .ZN(n7330) );
  OAI21_X1 U9521 ( .B1(n11348), .B2(n7335), .A(n7334), .ZN(n11413) );
  NAND2_X1 U9522 ( .A1(n11348), .A2(n7334), .ZN(n7333) );
  NAND2_X1 U9523 ( .A1(n7743), .A2(n7532), .ZN(n7977) );
  INV_X1 U9524 ( .A(n7535), .ZN(n7340) );
  NAND2_X1 U9525 ( .A1(n7678), .A2(n7342), .ZN(n7341) );
  NAND2_X1 U9526 ( .A1(n7483), .A2(n7482), .ZN(n7801) );
  NAND2_X1 U9527 ( .A1(n7350), .A2(n7354), .ZN(n7491) );
  NAND2_X1 U9528 ( .A1(n7483), .A2(n7351), .ZN(n7350) );
  INV_X1 U9529 ( .A(n7361), .ZN(n13957) );
  OAI211_X1 U9530 ( .C1(n7911), .C2(n7366), .A(n7367), .B(n6435), .ZN(n11871)
         );
  NOR2_X1 U9531 ( .A1(n9780), .A2(n7384), .ZN(n7383) );
  INV_X1 U9532 ( .A(n7386), .ZN(n10775) );
  OAI211_X1 U9533 ( .C1(n13698), .C2(n7392), .A(n7389), .B(n7387), .ZN(n12242)
         );
  NAND2_X1 U9534 ( .A1(n13698), .A2(n7388), .ZN(n7387) );
  NAND2_X1 U9535 ( .A1(n13698), .A2(n13699), .ZN(n7394) );
  INV_X1 U9536 ( .A(n7406), .ZN(n11424) );
  NAND2_X1 U9537 ( .A1(n12249), .A2(n12248), .ZN(n12259) );
  NAND2_X1 U9538 ( .A1(n14096), .A2(n12073), .ZN(n11533) );
  NAND2_X2 U9539 ( .A1(n12163), .A2(n11972), .ZN(n12037) );
  OR2_X2 U9540 ( .A1(n12740), .A2(n8513), .ZN(n8515) );
  NAND2_X1 U9541 ( .A1(n12144), .A2(n12143), .ZN(n12145) );
  OAI21_X1 U9542 ( .B1(n8670), .B2(n8669), .A(n10109), .ZN(n9440) );
  AOI21_X1 U9543 ( .B1(n10109), .B2(n8660), .A(n8659), .ZN(n12966) );
  XNOR2_X1 U9544 ( .A(n8595), .B(n8594), .ZN(n8616) );
  XNOR2_X1 U9545 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8176) );
  NAND2_X1 U9546 ( .A1(n8016), .A2(n7416), .ZN(n8018) );
  NAND2_X1 U9547 ( .A1(n6515), .A2(n9218), .ZN(n9222) );
  XNOR2_X2 U9548 ( .A(n8177), .B(n8178), .ZN(n10311) );
  NAND2_X1 U9549 ( .A1(n8689), .A2(n8688), .ZN(n8696) );
  OAI21_X1 U9550 ( .B1(n10235), .B2(n9167), .A(n9158), .ZN(n9163) );
  OAI211_X1 U9551 ( .C1(n8240), .C2(SI_2_), .A(n8200), .B(n8199), .ZN(n15077)
         );
  CLKBUF_X1 U9552 ( .A(n8033), .Z(n9869) );
  NAND2_X1 U9553 ( .A1(n12974), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U9554 ( .A1(n9431), .A2(n9430), .ZN(n9432) );
  AOI21_X2 U9555 ( .B1(n9548), .B2(n9547), .A(n7409), .ZN(n11223) );
  AOI21_X1 U9556 ( .B1(n11956), .B2(n11955), .A(n13088), .ZN(n11962) );
  NAND2_X1 U9557 ( .A1(n9701), .A2(n9948), .ZN(n9946) );
  AND2_X1 U9558 ( .A1(n9546), .A2(n9545), .ZN(n7409) );
  OR2_X1 U9559 ( .A1(n9759), .A2(n9758), .ZN(n7410) );
  OR2_X1 U9560 ( .A1(n12250), .A2(n12743), .ZN(n7411) );
  AND2_X1 U9561 ( .A1(n7977), .A2(n7978), .ZN(n7412) );
  AND2_X2 U9562 ( .A1(n8924), .A2(n8923), .ZN(n14857) );
  INV_X1 U9563 ( .A(n13497), .ZN(n11336) );
  AND2_X1 U9564 ( .A1(n8924), .A2(n14834), .ZN(n14457) );
  INV_X1 U9565 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10744) );
  INV_X1 U9566 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8133) );
  AND2_X1 U9567 ( .A1(n7470), .A2(n7469), .ZN(n7413) );
  INV_X1 U9568 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U9569 ( .A1(n14562), .A2(n14561), .ZN(n14092) );
  INV_X1 U9570 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7546) );
  INV_X1 U9571 ( .A(n9416), .ZN(n8695) );
  AND2_X1 U9572 ( .A1(n7487), .A2(n7486), .ZN(n7415) );
  OR2_X1 U9573 ( .A1(n13505), .A2(n11607), .ZN(n7416) );
  INV_X1 U9574 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10424) );
  AND2_X1 U9575 ( .A1(n9259), .A2(n9256), .ZN(n7417) );
  INV_X1 U9576 ( .A(n13199), .ZN(n8925) );
  XOR2_X1 U9577 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n7418) );
  AND2_X1 U9578 ( .A1(n12004), .A2(n12003), .ZN(n7419) );
  OR2_X1 U9579 ( .A1(n9222), .A2(n9221), .ZN(n7420) );
  INV_X1 U9580 ( .A(n9728), .ZN(n11746) );
  INV_X1 U9581 ( .A(n15159), .ZN(n9457) );
  INV_X2 U9582 ( .A(n15142), .ZN(n15143) );
  INV_X1 U9583 ( .A(n11506), .ZN(n8625) );
  INV_X1 U9584 ( .A(n12757), .ZN(n8635) );
  AND2_X1 U9585 ( .A1(n12258), .A2(n12257), .ZN(n7421) );
  AOI21_X1 U9586 ( .B1(n10243), .B2(n9153), .A(n9500), .ZN(n9154) );
  NAND2_X1 U9587 ( .A1(n9160), .A2(n9159), .ZN(n9162) );
  NAND2_X1 U9588 ( .A1(n12010), .A2(n12009), .ZN(n12014) );
  NAND2_X1 U9589 ( .A1(n9192), .A2(n9191), .ZN(n9198) );
  OAI21_X1 U9590 ( .B1(n10831), .B2(n9177), .A(n9210), .ZN(n9211) );
  OAI21_X1 U9591 ( .B1(n10912), .B2(n9369), .A(n9223), .ZN(n9224) );
  AOI21_X1 U9592 ( .B1(n13246), .B2(n9369), .A(n9324), .ZN(n9327) );
  OR2_X1 U9593 ( .A1(n11966), .A2(n12226), .ZN(n11968) );
  AOI21_X1 U9594 ( .B1(n9388), .B2(n9369), .A(n9362), .ZN(n9381) );
  INV_X1 U9595 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7533) );
  INV_X1 U9596 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9482) );
  INV_X1 U9597 ( .A(n12782), .ZN(n8474) );
  AND2_X1 U9598 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n7550) );
  INV_X1 U9599 ( .A(n10263), .ZN(n9393) );
  INV_X1 U9600 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9479) );
  AND2_X1 U9601 ( .A1(n8575), .A2(n8143), .ZN(n8164) );
  NOR2_X1 U9602 ( .A1(n8544), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8562) );
  INV_X1 U9603 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8419) );
  NOR2_X1 U9604 ( .A1(n9381), .A2(n9382), .ZN(n9383) );
  INV_X1 U9605 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7807) );
  AND2_X1 U9606 ( .A1(n7947), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7963) );
  INV_X1 U9607 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7859) );
  INV_X1 U9608 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7715) );
  INV_X1 U9609 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7650) );
  INV_X1 U9610 ( .A(n11818), .ZN(n11816) );
  OR2_X1 U9611 ( .A1(n14304), .A2(n11661), .ZN(n11299) );
  INV_X1 U9612 ( .A(P1_B_REG_SCAN_IN), .ZN(n9761) );
  NAND2_X1 U9613 ( .A1(n9491), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9481) );
  INV_X1 U9614 ( .A(SI_16_), .ZN(n8423) );
  INV_X1 U9615 ( .A(SI_11_), .ZN(n8345) );
  INV_X1 U9616 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U9617 ( .A1(n8164), .A2(n8144), .ZN(n8166) );
  AND2_X1 U9618 ( .A1(n8562), .A2(n8561), .ZN(n8575) );
  NAND2_X1 U9619 ( .A1(n8454), .A2(n8453), .ZN(n8468) );
  INV_X1 U9620 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8231) );
  NOR2_X1 U9621 ( .A1(n12265), .A2(n15044), .ZN(n8614) );
  AND2_X1 U9622 ( .A1(n8675), .A2(n9078), .ZN(n10426) );
  INV_X1 U9623 ( .A(n9610), .ZN(n9608) );
  AND2_X1 U9624 ( .A1(n7858), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7885) );
  INV_X1 U9625 ( .A(n12247), .ZN(n7548) );
  INV_X1 U9626 ( .A(n7930), .ZN(n7551) );
  INV_X1 U9627 ( .A(n13110), .ZN(n7922) );
  OR2_X1 U9628 ( .A1(n7701), .A2(n7700), .ZN(n7716) );
  INV_X1 U9629 ( .A(n9406), .ZN(n7799) );
  INV_X1 U9630 ( .A(n10266), .ZN(n7605) );
  XNOR2_X1 U9631 ( .A(n13129), .B(n10554), .ZN(n7986) );
  AND2_X1 U9632 ( .A1(n14461), .A2(n14458), .ZN(n11728) );
  INV_X1 U9633 ( .A(n13612), .ZN(n11827) );
  OR2_X1 U9634 ( .A1(n11919), .A2(n11940), .ZN(n13909) );
  OR2_X1 U9635 ( .A1(n11887), .A2(n11886), .ZN(n11905) );
  NAND2_X1 U9636 ( .A1(n11816), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11836) );
  OR2_X1 U9637 ( .A1(n11016), .A2(n11015), .ZN(n11447) );
  INV_X1 U9638 ( .A(n11835), .ZN(n11773) );
  INV_X1 U9639 ( .A(n14481), .ZN(n11542) );
  INV_X1 U9640 ( .A(n13903), .ZN(n14100) );
  INV_X1 U9641 ( .A(n9354), .ZN(n9346) );
  INV_X1 U9642 ( .A(n10582), .ZN(n10583) );
  NAND2_X1 U9643 ( .A1(n8892), .A2(n14768), .ZN(n8893) );
  NOR2_X1 U9644 ( .A1(n8482), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8495) );
  OR2_X1 U9645 ( .A1(n8249), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8265) );
  INV_X1 U9646 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n14891) );
  INV_X1 U9647 ( .A(n14865), .ZN(n14987) );
  INV_X1 U9648 ( .A(n12766), .ZN(n12792) );
  OR2_X1 U9649 ( .A1(n8332), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U9650 ( .A1(n15070), .A2(n14410), .ZN(n12826) );
  AND2_X1 U9651 ( .A1(n12968), .A2(n12966), .ZN(n9443) );
  OR2_X1 U9652 ( .A1(n8808), .A2(n9450), .ZN(n15044) );
  AND2_X1 U9653 ( .A1(n9451), .A2(n8645), .ZN(n15094) );
  INV_X1 U9654 ( .A(n15081), .ZN(n15046) );
  INV_X1 U9655 ( .A(SI_24_), .ZN(n12683) );
  INV_X1 U9656 ( .A(SI_12_), .ZN(n14271) );
  NAND2_X1 U9657 ( .A1(n7912), .A2(n6390), .ZN(n7914) );
  NOR2_X1 U9658 ( .A1(n7916), .A2(n9643), .ZN(n7931) );
  AND2_X1 U9659 ( .A1(n7885), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7898) );
  OR2_X1 U9660 ( .A1(n10088), .A2(n10087), .ZN(n14739) );
  AND2_X1 U9661 ( .A1(n9887), .A2(n9870), .ZN(n9900) );
  XNOR2_X1 U9662 ( .A(n13444), .B(n13106), .ZN(n13206) );
  INV_X1 U9663 ( .A(n9413), .ZN(n13239) );
  INV_X1 U9664 ( .A(n13117), .ZN(n11605) );
  OR2_X1 U9665 ( .A1(n8698), .A2(n8697), .ZN(n9631) );
  INV_X1 U9666 ( .A(n13121), .ZN(n10912) );
  INV_X1 U9667 ( .A(n9408), .ZN(n13389) );
  INV_X1 U9668 ( .A(n9498), .ZN(n13420) );
  INV_X1 U9669 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11302) );
  OR2_X1 U9670 ( .A1(n11778), .A2(n11777), .ZN(n11798) );
  NAND2_X1 U9671 ( .A1(n11252), .A2(n11254), .ZN(n11255) );
  OR2_X1 U9672 ( .A1(n11836), .A2(n13675), .ZN(n11856) );
  INV_X1 U9673 ( .A(n6415), .ZN(n9792) );
  AND2_X1 U9674 ( .A1(n13909), .A2(n11920), .ZN(n13937) );
  INV_X1 U9675 ( .A(n9744), .ZN(n11933) );
  INV_X1 U9676 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10980) );
  NAND2_X1 U9677 ( .A1(n14250), .A2(n10409), .ZN(n11979) );
  INV_X1 U9678 ( .A(n12200), .ZN(n13882) );
  NAND2_X1 U9679 ( .A1(n14591), .A2(n14559), .ZN(n10399) );
  INV_X2 U9680 ( .A(n11721), .ZN(n12232) );
  INV_X1 U9681 ( .A(n13885), .ZN(n14075) );
  OAI21_X1 U9682 ( .B1(n10405), .B2(P1_D_REG_1__SCAN_IN), .A(n10082), .ZN(
        n10858) );
  INV_X1 U9683 ( .A(n7480), .ZN(n7783) );
  INV_X1 U9684 ( .A(n12564), .ZN(n12731) );
  AND2_X1 U9685 ( .A1(n8553), .A2(n8552), .ZN(n9084) );
  INV_X1 U9686 ( .A(n15052), .ZN(n15089) );
  NOR2_X1 U9687 ( .A1(n8358), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8375) );
  INV_X1 U9688 ( .A(n11026), .ZN(n11023) );
  INV_X1 U9689 ( .A(n11047), .ZN(n15070) );
  NOR2_X1 U9690 ( .A1(n15159), .A2(n9459), .ZN(n9460) );
  NOR2_X1 U9691 ( .A1(n9444), .A2(n9443), .ZN(n10630) );
  NAND2_X1 U9692 ( .A1(n15094), .A2(n12839), .ZN(n15136) );
  INV_X1 U9693 ( .A(n12839), .ZN(n15140) );
  INV_X1 U9694 ( .A(n15076), .ZN(n14410) );
  NOR2_X1 U9695 ( .A1(n10109), .A2(n10108), .ZN(n10111) );
  INV_X1 U9696 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12969) );
  INV_X1 U9697 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8290) );
  INV_X1 U9698 ( .A(n13088), .ZN(n13093) );
  INV_X1 U9699 ( .A(n11585), .ZN(n9434) );
  AND2_X1 U9700 ( .A1(n14741), .A2(n11372), .ZN(n14756) );
  OR2_X1 U9701 ( .A1(n9867), .A2(n9866), .ZN(n9887) );
  AOI21_X1 U9702 ( .B1(n13436), .B2(n13422), .A(n8721), .ZN(n8722) );
  INV_X1 U9703 ( .A(n14428), .ZN(n14440) );
  NAND2_X1 U9704 ( .A1(n9798), .A2(n10859), .ZN(n13712) );
  INV_X1 U9705 ( .A(n13712), .ZN(n14472) );
  INV_X1 U9706 ( .A(n13705), .ZN(n14470) );
  OR2_X1 U9707 ( .A1(n13992), .A2(n9744), .ZN(n11862) );
  INV_X1 U9708 ( .A(n14533), .ZN(n13841) );
  AND2_X1 U9709 ( .A1(n10042), .A2(n10041), .ZN(n13846) );
  INV_X1 U9710 ( .A(n13890), .ZN(n14010) );
  INV_X1 U9711 ( .A(n12199), .ZN(n11541) );
  INV_X1 U9712 ( .A(n14652), .ZN(n14686) );
  INV_X1 U9713 ( .A(n14644), .ZN(n14683) );
  AND2_X1 U9714 ( .A1(n10407), .A2(n10406), .ZN(n10860) );
  OR2_X1 U9715 ( .A1(n9760), .A2(n9775), .ZN(n10404) );
  AND2_X1 U9716 ( .A1(n10299), .A2(n10298), .ZN(n14984) );
  NOR2_X1 U9717 ( .A1(n8816), .A2(n8815), .ZN(n8817) );
  INV_X1 U9718 ( .A(n12392), .ZN(n11503) );
  AND2_X1 U9719 ( .A1(n8949), .A2(n8611), .ZN(n10746) );
  NAND2_X1 U9720 ( .A1(n8541), .A2(n8540), .ZN(n12564) );
  INV_X1 U9721 ( .A(n14385), .ZN(n14997) );
  NAND2_X1 U9722 ( .A1(n10631), .A2(n15079), .ZN(n15078) );
  NAND2_X1 U9723 ( .A1(n10632), .A2(n15078), .ZN(n15109) );
  AND2_X2 U9724 ( .A1(n10630), .A2(n9456), .ZN(n15159) );
  INV_X1 U9725 ( .A(n12338), .ZN(n12936) );
  AND2_X1 U9726 ( .A1(n8683), .A2(n8682), .ZN(n15142) );
  NAND2_X1 U9727 ( .A1(n15143), .A2(n14410), .ZN(n12965) );
  INV_X1 U9728 ( .A(n9144), .ZN(n11248) );
  INV_X1 U9729 ( .A(SI_18_), .ZN(n10637) );
  INV_X1 U9730 ( .A(n12455), .ZN(n14931) );
  INV_X1 U9731 ( .A(n14287), .ZN(n14275) );
  INV_X1 U9732 ( .A(n11360), .ZN(n14444) );
  INV_X1 U9733 ( .A(n11337), .ZN(n11333) );
  INV_X1 U9734 ( .A(n13086), .ZN(n13102) );
  OR2_X1 U9735 ( .A1(n7849), .A2(n7848), .ZN(n13113) );
  INV_X1 U9736 ( .A(n14776), .ZN(n14816) );
  NAND2_X1 U9737 ( .A1(n9887), .A2(n9868), .ZN(n14807) );
  INV_X1 U9738 ( .A(n14773), .ZN(n14827) );
  AND2_X1 U9739 ( .A1(n8701), .A2(n13412), .ZN(n13384) );
  NAND2_X1 U9740 ( .A1(n13427), .A2(n8703), .ZN(n13425) );
  NAND2_X1 U9741 ( .A1(n14857), .A2(n13506), .ZN(n13497) );
  INV_X1 U9742 ( .A(n13299), .ZN(n13532) );
  INV_X1 U9743 ( .A(n14457), .ZN(n14450) );
  INV_X1 U9744 ( .A(n14450), .ZN(n14854) );
  INV_X1 U9745 ( .A(n14831), .ZN(n14832) );
  AND2_X1 U9746 ( .A1(n9633), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14835) );
  INV_X1 U9747 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13574) );
  INV_X1 U9748 ( .A(n14135), .ZN(n13939) );
  NAND2_X1 U9749 ( .A1(n9784), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14479) );
  INV_X1 U9750 ( .A(n14475), .ZN(n13718) );
  INV_X1 U9751 ( .A(n13682), .ZN(n13887) );
  OR2_X1 U9752 ( .A1(n10037), .A2(n13745), .ZN(n14533) );
  INV_X1 U9753 ( .A(n14595), .ZN(n14109) );
  INV_X1 U9754 ( .A(n14063), .ZN(n13930) );
  INV_X1 U9755 ( .A(n14709), .ZN(n14706) );
  AND4_X1 U9756 ( .A1(n14487), .A2(n14486), .A3(n14485), .A4(n14484), .ZN(
        n14505) );
  INV_X1 U9757 ( .A(n14693), .ZN(n14691) );
  INV_X1 U9758 ( .A(n10081), .ZN(n9948) );
  NAND2_X1 U9759 ( .A1(n10405), .A2(n9947), .ZN(n14603) );
  INV_X1 U9760 ( .A(n11976), .ZN(n14250) );
  INV_X1 U9761 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n12704) );
  XNOR2_X1 U9762 ( .A(n8867), .B(n8866), .ZN(n14282) );
  INV_X2 U9763 ( .A(n12399), .ZN(P3_U3897) );
  OAI21_X1 U9764 ( .B1(n9458), .B2(n15142), .A(n8687), .ZN(P3_U3456) );
  AND2_X1 U9765 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9866), .ZN(P2_U3947) );
  OAI21_X1 U9766 ( .B1(n8930), .B2(n14450), .A(n8084), .ZN(P2_U3495) );
  INV_X1 U9767 ( .A(n13732), .ZN(P1_U4016) );
  INV_X1 U9768 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9846) );
  AND2_X1 U9769 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U9770 ( .A1(n7432), .A2(n7425), .ZN(n7574) );
  AND2_X1 U9771 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7426) );
  NAND2_X1 U9772 ( .A1(n7431), .A2(n7426), .ZN(n9731) );
  NAND2_X1 U9773 ( .A1(n7574), .A2(n9731), .ZN(n7585) );
  NAND2_X1 U9774 ( .A1(n7586), .A2(n7585), .ZN(n7430) );
  INV_X1 U9775 ( .A(n7427), .ZN(n7428) );
  NAND2_X1 U9776 ( .A1(n7428), .A2(SI_1_), .ZN(n7429) );
  NAND2_X1 U9777 ( .A1(n7430), .A2(n7429), .ZN(n7594) );
  INV_X1 U9778 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9825) );
  INV_X1 U9779 ( .A(n7433), .ZN(n7434) );
  NAND2_X1 U9780 ( .A1(n7434), .A2(SI_2_), .ZN(n7435) );
  INV_X1 U9781 ( .A(n7614), .ZN(n7438) );
  NAND2_X1 U9782 ( .A1(n7615), .A2(n7438), .ZN(n7441) );
  NAND2_X1 U9783 ( .A1(n7439), .A2(SI_3_), .ZN(n7440) );
  MUX2_X1 U9784 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7476), .Z(n7443) );
  XNOR2_X1 U9785 ( .A(n7443), .B(SI_4_), .ZN(n7624) );
  INV_X1 U9786 ( .A(n7624), .ZN(n7442) );
  NAND2_X1 U9787 ( .A1(n7443), .A2(SI_4_), .ZN(n7444) );
  MUX2_X1 U9788 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7476), .Z(n7446) );
  XNOR2_X1 U9789 ( .A(n7446), .B(SI_5_), .ZN(n7632) );
  INV_X1 U9790 ( .A(n7632), .ZN(n7445) );
  NAND2_X1 U9791 ( .A1(n7446), .A2(SI_5_), .ZN(n7447) );
  MUX2_X1 U9792 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7476), .Z(n7449) );
  XNOR2_X1 U9793 ( .A(n7449), .B(SI_6_), .ZN(n7647) );
  INV_X1 U9794 ( .A(n7647), .ZN(n7448) );
  XNOR2_X1 U9795 ( .A(n7451), .B(SI_7_), .ZN(n7659) );
  INV_X1 U9796 ( .A(n7659), .ZN(n7450) );
  NAND2_X1 U9797 ( .A1(n7451), .A2(SI_7_), .ZN(n7452) );
  MUX2_X1 U9798 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n9828), .Z(n7455) );
  NAND2_X1 U9799 ( .A1(n7455), .A2(SI_8_), .ZN(n7456) );
  MUX2_X1 U9800 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n9828), .Z(n7458) );
  INV_X1 U9801 ( .A(n7690), .ZN(n7457) );
  MUX2_X1 U9802 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n9828), .Z(n7460) );
  XNOR2_X1 U9803 ( .A(n7460), .B(SI_10_), .ZN(n7709) );
  INV_X1 U9804 ( .A(n7709), .ZN(n7459) );
  NAND2_X1 U9805 ( .A1(n7710), .A2(n7459), .ZN(n7462) );
  NAND2_X1 U9806 ( .A1(n7460), .A2(SI_10_), .ZN(n7461) );
  MUX2_X1 U9807 ( .A(n10102), .B(n10107), .S(n9812), .Z(n7463) );
  NAND2_X1 U9808 ( .A1(n7463), .A2(n8345), .ZN(n7466) );
  INV_X1 U9809 ( .A(n7463), .ZN(n7464) );
  NAND2_X1 U9810 ( .A1(n7464), .A2(SI_11_), .ZN(n7465) );
  NAND2_X1 U9811 ( .A1(n7466), .A2(n7465), .ZN(n7727) );
  MUX2_X1 U9812 ( .A(n10189), .B(n6711), .S(n9828), .Z(n7467) );
  NAND2_X1 U9813 ( .A1(n7467), .A2(n14271), .ZN(n7470) );
  INV_X1 U9814 ( .A(n7467), .ZN(n7468) );
  NAND2_X1 U9815 ( .A1(n7468), .A2(SI_12_), .ZN(n7469) );
  MUX2_X1 U9816 ( .A(n10251), .B(n11285), .S(n9812), .Z(n7472) );
  INV_X1 U9817 ( .A(n7472), .ZN(n7473) );
  NAND2_X1 U9818 ( .A1(n7473), .A2(SI_13_), .ZN(n7474) );
  MUX2_X1 U9819 ( .A(n10443), .B(n6630), .S(n9812), .Z(n7480) );
  MUX2_X1 U9820 ( .A(n12681), .B(n6650), .S(n9812), .Z(n7477) );
  NAND2_X1 U9821 ( .A1(n7477), .A2(n8403), .ZN(n7482) );
  INV_X1 U9822 ( .A(n7477), .ZN(n7478) );
  NAND2_X1 U9823 ( .A1(n7478), .A2(SI_15_), .ZN(n7479) );
  NAND2_X1 U9824 ( .A1(n7482), .A2(n7479), .ZN(n7785) );
  NOR2_X1 U9825 ( .A1(n7480), .A2(n8386), .ZN(n7481) );
  MUX2_X1 U9826 ( .A(n10424), .B(n12704), .S(n9828), .Z(n7484) );
  INV_X1 U9827 ( .A(n7484), .ZN(n7485) );
  NAND2_X1 U9828 ( .A1(n7485), .A2(SI_16_), .ZN(n7486) );
  MUX2_X1 U9829 ( .A(n10589), .B(n6632), .S(n9812), .Z(n7814) );
  INV_X1 U9830 ( .A(n7814), .ZN(n7488) );
  NAND2_X1 U9831 ( .A1(n7488), .A2(SI_17_), .ZN(n7489) );
  NAND2_X1 U9832 ( .A1(n7814), .A2(n8449), .ZN(n7490) );
  MUX2_X1 U9833 ( .A(n10701), .B(n6707), .S(n9828), .Z(n7836) );
  MUX2_X1 U9834 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n9812), .Z(n7494) );
  XNOR2_X1 U9835 ( .A(n7494), .B(SI_19_), .ZN(n7851) );
  INV_X1 U9836 ( .A(n7494), .ZN(n7495) );
  INV_X1 U9837 ( .A(SI_19_), .ZN(n10690) );
  NAND2_X1 U9838 ( .A1(n7495), .A2(n10690), .ZN(n7496) );
  MUX2_X1 U9839 ( .A(n12660), .B(n7077), .S(n9812), .Z(n7865) );
  MUX2_X1 U9840 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n9812), .Z(n7500) );
  INV_X1 U9841 ( .A(n7500), .ZN(n7501) );
  INV_X1 U9842 ( .A(SI_21_), .ZN(n12626) );
  NAND2_X1 U9843 ( .A1(n7501), .A2(n12626), .ZN(n7502) );
  INV_X1 U9844 ( .A(n7504), .ZN(n7506) );
  INV_X1 U9845 ( .A(SI_22_), .ZN(n7505) );
  INV_X1 U9846 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8085) );
  MUX2_X1 U9847 ( .A(n11470), .B(n8085), .S(n9828), .Z(n7893) );
  INV_X1 U9848 ( .A(n7893), .ZN(n7508) );
  INV_X1 U9849 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11851) );
  MUX2_X1 U9850 ( .A(n13574), .B(n14246), .S(n9812), .Z(n7513) );
  NAND2_X1 U9851 ( .A1(n7513), .A2(n12683), .ZN(n7564) );
  INV_X1 U9852 ( .A(n7564), .ZN(n7519) );
  INV_X1 U9853 ( .A(n7510), .ZN(n7511) );
  MUX2_X1 U9854 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n9812), .Z(n7520) );
  XNOR2_X1 U9855 ( .A(n7520), .B(SI_25_), .ZN(n7926) );
  INV_X1 U9856 ( .A(n7926), .ZN(n7515) );
  INV_X1 U9857 ( .A(n7513), .ZN(n7514) );
  NAND2_X1 U9858 ( .A1(n7514), .A2(SI_24_), .ZN(n7924) );
  NAND2_X1 U9859 ( .A1(n7515), .A2(n7924), .ZN(n7516) );
  INV_X1 U9860 ( .A(n7520), .ZN(n7521) );
  INV_X1 U9861 ( .A(SI_25_), .ZN(n12993) );
  NAND2_X1 U9862 ( .A1(n7521), .A2(n12993), .ZN(n7522) );
  MUX2_X1 U9863 ( .A(n13566), .B(n6709), .S(n9812), .Z(n7937) );
  XNOR2_X1 U9864 ( .A(n7937), .B(SI_26_), .ZN(n7523) );
  AND2_X2 U9865 ( .A1(n7590), .A2(n7591), .ZN(n7612) );
  NOR2_X1 U9866 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7527) );
  NOR2_X1 U9867 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7526) );
  AND2_X1 U9868 ( .A1(n7527), .A2(n7526), .ZN(n7528) );
  NOR2_X1 U9869 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7530) );
  NOR2_X1 U9870 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7529) );
  NAND3_X1 U9871 ( .A1(n7819), .A2(n7530), .A3(n7529), .ZN(n7974) );
  NAND2_X1 U9872 ( .A1(n7818), .A2(n12614), .ZN(n7531) );
  NOR2_X2 U9873 ( .A1(n7974), .A2(n7531), .ZN(n7532) );
  NAND4_X1 U9874 ( .A1(n8063), .A2(n7981), .A3(n7534), .A4(n7533), .ZN(n7535)
         );
  NAND2_X1 U9875 ( .A1(n13565), .A2(n7626), .ZN(n7543) );
  OR2_X1 U9876 ( .A1(n6410), .A2(n13566), .ZN(n7542) );
  NAND2_X1 U9877 ( .A1(n7545), .A2(n7546), .ZN(n13551) );
  NAND2_X1 U9878 ( .A1(n9351), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7556) );
  INV_X1 U9879 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n13451) );
  OR2_X1 U9880 ( .A1(n7577), .A2(n13451), .ZN(n7555) );
  NAND2_X1 U9881 ( .A1(n7619), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U9882 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n7549) );
  NOR2_X1 U9883 ( .A1(n7669), .A2(n7549), .ZN(n7670) );
  NAND2_X1 U9884 ( .A1(n7670), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7701) );
  INV_X1 U9885 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U9886 ( .A1(n7736), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7775) );
  INV_X1 U9887 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7774) );
  INV_X1 U9888 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U9889 ( .A1(n7806), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7845) );
  INV_X1 U9890 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U9891 ( .A1(n7898), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n7899) );
  INV_X1 U9892 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9643) );
  NAND2_X1 U9893 ( .A1(n7931), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U9894 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n7551), .ZN(n7949) );
  OAI21_X1 U9895 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n7551), .A(n7949), .ZN(
        n13224) );
  OR2_X1 U9896 ( .A1(n8036), .A2(n13224), .ZN(n7554) );
  INV_X1 U9897 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13225) );
  OR2_X1 U9898 ( .A1(n8038), .A2(n13225), .ZN(n7553) );
  NAND4_X1 U9899 ( .A1(n7556), .A2(n7555), .A3(n7554), .A4(n7553), .ZN(n13107)
         );
  NAND2_X1 U9900 ( .A1(n9351), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7563) );
  INV_X1 U9901 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n7557) );
  OR2_X1 U9902 ( .A1(n7577), .A2(n7557), .ZN(n7562) );
  INV_X1 U9903 ( .A(n7916), .ZN(n7559) );
  INV_X1 U9904 ( .A(n7931), .ZN(n7558) );
  OAI21_X1 U9905 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n7559), .A(n7558), .ZN(
        n13264) );
  OR2_X1 U9906 ( .A1(n8036), .A2(n13264), .ZN(n7561) );
  INV_X1 U9907 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13265) );
  OR2_X1 U9908 ( .A1(n8038), .A2(n13265), .ZN(n7560) );
  NAND4_X1 U9909 ( .A1(n7563), .A2(n7562), .A3(n7561), .A4(n7560), .ZN(n13109)
         );
  AND2_X1 U9910 ( .A1(n7564), .A2(n7924), .ZN(n7565) );
  OR2_X1 U9911 ( .A1(n6410), .A2(n13574), .ZN(n7566) );
  NAND2_X1 U9912 ( .A1(n7862), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7572) );
  INV_X1 U9913 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10246) );
  INV_X1 U9914 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U9915 ( .A1(n7638), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7569) );
  NAND4_X1 U9916 ( .A1(n7572), .A2(n7571), .A3(n7570), .A4(n7569), .ZN(n9157)
         );
  INV_X1 U9917 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9931) );
  INV_X1 U9918 ( .A(SI_0_), .ZN(n8189) );
  INV_X1 U9919 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8086) );
  OAI21_X1 U9920 ( .B1(n9812), .B2(n8189), .A(n8086), .ZN(n7573) );
  NAND2_X1 U9921 ( .A1(n7574), .A2(n7573), .ZN(n13577) );
  INV_X1 U9922 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7575) );
  OR2_X1 U9923 ( .A1(n7576), .A2(n7575), .ZN(n7582) );
  INV_X1 U9924 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9871) );
  INV_X1 U9925 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10536) );
  OR2_X1 U9926 ( .A1(n7599), .A2(n10536), .ZN(n7580) );
  INV_X1 U9927 ( .A(n7578), .ZN(n7875) );
  NAND4_X2 U9928 ( .A1(n7582), .A2(n7581), .A3(n7580), .A4(n7579), .ZN(n13129)
         );
  INV_X1 U9929 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U9930 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7583) );
  XNOR2_X1 U9931 ( .A(n7584), .B(n7583), .ZN(n9929) );
  XNOR2_X1 U9932 ( .A(n7586), .B(n7585), .ZN(n9845) );
  NAND2_X1 U9933 ( .A1(n10231), .A2(n7986), .ZN(n10230) );
  OR2_X1 U9934 ( .A1(n13129), .A2(n10238), .ZN(n7588) );
  NAND2_X1 U9935 ( .A1(n10230), .A2(n7588), .ZN(n10259) );
  OR2_X1 U9936 ( .A1(n7590), .A2(n7980), .ZN(n7592) );
  XNOR2_X1 U9937 ( .A(n7592), .B(n7591), .ZN(n13136) );
  XNOR2_X1 U9938 ( .A(n7593), .B(n7594), .ZN(n9829) );
  OR2_X1 U9939 ( .A1(n9829), .A2(n7595), .ZN(n7598) );
  OR2_X1 U9940 ( .A1(n7596), .A2(n9825), .ZN(n7597) );
  NAND2_X1 U9941 ( .A1(n7862), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7604) );
  INV_X1 U9942 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10545) );
  OR2_X1 U9943 ( .A1(n7599), .A2(n10545), .ZN(n7603) );
  INV_X1 U9944 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9888) );
  OR2_X1 U9945 ( .A1(n7578), .A2(n9888), .ZN(n7602) );
  INV_X1 U9946 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7600) );
  OR2_X1 U9947 ( .A1(n7576), .A2(n7600), .ZN(n7601) );
  NAND2_X1 U9948 ( .A1(n10259), .A2(n10263), .ZN(n10258) );
  OR2_X1 U9949 ( .A1(n9166), .A2(n10266), .ZN(n7606) );
  NAND2_X1 U9950 ( .A1(n10258), .A2(n7606), .ZN(n10364) );
  NAND2_X1 U9951 ( .A1(n7862), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7611) );
  OR2_X1 U9952 ( .A1(n7599), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7610) );
  INV_X1 U9953 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10462) );
  OR2_X1 U9954 ( .A1(n7578), .A2(n10462), .ZN(n7609) );
  INV_X1 U9955 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7607) );
  OR2_X1 U9956 ( .A1(n7576), .A2(n7607), .ZN(n7608) );
  OR2_X1 U9957 ( .A1(n7612), .A2(n7980), .ZN(n7613) );
  XNOR2_X1 U9958 ( .A(n7613), .B(n7627), .ZN(n13154) );
  XNOR2_X1 U9959 ( .A(n7615), .B(n7614), .ZN(n9826) );
  NAND2_X1 U9960 ( .A1(n7626), .A2(n9826), .ZN(n7617) );
  OR2_X1 U9961 ( .A1(n6410), .A2(n9827), .ZN(n7616) );
  INV_X1 U9962 ( .A(n6398), .ZN(n10563) );
  NAND2_X1 U9963 ( .A1(n10364), .A2(n10366), .ZN(n10363) );
  OR2_X1 U9964 ( .A1(n13128), .A2(n6399), .ZN(n7618) );
  NAND2_X1 U9965 ( .A1(n10363), .A2(n7618), .ZN(n10445) );
  INV_X1 U9966 ( .A(n7576), .ZN(n7638) );
  NAND2_X1 U9967 ( .A1(n7638), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7623) );
  INV_X1 U9968 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9880) );
  OR2_X1 U9969 ( .A1(n7577), .A2(n9880), .ZN(n7622) );
  INV_X1 U9970 ( .A(n7619), .ZN(n7640) );
  OAI21_X1 U9971 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7640), .ZN(n10454) );
  OR2_X1 U9972 ( .A1(n7599), .A2(n10454), .ZN(n7621) );
  INV_X1 U9973 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10451) );
  OR2_X1 U9974 ( .A1(n7578), .A2(n10451), .ZN(n7620) );
  NAND4_X1 U9975 ( .A1(n7623), .A2(n7622), .A3(n7621), .A4(n7620), .ZN(n13127)
         );
  XNOR2_X1 U9976 ( .A(n7625), .B(n7624), .ZN(n10776) );
  NAND2_X1 U9977 ( .A1(n10776), .A2(n6389), .ZN(n7630) );
  NAND2_X1 U9978 ( .A1(n7612), .A2(n7627), .ZN(n7634) );
  NAND2_X1 U9979 ( .A1(n7634), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7628) );
  XNOR2_X1 U9980 ( .A(n7628), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9897) );
  AOI22_X1 U9981 ( .A1(n7855), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7854), .B2(
        n9897), .ZN(n7629) );
  NAND2_X1 U9982 ( .A1(n7630), .A2(n7629), .ZN(n10471) );
  NAND2_X1 U9983 ( .A1(n10445), .A2(n10446), .ZN(n10444) );
  OR2_X1 U9984 ( .A1(n13127), .A2(n10471), .ZN(n7631) );
  NAND2_X1 U9985 ( .A1(n10444), .A2(n7631), .ZN(n10593) );
  XNOR2_X1 U9986 ( .A(n7633), .B(n7632), .ZN(n10803) );
  NAND2_X1 U9987 ( .A1(n10803), .A2(n6390), .ZN(n7637) );
  NAND2_X1 U9988 ( .A1(n7649), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7635) );
  XNOR2_X1 U9989 ( .A(n7635), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U9990 ( .A1(n7855), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7854), .B2(
        n9915), .ZN(n7636) );
  NAND2_X1 U9991 ( .A1(n7638), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7645) );
  INV_X1 U9992 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9881) );
  OR2_X1 U9993 ( .A1(n7577), .A2(n9881), .ZN(n7644) );
  INV_X1 U9994 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7639) );
  NAND2_X1 U9995 ( .A1(n7640), .A2(n7639), .ZN(n7641) );
  NAND2_X1 U9996 ( .A1(n7669), .A2(n7641), .ZN(n10602) );
  OR2_X1 U9997 ( .A1(n8036), .A2(n10602), .ZN(n7643) );
  INV_X1 U9998 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10599) );
  OR2_X1 U9999 ( .A1(n8038), .A2(n10599), .ZN(n7642) );
  NAND4_X1 U10000 ( .A1(n7645), .A2(n7644), .A3(n7643), .A4(n7642), .ZN(n13126) );
  OR2_X1 U10001 ( .A1(n10623), .A2(n13126), .ZN(n7646) );
  XNOR2_X1 U10002 ( .A(n7648), .B(n7647), .ZN(n10951) );
  NAND2_X1 U10003 ( .A1(n10951), .A2(n6390), .ZN(n7654) );
  INV_X1 U10004 ( .A(n7649), .ZN(n7651) );
  NAND2_X1 U10005 ( .A1(n7651), .A2(n7650), .ZN(n7661) );
  NAND2_X1 U10006 ( .A1(n7661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7652) );
  XNOR2_X1 U10007 ( .A(n7652), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U10008 ( .A1(n7855), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7854), .B2(
        n9960), .ZN(n7653) );
  NAND2_X1 U10009 ( .A1(n9351), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7658) );
  INV_X1 U10010 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9908) );
  OR2_X1 U10011 ( .A1(n7577), .A2(n9908), .ZN(n7657) );
  INV_X1 U10012 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7668) );
  XNOR2_X1 U10013 ( .A(n7669), .B(n7668), .ZN(n10672) );
  OR2_X1 U10014 ( .A1(n8036), .A2(n10672), .ZN(n7656) );
  INV_X1 U10015 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10670) );
  OR2_X1 U10016 ( .A1(n7578), .A2(n10670), .ZN(n7655) );
  NAND4_X1 U10017 ( .A1(n7658), .A2(n7657), .A3(n7656), .A4(n7655), .ZN(n13125) );
  XNOR2_X1 U10018 ( .A(n10698), .B(n13125), .ZN(n9396) );
  XNOR2_X1 U10019 ( .A(n7660), .B(n7659), .ZN(n10962) );
  NAND2_X1 U10020 ( .A1(n10962), .A2(n6389), .ZN(n7666) );
  INV_X1 U10021 ( .A(n7661), .ZN(n7663) );
  INV_X1 U10022 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U10023 ( .A1(n7663), .A2(n7662), .ZN(n7679) );
  NAND2_X1 U10024 ( .A1(n7679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7664) );
  XNOR2_X1 U10025 ( .A(n7664), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13171) );
  AOI22_X1 U10026 ( .A1(n7855), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7854), .B2(
        n13171), .ZN(n7665) );
  NAND2_X1 U10027 ( .A1(n9351), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7675) );
  INV_X1 U10028 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9961) );
  OR2_X1 U10029 ( .A1(n7577), .A2(n9961), .ZN(n7674) );
  INV_X1 U10030 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7667) );
  OAI21_X1 U10031 ( .B1(n7669), .B2(n7668), .A(n7667), .ZN(n7671) );
  INV_X1 U10032 ( .A(n7670), .ZN(n7683) );
  NAND2_X1 U10033 ( .A1(n7671), .A2(n7683), .ZN(n10760) );
  OR2_X1 U10034 ( .A1(n8036), .A2(n10760), .ZN(n7673) );
  INV_X1 U10035 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10711) );
  OR2_X1 U10036 ( .A1(n8038), .A2(n10711), .ZN(n7672) );
  NAND4_X1 U10037 ( .A1(n7675), .A2(n7674), .A3(n7673), .A4(n7672), .ZN(n13124) );
  XNOR2_X1 U10038 ( .A(n10766), .B(n13124), .ZN(n9398) );
  OR2_X1 U10039 ( .A1(n10766), .A2(n13124), .ZN(n7676) );
  NAND2_X1 U10040 ( .A1(n11081), .A2(n6390), .ZN(n7682) );
  NAND2_X1 U10041 ( .A1(n7692), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7680) );
  XNOR2_X1 U10042 ( .A(n7680), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U10043 ( .A1(n7855), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7854), .B2(
        n9981), .ZN(n7681) );
  NAND2_X1 U10044 ( .A1(n9351), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7688) );
  INV_X1 U10045 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9965) );
  OR2_X1 U10046 ( .A1(n7577), .A2(n9965), .ZN(n7687) );
  INV_X1 U10047 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n12615) );
  NAND2_X1 U10048 ( .A1(n7683), .A2(n12615), .ZN(n7684) );
  NAND2_X1 U10049 ( .A1(n7701), .A2(n7684), .ZN(n10854) );
  OR2_X1 U10050 ( .A1(n8036), .A2(n10854), .ZN(n7686) );
  INV_X1 U10051 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9954) );
  OR2_X1 U10052 ( .A1(n8038), .A2(n9954), .ZN(n7685) );
  NAND4_X1 U10053 ( .A1(n7688), .A2(n7687), .A3(n7686), .A4(n7685), .ZN(n13123) );
  INV_X1 U10054 ( .A(n13123), .ZN(n10831) );
  XNOR2_X1 U10055 ( .A(n10853), .B(n10831), .ZN(n9400) );
  INV_X1 U10056 ( .A(n9400), .ZN(n10843) );
  NAND2_X1 U10057 ( .A1(n10853), .A2(n13123), .ZN(n7689) );
  XNOR2_X1 U10058 ( .A(n7691), .B(n7690), .ZN(n11086) );
  NAND2_X1 U10059 ( .A1(n11086), .A2(n6390), .ZN(n7699) );
  INV_X1 U10060 ( .A(n7692), .ZN(n7694) );
  INV_X1 U10061 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U10062 ( .A1(n7694), .A2(n7693), .ZN(n7696) );
  NAND2_X1 U10063 ( .A1(n7696), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7695) );
  MUX2_X1 U10064 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7695), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7697) );
  AOI22_X1 U10065 ( .A1(n7855), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7854), .B2(
        n9984), .ZN(n7698) );
  NAND2_X1 U10066 ( .A1(n9351), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7706) );
  INV_X1 U10067 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9976) );
  OR2_X1 U10068 ( .A1(n7577), .A2(n9976), .ZN(n7705) );
  NAND2_X1 U10069 ( .A1(n7701), .A2(n7700), .ZN(n7702) );
  NAND2_X1 U10070 ( .A1(n7716), .A2(n7702), .ZN(n10911) );
  OR2_X1 U10071 ( .A1(n8036), .A2(n10911), .ZN(n7704) );
  INV_X1 U10072 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10835) );
  OR2_X1 U10073 ( .A1(n8038), .A2(n10835), .ZN(n7703) );
  NAND4_X1 U10074 ( .A1(n7706), .A2(n7705), .A3(n7704), .A4(n7703), .ZN(n13122) );
  XNOR2_X1 U10075 ( .A(n11003), .B(n10937), .ZN(n10829) );
  NAND2_X1 U10076 ( .A1(n10828), .A2(n10829), .ZN(n7708) );
  NAND2_X1 U10077 ( .A1(n11003), .A2(n13122), .ZN(n7707) );
  NAND2_X1 U10078 ( .A1(n7708), .A2(n7707), .ZN(n10934) );
  XNOR2_X1 U10079 ( .A(n7710), .B(n7709), .ZN(n11164) );
  NAND2_X1 U10080 ( .A1(n11164), .A2(n6390), .ZN(n7713) );
  NAND2_X1 U10081 ( .A1(n7729), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7711) );
  XNOR2_X1 U10082 ( .A(n7711), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U10083 ( .A1(n7855), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10090), 
        .B2(n7854), .ZN(n7712) );
  NAND2_X1 U10084 ( .A1(n9351), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7721) );
  INV_X1 U10085 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9978) );
  OR2_X1 U10086 ( .A1(n7577), .A2(n9978), .ZN(n7720) );
  INV_X1 U10087 ( .A(n7714), .ZN(n7735) );
  NAND2_X1 U10088 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  NAND2_X1 U10089 ( .A1(n7735), .A2(n7717), .ZN(n10941) );
  OR2_X1 U10090 ( .A1(n8036), .A2(n10941), .ZN(n7719) );
  INV_X1 U10091 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10942) );
  OR2_X1 U10092 ( .A1(n8038), .A2(n10942), .ZN(n7718) );
  NAND4_X1 U10093 ( .A1(n7721), .A2(n7720), .A3(n7719), .A4(n7718), .ZN(n13121) );
  XNOR2_X1 U10094 ( .A(n10945), .B(n10912), .ZN(n10935) );
  NAND2_X1 U10095 ( .A1(n10945), .A2(n13121), .ZN(n7722) );
  NAND2_X1 U10096 ( .A1(n9351), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7726) );
  INV_X1 U10097 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10091) );
  OR2_X1 U10098 ( .A1(n7577), .A2(n10091), .ZN(n7725) );
  INV_X1 U10099 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7734) );
  XNOR2_X1 U10100 ( .A(n7735), .B(n7734), .ZN(n11240) );
  OR2_X1 U10101 ( .A1(n8036), .A2(n11240), .ZN(n7724) );
  INV_X1 U10102 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11241) );
  OR2_X1 U10103 ( .A1(n8038), .A2(n11241), .ZN(n7723) );
  NAND4_X1 U10104 ( .A1(n7726), .A2(n7725), .A3(n7724), .A4(n7723), .ZN(n13120) );
  XNOR2_X1 U10105 ( .A(n7728), .B(n7727), .ZN(n11171) );
  NAND2_X1 U10106 ( .A1(n11171), .A2(n6390), .ZN(n7732) );
  OAI21_X1 U10107 ( .B1(n7729), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7730) );
  XNOR2_X1 U10108 ( .A(n7730), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U10109 ( .A1(n7854), .A2(n11384), .B1(n7855), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U10110 ( .A1(n9351), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7741) );
  INV_X1 U10111 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11387) );
  OR2_X1 U10112 ( .A1(n7577), .A2(n11387), .ZN(n7740) );
  INV_X1 U10113 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7733) );
  OAI21_X1 U10114 ( .B1(n7735), .B2(n7734), .A(n7733), .ZN(n7737) );
  INV_X1 U10115 ( .A(n7736), .ZN(n7748) );
  NAND2_X1 U10116 ( .A1(n7737), .A2(n7748), .ZN(n11355) );
  OR2_X1 U10117 ( .A1(n8036), .A2(n11355), .ZN(n7739) );
  INV_X1 U10118 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11356) );
  OR2_X1 U10119 ( .A1(n7578), .A2(n11356), .ZN(n7738) );
  NAND4_X1 U10120 ( .A1(n7741), .A2(n7740), .A3(n7739), .A4(n7738), .ZN(n13119) );
  XNOR2_X1 U10121 ( .A(n7742), .B(n7413), .ZN(n11277) );
  NAND2_X1 U10122 ( .A1(n11277), .A2(n6390), .ZN(n7746) );
  XNOR2_X1 U10123 ( .A(n7744), .B(P2_IR_REG_12__SCAN_IN), .ZN(n14742) );
  AOI22_X1 U10124 ( .A1(n7855), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7854), 
        .B2(n14742), .ZN(n7745) );
  NAND2_X1 U10125 ( .A1(n9351), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7753) );
  INV_X1 U10126 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11390) );
  OR2_X1 U10127 ( .A1(n7577), .A2(n11390), .ZN(n7752) );
  INV_X1 U10128 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7747) );
  NAND2_X1 U10129 ( .A1(n7748), .A2(n7747), .ZN(n7749) );
  NAND2_X1 U10130 ( .A1(n7775), .A2(n7749), .ZN(n11414) );
  OR2_X1 U10131 ( .A1(n8036), .A2(n11414), .ZN(n7751) );
  INV_X1 U10132 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11415) );
  OR2_X1 U10133 ( .A1(n8038), .A2(n11415), .ZN(n7750) );
  NAND4_X1 U10134 ( .A1(n7753), .A2(n7752), .A3(n7751), .A4(n7750), .ZN(n13118) );
  XNOR2_X1 U10135 ( .A(n7754), .B(n6443), .ZN(n11284) );
  NAND2_X1 U10136 ( .A1(n11284), .A2(n6390), .ZN(n7758) );
  INV_X1 U10137 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U10138 ( .A1(n7766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7756) );
  XNOR2_X1 U10139 ( .A(n7756), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U10140 ( .A1(n7855), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7854), 
        .B2(n11389), .ZN(n7757) );
  INV_X1 U10141 ( .A(n11420), .ZN(n14438) );
  NAND2_X1 U10142 ( .A1(n7759), .A2(n14438), .ZN(n7763) );
  INV_X1 U10143 ( .A(n11413), .ZN(n7761) );
  INV_X1 U10144 ( .A(n13118), .ZN(n7760) );
  NAND2_X1 U10145 ( .A1(n7761), .A2(n7760), .ZN(n7762) );
  NAND2_X1 U10146 ( .A1(n7763), .A2(n7762), .ZN(n11491) );
  NAND2_X1 U10147 ( .A1(n7764), .A2(n8386), .ZN(n7782) );
  NAND2_X1 U10148 ( .A1(n7782), .A2(n7765), .ZN(n7784) );
  XNOR2_X1 U10149 ( .A(n7784), .B(n7783), .ZN(n11516) );
  NAND2_X1 U10150 ( .A1(n11516), .A2(n6390), .ZN(n7772) );
  INV_X1 U10151 ( .A(n7766), .ZN(n7768) );
  NAND2_X1 U10152 ( .A1(n7768), .A2(n7767), .ZN(n7975) );
  NAND2_X1 U10153 ( .A1(n7975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7769) );
  XNOR2_X1 U10154 ( .A(n7769), .B(n7817), .ZN(n14772) );
  INV_X1 U10155 ( .A(n14772), .ZN(n7770) );
  AOI22_X1 U10156 ( .A1(n7855), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7854), 
        .B2(n7770), .ZN(n7771) );
  NAND2_X1 U10157 ( .A1(n9351), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7780) );
  INV_X1 U10158 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7773) );
  OR2_X1 U10159 ( .A1(n7577), .A2(n7773), .ZN(n7779) );
  NAND2_X1 U10160 ( .A1(n7775), .A2(n7774), .ZN(n7776) );
  NAND2_X1 U10161 ( .A1(n7793), .A2(n7776), .ZN(n11561) );
  OR2_X1 U10162 ( .A1(n8036), .A2(n11561), .ZN(n7778) );
  INV_X1 U10163 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11485) );
  OR2_X1 U10164 ( .A1(n8038), .A2(n11485), .ZN(n7777) );
  NAND4_X1 U10165 ( .A1(n7780), .A2(n7779), .A3(n7778), .A4(n7777), .ZN(n13117) );
  XNOR2_X1 U10166 ( .A(n11490), .B(n11605), .ZN(n9405) );
  NAND2_X1 U10167 ( .A1(n11490), .A2(n13117), .ZN(n7781) );
  INV_X1 U10168 ( .A(n7785), .ZN(n7786) );
  NAND2_X1 U10169 ( .A1(n11520), .A2(n7626), .ZN(n7791) );
  INV_X1 U10170 ( .A(n7975), .ZN(n7788) );
  NAND2_X1 U10171 ( .A1(n7788), .A2(n7817), .ZN(n7802) );
  NAND2_X1 U10172 ( .A1(n7802), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7789) );
  XNOR2_X1 U10173 ( .A(n7789), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14774) );
  AOI22_X1 U10174 ( .A1(n7855), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7854), 
        .B2(n14774), .ZN(n7790) );
  NAND2_X1 U10175 ( .A1(n9351), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7798) );
  INV_X1 U10176 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7792) );
  OR2_X1 U10177 ( .A1(n7577), .A2(n7792), .ZN(n7797) );
  NAND2_X1 U10178 ( .A1(n7793), .A2(n11604), .ZN(n7794) );
  NAND2_X1 U10179 ( .A1(n7808), .A2(n7794), .ZN(n11606) );
  OR2_X1 U10180 ( .A1(n8036), .A2(n11606), .ZN(n7796) );
  INV_X1 U10181 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11594) );
  OR2_X1 U10182 ( .A1(n7578), .A2(n11594), .ZN(n7795) );
  NAND4_X1 U10183 ( .A1(n7798), .A2(n7797), .A3(n7796), .A4(n7795), .ZN(n13116) );
  XNOR2_X1 U10184 ( .A(n11610), .B(n13116), .ZN(n9406) );
  OR2_X1 U10185 ( .A1(n11610), .A2(n13116), .ZN(n7800) );
  XNOR2_X1 U10186 ( .A(n7801), .B(n7415), .ZN(n11686) );
  NAND2_X1 U10187 ( .A1(n11686), .A2(n6390), .ZN(n7805) );
  OAI21_X1 U10188 ( .B1(n7802), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7803) );
  XNOR2_X1 U10189 ( .A(n7803), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U10190 ( .A1(n7855), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7854), 
        .B2(n11383), .ZN(n7804) );
  NAND2_X1 U10191 ( .A1(n9351), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7813) );
  INV_X1 U10192 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11396) );
  OR2_X1 U10193 ( .A1(n7577), .A2(n11396), .ZN(n7812) );
  INV_X1 U10194 ( .A(n7806), .ZN(n7829) );
  NAND2_X1 U10195 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  NAND2_X1 U10196 ( .A1(n7829), .A2(n7809), .ZN(n13413) );
  OR2_X1 U10197 ( .A1(n8036), .A2(n13413), .ZN(n7811) );
  INV_X1 U10198 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13414) );
  OR2_X1 U10199 ( .A1(n8038), .A2(n13414), .ZN(n7810) );
  NAND4_X1 U10200 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n13115) );
  XNOR2_X1 U10201 ( .A(n13505), .B(n13115), .ZN(n13401) );
  INV_X1 U10202 ( .A(n13401), .ZN(n13411) );
  XNOR2_X1 U10203 ( .A(n7814), .B(SI_17_), .ZN(n7815) );
  XNOR2_X1 U10204 ( .A(n7816), .B(n7815), .ZN(n11742) );
  NAND2_X1 U10205 ( .A1(n11742), .A2(n7626), .ZN(n7827) );
  AND3_X1 U10206 ( .A1(n7819), .A2(n7818), .A3(n7817), .ZN(n7820) );
  NAND2_X1 U10207 ( .A1(n7822), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7821) );
  MUX2_X1 U10208 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7821), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7825) );
  AND2_X1 U10209 ( .A1(n7825), .A2(n7840), .ZN(n11382) );
  AOI22_X1 U10210 ( .A1(n7855), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7854), 
        .B2(n11382), .ZN(n7826) );
  NAND2_X1 U10211 ( .A1(n9351), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7834) );
  INV_X1 U10212 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11397) );
  OR2_X1 U10213 ( .A1(n7577), .A2(n11397), .ZN(n7833) );
  INV_X1 U10214 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U10215 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  NAND2_X1 U10216 ( .A1(n7845), .A2(n7830), .ZN(n13391) );
  OR2_X1 U10217 ( .A1(n8036), .A2(n13391), .ZN(n7832) );
  INV_X1 U10218 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13392) );
  OR2_X1 U10219 ( .A1(n8038), .A2(n13392), .ZN(n7831) );
  NAND4_X1 U10220 ( .A1(n7834), .A2(n7833), .A3(n7832), .A4(n7831), .ZN(n13114) );
  XNOR2_X1 U10221 ( .A(n13500), .B(n13114), .ZN(n9408) );
  NAND2_X1 U10222 ( .A1(n13390), .A2(n13389), .ZN(n13388) );
  NAND2_X1 U10223 ( .A1(n13500), .A2(n13114), .ZN(n7835) );
  NAND2_X1 U10224 ( .A1(n13388), .A2(n7835), .ZN(n13372) );
  NAND2_X1 U10225 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  NAND2_X1 U10226 ( .A1(n7839), .A2(n7838), .ZN(n11753) );
  OR2_X1 U10227 ( .A1(n11753), .A2(n7595), .ZN(n7843) );
  NAND2_X1 U10228 ( .A1(n7840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7841) );
  XNOR2_X1 U10229 ( .A(n7841), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14818) );
  AOI22_X1 U10230 ( .A1(n7855), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7854), 
        .B2(n14818), .ZN(n7842) );
  NAND2_X1 U10231 ( .A1(n7845), .A2(n7844), .ZN(n7846) );
  NAND2_X1 U10232 ( .A1(n7860), .A2(n7846), .ZN(n13377) );
  NAND2_X1 U10233 ( .A1(n9351), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7847) );
  OAI21_X1 U10234 ( .B1(n13377), .B2(n8036), .A(n7847), .ZN(n7849) );
  INV_X1 U10235 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13495) );
  INV_X1 U10236 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13378) );
  OAI22_X1 U10237 ( .A1(n7577), .A2(n13495), .B1(n8038), .B2(n13378), .ZN(
        n7848) );
  INV_X1 U10238 ( .A(n13113), .ZN(n13349) );
  XNOR2_X1 U10239 ( .A(n13375), .B(n13349), .ZN(n9410) );
  OR2_X1 U10240 ( .A1(n13375), .A2(n13113), .ZN(n7850) );
  XNOR2_X1 U10241 ( .A(n7852), .B(n7851), .ZN(n11772) );
  NAND2_X1 U10242 ( .A1(n11772), .A2(n6390), .ZN(n7857) );
  AOI22_X1 U10243 ( .A1(n7855), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9423), 
        .B2(n7854), .ZN(n7856) );
  INV_X1 U10244 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13362) );
  INV_X1 U10245 ( .A(n7858), .ZN(n7872) );
  NAND2_X1 U10246 ( .A1(n7860), .A2(n7859), .ZN(n7861) );
  NAND2_X1 U10247 ( .A1(n7872), .A2(n7861), .ZN(n13361) );
  OR2_X1 U10248 ( .A1(n13361), .A2(n8036), .ZN(n7864) );
  AOI22_X1 U10249 ( .A1(n7887), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9351), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n7863) );
  OAI211_X1 U10250 ( .C1(n8038), .C2(n13362), .A(n7864), .B(n7863), .ZN(n13112) );
  INV_X1 U10251 ( .A(n13112), .ZN(n13333) );
  NAND2_X1 U10252 ( .A1(n7866), .A2(n7865), .ZN(n7867) );
  NAND2_X1 U10253 ( .A1(n7868), .A2(n7867), .ZN(n11794) );
  OR2_X1 U10254 ( .A1(n11794), .A2(n7595), .ZN(n7870) );
  OR2_X1 U10255 ( .A1(n6410), .A2(n12660), .ZN(n7869) );
  INV_X1 U10256 ( .A(n7885), .ZN(n7874) );
  INV_X1 U10257 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10258 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  NAND2_X1 U10259 ( .A1(n7874), .A2(n7873), .ZN(n13338) );
  AOI22_X1 U10260 ( .A1(n7887), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n7875), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U10261 ( .A1(n9351), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7876) );
  OAI211_X1 U10262 ( .C1(n13338), .C2(n8036), .A(n7877), .B(n7876), .ZN(n13310) );
  INV_X1 U10263 ( .A(n13310), .ZN(n13350) );
  NAND2_X1 U10264 ( .A1(n13540), .A2(n13350), .ZN(n7878) );
  OR2_X1 U10265 ( .A1(n7880), .A2(n7879), .ZN(n7881) );
  AND2_X1 U10266 ( .A1(n7882), .A2(n7881), .ZN(n11812) );
  NAND2_X1 U10267 ( .A1(n11812), .A2(n6390), .ZN(n7884) );
  OR2_X1 U10268 ( .A1(n6410), .A2(n11326), .ZN(n7883) );
  NOR2_X1 U10269 ( .A1(n7885), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7886) );
  OR2_X1 U10270 ( .A1(n7898), .A2(n7886), .ZN(n13321) );
  INV_X1 U10271 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U10272 ( .A1(n9351), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U10273 ( .A1(n7887), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7888) );
  OAI211_X1 U10274 ( .C1(n13320), .C2(n8038), .A(n7889), .B(n7888), .ZN(n7890)
         );
  INV_X1 U10275 ( .A(n7890), .ZN(n7891) );
  OAI21_X1 U10276 ( .B1(n13321), .B2(n8036), .A(n7891), .ZN(n13111) );
  XNOR2_X1 U10277 ( .A(n13319), .B(n13111), .ZN(n13307) );
  INV_X1 U10278 ( .A(n13307), .ZN(n13316) );
  OR2_X1 U10279 ( .A1(n13319), .A2(n13111), .ZN(n7892) );
  NAND2_X1 U10280 ( .A1(n11833), .A2(n7893), .ZN(n7894) );
  AND2_X1 U10281 ( .A1(n7895), .A2(n7894), .ZN(n11469) );
  NAND2_X1 U10282 ( .A1(n11469), .A2(n7626), .ZN(n7897) );
  OR2_X1 U10283 ( .A1(n6410), .A2(n11470), .ZN(n7896) );
  OR2_X1 U10284 ( .A1(n7898), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n7900) );
  AND2_X1 U10285 ( .A1(n7900), .A2(n7899), .ZN(n13302) );
  INV_X1 U10286 ( .A(n8036), .ZN(n7901) );
  NAND2_X1 U10287 ( .A1(n13302), .A2(n7901), .ZN(n7907) );
  INV_X1 U10288 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U10289 ( .A1(n9351), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U10290 ( .A1(n7875), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7902) );
  OAI211_X1 U10291 ( .C1(n7577), .C2(n7904), .A(n7903), .B(n7902), .ZN(n7905)
         );
  INV_X1 U10292 ( .A(n7905), .ZN(n7906) );
  NAND2_X1 U10293 ( .A1(n7907), .A2(n7906), .ZN(n13313) );
  XNOR2_X1 U10294 ( .A(n13299), .B(n13313), .ZN(n13293) );
  NAND2_X1 U10295 ( .A1(n13299), .A2(n13313), .ZN(n7908) );
  INV_X1 U10296 ( .A(n11850), .ZN(n7912) );
  OR2_X1 U10297 ( .A1(n6410), .A2(n8118), .ZN(n7913) );
  NAND2_X1 U10298 ( .A1(n9351), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7921) );
  INV_X1 U10299 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n7915) );
  OR2_X1 U10300 ( .A1(n7577), .A2(n7915), .ZN(n7920) );
  OAI21_X1 U10301 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n7917), .A(n7916), .ZN(
        n13286) );
  OR2_X1 U10302 ( .A1(n7599), .A2(n13286), .ZN(n7919) );
  INV_X1 U10303 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13280) );
  OR2_X1 U10304 ( .A1(n8038), .A2(n13280), .ZN(n7918) );
  NAND4_X1 U10305 ( .A1(n7921), .A2(n7920), .A3(n7919), .A4(n7918), .ZN(n13110) );
  NAND2_X1 U10306 ( .A1(n13281), .A2(n7922), .ZN(n7923) );
  NAND2_X1 U10307 ( .A1(n13568), .A2(n6389), .ZN(n7929) );
  INV_X1 U10308 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13569) );
  OR2_X1 U10309 ( .A1(n6410), .A2(n13569), .ZN(n7928) );
  NAND2_X1 U10310 ( .A1(n9351), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7935) );
  INV_X1 U10311 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13456) );
  OR2_X1 U10312 ( .A1(n7577), .A2(n13456), .ZN(n7934) );
  OAI21_X1 U10313 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n7931), .A(n7930), .ZN(
        n13247) );
  OR2_X1 U10314 ( .A1(n8036), .A2(n13247), .ZN(n7933) );
  INV_X1 U10315 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13248) );
  OR2_X1 U10316 ( .A1(n8038), .A2(n13248), .ZN(n7932) );
  NAND4_X1 U10317 ( .A1(n7935), .A2(n7934), .A3(n7933), .A4(n7932), .ZN(n13108) );
  NOR2_X1 U10318 ( .A1(n13246), .A2(n13108), .ZN(n7936) );
  INV_X1 U10319 ( .A(n7937), .ZN(n7938) );
  NAND2_X1 U10320 ( .A1(n7938), .A2(SI_26_), .ZN(n7939) );
  MUX2_X1 U10321 ( .A(n13563), .B(n7103), .S(n9812), .Z(n7941) );
  INV_X1 U10322 ( .A(SI_27_), .ZN(n12986) );
  NAND2_X1 U10323 ( .A1(n7941), .A2(n12986), .ZN(n7955) );
  INV_X1 U10324 ( .A(n7941), .ZN(n7942) );
  NAND2_X1 U10325 ( .A1(n7942), .A2(SI_27_), .ZN(n7943) );
  NAND2_X1 U10326 ( .A1(n7955), .A2(n7943), .ZN(n7956) );
  NAND2_X1 U10327 ( .A1(n13562), .A2(n6390), .ZN(n7945) );
  OR2_X1 U10328 ( .A1(n6410), .A2(n13563), .ZN(n7944) );
  NAND2_X2 U10329 ( .A1(n7945), .A2(n7944), .ZN(n13444) );
  NAND2_X1 U10330 ( .A1(n9351), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7954) );
  INV_X1 U10331 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7946) );
  OR2_X1 U10332 ( .A1(n7577), .A2(n7946), .ZN(n7953) );
  INV_X1 U10333 ( .A(n7949), .ZN(n7947) );
  INV_X1 U10334 ( .A(n7963), .ZN(n7965) );
  INV_X1 U10335 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U10336 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  NAND2_X1 U10337 ( .A1(n7965), .A2(n7950), .ZN(n13212) );
  OR2_X1 U10338 ( .A1(n8036), .A2(n13212), .ZN(n7952) );
  INV_X1 U10339 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13213) );
  OR2_X1 U10340 ( .A1(n8038), .A2(n13213), .ZN(n7951) );
  NAND4_X1 U10341 ( .A1(n7954), .A2(n7953), .A3(n7952), .A4(n7951), .ZN(n13106) );
  INV_X1 U10342 ( .A(n13206), .ZN(n13210) );
  INV_X1 U10343 ( .A(n13444), .ZN(n13215) );
  INV_X1 U10344 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13560) );
  MUX2_X1 U10345 ( .A(n13560), .B(n14236), .S(n9828), .Z(n7958) );
  INV_X1 U10346 ( .A(SI_28_), .ZN(n12983) );
  NAND2_X1 U10347 ( .A1(n7958), .A2(n12983), .ZN(n8692) );
  INV_X1 U10348 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U10349 ( .A1(n7959), .A2(SI_28_), .ZN(n7960) );
  NAND2_X1 U10350 ( .A1(n14235), .A2(n6390), .ZN(n7962) );
  OR2_X1 U10351 ( .A1(n6410), .A2(n13560), .ZN(n7961) );
  NAND2_X1 U10352 ( .A1(n9351), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7970) );
  INV_X1 U10353 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8926) );
  OR2_X1 U10354 ( .A1(n7577), .A2(n8926), .ZN(n7969) );
  NAND2_X1 U10355 ( .A1(n7963), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8718) );
  INV_X1 U10356 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10357 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  NAND2_X1 U10358 ( .A1(n8718), .A2(n7966), .ZN(n13193) );
  OR2_X1 U10359 ( .A1(n7599), .A2(n13193), .ZN(n7968) );
  INV_X1 U10360 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13197) );
  OR2_X1 U10361 ( .A1(n8038), .A2(n13197), .ZN(n7967) );
  NAND4_X1 U10362 ( .A1(n7970), .A2(n7969), .A3(n7968), .A4(n7967), .ZN(n13105) );
  NAND2_X1 U10363 ( .A1(n13199), .A2(n13105), .ZN(n8688) );
  OR2_X1 U10364 ( .A1(n13199), .A2(n13105), .ZN(n7971) );
  NAND2_X1 U10365 ( .A1(n8688), .A2(n7971), .ZN(n9415) );
  INV_X1 U10366 ( .A(n9415), .ZN(n7972) );
  OAI21_X1 U10367 ( .B1(n7973), .B2(n7972), .A(n8689), .ZN(n13196) );
  OAI21_X1 U10368 ( .B1(n7975), .B2(n7974), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7976) );
  NAND2_X1 U10369 ( .A1(n7980), .A2(n12614), .ZN(n7978) );
  NAND2_X2 U10370 ( .A1(n7979), .A2(n7412), .ZN(n11059) );
  NAND2_X1 U10371 ( .A1(n7982), .A2(n7981), .ZN(n8062) );
  INV_X1 U10372 ( .A(n9151), .ZN(n10254) );
  NAND2_X1 U10373 ( .A1(n7977), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7983) );
  XNOR2_X2 U10374 ( .A(n7983), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9428) );
  XNOR2_X1 U10375 ( .A(n9500), .B(n9436), .ZN(n7984) );
  INV_X1 U10376 ( .A(n13267), .ZN(n13461) );
  NAND2_X1 U10377 ( .A1(n7587), .A2(n10014), .ZN(n10260) );
  INV_X1 U10378 ( .A(n10766), .ZN(n10723) );
  INV_X1 U10379 ( .A(n10853), .ZN(n14842) );
  NAND2_X1 U10380 ( .A1(n10849), .A2(n14842), .ZN(n10850) );
  OR2_X2 U10381 ( .A1(n11416), .A2(n11420), .ZN(n11486) );
  OR2_X2 U10382 ( .A1(n11486), .A2(n11490), .ZN(n11595) );
  INV_X1 U10383 ( .A(n13505), .ZN(n13417) );
  NAND2_X1 U10384 ( .A1(n13544), .A2(n13374), .ZN(n13357) );
  NAND2_X1 U10385 ( .A1(n13461), .A2(n13279), .ZN(n13262) );
  OR2_X2 U10386 ( .A1(n13262), .A2(n13246), .ZN(n13244) );
  NOR2_X2 U10387 ( .A1(n9436), .A2(n9428), .ZN(n10242) );
  OAI21_X1 U10388 ( .B1(n13216), .B2(n8925), .A(n13420), .ZN(n7985) );
  OAI21_X1 U10389 ( .B1(n13196), .B2(n14428), .A(n13201), .ZN(n8045) );
  INV_X1 U10390 ( .A(n9157), .ZN(n7987) );
  NAND2_X1 U10391 ( .A1(n7987), .A2(n10243), .ZN(n10235) );
  INV_X1 U10392 ( .A(n10235), .ZN(n7988) );
  NAND2_X1 U10393 ( .A1(n9394), .A2(n7988), .ZN(n10233) );
  OR2_X1 U10394 ( .A1(n13129), .A2(n10554), .ZN(n7989) );
  NAND2_X1 U10395 ( .A1(n10233), .A2(n7989), .ZN(n10262) );
  NAND2_X1 U10396 ( .A1(n10262), .A2(n9393), .ZN(n7991) );
  OR2_X1 U10397 ( .A1(n9166), .A2(n7605), .ZN(n7990) );
  NAND2_X1 U10398 ( .A1(n7991), .A2(n7990), .ZN(n10367) );
  INV_X1 U10399 ( .A(n10366), .ZN(n7992) );
  NAND2_X1 U10400 ( .A1(n10367), .A2(n7992), .ZN(n7994) );
  OR2_X1 U10401 ( .A1(n13128), .A2(n10563), .ZN(n7993) );
  NAND2_X1 U10402 ( .A1(n7994), .A2(n7993), .ZN(n10447) );
  INV_X1 U10403 ( .A(n10446), .ZN(n7995) );
  NAND2_X1 U10404 ( .A1(n10447), .A2(n7995), .ZN(n7997) );
  OR2_X1 U10405 ( .A1(n13127), .A2(n10559), .ZN(n7996) );
  NAND2_X1 U10406 ( .A1(n7997), .A2(n7996), .ZN(n10595) );
  INV_X1 U10407 ( .A(n13126), .ZN(n7998) );
  NAND2_X1 U10408 ( .A1(n7998), .A2(n10623), .ZN(n7999) );
  INV_X1 U10409 ( .A(n13125), .ZN(n9194) );
  INV_X1 U10410 ( .A(n13124), .ZN(n10752) );
  AND2_X1 U10411 ( .A1(n10766), .A2(n10752), .ZN(n8000) );
  NAND2_X1 U10412 ( .A1(n10844), .A2(n10843), .ZN(n8002) );
  OR2_X1 U10413 ( .A1(n10853), .A2(n10831), .ZN(n8001) );
  NAND2_X1 U10414 ( .A1(n8002), .A2(n8001), .ZN(n10830) );
  INV_X1 U10415 ( .A(n10829), .ZN(n8003) );
  NAND2_X1 U10416 ( .A1(n10830), .A2(n8003), .ZN(n8005) );
  OR2_X1 U10417 ( .A1(n11003), .A2(n10937), .ZN(n8004) );
  NAND2_X1 U10418 ( .A1(n8005), .A2(n8004), .ZN(n10936) );
  INV_X1 U10419 ( .A(n10935), .ZN(n8006) );
  NAND2_X1 U10420 ( .A1(n10936), .A2(n8006), .ZN(n8008) );
  OR2_X1 U10421 ( .A1(n10945), .A2(n10912), .ZN(n8007) );
  INV_X1 U10422 ( .A(n13120), .ZN(n11351) );
  NAND2_X1 U10423 ( .A1(n11337), .A2(n11351), .ZN(n8010) );
  OR2_X1 U10424 ( .A1(n11337), .A2(n11351), .ZN(n8009) );
  NAND2_X1 U10425 ( .A1(n8010), .A2(n8009), .ZN(n11234) );
  OR2_X1 U10426 ( .A1(n11360), .A2(n11225), .ZN(n8011) );
  NAND2_X1 U10427 ( .A1(n11360), .A2(n11225), .ZN(n8012) );
  NAND2_X1 U10428 ( .A1(n8013), .A2(n8012), .ZN(n11409) );
  OR2_X1 U10429 ( .A1(n11420), .A2(n7760), .ZN(n9402) );
  NAND2_X1 U10430 ( .A1(n11409), .A2(n9402), .ZN(n8014) );
  NAND2_X1 U10431 ( .A1(n11420), .A2(n7760), .ZN(n9401) );
  NAND2_X1 U10432 ( .A1(n8014), .A2(n9401), .ZN(n11483) );
  NAND2_X1 U10433 ( .A1(n11490), .A2(n11605), .ZN(n8015) );
  INV_X1 U10434 ( .A(n13116), .ZN(n13403) );
  INV_X1 U10435 ( .A(n13402), .ZN(n8016) );
  INV_X1 U10436 ( .A(n13115), .ZN(n11607) );
  NAND2_X1 U10437 ( .A1(n13505), .A2(n11607), .ZN(n8017) );
  NAND2_X1 U10438 ( .A1(n8018), .A2(n8017), .ZN(n13385) );
  INV_X1 U10439 ( .A(n13114), .ZN(n13407) );
  AND2_X1 U10440 ( .A1(n13500), .A2(n13407), .ZN(n8020) );
  OR2_X1 U10441 ( .A1(n13500), .A2(n13407), .ZN(n8019) );
  NOR2_X1 U10442 ( .A1(n13375), .A2(n13349), .ZN(n8021) );
  NAND2_X1 U10443 ( .A1(n13375), .A2(n13349), .ZN(n8022) );
  AND2_X1 U10444 ( .A1(n13360), .A2(n13333), .ZN(n8023) );
  INV_X1 U10445 ( .A(n13330), .ZN(n8026) );
  NAND2_X1 U10446 ( .A1(n13540), .A2(n13310), .ZN(n8024) );
  NAND2_X1 U10447 ( .A1(n13337), .A2(n13350), .ZN(n8027) );
  NAND2_X1 U10448 ( .A1(n8024), .A2(n8027), .ZN(n13331) );
  NAND2_X1 U10449 ( .A1(n8026), .A2(n8025), .ZN(n13328) );
  NAND2_X1 U10450 ( .A1(n13328), .A2(n8027), .ZN(n13308) );
  INV_X1 U10451 ( .A(n13111), .ZN(n13334) );
  OR2_X1 U10452 ( .A1(n13319), .A2(n13334), .ZN(n8028) );
  NOR2_X1 U10453 ( .A1(n13255), .A2(n13256), .ZN(n13254) );
  XNOR2_X1 U10454 ( .A(n13246), .B(n13108), .ZN(n9413) );
  OR2_X1 U10455 ( .A1(n13229), .A2(n13243), .ZN(n9390) );
  INV_X1 U10456 ( .A(n9390), .ZN(n8030) );
  NAND2_X1 U10457 ( .A1(n13229), .A2(n13243), .ZN(n9389) );
  INV_X1 U10458 ( .A(n9428), .ZN(n11328) );
  NAND2_X1 U10459 ( .A1(n9436), .A2(n9423), .ZN(n8031) );
  OAI21_X2 U10460 ( .B1(n11059), .B2(n11328), .A(n8031), .ZN(n13352) );
  OAI211_X1 U10461 ( .C1(n8032), .C2(n9415), .A(n8705), .B(n13352), .ZN(n8044)
         );
  INV_X1 U10462 ( .A(n9869), .ZN(n8034) );
  NAND2_X1 U10463 ( .A1(n9351), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8042) );
  INV_X1 U10464 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8035) );
  OR2_X1 U10465 ( .A1(n7577), .A2(n8035), .ZN(n8041) );
  OR2_X1 U10466 ( .A1(n8036), .A2(n8718), .ZN(n8040) );
  INV_X1 U10467 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8037) );
  OR2_X1 U10468 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  AND4_X1 U10469 ( .A1(n8042), .A2(n8041), .A3(n8040), .A4(n8039), .ZN(n9363)
         );
  NAND2_X1 U10470 ( .A1(n9869), .A2(n9864), .ZN(n13408) );
  OAI22_X1 U10471 ( .A1(n13223), .A2(n13404), .B1(n9363), .B2(n13408), .ZN(
        n13030) );
  INV_X1 U10472 ( .A(n13030), .ZN(n8043) );
  NAND2_X1 U10473 ( .A1(n8044), .A2(n8043), .ZN(n13194) );
  NOR2_X1 U10474 ( .A1(n8045), .A2(n13194), .ZN(n8930) );
  OAI21_X1 U10475 ( .B1(n8062), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8046) );
  MUX2_X1 U10476 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8046), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8048) );
  INV_X1 U10477 ( .A(n8047), .ZN(n8049) );
  INV_X1 U10478 ( .A(P2_B_REG_SCAN_IN), .ZN(n8710) );
  XNOR2_X1 U10479 ( .A(n13571), .B(n8710), .ZN(n8053) );
  NAND2_X1 U10480 ( .A1(n8049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8050) );
  MUX2_X1 U10481 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8050), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8052) );
  NAND2_X1 U10482 ( .A1(n8047), .A2(n8051), .ZN(n8054) );
  NAND2_X1 U10483 ( .A1(n8052), .A2(n8054), .ZN(n13570) );
  NAND2_X1 U10484 ( .A1(n8053), .A2(n13570), .ZN(n8058) );
  NAND2_X1 U10485 ( .A1(n8054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8055) );
  MUX2_X1 U10486 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8055), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8057) );
  NAND2_X1 U10487 ( .A1(n8057), .A2(n8056), .ZN(n13567) );
  INV_X1 U10488 ( .A(n13567), .ZN(n8078) );
  AND2_X1 U10489 ( .A1(n8058), .A2(n8078), .ZN(n14829) );
  INV_X1 U10490 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14838) );
  NAND2_X1 U10491 ( .A1(n14829), .A2(n14838), .ZN(n8060) );
  NAND2_X1 U10492 ( .A1(n13567), .A2(n13570), .ZN(n8059) );
  NAND2_X1 U10493 ( .A1(n8060), .A2(n8059), .ZN(n8698) );
  NOR2_X1 U10494 ( .A1(n13567), .A2(n13570), .ZN(n8061) );
  NAND2_X1 U10495 ( .A1(n8061), .A2(n13571), .ZN(n9464) );
  NAND2_X1 U10496 ( .A1(n8062), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8064) );
  XNOR2_X1 U10497 ( .A(n8064), .B(n8063), .ZN(n9863) );
  AND2_X1 U10498 ( .A1(n9464), .A2(n9863), .ZN(n9633) );
  AND2_X1 U10499 ( .A1(n8698), .A2(n14835), .ZN(n14836) );
  NOR4_X1 U10500 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8068) );
  NOR4_X1 U10501 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8067) );
  NOR4_X1 U10502 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8066) );
  NOR4_X1 U10503 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8065) );
  AND4_X1 U10504 ( .A1(n8068), .A2(n8067), .A3(n8066), .A4(n8065), .ZN(n8074)
         );
  NOR2_X1 U10505 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n8072) );
  NOR4_X1 U10506 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n8071) );
  NOR4_X1 U10507 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8070) );
  NOR4_X1 U10508 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n8069) );
  AND4_X1 U10509 ( .A1(n8072), .A2(n8071), .A3(n8070), .A4(n8069), .ZN(n8073)
         );
  NAND2_X1 U10510 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  AND2_X1 U10511 ( .A1(n14829), .A2(n8075), .ZN(n8697) );
  NAND2_X1 U10512 ( .A1(n10242), .A2(n10245), .ZN(n9630) );
  NAND2_X1 U10513 ( .A1(n9864), .A2(n9627), .ZN(n9632) );
  NAND2_X1 U10514 ( .A1(n9630), .A2(n9632), .ZN(n8076) );
  NOR2_X1 U10515 ( .A1(n8697), .A2(n8076), .ZN(n8077) );
  AND2_X1 U10516 ( .A1(n14836), .A2(n8077), .ZN(n8924) );
  INV_X1 U10517 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14833) );
  NAND2_X1 U10518 ( .A1(n14829), .A2(n14833), .ZN(n8080) );
  OR2_X1 U10519 ( .A1(n13571), .A2(n8078), .ZN(n8079) );
  NAND2_X1 U10520 ( .A1(n8080), .A2(n8079), .ZN(n14834) );
  INV_X1 U10521 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8082) );
  NOR2_X1 U10522 ( .A1(n14457), .A2(n8082), .ZN(n8083) );
  AOI22_X1 U10523 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13566), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n6709), .ZN(n8569) );
  AOI22_X1 U10524 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n8118), .B2(n11851), .ZN(n8532) );
  AOI22_X1 U10525 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n11470), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n8085), .ZN(n8516) );
  AOI22_X1 U10526 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n12660), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n7077), .ZN(n8489) );
  AOI22_X1 U10527 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n10701), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n6707), .ZN(n8461) );
  AOI22_X1 U10528 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10589), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n6632), .ZN(n8441) );
  AOI22_X1 U10529 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n12681), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n6650), .ZN(n8397) );
  XNOR2_X1 U10530 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8382) );
  NAND2_X1 U10531 ( .A1(n12631), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8087) );
  AND2_X1 U10532 ( .A1(n9825), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U10533 ( .A1(n9827), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U10534 ( .A1(n9848), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10535 ( .A1(n8090), .A2(n8089), .ZN(n8209) );
  XNOR2_X1 U10536 ( .A(n8091), .B(P1_DATAO_REG_4__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U10537 ( .A1(n8091), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10538 ( .A1(n9834), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U10539 ( .A1(n8094), .A2(n8093), .ZN(n8241) );
  NAND2_X1 U10540 ( .A1(n9838), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10541 ( .A1(n9844), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U10542 ( .A1(n8097), .A2(n8096), .ZN(n8273) );
  XNOR2_X1 U10543 ( .A(n9852), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U10544 ( .A1(n9852), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U10545 ( .A1(n9943), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U10546 ( .A1(n8102), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U10547 ( .A1(n10102), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10548 ( .A1(n10107), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U10549 ( .A1(n8106), .A2(n8105), .ZN(n8339) );
  XNOR2_X1 U10550 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8352) );
  NAND2_X1 U10551 ( .A1(n11285), .A2(n8108), .ZN(n8109) );
  AOI22_X1 U10552 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n10424), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n12704), .ZN(n8412) );
  INV_X1 U10553 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U10554 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n10744), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n12228), .ZN(n8475) );
  INV_X1 U10555 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U10556 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(
        P1_DATAO_REG_21__SCAN_IN), .B1(n11326), .B2(n11813), .ZN(n8502) );
  NOR2_X1 U10557 ( .A1(n8532), .A2(n8531), .ZN(n8117) );
  NOR2_X1 U10558 ( .A1(n8119), .A2(n14246), .ZN(n8120) );
  AOI22_X1 U10559 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13569), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n6685), .ZN(n8556) );
  AOI22_X1 U10560 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(
        P2_DATAO_REG_28__SCAN_IN), .B1(n14236), .B2(n13560), .ZN(n8122) );
  NOR2_X1 U10561 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8136) );
  NAND2_X1 U10562 ( .A1(n12980), .A2(n8587), .ZN(n8142) );
  OR2_X1 U10563 ( .A1(n8572), .A2(n12983), .ZN(n8141) );
  NOR2_X1 U10564 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8232) );
  NAND2_X1 U10565 ( .A1(n8232), .A2(n8231), .ZN(n8249) );
  NAND2_X1 U10566 ( .A1(n8375), .A2(n12350), .ZN(n8390) );
  INV_X1 U10567 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12326) );
  INV_X1 U10568 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8453) );
  INV_X1 U10569 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8494) );
  INV_X1 U10570 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8506) );
  INV_X1 U10571 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8561) );
  INV_X1 U10572 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n8143) );
  INV_X1 U10573 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8144) );
  INV_X1 U10574 ( .A(n8166), .ZN(n8146) );
  INV_X1 U10575 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10576 ( .A1(n8146), .A2(n8145), .ZN(n12493) );
  NAND2_X1 U10577 ( .A1(n8166), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U10578 ( .A1(n12493), .A2(n8147), .ZN(n12506) );
  INV_X1 U10579 ( .A(n8152), .ZN(n8155) );
  INV_X1 U10580 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8158) );
  INV_X1 U10581 ( .A(n8153), .ZN(n8154) );
  NAND2_X2 U10582 ( .A1(n8154), .A2(n8152), .ZN(n8509) );
  AND2_X2 U10583 ( .A1(n8152), .A2(n8153), .ZN(n8588) );
  NAND2_X1 U10584 ( .A1(n8523), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10585 ( .A1(n8606), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8156) );
  OAI211_X1 U10586 ( .C1(n8158), .C2(n8946), .A(n8157), .B(n8156), .ZN(n8159)
         );
  AOI21_X1 U10587 ( .B1(n12506), .B2(n8547), .A(n8159), .ZN(n12265) );
  INV_X1 U10588 ( .A(n12265), .ZN(n12516) );
  NAND2_X1 U10589 ( .A1(n12984), .A2(n8587), .ZN(n8163) );
  OR2_X1 U10590 ( .A1(n8572), .A2(n12986), .ZN(n8162) );
  INV_X1 U10591 ( .A(n8164), .ZN(n8578) );
  NAND2_X1 U10592 ( .A1(n8578), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10593 ( .A1(n8166), .A2(n8165), .ZN(n12525) );
  INV_X1 U10594 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12913) );
  NAND2_X1 U10595 ( .A1(n8523), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10596 ( .A1(n8606), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8167) );
  OAI211_X1 U10597 ( .C1(n12913), .C2(n8946), .A(n8168), .B(n8167), .ZN(n8169)
         );
  INV_X1 U10598 ( .A(n12536), .ZN(n12397) );
  NAND2_X1 U10599 ( .A1(n6412), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U10600 ( .A1(n8588), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8173) );
  INV_X1 U10601 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8170) );
  XNOR2_X1 U10602 ( .A(n8176), .B(n8187), .ZN(n9819) );
  NAND2_X1 U10603 ( .A1(n8175), .A2(n9819), .ZN(n8181) );
  INV_X1 U10604 ( .A(SI_1_), .ZN(n9821) );
  OR2_X1 U10605 ( .A1(n8240), .A2(n9821), .ZN(n8180) );
  INV_X1 U10606 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8178) );
  OR2_X1 U10607 ( .A1(n10290), .A2(n10311), .ZN(n8179) );
  AND3_X2 U10608 ( .A1(n8181), .A2(n8180), .A3(n8179), .ZN(n12908) );
  NAND2_X1 U10609 ( .A1(n6412), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10610 ( .A1(n8588), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8183) );
  INV_X1 U10611 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10585) );
  INV_X1 U10612 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9729) );
  AND2_X1 U10613 ( .A1(n9729), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8186) );
  NOR2_X1 U10614 ( .A1(n8187), .A2(n8186), .ZN(n8188) );
  MUX2_X1 U10615 ( .A(n8189), .B(n8188), .S(n9828), .Z(n9803) );
  MUX2_X1 U10616 ( .A(n8190), .B(n9803), .S(n10290), .Z(n10588) );
  NAND2_X1 U10617 ( .A1(n15088), .A2(n15086), .ZN(n8201) );
  NAND2_X1 U10618 ( .A1(n6412), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10619 ( .A1(n8588), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8193) );
  INV_X1 U10620 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8191) );
  OR2_X1 U10621 ( .A1(n8509), .A2(n8191), .ZN(n8192) );
  NAND4_X2 U10622 ( .A1(n8195), .A2(n8194), .A3(n8193), .A4(n8192), .ZN(n15061) );
  XNOR2_X1 U10623 ( .A(n9825), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n8196) );
  XNOR2_X1 U10624 ( .A(n8197), .B(n8196), .ZN(n9807) );
  NAND2_X1 U10625 ( .A1(n8175), .A2(n9807), .ZN(n8200) );
  OR2_X1 U10626 ( .A1(n10290), .A2(n10351), .ZN(n8199) );
  NAND2_X1 U10627 ( .A1(n15061), .A2(n15077), .ZN(n8981) );
  INV_X1 U10628 ( .A(n15087), .ZN(n15074) );
  NAND2_X1 U10629 ( .A1(n8201), .A2(n15074), .ZN(n15085) );
  OR2_X1 U10630 ( .A1(n15061), .A2(n6601), .ZN(n8202) );
  NAND2_X1 U10631 ( .A1(n15085), .A2(n8202), .ZN(n15062) );
  INV_X1 U10632 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10633 ( .A1(n6412), .A2(n8203), .ZN(n8208) );
  NAND2_X1 U10634 ( .A1(n8588), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8207) );
  INV_X1 U10635 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8204) );
  OR2_X1 U10636 ( .A1(n8509), .A2(n8204), .ZN(n8205) );
  INV_X1 U10637 ( .A(n8209), .ZN(n8210) );
  XNOR2_X1 U10638 ( .A(n8211), .B(n8210), .ZN(n9805) );
  NAND2_X1 U10639 ( .A1(n6411), .A2(n9805), .ZN(n8215) );
  OR2_X1 U10640 ( .A1(n8212), .A2(n8416), .ZN(n8213) );
  XNOR2_X1 U10641 ( .A(n8213), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10330) );
  OR2_X1 U10642 ( .A1(n6675), .A2(n10330), .ZN(n8214) );
  OAI211_X1 U10643 ( .C1(n8572), .C2(SI_3_), .A(n8215), .B(n8214), .ZN(n15069)
         );
  NAND2_X1 U10644 ( .A1(n15082), .A2(n15069), .ZN(n8989) );
  OR2_X1 U10645 ( .A1(n15062), .A2(n15059), .ZN(n15063) );
  INV_X1 U10646 ( .A(n15069), .ZN(n10681) );
  NAND2_X1 U10647 ( .A1(n15082), .A2(n10681), .ZN(n8216) );
  AND2_X1 U10648 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8217) );
  NOR2_X1 U10649 ( .A1(n8232), .A2(n8217), .ZN(n15057) );
  INV_X1 U10650 ( .A(n15057), .ZN(n10796) );
  NAND2_X1 U10651 ( .A1(n8547), .A2(n10796), .ZN(n8222) );
  NAND2_X1 U10652 ( .A1(n8588), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U10653 ( .A1(n6419), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8220) );
  INV_X1 U10654 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8218) );
  OR2_X1 U10655 ( .A1(n8509), .A2(n8218), .ZN(n8219) );
  NAND4_X1 U10656 ( .A1(n8222), .A2(n8221), .A3(n8220), .A4(n8219), .ZN(n15060) );
  XNOR2_X1 U10657 ( .A(n6576), .B(n8223), .ZN(n9811) );
  NAND2_X1 U10658 ( .A1(n6411), .A2(n9811), .ZN(n8228) );
  NAND2_X1 U10659 ( .A1(n8212), .A2(n8225), .ZN(n8244) );
  NAND2_X1 U10660 ( .A1(n8244), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8226) );
  XNOR2_X1 U10661 ( .A(n8226), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10498) );
  OR2_X1 U10662 ( .A1(n6413), .A2(n10498), .ZN(n8227) );
  OAI211_X1 U10663 ( .C1(n8572), .C2(SI_4_), .A(n8228), .B(n8227), .ZN(n15039)
         );
  INV_X1 U10664 ( .A(n15039), .ZN(n8229) );
  INV_X1 U10665 ( .A(n15043), .ZN(n15041) );
  AND2_X1 U10666 ( .A1(n15060), .A2(n8229), .ZN(n8230) );
  AOI21_X1 U10667 ( .B1(n15040), .B2(n15041), .A(n8230), .ZN(n15027) );
  NAND2_X1 U10668 ( .A1(n8606), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10669 ( .A1(n8588), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8238) );
  OR2_X1 U10670 ( .A1(n8232), .A2(n8231), .ZN(n8233) );
  NAND2_X1 U10671 ( .A1(n8249), .A2(n8233), .ZN(n15035) );
  NAND2_X1 U10672 ( .A1(n8547), .A2(n15035), .ZN(n8237) );
  INV_X1 U10673 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8235) );
  INV_X1 U10674 ( .A(n8241), .ZN(n8242) );
  XNOR2_X1 U10675 ( .A(n8243), .B(n8242), .ZN(n9809) );
  NAND2_X1 U10676 ( .A1(n8587), .A2(n9809), .ZN(n8247) );
  NAND2_X1 U10677 ( .A1(n8258), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8245) );
  XNOR2_X1 U10678 ( .A(n8245), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10499) );
  OR2_X1 U10679 ( .A1(n6413), .A2(n10499), .ZN(n8246) );
  OAI211_X1 U10680 ( .C1(n8572), .C2(SI_5_), .A(n8247), .B(n8246), .ZN(n15034)
         );
  OR2_X1 U10681 ( .A1(n11052), .A2(n15034), .ZN(n8996) );
  NAND2_X1 U10682 ( .A1(n11052), .A2(n15034), .ZN(n8997) );
  NAND2_X1 U10683 ( .A1(n8996), .A2(n8997), .ZN(n15026) );
  INV_X1 U10684 ( .A(n15034), .ZN(n10900) );
  OR2_X1 U10685 ( .A1(n11052), .A2(n10900), .ZN(n8248) );
  NAND2_X1 U10686 ( .A1(n8588), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8255) );
  NAND2_X1 U10687 ( .A1(n8606), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U10688 ( .A1(n8249), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U10689 ( .A1(n8265), .A2(n8250), .ZN(n10925) );
  NAND2_X1 U10690 ( .A1(n8547), .A2(n10925), .ZN(n8253) );
  INV_X1 U10691 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8251) );
  OR2_X1 U10692 ( .A1(n8509), .A2(n8251), .ZN(n8252) );
  NAND4_X1 U10693 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n8252), .ZN(n11027) );
  XNOR2_X1 U10694 ( .A(n8257), .B(n8256), .ZN(n9816) );
  NAND2_X1 U10695 ( .A1(n8587), .A2(n9816), .ZN(n8262) );
  INV_X1 U10696 ( .A(SI_6_), .ZN(n9818) );
  OR2_X1 U10697 ( .A1(n8572), .A2(n9818), .ZN(n8261) );
  OR2_X1 U10698 ( .A1(n8275), .A2(n8416), .ZN(n8259) );
  XNOR2_X1 U10699 ( .A(n8259), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10520) );
  OR2_X1 U10700 ( .A1(n6413), .A2(n10525), .ZN(n8260) );
  NAND2_X1 U10701 ( .A1(n11027), .A2(n10929), .ZN(n9001) );
  INV_X1 U10702 ( .A(n11048), .ZN(n8263) );
  INV_X1 U10703 ( .A(n10929), .ZN(n11045) );
  NAND2_X1 U10704 ( .A1(n11027), .A2(n11045), .ZN(n8264) );
  NAND2_X1 U10705 ( .A1(n11051), .A2(n8264), .ZN(n11025) );
  NAND2_X1 U10706 ( .A1(n8606), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8271) );
  AND2_X1 U10707 ( .A1(n8265), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8266) );
  OR2_X1 U10708 ( .A1(n8266), .A2(n8281), .ZN(n11034) );
  NAND2_X1 U10709 ( .A1(n8547), .A2(n11034), .ZN(n8270) );
  NAND2_X1 U10710 ( .A1(n8523), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8269) );
  INV_X1 U10711 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8267) );
  OR2_X1 U10712 ( .A1(n8509), .A2(n8267), .ZN(n8268) );
  NAND4_X1 U10713 ( .A1(n8271), .A2(n8270), .A3(n8269), .A4(n8268), .ZN(n12410) );
  XNOR2_X1 U10714 ( .A(n8273), .B(n8272), .ZN(n9823) );
  NAND2_X1 U10715 ( .A1(n8587), .A2(n9823), .ZN(n8278) );
  OR2_X1 U10716 ( .A1(n8291), .A2(n8416), .ZN(n8276) );
  XNOR2_X1 U10717 ( .A(n8276), .B(n8290), .ZN(n10644) );
  INV_X1 U10718 ( .A(n10644), .ZN(n10652) );
  OR2_X1 U10719 ( .A1(n6413), .A2(n10652), .ZN(n8277) );
  OAI211_X1 U10720 ( .C1(n8572), .C2(SI_7_), .A(n8278), .B(n8277), .ZN(n11038)
         );
  OR2_X1 U10721 ( .A1(n12410), .A2(n11038), .ZN(n9008) );
  NAND2_X1 U10722 ( .A1(n12410), .A2(n11038), .ZN(n9007) );
  INV_X1 U10723 ( .A(n11038), .ZN(n8745) );
  NAND2_X1 U10724 ( .A1(n12410), .A2(n8745), .ZN(n8279) );
  NAND2_X1 U10725 ( .A1(n8588), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U10726 ( .A1(n8606), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8286) );
  NOR2_X1 U10727 ( .A1(n8281), .A2(n8280), .ZN(n8282) );
  OR2_X1 U10728 ( .A1(n8300), .A2(n8282), .ZN(n15011) );
  NAND2_X1 U10729 ( .A1(n8547), .A2(n15011), .ZN(n8285) );
  INV_X1 U10730 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8283) );
  OR2_X1 U10731 ( .A1(n8946), .A2(n8283), .ZN(n8284) );
  NAND4_X1 U10732 ( .A1(n8287), .A2(n8286), .A3(n8285), .A4(n8284), .ZN(n12409) );
  XNOR2_X1 U10733 ( .A(n9860), .B(P1_DATAO_REG_8__SCAN_IN), .ZN(n8288) );
  XNOR2_X1 U10734 ( .A(n8289), .B(n8288), .ZN(n9813) );
  NAND2_X1 U10735 ( .A1(n8587), .A2(n9813), .ZN(n8298) );
  NOR2_X1 U10736 ( .A1(n8294), .A2(n8416), .ZN(n8292) );
  MUX2_X1 U10737 ( .A(n8416), .B(n8292), .S(P3_IR_REG_8__SCAN_IN), .Z(n8293)
         );
  INV_X1 U10738 ( .A(n8293), .ZN(n8295) );
  NAND2_X1 U10739 ( .A1(n8294), .A2(n12632), .ZN(n8310) );
  NAND2_X1 U10740 ( .A1(n8295), .A2(n8310), .ZN(n12442) );
  OR2_X1 U10741 ( .A1(n6413), .A2(n12442), .ZN(n8297) );
  INV_X1 U10742 ( .A(SI_8_), .ZN(n9814) );
  OR2_X1 U10743 ( .A1(n8572), .A2(n9814), .ZN(n8296) );
  NAND2_X1 U10744 ( .A1(n12409), .A2(n15010), .ZN(n9014) );
  NAND2_X1 U10745 ( .A1(n9015), .A2(n9014), .ZN(n9011) );
  INV_X1 U10746 ( .A(n15010), .ZN(n8749) );
  OR2_X1 U10747 ( .A1(n8749), .A2(n12409), .ZN(n8299) );
  NAND2_X1 U10748 ( .A1(n8523), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U10749 ( .A1(n8606), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8305) );
  OR2_X1 U10750 ( .A1(n8300), .A2(n14891), .ZN(n8301) );
  NAND2_X1 U10751 ( .A1(n8316), .A2(n8301), .ZN(n11466) );
  NAND2_X1 U10752 ( .A1(n8547), .A2(n11466), .ZN(n8304) );
  INV_X1 U10753 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8302) );
  OR2_X1 U10754 ( .A1(n8509), .A2(n8302), .ZN(n8303) );
  NAND4_X1 U10755 ( .A1(n8306), .A2(n8305), .A3(n8304), .A4(n8303), .ZN(n12408) );
  XNOR2_X1 U10756 ( .A(n9945), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n8307) );
  XNOR2_X1 U10757 ( .A(n8308), .B(n8307), .ZN(n14262) );
  NAND2_X1 U10758 ( .A1(n8587), .A2(n14262), .ZN(n8313) );
  NAND2_X1 U10759 ( .A1(n8310), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8309) );
  MUX2_X1 U10760 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8309), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8311) );
  NAND2_X1 U10761 ( .A1(n8311), .A2(n8343), .ZN(n14896) );
  OR2_X1 U10762 ( .A1(n6413), .A2(n12446), .ZN(n8312) );
  OAI211_X1 U10763 ( .C1(n8572), .C2(SI_9_), .A(n8313), .B(n8312), .ZN(n11463)
         );
  INV_X1 U10764 ( .A(n11463), .ZN(n8315) );
  NAND2_X1 U10765 ( .A1(n12408), .A2(n8315), .ZN(n8314) );
  NAND2_X1 U10766 ( .A1(n8606), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10767 ( .A1(n8316), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8317) );
  AND2_X1 U10768 ( .A1(n8332), .A2(n8317), .ZN(n15009) );
  INV_X1 U10769 ( .A(n15009), .ZN(n8318) );
  NAND2_X1 U10770 ( .A1(n8547), .A2(n8318), .ZN(n8322) );
  NAND2_X1 U10771 ( .A1(n8523), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8321) );
  INV_X1 U10772 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8319) );
  OR2_X1 U10773 ( .A1(n8946), .A2(n8319), .ZN(n8320) );
  NAND4_X1 U10774 ( .A1(n8323), .A2(n8322), .A3(n8321), .A4(n8320), .ZN(n11461) );
  XNOR2_X1 U10775 ( .A(n8325), .B(n8324), .ZN(n14266) );
  NAND2_X1 U10776 ( .A1(n14266), .A2(n8587), .ZN(n8330) );
  NAND2_X1 U10777 ( .A1(n8343), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8327) );
  INV_X1 U10778 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8326) );
  OAI22_X1 U10779 ( .A1(n8572), .A2(SI_10_), .B1(n12451), .B2(n6413), .ZN(
        n8328) );
  INV_X1 U10780 ( .A(n8328), .ZN(n8329) );
  NAND2_X1 U10781 ( .A1(n11461), .A2(n11499), .ZN(n8331) );
  NAND2_X1 U10782 ( .A1(n11508), .A2(n8331), .ZN(n11475) );
  INV_X1 U10783 ( .A(n11475), .ZN(n11473) );
  INV_X1 U10784 ( .A(n11499), .ZN(n15002) );
  NAND2_X1 U10785 ( .A1(n8523), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10786 ( .A1(n8606), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10787 ( .A1(n8332), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U10788 ( .A1(n8358), .A2(n8333), .ZN(n11619) );
  NAND2_X1 U10789 ( .A1(n8547), .A2(n11619), .ZN(n8336) );
  INV_X1 U10790 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8334) );
  OR2_X1 U10791 ( .A1(n8946), .A2(n8334), .ZN(n8335) );
  NAND4_X1 U10792 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(n12407) );
  INV_X1 U10793 ( .A(n12407), .ZN(n11680) );
  NAND2_X1 U10794 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  NAND2_X1 U10795 ( .A1(n8342), .A2(n8341), .ZN(n14269) );
  NAND2_X1 U10796 ( .A1(n14269), .A2(n8587), .ZN(n8348) );
  OAI21_X1 U10797 ( .B1(n8343), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8344) );
  XNOR2_X1 U10798 ( .A(n8344), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12455) );
  OAI22_X1 U10799 ( .A1(n8572), .A2(n8345), .B1(n6413), .B2(n14931), .ZN(n8346) );
  INV_X1 U10800 ( .A(n8346), .ZN(n8347) );
  NAND2_X1 U10801 ( .A1(n11680), .A2(n14413), .ZN(n8349) );
  INV_X1 U10802 ( .A(n14413), .ZN(n8626) );
  NAND2_X1 U10803 ( .A1(n8626), .A2(n12407), .ZN(n8350) );
  XNOR2_X1 U10804 ( .A(n6527), .B(n8352), .ZN(n14272) );
  NAND2_X1 U10805 ( .A1(n14272), .A2(n8587), .ZN(n8357) );
  NAND2_X1 U10806 ( .A1(n8353), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8354) );
  INV_X1 U10807 ( .A(n14949), .ZN(n12433) );
  OAI22_X1 U10808 ( .A1(n8572), .A2(SI_12_), .B1(n12433), .B2(n6413), .ZN(
        n8355) );
  INV_X1 U10809 ( .A(n8355), .ZN(n8356) );
  NAND2_X1 U10810 ( .A1(n8606), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8364) );
  AND2_X1 U10811 ( .A1(n8358), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8359) );
  NOR2_X1 U10812 ( .A1(n8375), .A2(n8359), .ZN(n14406) );
  INV_X1 U10813 ( .A(n14406), .ZN(n11637) );
  NAND2_X1 U10814 ( .A1(n8547), .A2(n11637), .ZN(n8363) );
  NAND2_X1 U10815 ( .A1(n8523), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8362) );
  INV_X1 U10816 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8360) );
  OR2_X1 U10817 ( .A1(n8946), .A2(n8360), .ZN(n8361) );
  NAND4_X1 U10818 ( .A1(n8364), .A2(n8363), .A3(n8362), .A4(n8361), .ZN(n12406) );
  INV_X1 U10819 ( .A(n12406), .ZN(n12352) );
  NOR2_X1 U10820 ( .A1(n11684), .A2(n12352), .ZN(n8365) );
  INV_X1 U10821 ( .A(n11684), .ZN(n14401) );
  XNOR2_X1 U10822 ( .A(n8366), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n14278) );
  NAND2_X1 U10823 ( .A1(n14278), .A2(n8587), .ZN(n8374) );
  NAND2_X1 U10824 ( .A1(n8367), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8368) );
  MUX2_X1 U10825 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8368), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8371) );
  INV_X1 U10826 ( .A(n8369), .ZN(n8370) );
  NAND2_X1 U10827 ( .A1(n8371), .A2(n8370), .ZN(n14967) );
  OAI22_X1 U10828 ( .A1(n8572), .A2(SI_13_), .B1(n12461), .B2(n6413), .ZN(
        n8372) );
  INV_X1 U10829 ( .A(n8372), .ZN(n8373) );
  NAND2_X1 U10830 ( .A1(n8588), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U10831 ( .A1(n8606), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8380) );
  OR2_X1 U10832 ( .A1(n8375), .A2(n12350), .ZN(n8376) );
  NAND2_X1 U10833 ( .A1(n8390), .A2(n8376), .ZN(n12355) );
  NAND2_X1 U10834 ( .A1(n8547), .A2(n12355), .ZN(n8379) );
  INV_X1 U10835 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n8377) );
  OR2_X1 U10836 ( .A1(n8946), .A2(n8377), .ZN(n8378) );
  NAND4_X1 U10837 ( .A1(n8381), .A2(n8380), .A3(n8379), .A4(n8378), .ZN(n12405) );
  NAND2_X1 U10838 ( .A1(n12964), .A2(n12405), .ZN(n9040) );
  INV_X1 U10839 ( .A(n12405), .ZN(n12273) );
  INV_X1 U10840 ( .A(n8382), .ZN(n8383) );
  XNOR2_X1 U10841 ( .A(n8384), .B(n8383), .ZN(n14283) );
  NAND2_X1 U10842 ( .A1(n14283), .A2(n8587), .ZN(n8389) );
  OR2_X1 U10843 ( .A1(n8369), .A2(n8416), .ZN(n8385) );
  XNOR2_X1 U10844 ( .A(n8385), .B(n8400), .ZN(n14986) );
  OAI22_X1 U10845 ( .A1(n8572), .A2(n8386), .B1(n6413), .B2(n14986), .ZN(n8387) );
  INV_X1 U10846 ( .A(n8387), .ZN(n8388) );
  NAND2_X1 U10847 ( .A1(n8389), .A2(n8388), .ZN(n11630) );
  NAND2_X1 U10848 ( .A1(n8523), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10849 ( .A1(n8606), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10850 ( .A1(n8390), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10851 ( .A1(n8407), .A2(n8391), .ZN(n12275) );
  NAND2_X1 U10852 ( .A1(n8547), .A2(n12275), .ZN(n8393) );
  INV_X1 U10853 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12957) );
  OR2_X1 U10854 ( .A1(n8509), .A2(n12957), .ZN(n8392) );
  NAND4_X1 U10855 ( .A1(n8395), .A2(n8394), .A3(n8393), .A4(n8392), .ZN(n12404) );
  OR2_X1 U10856 ( .A1(n11630), .A2(n12819), .ZN(n9045) );
  NAND2_X1 U10857 ( .A1(n11630), .A2(n12819), .ZN(n9044) );
  INV_X1 U10858 ( .A(n11628), .ZN(n11624) );
  NAND2_X1 U10859 ( .A1(n11625), .A2(n11624), .ZN(n11623) );
  NAND2_X1 U10860 ( .A1(n11630), .A2(n12404), .ZN(n8396) );
  NAND2_X1 U10861 ( .A1(n11623), .A2(n8396), .ZN(n12817) );
  INV_X1 U10862 ( .A(n8397), .ZN(n8398) );
  XNOR2_X1 U10863 ( .A(n8399), .B(n8398), .ZN(n14285) );
  NAND2_X1 U10864 ( .A1(n14285), .A2(n8587), .ZN(n8406) );
  NAND2_X1 U10865 ( .A1(n8369), .A2(n8400), .ZN(n8401) );
  NAND2_X1 U10866 ( .A1(n8401), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8402) );
  XNOR2_X1 U10867 ( .A(n8402), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12469) );
  OAI22_X1 U10868 ( .A1(n8572), .A2(n8403), .B1(n6675), .B2(n14331), .ZN(n8404) );
  INV_X1 U10869 ( .A(n8404), .ZN(n8405) );
  NAND2_X1 U10870 ( .A1(n8523), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U10871 ( .A1(n8606), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8410) );
  XNOR2_X1 U10872 ( .A(n8407), .B(P3_REG3_REG_15__SCAN_IN), .ZN(n12824) );
  NAND2_X1 U10873 ( .A1(n8547), .A2(n12824), .ZN(n8409) );
  INV_X1 U10874 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12954) );
  OR2_X1 U10875 ( .A1(n8509), .A2(n12954), .ZN(n8408) );
  NAND4_X1 U10876 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), .ZN(n12403) );
  OR2_X1 U10877 ( .A1(n12384), .A2(n12403), .ZN(n12801) );
  INV_X1 U10878 ( .A(n8412), .ZN(n8413) );
  XNOR2_X1 U10879 ( .A(n8414), .B(n8413), .ZN(n14289) );
  NAND2_X1 U10880 ( .A1(n14289), .A2(n8587), .ZN(n8426) );
  NOR2_X1 U10881 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n8415) );
  NOR2_X1 U10882 ( .A1(n8420), .A2(n8416), .ZN(n8417) );
  MUX2_X1 U10883 ( .A(n8416), .B(n8417), .S(P3_IR_REG_16__SCAN_IN), .Z(n8418)
         );
  INV_X1 U10884 ( .A(n8418), .ZN(n8422) );
  INV_X1 U10885 ( .A(n8447), .ZN(n8421) );
  AND2_X1 U10886 ( .A1(n8422), .A2(n8421), .ZN(n12471) );
  OAI22_X1 U10887 ( .A1(n8572), .A2(n8423), .B1(n6675), .B2(n14349), .ZN(n8424) );
  INV_X1 U10888 ( .A(n8424), .ZN(n8425) );
  NAND2_X1 U10889 ( .A1(n8588), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U10890 ( .A1(n8606), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8431) );
  NOR2_X1 U10891 ( .A1(n8427), .A2(n12326), .ZN(n8428) );
  OR2_X1 U10892 ( .A1(n8454), .A2(n8428), .ZN(n12812) );
  NAND2_X1 U10893 ( .A1(n8547), .A2(n12812), .ZN(n8430) );
  INV_X1 U10894 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12950) );
  OR2_X1 U10895 ( .A1(n8946), .A2(n12950), .ZN(n8429) );
  NAND4_X1 U10896 ( .A1(n8432), .A2(n8431), .A3(n8430), .A4(n8429), .ZN(n12402) );
  NAND2_X1 U10897 ( .A1(n12322), .A2(n12402), .ZN(n8436) );
  INV_X1 U10898 ( .A(n8436), .ZN(n8433) );
  OR2_X1 U10899 ( .A1(n12322), .A2(n12820), .ZN(n9058) );
  NAND2_X1 U10900 ( .A1(n12322), .A2(n12820), .ZN(n9054) );
  AND2_X1 U10901 ( .A1(n12801), .A2(n8435), .ZN(n8434) );
  NAND2_X1 U10902 ( .A1(n12817), .A2(n8434), .ZN(n8440) );
  INV_X1 U10903 ( .A(n8435), .ZN(n8438) );
  NAND2_X1 U10904 ( .A1(n12384), .A2(n12403), .ZN(n12802) );
  AND2_X1 U10905 ( .A1(n12802), .A2(n8436), .ZN(n8437) );
  OR2_X1 U10906 ( .A1(n8438), .A2(n8437), .ZN(n8439) );
  NAND2_X1 U10907 ( .A1(n8440), .A2(n8439), .ZN(n12789) );
  INV_X1 U10908 ( .A(n8441), .ZN(n8442) );
  XNOR2_X1 U10909 ( .A(n8443), .B(n8442), .ZN(n10396) );
  NAND2_X1 U10910 ( .A1(n10396), .A2(n8587), .ZN(n8452) );
  NOR2_X1 U10911 ( .A1(n8447), .A2(n8416), .ZN(n8444) );
  MUX2_X1 U10912 ( .A(n8416), .B(n8444), .S(P3_IR_REG_17__SCAN_IN), .Z(n8445)
         );
  INV_X1 U10913 ( .A(n8445), .ZN(n8448) );
  AND2_X1 U10914 ( .A1(n8448), .A2(n8477), .ZN(n14361) );
  OAI22_X1 U10915 ( .A1(n8572), .A2(n8449), .B1(n6413), .B2(n12474), .ZN(n8450) );
  INV_X1 U10916 ( .A(n8450), .ZN(n8451) );
  NAND2_X1 U10917 ( .A1(n8523), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U10918 ( .A1(n8606), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8458) );
  OR2_X1 U10919 ( .A1(n8454), .A2(n8453), .ZN(n8455) );
  NAND2_X1 U10920 ( .A1(n8468), .A2(n8455), .ZN(n12796) );
  NAND2_X1 U10921 ( .A1(n8547), .A2(n12796), .ZN(n8457) );
  INV_X1 U10922 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12946) );
  OR2_X1 U10923 ( .A1(n8509), .A2(n12946), .ZN(n8456) );
  NAND4_X1 U10924 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n12401) );
  OR2_X1 U10925 ( .A1(n12795), .A2(n12808), .ZN(n8966) );
  NAND2_X1 U10926 ( .A1(n12795), .A2(n12808), .ZN(n8967) );
  NAND2_X1 U10927 ( .A1(n12795), .A2(n12401), .ZN(n8460) );
  INV_X1 U10928 ( .A(n8461), .ZN(n8462) );
  XNOR2_X1 U10929 ( .A(n8463), .B(n8462), .ZN(n10636) );
  NAND2_X1 U10930 ( .A1(n10636), .A2(n8587), .ZN(n8467) );
  NAND2_X1 U10931 ( .A1(n8477), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8464) );
  XNOR2_X1 U10932 ( .A(n8464), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14376) );
  OAI22_X1 U10933 ( .A1(n8572), .A2(n10637), .B1(n6675), .B2(n12477), .ZN(
        n8465) );
  INV_X1 U10934 ( .A(n8465), .ZN(n8466) );
  NAND2_X1 U10935 ( .A1(n8606), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10936 ( .A1(n8468), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U10937 ( .A1(n8482), .A2(n8469), .ZN(n12784) );
  NAND2_X1 U10938 ( .A1(n8547), .A2(n12784), .ZN(n8472) );
  NAND2_X1 U10939 ( .A1(n8523), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8471) );
  INV_X1 U10940 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12942) );
  OR2_X1 U10941 ( .A1(n8946), .A2(n12942), .ZN(n8470) );
  NAND4_X1 U10942 ( .A1(n8473), .A2(n8472), .A3(n8471), .A4(n8470), .ZN(n12766) );
  NAND2_X1 U10943 ( .A1(n12364), .A2(n12792), .ZN(n9063) );
  XNOR2_X1 U10944 ( .A(n8476), .B(n8475), .ZN(n10689) );
  NAND2_X1 U10945 ( .A1(n10689), .A2(n8587), .ZN(n8481) );
  OAI22_X1 U10946 ( .A1(n8572), .A2(SI_19_), .B1(n6403), .B2(n6413), .ZN(n8479) );
  INV_X1 U10947 ( .A(n8479), .ZN(n8480) );
  AND2_X1 U10948 ( .A1(n8482), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8483) );
  OR2_X1 U10949 ( .A1(n8483), .A2(n8495), .ZN(n12773) );
  NAND2_X1 U10950 ( .A1(n12773), .A2(n8547), .ZN(n8486) );
  AOI22_X1 U10951 ( .A1(n8605), .A2(P3_REG0_REG_19__SCAN_IN), .B1(n8606), .B2(
        P3_REG2_REG_19__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U10952 ( .A1(n8523), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8484) );
  NOR2_X1 U10953 ( .A1(n12940), .A2(n12781), .ZN(n9069) );
  INV_X1 U10954 ( .A(n9069), .ZN(n8488) );
  NAND2_X1 U10955 ( .A1(n12940), .A2(n12781), .ZN(n9062) );
  OR2_X1 U10956 ( .A1(n12364), .A2(n12766), .ZN(n12765) );
  AND2_X1 U10957 ( .A1(n12771), .A2(n12765), .ZN(n8487) );
  NAND2_X1 U10958 ( .A1(n12764), .A2(n8487), .ZN(n12763) );
  NAND2_X1 U10959 ( .A1(n12763), .A2(n8488), .ZN(n12752) );
  INV_X1 U10960 ( .A(n8489), .ZN(n8490) );
  XNOR2_X1 U10961 ( .A(n8491), .B(n8490), .ZN(n10768) );
  NAND2_X1 U10962 ( .A1(n10768), .A2(n8587), .ZN(n8493) );
  OR2_X1 U10963 ( .A1(n8572), .A2(n10770), .ZN(n8492) );
  NOR2_X1 U10964 ( .A1(n8495), .A2(n8494), .ZN(n8496) );
  OR2_X1 U10965 ( .A1(n8507), .A2(n8496), .ZN(n12758) );
  NAND2_X1 U10966 ( .A1(n12758), .A2(n8547), .ZN(n8499) );
  AOI22_X1 U10967 ( .A1(n8606), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n8523), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n8498) );
  INV_X1 U10968 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12934) );
  OR2_X1 U10969 ( .A1(n8946), .A2(n12934), .ZN(n8497) );
  NAND2_X1 U10970 ( .A1(n12338), .A2(n12742), .ZN(n9072) );
  NAND2_X1 U10971 ( .A1(n9071), .A2(n9072), .ZN(n12757) );
  NAND2_X1 U10972 ( .A1(n12752), .A2(n12757), .ZN(n8501) );
  NAND2_X1 U10973 ( .A1(n12338), .A2(n12767), .ZN(n8500) );
  NAND2_X1 U10974 ( .A1(n8501), .A2(n8500), .ZN(n12740) );
  XNOR2_X1 U10975 ( .A(n8503), .B(n8502), .ZN(n10905) );
  NAND2_X1 U10976 ( .A1(n10905), .A2(n8587), .ZN(n8505) );
  OR2_X1 U10977 ( .A1(n8572), .A2(n12626), .ZN(n8504) );
  OR2_X1 U10978 ( .A1(n8507), .A2(n8506), .ZN(n8508) );
  NAND2_X1 U10979 ( .A1(n8521), .A2(n8508), .ZN(n12747) );
  NAND2_X1 U10980 ( .A1(n12747), .A2(n8547), .ZN(n8512) );
  AOI22_X1 U10981 ( .A1(n8606), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n8523), .B2(
        P3_REG1_REG_21__SCAN_IN), .ZN(n8511) );
  INV_X1 U10982 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12930) );
  OR2_X1 U10983 ( .A1(n8946), .A2(n12930), .ZN(n8510) );
  INV_X1 U10984 ( .A(n12754), .ZN(n12398) );
  AND2_X1 U10985 ( .A1(n12746), .A2(n12398), .ZN(n8513) );
  OR2_X1 U10986 ( .A1(n12746), .A2(n12398), .ZN(n8514) );
  INV_X1 U10987 ( .A(n8516), .ZN(n8517) );
  XNOR2_X1 U10988 ( .A(n8518), .B(n8517), .ZN(n11006) );
  NAND2_X1 U10989 ( .A1(n11006), .A2(n6411), .ZN(n8520) );
  OR2_X1 U10990 ( .A1(n8572), .A2(n7505), .ZN(n8519) );
  NAND2_X1 U10991 ( .A1(n8521), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U10992 ( .A1(n8535), .A2(n8522), .ZN(n12735) );
  NAND2_X1 U10993 ( .A1(n12735), .A2(n8547), .ZN(n8528) );
  INV_X1 U10994 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12926) );
  NAND2_X1 U10995 ( .A1(n8523), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U10996 ( .A1(n8606), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8524) );
  OAI211_X1 U10997 ( .C1(n12926), .C2(n8946), .A(n8525), .B(n8524), .ZN(n8526)
         );
  INV_X1 U10998 ( .A(n8526), .ZN(n8527) );
  NOR2_X1 U10999 ( .A1(n12734), .A2(n12581), .ZN(n8530) );
  NAND2_X1 U11000 ( .A1(n12734), .A2(n12581), .ZN(n8529) );
  XNOR2_X1 U11001 ( .A(n8532), .B(n8531), .ZN(n11247) );
  NAND2_X1 U11002 ( .A1(n11247), .A2(n6411), .ZN(n8534) );
  INV_X1 U11003 ( .A(SI_23_), .ZN(n11250) );
  OR2_X1 U11004 ( .A1(n8572), .A2(n11250), .ZN(n8533) );
  NAND2_X1 U11005 ( .A1(n8535), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U11006 ( .A1(n8544), .A2(n8536), .ZN(n12587) );
  NAND2_X1 U11007 ( .A1(n12587), .A2(n8547), .ZN(n8541) );
  INV_X1 U11008 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12922) );
  NAND2_X1 U11009 ( .A1(n8606), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U11010 ( .A1(n8523), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8537) );
  OAI211_X1 U11011 ( .C1(n12922), .C2(n8946), .A(n8538), .B(n8537), .ZN(n8539)
         );
  INV_X1 U11012 ( .A(n8539), .ZN(n8540) );
  NAND2_X1 U11013 ( .A1(n12924), .A2(n12564), .ZN(n8962) );
  INV_X1 U11014 ( .A(n12924), .ZN(n12282) );
  NAND2_X1 U11015 ( .A1(n12282), .A2(n12731), .ZN(n8961) );
  NAND2_X1 U11016 ( .A1(n8962), .A2(n8961), .ZN(n9132) );
  INV_X1 U11017 ( .A(n12560), .ZN(n8555) );
  NOR2_X1 U11018 ( .A1(n8572), .A2(n12683), .ZN(n8543) );
  INV_X1 U11019 ( .A(n6392), .ZN(n12849) );
  INV_X1 U11020 ( .A(n8562), .ZN(n8546) );
  NAND2_X1 U11021 ( .A1(n8544), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U11022 ( .A1(n8546), .A2(n8545), .ZN(n12570) );
  NAND2_X1 U11023 ( .A1(n12570), .A2(n8547), .ZN(n8553) );
  INV_X1 U11024 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U11025 ( .A1(n8606), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U11026 ( .A1(n8523), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8548) );
  OAI211_X1 U11027 ( .C1(n8946), .C2(n8550), .A(n8549), .B(n8548), .ZN(n8551)
         );
  INV_X1 U11028 ( .A(n8551), .ZN(n8552) );
  NAND2_X1 U11029 ( .A1(n12849), .A2(n12582), .ZN(n8638) );
  NAND2_X1 U11030 ( .A1(n6392), .A2(n9084), .ZN(n9085) );
  INV_X1 U11031 ( .A(n9085), .ZN(n8554) );
  AOI21_X2 U11032 ( .B1(n8555), .B2(n8638), .A(n8554), .ZN(n12549) );
  INV_X1 U11033 ( .A(n8556), .ZN(n8557) );
  XNOR2_X1 U11034 ( .A(n8558), .B(n8557), .ZN(n12991) );
  NAND2_X1 U11035 ( .A1(n12991), .A2(n6411), .ZN(n8560) );
  OR2_X1 U11036 ( .A1(n8572), .A2(n12993), .ZN(n8559) );
  NOR2_X1 U11037 ( .A1(n8562), .A2(n8561), .ZN(n8563) );
  OR2_X1 U11038 ( .A1(n8575), .A2(n8563), .ZN(n12555) );
  INV_X1 U11039 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U11040 ( .A1(n8523), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U11041 ( .A1(n8606), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8564) );
  OAI211_X1 U11042 ( .C1(n8566), .C2(n8946), .A(n8565), .B(n8564), .ZN(n8567)
         );
  OR2_X1 U11043 ( .A1(n12845), .A2(n12535), .ZN(n8957) );
  NAND2_X1 U11044 ( .A1(n12845), .A2(n12535), .ZN(n8641) );
  NAND2_X1 U11045 ( .A1(n12549), .A2(n12548), .ZN(n12547) );
  INV_X1 U11046 ( .A(n12535), .ZN(n12565) );
  NAND2_X1 U11047 ( .A1(n12845), .A2(n12565), .ZN(n8568) );
  INV_X1 U11048 ( .A(n8569), .ZN(n8570) );
  XNOR2_X1 U11049 ( .A(n8571), .B(n8570), .ZN(n12987) );
  NAND2_X1 U11050 ( .A1(n12987), .A2(n6411), .ZN(n8574) );
  INV_X1 U11051 ( .A(SI_26_), .ZN(n12989) );
  OR2_X1 U11052 ( .A1(n8572), .A2(n12989), .ZN(n8573) );
  INV_X1 U11053 ( .A(n8575), .ZN(n8576) );
  NAND2_X1 U11054 ( .A1(n8576), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U11055 ( .A1(n8578), .A2(n8577), .ZN(n12540) );
  NAND2_X1 U11056 ( .A1(n12540), .A2(n8547), .ZN(n8583) );
  INV_X1 U11057 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12917) );
  NAND2_X1 U11058 ( .A1(n8606), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U11059 ( .A1(n8523), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8579) );
  OAI211_X1 U11060 ( .C1(n12917), .C2(n8946), .A(n8580), .B(n8579), .ZN(n8581)
         );
  INV_X1 U11061 ( .A(n8581), .ZN(n8582) );
  INV_X1 U11062 ( .A(n12550), .ZN(n12318) );
  NAND2_X1 U11063 ( .A1(n12838), .A2(n12318), .ZN(n8584) );
  NAND2_X1 U11064 ( .A1(n12524), .A2(n12536), .ZN(n9092) );
  AND2_X2 U11065 ( .A1(n9094), .A2(n9092), .ZN(n12511) );
  NAND2_X1 U11066 ( .A1(n12519), .A2(n12518), .ZN(n12517) );
  OAI21_X1 U11067 ( .B1(n12524), .B2(n12397), .A(n12517), .ZN(n12501) );
  NAND2_X1 U11068 ( .A1(n12830), .A2(n12265), .ZN(n8642) );
  AND2_X2 U11069 ( .A1(n9100), .A2(n8642), .ZN(n12504) );
  INV_X1 U11070 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U11071 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(
        P2_DATAO_REG_29__SCAN_IN), .B1(n12148), .B2(n11944), .ZN(n8932) );
  INV_X1 U11072 ( .A(SI_29_), .ZN(n12976) );
  NOR2_X1 U11073 ( .A1(n8240), .A2(n12976), .ZN(n8586) );
  INV_X1 U11074 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U11075 ( .A1(n8606), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U11076 ( .A1(n8588), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8589) );
  OAI211_X1 U11077 ( .C1(n8946), .C2(n8684), .A(n8590), .B(n8589), .ZN(n8591)
         );
  INV_X1 U11078 ( .A(n8591), .ZN(n8592) );
  NAND2_X1 U11079 ( .A1(n8949), .A2(n8592), .ZN(n12503) );
  NAND2_X1 U11080 ( .A1(n12494), .A2(n12503), .ZN(n9104) );
  INV_X1 U11081 ( .A(n12494), .ZN(n8593) );
  INV_X1 U11082 ( .A(n12503), .ZN(n12301) );
  NAND2_X1 U11083 ( .A1(n9104), .A2(n8950), .ZN(n9103) );
  INV_X1 U11084 ( .A(n9103), .ZN(n8594) );
  NAND2_X1 U11085 ( .A1(n8646), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U11086 ( .A1(n6403), .A2(n11007), .ZN(n8676) );
  NAND2_X1 U11087 ( .A1(n8596), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8600) );
  XNOR2_X2 U11088 ( .A(n8600), .B(P3_IR_REG_21__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U11089 ( .A1(n8601), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8602) );
  INV_X1 U11090 ( .A(n10771), .ZN(n8724) );
  NAND2_X1 U11091 ( .A1(n9117), .A2(n8724), .ZN(n8603) );
  INV_X1 U11092 ( .A(n10285), .ZN(n10291) );
  NAND2_X1 U11093 ( .A1(n10291), .A2(n12480), .ZN(n10292) );
  NAND2_X1 U11094 ( .A1(n10292), .A2(n6675), .ZN(n8808) );
  NAND2_X2 U11095 ( .A1(n11007), .A2(n9117), .ZN(n9450) );
  INV_X1 U11096 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14412) );
  NAND2_X1 U11097 ( .A1(n8605), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U11098 ( .A1(n8606), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8607) );
  OAI211_X1 U11099 ( .C1(n8609), .C2(n14412), .A(n8608), .B(n8607), .ZN(n8610)
         );
  INV_X1 U11100 ( .A(n8610), .ZN(n8611) );
  INV_X1 U11101 ( .A(P3_B_REG_SCAN_IN), .ZN(n8612) );
  OAI21_X1 U11102 ( .B1(n10285), .B2(n8612), .A(n15081), .ZN(n14393) );
  NOR2_X1 U11103 ( .A1(n10746), .A2(n14393), .ZN(n8613) );
  OAI21_X2 U11104 ( .B1(n8616), .B2(n15052), .A(n8615), .ZN(n12492) );
  NOR2_X1 U11105 ( .A1(n12746), .A2(n12754), .ZN(n8964) );
  NAND2_X1 U11106 ( .A1(n15075), .A2(n15087), .ZN(n8617) );
  NAND2_X1 U11107 ( .A1(n8617), .A2(n8985), .ZN(n15058) );
  NAND2_X1 U11108 ( .A1(n15058), .A2(n15059), .ZN(n8618) );
  NAND2_X1 U11109 ( .A1(n8618), .A2(n8987), .ZN(n15042) );
  NAND2_X1 U11110 ( .A1(n15042), .A2(n15043), .ZN(n8620) );
  NOR2_X1 U11111 ( .A1(n15060), .A2(n15039), .ZN(n8990) );
  INV_X1 U11112 ( .A(n8990), .ZN(n8619) );
  INV_X1 U11113 ( .A(n15026), .ZN(n9123) );
  NAND2_X1 U11114 ( .A1(n15024), .A2(n9123), .ZN(n8621) );
  NAND2_X1 U11115 ( .A1(n11044), .A2(n11048), .ZN(n8622) );
  NAND2_X1 U11116 ( .A1(n8622), .A2(n9002), .ZN(n11022) );
  NAND2_X1 U11117 ( .A1(n11022), .A2(n11026), .ZN(n8623) );
  NAND2_X1 U11118 ( .A1(n15019), .A2(n15018), .ZN(n8624) );
  NAND2_X1 U11119 ( .A1(n8624), .A2(n9015), .ZN(n11315) );
  OR2_X1 U11120 ( .A1(n12408), .A2(n11463), .ZN(n9018) );
  INV_X1 U11121 ( .A(n9018), .ZN(n9023) );
  NAND2_X1 U11122 ( .A1(n12408), .A2(n11463), .ZN(n9022) );
  XNOR2_X1 U11123 ( .A(n14413), .B(n12407), .ZN(n11506) );
  INV_X1 U11124 ( .A(n11508), .ZN(n8628) );
  AND2_X1 U11125 ( .A1(n11680), .A2(n8626), .ZN(n8627) );
  AOI21_X1 U11126 ( .B1(n8625), .B2(n8628), .A(n8627), .ZN(n9030) );
  OR2_X1 U11127 ( .A1(n11684), .A2(n12406), .ZN(n9037) );
  NAND2_X1 U11128 ( .A1(n11684), .A2(n12406), .ZN(n9035) );
  NAND2_X1 U11129 ( .A1(n11676), .A2(n11677), .ZN(n11675) );
  NAND2_X1 U11130 ( .A1(n11675), .A2(n9037), .ZN(n11577) );
  NAND2_X1 U11131 ( .A1(n11579), .A2(n9041), .ZN(n11629) );
  NAND2_X1 U11132 ( .A1(n11629), .A2(n11628), .ZN(n8629) );
  INV_X1 U11133 ( .A(n12403), .ZN(n12807) );
  OR2_X1 U11134 ( .A1(n12384), .A2(n12807), .ZN(n9048) );
  NAND2_X1 U11135 ( .A1(n12384), .A2(n12807), .ZN(n9052) );
  NAND2_X1 U11136 ( .A1(n12794), .A2(n12793), .ZN(n8630) );
  INV_X1 U11137 ( .A(n12772), .ZN(n8632) );
  INV_X1 U11138 ( .A(n12771), .ZN(n8631) );
  INV_X1 U11139 ( .A(n12940), .ZN(n8633) );
  NAND2_X1 U11140 ( .A1(n8633), .A2(n12781), .ZN(n8634) );
  AND2_X1 U11141 ( .A1(n12746), .A2(n12754), .ZN(n8963) );
  INV_X1 U11142 ( .A(n8963), .ZN(n8636) );
  XNOR2_X1 U11143 ( .A(n12734), .B(n12581), .ZN(n12732) );
  AND2_X1 U11144 ( .A1(n12734), .A2(n12743), .ZN(n8637) );
  INV_X1 U11145 ( .A(n12561), .ZN(n12563) );
  NAND2_X1 U11146 ( .A1(n12849), .A2(n9084), .ZN(n8640) );
  INV_X1 U11147 ( .A(n8641), .ZN(n8959) );
  NAND2_X1 U11148 ( .A1(n12380), .A2(n12318), .ZN(n9091) );
  AND2_X2 U11149 ( .A1(n12512), .A2(n9091), .ZN(n12533) );
  NAND3_X1 U11150 ( .A1(n12511), .A2(n12512), .A3(n12530), .ZN(n12513) );
  INV_X1 U11151 ( .A(n8642), .ZN(n9102) );
  AOI21_X2 U11152 ( .B1(n12505), .B2(n9100), .A(n9102), .ZN(n8952) );
  XNOR2_X1 U11153 ( .A(n9103), .B(n8952), .ZN(n12491) );
  NAND2_X1 U11154 ( .A1(n9116), .A2(n8676), .ZN(n9445) );
  INV_X1 U11155 ( .A(n11007), .ZN(n9447) );
  OR2_X1 U11156 ( .A1(n9445), .A2(n9447), .ZN(n9451) );
  INV_X1 U11157 ( .A(n9116), .ZN(n8675) );
  OR2_X1 U11158 ( .A1(n9117), .A2(n8724), .ZN(n9446) );
  XNOR2_X1 U11159 ( .A(n11007), .B(n9446), .ZN(n8644) );
  OR2_X1 U11160 ( .A1(n6403), .A2(n9117), .ZN(n8643) );
  NAND2_X1 U11161 ( .A1(n8644), .A2(n8643), .ZN(n8798) );
  NAND3_X1 U11162 ( .A1(n8675), .A2(n8798), .A3(n15076), .ZN(n8645) );
  OR2_X1 U11163 ( .A1(n15101), .A2(n11007), .ZN(n12839) );
  NOR2_X2 U11164 ( .A1(n12492), .A2(n7422), .ZN(n9458) );
  NAND2_X2 U11165 ( .A1(n6442), .A2(n8650), .ZN(n11567) );
  XNOR2_X1 U11166 ( .A(n11567), .B(P3_B_REG_SCAN_IN), .ZN(n8658) );
  NAND2_X1 U11167 ( .A1(n6442), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8651) );
  MUX2_X1 U11168 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8651), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8653) );
  INV_X1 U11169 ( .A(n8652), .ZN(n8654) );
  INV_X1 U11170 ( .A(n12990), .ZN(n8657) );
  INV_X1 U11171 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8660) );
  NOR2_X1 U11172 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .ZN(
        n8664) );
  NOR4_X1 U11173 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8663) );
  NOR4_X1 U11174 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n8662) );
  NOR4_X1 U11175 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8661) );
  NAND4_X1 U11176 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), .ZN(n8670)
         );
  NOR4_X1 U11177 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8668) );
  NOR4_X1 U11178 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8667) );
  NOR4_X1 U11179 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8666) );
  NOR4_X1 U11180 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8665) );
  NAND4_X1 U11181 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8665), .ZN(n8669)
         );
  NAND2_X1 U11182 ( .A1(n9443), .A2(n9440), .ZN(n8799) );
  INV_X1 U11183 ( .A(n12994), .ZN(n8672) );
  NOR2_X1 U11184 ( .A1(n11567), .A2(n12990), .ZN(n8671) );
  NAND2_X1 U11185 ( .A1(n8672), .A2(n8671), .ZN(n9497) );
  NAND2_X1 U11186 ( .A1(n6560), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8673) );
  INV_X1 U11187 ( .A(n10288), .ZN(n8674) );
  NAND2_X1 U11188 ( .A1(n10286), .A2(n10426), .ZN(n9147) );
  OR3_X1 U11189 ( .A1(n8676), .A2(n9117), .A3(n10771), .ZN(n8802) );
  INV_X1 U11190 ( .A(n8802), .ZN(n8792) );
  NAND2_X1 U11191 ( .A1(n10286), .A2(n8792), .ZN(n8677) );
  AND2_X1 U11192 ( .A1(n9147), .A2(n8677), .ZN(n8678) );
  OR2_X1 U11193 ( .A1(n8799), .A2(n8678), .ZN(n8683) );
  INV_X1 U11194 ( .A(n12968), .ZN(n8680) );
  INV_X1 U11195 ( .A(n12966), .ZN(n8679) );
  AND2_X1 U11196 ( .A1(n8680), .A2(n8679), .ZN(n9442) );
  AND2_X1 U11197 ( .A1(n10286), .A2(n8798), .ZN(n8681) );
  NAND2_X1 U11198 ( .A1(n8811), .A2(n8681), .ZN(n8682) );
  INV_X1 U11199 ( .A(n12965), .ZN(n8686) );
  NOR2_X1 U11200 ( .A1(n15143), .A2(n8684), .ZN(n8685) );
  AOI21_X1 U11201 ( .B1(n8593), .B2(n8686), .A(n8685), .ZN(n8687) );
  MUX2_X1 U11202 ( .A(n11944), .B(n12148), .S(n9812), .Z(n9342) );
  NAND2_X1 U11203 ( .A1(n12147), .A2(n7626), .ZN(n8694) );
  OR2_X1 U11204 ( .A1(n6410), .A2(n11944), .ZN(n8693) );
  INV_X1 U11205 ( .A(n9363), .ZN(n13104) );
  XNOR2_X1 U11206 ( .A(n13437), .B(n13104), .ZN(n9416) );
  NAND3_X1 U11207 ( .A1(n14834), .A2(n14835), .A3(n9632), .ZN(n8699) );
  OR2_X1 U11208 ( .A1(n9631), .A2(n8699), .ZN(n8701) );
  INV_X1 U11209 ( .A(n9630), .ZN(n8700) );
  INV_X1 U11210 ( .A(n9500), .ZN(n8702) );
  NAND2_X1 U11211 ( .A1(n8702), .A2(n9423), .ZN(n10240) );
  NAND2_X1 U11212 ( .A1(n13355), .A2(n10240), .ZN(n8703) );
  INV_X1 U11213 ( .A(n13105), .ZN(n11957) );
  NAND2_X1 U11214 ( .A1(n8925), .A2(n13105), .ZN(n8704) );
  NAND2_X1 U11215 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  XNOR2_X1 U11216 ( .A(n8706), .B(n8695), .ZN(n8707) );
  INV_X1 U11217 ( .A(n13404), .ZN(n13311) );
  INV_X1 U11218 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U11219 ( .A1(n7875), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U11220 ( .A1(n9351), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8708) );
  OAI211_X1 U11221 ( .C1(n7577), .C2(n13434), .A(n8709), .B(n8708), .ZN(n13103) );
  NOR2_X1 U11222 ( .A1(n13564), .A2(n8710), .ZN(n8711) );
  NOR2_X1 U11223 ( .A1(n13408), .A2(n8711), .ZN(n13182) );
  AND2_X1 U11224 ( .A1(n13103), .A2(n13182), .ZN(n8712) );
  AOI21_X1 U11225 ( .B1(n13105), .B2(n13311), .A(n8712), .ZN(n8713) );
  INV_X1 U11226 ( .A(n8714), .ZN(n8715) );
  NAND2_X1 U11227 ( .A1(n13437), .A2(n8715), .ZN(n8716) );
  INV_X2 U11228 ( .A(n13384), .ZN(n13427) );
  AND2_X2 U11229 ( .A1(n13427), .A2(n11405), .ZN(n13422) );
  INV_X1 U11230 ( .A(n11059), .ZN(n9392) );
  NAND2_X1 U11231 ( .A1(n10242), .A2(n9392), .ZN(n9626) );
  INV_X1 U11232 ( .A(n9626), .ZN(n8717) );
  NOR2_X1 U11233 ( .A1(n13412), .A2(n8718), .ZN(n8719) );
  AOI21_X1 U11234 ( .B1(n13384), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8719), .ZN(
        n8720) );
  OAI21_X1 U11235 ( .B1(n9364), .B2(n13376), .A(n8720), .ZN(n8721) );
  NAND2_X1 U11236 ( .A1(n6463), .A2(n8723), .ZN(P2_U3236) );
  NAND3_X1 U11237 ( .A1(n8764), .A2(n6695), .A3(n15083), .ZN(n8728) );
  INV_X1 U11238 ( .A(n12900), .ZN(n8729) );
  AOI21_X1 U11239 ( .B1(n6401), .B2(n8730), .A(n8729), .ZN(n8731) );
  NAND2_X1 U11240 ( .A1(n9649), .A2(n8732), .ZN(n9659) );
  XNOR2_X1 U11241 ( .A(n6402), .B(n6601), .ZN(n8733) );
  XNOR2_X1 U11242 ( .A(n8733), .B(n15061), .ZN(n9660) );
  NAND2_X1 U11243 ( .A1(n9659), .A2(n9660), .ZN(n9658) );
  INV_X1 U11244 ( .A(n15061), .ZN(n9652) );
  NAND2_X1 U11245 ( .A1(n8733), .A2(n9652), .ZN(n8734) );
  INV_X1 U11246 ( .A(n8735), .ZN(n8736) );
  NAND2_X1 U11247 ( .A1(n8736), .A2(n15082), .ZN(n8737) );
  XNOR2_X1 U11248 ( .A(n6401), .B(n15039), .ZN(n8738) );
  XNOR2_X1 U11249 ( .A(n8738), .B(n15060), .ZN(n10793) );
  INV_X1 U11250 ( .A(n8738), .ZN(n8739) );
  INV_X1 U11251 ( .A(n15060), .ZN(n15029) );
  XNOR2_X1 U11252 ( .A(n6401), .B(n10900), .ZN(n8740) );
  XNOR2_X1 U11253 ( .A(n8740), .B(n11052), .ZN(n10899) );
  INV_X1 U11254 ( .A(n11052), .ZN(n15047) );
  AND2_X1 U11255 ( .A1(n8740), .A2(n15047), .ZN(n8741) );
  XNOR2_X1 U11256 ( .A(n6402), .B(n11045), .ZN(n8742) );
  XNOR2_X1 U11257 ( .A(n8742), .B(n11027), .ZN(n10927) );
  NAND2_X1 U11258 ( .A1(n10928), .A2(n10927), .ZN(n10926) );
  INV_X1 U11259 ( .A(n8742), .ZN(n8743) );
  NAND2_X1 U11260 ( .A1(n8743), .A2(n11027), .ZN(n8744) );
  NAND2_X1 U11261 ( .A1(n10926), .A2(n8744), .ZN(n11037) );
  XNOR2_X1 U11262 ( .A(n6402), .B(n8745), .ZN(n8746) );
  XNOR2_X1 U11263 ( .A(n8746), .B(n12410), .ZN(n11036) );
  INV_X1 U11264 ( .A(n8746), .ZN(n8747) );
  NAND2_X1 U11265 ( .A1(n8747), .A2(n12410), .ZN(n8748) );
  NAND2_X1 U11266 ( .A1(n11035), .A2(n8748), .ZN(n11267) );
  XNOR2_X1 U11267 ( .A(n6402), .B(n8749), .ZN(n8750) );
  XNOR2_X1 U11268 ( .A(n8750), .B(n12409), .ZN(n11266) );
  NAND2_X1 U11269 ( .A1(n11267), .A2(n11266), .ZN(n11265) );
  INV_X1 U11270 ( .A(n8750), .ZN(n8751) );
  NAND2_X1 U11271 ( .A1(n8751), .A2(n12409), .ZN(n8752) );
  XNOR2_X1 U11272 ( .A(n6401), .B(n11463), .ZN(n8753) );
  XNOR2_X1 U11273 ( .A(n8753), .B(n12408), .ZN(n11460) );
  OR2_X2 U11274 ( .A1(n11459), .A2(n11460), .ZN(n11457) );
  INV_X1 U11275 ( .A(n8753), .ZN(n8754) );
  INV_X1 U11276 ( .A(n12408), .ZN(n15017) );
  NAND2_X1 U11277 ( .A1(n8754), .A2(n15017), .ZN(n8755) );
  XNOR2_X1 U11278 ( .A(n6402), .B(n11499), .ZN(n8756) );
  XNOR2_X1 U11279 ( .A(n8756), .B(n11461), .ZN(n11495) );
  NAND2_X1 U11280 ( .A1(n8756), .A2(n11461), .ZN(n8757) );
  XNOR2_X1 U11281 ( .A(n6401), .B(n14413), .ZN(n8758) );
  NAND2_X1 U11282 ( .A1(n11614), .A2(n12407), .ZN(n8760) );
  NAND2_X1 U11283 ( .A1(n8759), .A2(n8758), .ZN(n11613) );
  XNOR2_X1 U11284 ( .A(n8764), .B(n11684), .ZN(n11634) );
  NAND2_X1 U11285 ( .A1(n11634), .A2(n12352), .ZN(n8761) );
  INV_X1 U11286 ( .A(n11634), .ZN(n8762) );
  NAND2_X1 U11287 ( .A1(n8762), .A2(n12406), .ZN(n8763) );
  XNOR2_X1 U11288 ( .A(n12964), .B(n8764), .ZN(n8765) );
  NAND2_X1 U11289 ( .A1(n8765), .A2(n12273), .ZN(n12346) );
  INV_X1 U11290 ( .A(n8765), .ZN(n8766) );
  NAND2_X1 U11291 ( .A1(n8766), .A2(n12405), .ZN(n12347) );
  XNOR2_X1 U11292 ( .A(n11630), .B(n6402), .ZN(n8767) );
  XNOR2_X1 U11293 ( .A(n8767), .B(n12404), .ZN(n12270) );
  INV_X1 U11294 ( .A(n8767), .ZN(n8768) );
  NAND2_X1 U11295 ( .A1(n8768), .A2(n12404), .ZN(n8769) );
  NAND2_X1 U11296 ( .A1(n12269), .A2(n8769), .ZN(n12387) );
  XNOR2_X1 U11297 ( .A(n12384), .B(n6402), .ZN(n8770) );
  XNOR2_X1 U11298 ( .A(n8770), .B(n12403), .ZN(n12386) );
  NAND2_X1 U11299 ( .A1(n12387), .A2(n12386), .ZN(n12385) );
  INV_X1 U11300 ( .A(n8770), .ZN(n8771) );
  NAND2_X1 U11301 ( .A1(n8771), .A2(n12403), .ZN(n8772) );
  NAND2_X1 U11302 ( .A1(n12385), .A2(n8772), .ZN(n12325) );
  XNOR2_X1 U11303 ( .A(n12322), .B(n6401), .ZN(n8773) );
  XNOR2_X1 U11304 ( .A(n8773), .B(n12402), .ZN(n12324) );
  INV_X1 U11305 ( .A(n8773), .ZN(n8774) );
  NAND2_X1 U11306 ( .A1(n8774), .A2(n12402), .ZN(n8775) );
  XNOR2_X1 U11307 ( .A(n12795), .B(n6401), .ZN(n8776) );
  XNOR2_X1 U11308 ( .A(n8776), .B(n12808), .ZN(n12332) );
  XNOR2_X1 U11309 ( .A(n12364), .B(n6402), .ZN(n8777) );
  XNOR2_X1 U11310 ( .A(n8777), .B(n12792), .ZN(n12365) );
  OR2_X2 U11311 ( .A1(n12366), .A2(n12365), .ZN(n12367) );
  INV_X1 U11312 ( .A(n8777), .ZN(n8778) );
  NAND2_X1 U11313 ( .A1(n8778), .A2(n12766), .ZN(n8779) );
  XNOR2_X1 U11314 ( .A(n12940), .B(n6401), .ZN(n8780) );
  XNOR2_X1 U11315 ( .A(n8780), .B(n12781), .ZN(n12286) );
  INV_X1 U11316 ( .A(n12781), .ZN(n12400) );
  NAND2_X1 U11317 ( .A1(n8780), .A2(n12400), .ZN(n8781) );
  NAND2_X1 U11318 ( .A1(n12285), .A2(n8781), .ZN(n12341) );
  XNOR2_X1 U11319 ( .A(n12338), .B(n6402), .ZN(n8782) );
  XNOR2_X1 U11320 ( .A(n8782), .B(n12767), .ZN(n12340) );
  NAND2_X1 U11321 ( .A1(n12341), .A2(n12340), .ZN(n12339) );
  INV_X1 U11322 ( .A(n8782), .ZN(n8783) );
  NAND2_X1 U11323 ( .A1(n8783), .A2(n12767), .ZN(n8784) );
  XNOR2_X1 U11324 ( .A(n12746), .B(n6401), .ZN(n8785) );
  XNOR2_X1 U11325 ( .A(n8785), .B(n12754), .ZN(n12308) );
  NAND2_X1 U11326 ( .A1(n8785), .A2(n12754), .ZN(n8786) );
  NAND2_X2 U11327 ( .A1(n12305), .A2(n8786), .ZN(n12249) );
  XNOR2_X1 U11328 ( .A(n12734), .B(n8764), .ZN(n8787) );
  INV_X1 U11329 ( .A(n8787), .ZN(n12250) );
  AND2_X1 U11330 ( .A1(n12249), .A2(n12250), .ZN(n8788) );
  XNOR2_X1 U11331 ( .A(n12924), .B(n6402), .ZN(n12253) );
  XNOR2_X1 U11332 ( .A(n8789), .B(n12253), .ZN(n12278) );
  OAI22_X1 U11333 ( .A1(n12278), .A2(n12564), .B1(n12253), .B2(n8789), .ZN(
        n8791) );
  XNOR2_X1 U11334 ( .A(n6392), .B(n6401), .ZN(n12252) );
  XNOR2_X1 U11335 ( .A(n12252), .B(n9084), .ZN(n8790) );
  XNOR2_X1 U11336 ( .A(n8791), .B(n8790), .ZN(n8796) );
  NAND2_X1 U11337 ( .A1(n8798), .A2(n15076), .ZN(n8794) );
  NAND2_X1 U11338 ( .A1(n8811), .A2(n8792), .ZN(n8793) );
  OAI21_X1 U11339 ( .B1(n8799), .B2(n8794), .A(n8793), .ZN(n8795) );
  NAND2_X1 U11340 ( .A1(n8796), .A2(n14861), .ZN(n8818) );
  NAND2_X1 U11341 ( .A1(n8799), .A2(n15101), .ZN(n8797) );
  NOR2_X1 U11342 ( .A1(n6392), .A2(n12395), .ZN(n8816) );
  NAND2_X1 U11343 ( .A1(n9116), .A2(n9078), .ZN(n10629) );
  AND2_X1 U11344 ( .A1(n9497), .A2(n10629), .ZN(n8801) );
  NAND2_X1 U11345 ( .A1(n8799), .A2(n8798), .ZN(n8800) );
  OAI211_X1 U11346 ( .C1(n8811), .C2(n8802), .A(n8801), .B(n8800), .ZN(n8803)
         );
  NAND2_X1 U11347 ( .A1(n8803), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8806) );
  AND2_X1 U11348 ( .A1(n10288), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9144) );
  OAI21_X1 U11349 ( .B1(n8811), .B2(n9147), .A(n11248), .ZN(n8804) );
  INV_X1 U11350 ( .A(n8804), .ZN(n8805) );
  NOR2_X1 U11351 ( .A1(n9147), .A2(n8808), .ZN(n8807) );
  NAND2_X1 U11352 ( .A1(n8811), .A2(n8807), .ZN(n12390) );
  NOR2_X1 U11353 ( .A1(n12731), .A2(n12390), .ZN(n8813) );
  INV_X1 U11354 ( .A(n8808), .ZN(n8809) );
  NOR2_X1 U11355 ( .A1(n9147), .A2(n8809), .ZN(n8810) );
  NAND2_X1 U11356 ( .A1(n8811), .A2(n8810), .ZN(n12378) );
  INV_X1 U11357 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12656) );
  OAI22_X1 U11358 ( .A1(n12535), .A2(n12378), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12656), .ZN(n8812) );
  AOI211_X1 U11359 ( .C1(n12570), .C2(n12392), .A(n8813), .B(n8812), .ZN(n8814) );
  INV_X1 U11360 ( .A(n8814), .ZN(n8815) );
  NAND2_X1 U11361 ( .A1(n8818), .A2(n8817), .ZN(P3_U3169) );
  INV_X1 U11362 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14797) );
  INV_X1 U11363 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10434) );
  XNOR2_X1 U11364 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n10434), .ZN(n8896) );
  INV_X1 U11365 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8841) );
  INV_X1 U11366 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n8839) );
  INV_X1 U11367 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n13820) );
  INV_X1 U11368 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10039) );
  INV_X1 U11369 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11370 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n12654), .ZN(n8850) );
  NOR2_X1 U11371 ( .A1(n8822), .A2(n10480), .ZN(n8824) );
  NOR2_X1 U11372 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n8856), .ZN(n8823) );
  INV_X1 U11373 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n8825) );
  INV_X1 U11374 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14887) );
  NOR2_X1 U11375 ( .A1(n8827), .A2(n14887), .ZN(n8829) );
  XNOR2_X1 U11376 ( .A(n13800), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n8868) );
  INV_X1 U11377 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n8830) );
  NOR2_X1 U11378 ( .A1(n8831), .A2(n8830), .ZN(n8833) );
  XOR2_X1 U11379 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n8831), .Z(n8871) );
  XNOR2_X1 U11380 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n8835), .ZN(n8873) );
  XNOR2_X1 U11381 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n10039), .ZN(n8844) );
  NOR2_X1 U11382 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n8836), .ZN(n8837) );
  XOR2_X1 U11383 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n8836), .Z(n8880) );
  XNOR2_X1 U11384 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n13820), .ZN(n8884) );
  XNOR2_X1 U11385 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n8839), .ZN(n8888) );
  AND2_X1 U11386 ( .A1(n8841), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n8840) );
  XOR2_X1 U11387 ( .A(n8896), .B(n8895), .Z(n14519) );
  XOR2_X1 U11388 ( .A(n8841), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n8843) );
  XOR2_X1 U11389 ( .A(n8843), .B(n8842), .Z(n14515) );
  INV_X1 U11390 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8887) );
  INV_X1 U11391 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8883) );
  XNOR2_X1 U11392 ( .A(n8845), .B(n8844), .ZN(n8879) );
  NOR2_X1 U11393 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n8858), .ZN(n8860) );
  INV_X1 U11394 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n8855) );
  XNOR2_X1 U11395 ( .A(n8847), .B(n8848), .ZN(n14259) );
  XNOR2_X1 U11396 ( .A(n8850), .B(n8849), .ZN(n8852) );
  NAND2_X1 U11397 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n8852), .ZN(n8853) );
  INV_X1 U11398 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15163) );
  OAI21_X1 U11399 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n12654), .A(n8850), .ZN(
        n8851) );
  INV_X1 U11400 ( .A(n8851), .ZN(n15164) );
  NOR2_X1 U11401 ( .A1(n15163), .A2(n15164), .ZN(n15173) );
  NAND2_X1 U11402 ( .A1(n14259), .A2(n14260), .ZN(n8854) );
  XNOR2_X1 U11403 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n8856), .ZN(n15169) );
  NOR2_X1 U11404 ( .A1(n15168), .A2(n15169), .ZN(n8857) );
  INV_X1 U11405 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15170) );
  NAND2_X1 U11406 ( .A1(n15168), .A2(n15169), .ZN(n15167) );
  OAI21_X1 U11407 ( .B1(n8857), .B2(n15170), .A(n15167), .ZN(n15161) );
  XNOR2_X1 U11408 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n8858), .ZN(n15160) );
  NOR2_X1 U11409 ( .A1(n15161), .A2(n15160), .ZN(n8859) );
  XNOR2_X1 U11410 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n8861), .ZN(n8862) );
  NOR2_X1 U11411 ( .A1(n8863), .A2(n8862), .ZN(n8864) );
  NAND2_X1 U11412 ( .A1(n8867), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8870) );
  INV_X1 U11413 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8866) );
  XNOR2_X1 U11414 ( .A(n8869), .B(n8868), .ZN(n14281) );
  XNOR2_X1 U11415 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8871), .ZN(n15165) );
  XNOR2_X1 U11416 ( .A(n8874), .B(n8873), .ZN(n8876) );
  NAND2_X1 U11417 ( .A1(n8875), .A2(n8876), .ZN(n8878) );
  NAND2_X1 U11418 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14291), .ZN(n8877) );
  INV_X1 U11419 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n8881) );
  XOR2_X1 U11420 ( .A(n8881), .B(n8880), .Z(n14294) );
  NAND2_X1 U11421 ( .A1(n14295), .A2(n14294), .ZN(n8882) );
  XNOR2_X1 U11422 ( .A(n8885), .B(n8884), .ZN(n14510) );
  XNOR2_X1 U11423 ( .A(n8889), .B(n8888), .ZN(n8891) );
  INV_X1 U11424 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14768) );
  INV_X1 U11425 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14545) );
  XOR2_X1 U11426 ( .A(n14545), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n8899) );
  INV_X1 U11427 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n8898) );
  XOR2_X1 U11428 ( .A(n8899), .B(n8903), .Z(n8900) );
  INV_X1 U11429 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n8909) );
  XOR2_X1 U11430 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n8909), .Z(n8905) );
  INV_X1 U11431 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U11432 ( .A1(n8902), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n8904) );
  XOR2_X1 U11433 ( .A(n8905), .B(n8908), .Z(n14527) );
  NAND2_X1 U11434 ( .A1(n14526), .A2(n14527), .ZN(n8906) );
  AOI21_X2 U11435 ( .B1(n14797), .B2(n8906), .A(n14525), .ZN(n14322) );
  OR2_X1 U11436 ( .A1(n8909), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8907) );
  AOI22_X1 U11437 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n8909), .B1(n8908), .B2(
        n8907), .ZN(n8910) );
  INV_X1 U11438 ( .A(n8910), .ZN(n8914) );
  XOR2_X1 U11439 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n8914), .Z(n8915) );
  XNOR2_X1 U11440 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n8915), .ZN(n14321) );
  NAND2_X1 U11441 ( .A1(n14322), .A2(n14321), .ZN(n8911) );
  INV_X1 U11442 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14811) );
  INV_X1 U11443 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n8921) );
  XOR2_X1 U11444 ( .A(n8921), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n8919) );
  XNOR2_X1 U11445 ( .A(n8918), .B(n8919), .ZN(n8916) );
  NAND2_X1 U11446 ( .A1(n8919), .A2(n8918), .ZN(n8920) );
  OAI21_X1 U11447 ( .B1(n8921), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n8920), .ZN(
        n8922) );
  INV_X1 U11448 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n12642) );
  INV_X1 U11449 ( .A(n14834), .ZN(n8923) );
  INV_X2 U11450 ( .A(n14857), .ZN(n8929) );
  NOR2_X1 U11451 ( .A1(n14857), .A2(n8926), .ZN(n8927) );
  OAI21_X1 U11452 ( .B1(n8930), .B2(n8929), .A(n8928), .ZN(P2_U3527) );
  INV_X1 U11453 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12246) );
  INV_X1 U11454 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14232) );
  OAI22_X1 U11455 ( .A1(n14232), .A2(n12246), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U11456 ( .A1(n8939), .A2(n8941), .ZN(n8933) );
  OAI21_X1 U11457 ( .B1(n12246), .B2(P2_DATAO_REG_30__SCAN_IN), .A(n8933), 
        .ZN(n8935) );
  INV_X1 U11458 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14231) );
  INV_X1 U11459 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13553) );
  AOI22_X1 U11460 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n14231), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n13553), .ZN(n8934) );
  XOR2_X1 U11461 ( .A(n8935), .B(n8934), .Z(n12970) );
  NAND2_X1 U11462 ( .A1(n12970), .A2(n8587), .ZN(n8938) );
  INV_X1 U11463 ( .A(n8240), .ZN(n8936) );
  NAND2_X1 U11464 ( .A1(n8936), .A2(SI_31_), .ZN(n8937) );
  INV_X1 U11465 ( .A(n8939), .ZN(n8940) );
  XNOR2_X1 U11466 ( .A(n8941), .B(n8940), .ZN(n12243) );
  NAND2_X1 U11467 ( .A1(n12243), .A2(n6411), .ZN(n8943) );
  INV_X1 U11468 ( .A(SI_30_), .ZN(n12658) );
  OR2_X1 U11469 ( .A1(n8240), .A2(n12658), .ZN(n8942) );
  INV_X1 U11470 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14418) );
  NAND2_X1 U11471 ( .A1(n8523), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8945) );
  NAND2_X1 U11472 ( .A1(n8606), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n8944) );
  OAI211_X1 U11473 ( .C1(n14418), .C2(n8946), .A(n8945), .B(n8944), .ZN(n8947)
         );
  INV_X1 U11474 ( .A(n8947), .ZN(n8948) );
  NOR2_X1 U11475 ( .A1(n6687), .A2(n14394), .ZN(n8955) );
  NAND2_X1 U11476 ( .A1(n14411), .A2(n10746), .ZN(n9107) );
  NAND2_X1 U11477 ( .A1(n9107), .A2(n8950), .ZN(n9109) );
  INV_X1 U11478 ( .A(n9109), .ZN(n8951) );
  INV_X1 U11479 ( .A(n14394), .ZN(n12396) );
  INV_X1 U11480 ( .A(n14411), .ZN(n8953) );
  INV_X1 U11481 ( .A(n9104), .ZN(n9137) );
  INV_X1 U11482 ( .A(n8957), .ZN(n8958) );
  MUX2_X1 U11483 ( .A(n8959), .B(n8958), .S(n9078), .Z(n8960) );
  INV_X1 U11484 ( .A(n8960), .ZN(n9090) );
  MUX2_X1 U11485 ( .A(n8962), .B(n8961), .S(n9450), .Z(n9083) );
  MUX2_X1 U11486 ( .A(n8964), .B(n8963), .S(n9450), .Z(n8965) );
  INV_X1 U11487 ( .A(n8965), .ZN(n9077) );
  XNOR2_X1 U11488 ( .A(n12746), .B(n12754), .ZN(n12745) );
  INV_X1 U11489 ( .A(n12745), .ZN(n9075) );
  MUX2_X1 U11490 ( .A(n12781), .B(n12940), .S(n9450), .Z(n9070) );
  NAND2_X1 U11491 ( .A1(n9057), .A2(n8966), .ZN(n8971) );
  INV_X1 U11492 ( .A(n8967), .ZN(n8968) );
  NAND2_X1 U11493 ( .A1(n9057), .A2(n8968), .ZN(n8969) );
  NAND2_X1 U11494 ( .A1(n8969), .A2(n9063), .ZN(n8970) );
  MUX2_X1 U11495 ( .A(n8971), .B(n8970), .S(n9450), .Z(n9067) );
  MUX2_X1 U11496 ( .A(n8974), .B(n8972), .S(n9450), .Z(n8980) );
  NAND2_X1 U11497 ( .A1(n9120), .A2(n11007), .ZN(n8977) );
  NAND2_X1 U11498 ( .A1(n9120), .A2(n9117), .ZN(n8975) );
  NAND3_X1 U11499 ( .A1(n8975), .A2(n8974), .A3(n9450), .ZN(n8976) );
  OAI21_X1 U11500 ( .B1(n8973), .B2(n8977), .A(n8976), .ZN(n8978) );
  OAI21_X1 U11501 ( .B1(n9117), .B2(n12905), .A(n8978), .ZN(n8979) );
  NAND3_X1 U11502 ( .A1(n8980), .A2(n15087), .A3(n8979), .ZN(n8984) );
  NAND2_X1 U11503 ( .A1(n8989), .A2(n8981), .ZN(n8982) );
  NAND2_X1 U11504 ( .A1(n8982), .A2(n9078), .ZN(n8983) );
  NAND2_X1 U11505 ( .A1(n8984), .A2(n8983), .ZN(n8988) );
  AOI21_X1 U11506 ( .B1(n8987), .B2(n8985), .A(n9078), .ZN(n8986) );
  AOI21_X1 U11507 ( .B1(n8988), .B2(n8987), .A(n8986), .ZN(n8995) );
  OAI21_X1 U11508 ( .B1(n9078), .B2(n8989), .A(n15043), .ZN(n8994) );
  AND2_X1 U11509 ( .A1(n15060), .A2(n15039), .ZN(n8991) );
  MUX2_X1 U11510 ( .A(n8991), .B(n8990), .S(n9450), .Z(n8992) );
  NOR2_X1 U11511 ( .A1(n8992), .A2(n15026), .ZN(n8993) );
  OAI21_X1 U11512 ( .B1(n8995), .B2(n8994), .A(n8993), .ZN(n9006) );
  NAND2_X1 U11513 ( .A1(n9002), .A2(n8996), .ZN(n8999) );
  NAND2_X1 U11514 ( .A1(n9001), .A2(n8997), .ZN(n8998) );
  MUX2_X1 U11515 ( .A(n8999), .B(n8998), .S(n9450), .Z(n9000) );
  INV_X1 U11516 ( .A(n9000), .ZN(n9005) );
  MUX2_X1 U11517 ( .A(n9002), .B(n9001), .S(n9078), .Z(n9003) );
  NAND2_X1 U11518 ( .A1(n9003), .A2(n11026), .ZN(n9004) );
  AOI21_X1 U11519 ( .B1(n9006), .B2(n9005), .A(n9004), .ZN(n9013) );
  INV_X1 U11520 ( .A(n9007), .ZN(n9010) );
  INV_X1 U11521 ( .A(n9008), .ZN(n9009) );
  MUX2_X1 U11522 ( .A(n9010), .B(n9009), .S(n9078), .Z(n9012) );
  OR3_X1 U11523 ( .A1(n9013), .A2(n9012), .A3(n9011), .ZN(n9021) );
  INV_X1 U11524 ( .A(n9014), .ZN(n9017) );
  INV_X1 U11525 ( .A(n9015), .ZN(n9016) );
  MUX2_X1 U11526 ( .A(n9017), .B(n9016), .S(n9450), .Z(n9019) );
  NAND2_X1 U11527 ( .A1(n9018), .A2(n9022), .ZN(n11316) );
  NOR2_X1 U11528 ( .A1(n9019), .A2(n11316), .ZN(n9020) );
  NAND2_X1 U11529 ( .A1(n9021), .A2(n9020), .ZN(n9027) );
  INV_X1 U11530 ( .A(n9022), .ZN(n9024) );
  MUX2_X1 U11531 ( .A(n9024), .B(n9023), .S(n9078), .Z(n9025) );
  NOR2_X1 U11532 ( .A1(n9025), .A2(n11475), .ZN(n9026) );
  NAND2_X1 U11533 ( .A1(n9027), .A2(n9026), .ZN(n9029) );
  NAND3_X1 U11534 ( .A1(n11461), .A2(n9078), .A3(n11499), .ZN(n9028) );
  AOI21_X1 U11535 ( .B1(n9029), .B2(n9028), .A(n11506), .ZN(n9032) );
  AOI21_X1 U11536 ( .B1(n9030), .B2(n9037), .A(n9078), .ZN(n9031) );
  OR2_X1 U11537 ( .A1(n9032), .A2(n9031), .ZN(n9036) );
  NAND2_X1 U11538 ( .A1(n14413), .A2(n12407), .ZN(n9033) );
  AOI21_X1 U11539 ( .B1(n9035), .B2(n9033), .A(n9450), .ZN(n9034) );
  AOI21_X1 U11540 ( .B1(n9036), .B2(n9035), .A(n9034), .ZN(n9039) );
  NOR2_X1 U11541 ( .A1(n9037), .A2(n9450), .ZN(n9038) );
  OAI21_X1 U11542 ( .B1(n9039), .B2(n9038), .A(n11576), .ZN(n9043) );
  MUX2_X1 U11543 ( .A(n9041), .B(n9040), .S(n9450), .Z(n9042) );
  NAND3_X1 U11544 ( .A1(n9043), .A2(n11628), .A3(n9042), .ZN(n9047) );
  MUX2_X1 U11545 ( .A(n9045), .B(n9044), .S(n9450), .Z(n9046) );
  NAND3_X1 U11546 ( .A1(n9047), .A2(n12822), .A3(n9046), .ZN(n9051) );
  NAND2_X1 U11547 ( .A1(n9058), .A2(n9048), .ZN(n9049) );
  NAND2_X1 U11548 ( .A1(n9049), .A2(n9450), .ZN(n9050) );
  NAND2_X1 U11549 ( .A1(n9051), .A2(n9050), .ZN(n9055) );
  AOI21_X1 U11550 ( .B1(n9054), .B2(n9052), .A(n9450), .ZN(n9053) );
  AOI21_X1 U11551 ( .B1(n9055), .B2(n9054), .A(n9053), .ZN(n9056) );
  NAND2_X1 U11552 ( .A1(n9057), .A2(n9056), .ZN(n9061) );
  INV_X1 U11553 ( .A(n9058), .ZN(n9059) );
  NAND2_X1 U11554 ( .A1(n9059), .A2(n9078), .ZN(n9060) );
  AOI21_X1 U11555 ( .B1(n9061), .B2(n9060), .A(n12790), .ZN(n9066) );
  NAND2_X1 U11556 ( .A1(n9070), .A2(n9062), .ZN(n9065) );
  OR2_X1 U11557 ( .A1(n9063), .A2(n9450), .ZN(n9064) );
  OAI211_X1 U11558 ( .C1(n9067), .C2(n9066), .A(n9065), .B(n9064), .ZN(n9068)
         );
  OAI211_X1 U11559 ( .C1(n9070), .C2(n9069), .A(n8635), .B(n9068), .ZN(n9074)
         );
  MUX2_X1 U11560 ( .A(n9072), .B(n9071), .S(n9450), .Z(n9073) );
  NAND3_X1 U11561 ( .A1(n9075), .A2(n9074), .A3(n9073), .ZN(n9076) );
  NAND3_X1 U11562 ( .A1(n12732), .A2(n9077), .A3(n9076), .ZN(n9081) );
  NAND3_X1 U11563 ( .A1(n12734), .A2(n12743), .A3(n9078), .ZN(n9080) );
  OR3_X1 U11564 ( .A1(n12734), .A2(n12743), .A3(n9078), .ZN(n9079) );
  NAND4_X1 U11565 ( .A1(n9081), .A2(n12578), .A3(n9080), .A4(n9079), .ZN(n9082) );
  AND2_X1 U11566 ( .A1(n9083), .A2(n9082), .ZN(n9087) );
  MUX2_X1 U11567 ( .A(n9084), .B(n6392), .S(n9450), .Z(n9086) );
  AOI22_X1 U11568 ( .A1(n12561), .A2(n9087), .B1(n9086), .B2(n9085), .ZN(n9088) );
  NAND2_X1 U11569 ( .A1(n9134), .A2(n9088), .ZN(n9089) );
  NAND3_X1 U11570 ( .A1(n12533), .A2(n9090), .A3(n9089), .ZN(n9099) );
  NAND2_X1 U11571 ( .A1(n9092), .A2(n9091), .ZN(n9093) );
  NAND2_X1 U11572 ( .A1(n9093), .A2(n9094), .ZN(n9098) );
  INV_X1 U11573 ( .A(n9094), .ZN(n9095) );
  AOI21_X1 U11574 ( .B1(n12511), .B2(n9096), .A(n9095), .ZN(n9097) );
  INV_X1 U11575 ( .A(n9100), .ZN(n9101) );
  NAND2_X1 U11576 ( .A1(n9140), .A2(n9104), .ZN(n9105) );
  NAND2_X1 U11577 ( .A1(n9105), .A2(n9450), .ZN(n9106) );
  NAND2_X1 U11578 ( .A1(n9108), .A2(n9107), .ZN(n9112) );
  AOI21_X1 U11579 ( .B1(n9109), .B2(n9140), .A(n9450), .ZN(n9110) );
  NAND2_X1 U11580 ( .A1(n9112), .A2(n9110), .ZN(n9111) );
  NAND2_X1 U11581 ( .A1(n14407), .A2(n14394), .ZN(n9139) );
  OAI211_X1 U11582 ( .C1(n9112), .C2(n9078), .A(n9111), .B(n9139), .ZN(n9114)
         );
  NAND2_X1 U11583 ( .A1(n9114), .A2(n9113), .ZN(n9115) );
  INV_X1 U11584 ( .A(n9119), .ZN(n9142) );
  INV_X1 U11585 ( .A(n12504), .ZN(n9138) );
  INV_X1 U11586 ( .A(n9120), .ZN(n9121) );
  NOR2_X1 U11587 ( .A1(n9122), .A2(n9121), .ZN(n14858) );
  NAND4_X1 U11588 ( .A1(n15087), .A2(n14858), .A3(n9123), .A4(n11026), .ZN(
        n9126) );
  INV_X1 U11589 ( .A(n8973), .ZN(n9124) );
  NAND4_X1 U11590 ( .A1(n9124), .A2(n15018), .A3(n15059), .A4(n11048), .ZN(
        n9125) );
  NOR4_X1 U11591 ( .A1(n9126), .A2(n9125), .A3(n15041), .A4(n11316), .ZN(n9127) );
  AND4_X1 U11592 ( .A1(n9127), .A2(n11473), .A3(n11677), .A4(n8625), .ZN(n9128) );
  NAND4_X1 U11593 ( .A1(n12822), .A2(n11628), .A3(n11576), .A4(n9128), .ZN(
        n9129) );
  NOR3_X1 U11594 ( .A1(n12771), .A2(n12804), .A3(n9129), .ZN(n9130) );
  NAND4_X1 U11595 ( .A1(n12782), .A2(n12793), .A3(n12732), .A4(n9130), .ZN(
        n9131) );
  NOR4_X1 U11596 ( .A1(n12745), .A2(n12757), .A3(n9132), .A4(n9131), .ZN(n9133) );
  NAND4_X1 U11597 ( .A1(n12511), .A2(n9134), .A3(n9133), .A4(n12561), .ZN(
        n9136) );
  INV_X1 U11598 ( .A(n12533), .ZN(n9135) );
  NOR4_X1 U11599 ( .A1(n9138), .A2(n9137), .A3(n9136), .A4(n9135), .ZN(n9141)
         );
  NAND4_X1 U11600 ( .A1(n9142), .A2(n9141), .A3(n9140), .A4(n9139), .ZN(n9143)
         );
  NAND2_X1 U11601 ( .A1(n10291), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12981) );
  NOR3_X1 U11602 ( .A1(n9147), .A2(n12480), .A3(n12981), .ZN(n9149) );
  OAI21_X1 U11603 ( .B1(n11248), .B2(n11007), .A(P3_B_REG_SCAN_IN), .ZN(n9148)
         );
  OR2_X1 U11604 ( .A1(n9149), .A2(n9148), .ZN(n9150) );
  AND2_X1 U11605 ( .A1(n11471), .A2(n9423), .ZN(n9153) );
  INV_X1 U11606 ( .A(n9153), .ZN(n9156) );
  NAND2_X1 U11607 ( .A1(n10245), .A2(n9436), .ZN(n9424) );
  AND2_X1 U11608 ( .A1(n9627), .A2(n9428), .ZN(n9152) );
  NAND2_X1 U11609 ( .A1(n9424), .A2(n9152), .ZN(n9360) );
  NAND3_X1 U11610 ( .A1(n9157), .A2(n9360), .A3(n10014), .ZN(n9155) );
  OAI211_X1 U11611 ( .C1(n9157), .C2(n9156), .A(n9155), .B(n9154), .ZN(n9158)
         );
  NAND2_X1 U11612 ( .A1(n13129), .A2(n9167), .ZN(n9160) );
  NAND2_X1 U11613 ( .A1(n10238), .A2(n9190), .ZN(n9159) );
  AOI22_X1 U11614 ( .A1(n13129), .A2(n9190), .B1(n10238), .B2(n9167), .ZN(
        n9161) );
  AOI21_X1 U11615 ( .B1(n9163), .B2(n9162), .A(n9161), .ZN(n9165) );
  NOR2_X1 U11616 ( .A1(n9163), .A2(n9162), .ZN(n9164) );
  NAND2_X1 U11617 ( .A1(n9166), .A2(n9177), .ZN(n9169) );
  NAND2_X1 U11618 ( .A1(n10266), .A2(n9167), .ZN(n9168) );
  NAND2_X1 U11619 ( .A1(n9169), .A2(n9168), .ZN(n9171) );
  AOI22_X1 U11620 ( .A1(n9166), .A2(n9167), .B1(n9190), .B2(n10266), .ZN(n9170) );
  AOI21_X1 U11621 ( .B1(n9172), .B2(n9171), .A(n9170), .ZN(n9174) );
  NOR2_X1 U11622 ( .A1(n9172), .A2(n9171), .ZN(n9173) );
  NAND2_X1 U11623 ( .A1(n13128), .A2(n9167), .ZN(n9176) );
  NAND2_X1 U11624 ( .A1(n6399), .A2(n9369), .ZN(n9175) );
  NAND2_X1 U11625 ( .A1(n9176), .A2(n9175), .ZN(n9180) );
  AOI22_X1 U11626 ( .A1(n13128), .A2(n9369), .B1(n9167), .B2(n6398), .ZN(n9178) );
  AOI21_X1 U11627 ( .B1(n9181), .B2(n9180), .A(n9178), .ZN(n9179) );
  INV_X1 U11628 ( .A(n9179), .ZN(n9182) );
  AOI22_X1 U11629 ( .A1(n13127), .A2(n9177), .B1(n9167), .B2(n10471), .ZN(
        n9185) );
  NAND2_X1 U11630 ( .A1(n13127), .A2(n9167), .ZN(n9183) );
  OAI21_X1 U11631 ( .B1(n9167), .B2(n10559), .A(n9183), .ZN(n9184) );
  NAND2_X1 U11632 ( .A1(n10623), .A2(n9369), .ZN(n9187) );
  NAND2_X1 U11633 ( .A1(n13126), .A2(n9167), .ZN(n9186) );
  NAND2_X1 U11634 ( .A1(n9187), .A2(n9186), .ZN(n9189) );
  AOI22_X1 U11635 ( .A1(n10623), .A2(n9167), .B1(n13126), .B2(n9369), .ZN(
        n9188) );
  NAND2_X1 U11636 ( .A1(n10698), .A2(n9167), .ZN(n9192) );
  NAND2_X1 U11637 ( .A1(n13125), .A2(n9369), .ZN(n9191) );
  NAND2_X1 U11638 ( .A1(n9197), .A2(n9198), .ZN(n9196) );
  NAND2_X1 U11639 ( .A1(n10698), .A2(n9369), .ZN(n9193) );
  OAI21_X1 U11640 ( .B1(n9194), .B2(n9369), .A(n9193), .ZN(n9195) );
  NAND2_X1 U11641 ( .A1(n9196), .A2(n9195), .ZN(n9202) );
  INV_X1 U11642 ( .A(n9197), .ZN(n9200) );
  INV_X1 U11643 ( .A(n9198), .ZN(n9199) );
  NAND2_X1 U11644 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  NAND2_X1 U11645 ( .A1(n9202), .A2(n9201), .ZN(n9207) );
  NAND2_X1 U11646 ( .A1(n10766), .A2(n9369), .ZN(n9204) );
  NAND2_X1 U11647 ( .A1(n13124), .A2(n9167), .ZN(n9203) );
  NAND2_X1 U11648 ( .A1(n9204), .A2(n9203), .ZN(n9206) );
  AOI22_X1 U11649 ( .A1(n10766), .A2(n9167), .B1(n9369), .B2(n13124), .ZN(
        n9205) );
  NAND2_X1 U11650 ( .A1(n10853), .A2(n9167), .ZN(n9209) );
  NAND2_X1 U11651 ( .A1(n13123), .A2(n9177), .ZN(n9208) );
  NAND2_X1 U11652 ( .A1(n10853), .A2(n9369), .ZN(n9210) );
  NAND2_X1 U11653 ( .A1(n11003), .A2(n9177), .ZN(n9213) );
  NAND2_X1 U11654 ( .A1(n13122), .A2(n9167), .ZN(n9212) );
  NAND2_X1 U11655 ( .A1(n9213), .A2(n9212), .ZN(n9215) );
  AOI22_X1 U11656 ( .A1(n11003), .A2(n9167), .B1(n9369), .B2(n13122), .ZN(
        n9214) );
  AOI21_X1 U11657 ( .B1(n9216), .B2(n9215), .A(n9214), .ZN(n9217) );
  INV_X1 U11658 ( .A(n9217), .ZN(n9218) );
  NAND2_X1 U11659 ( .A1(n10945), .A2(n9167), .ZN(n9220) );
  NAND2_X1 U11660 ( .A1(n13121), .A2(n9369), .ZN(n9219) );
  NAND2_X1 U11661 ( .A1(n9220), .A2(n9219), .ZN(n9221) );
  NAND2_X1 U11662 ( .A1(n9222), .A2(n9221), .ZN(n9225) );
  NAND2_X1 U11663 ( .A1(n10945), .A2(n9177), .ZN(n9223) );
  NAND2_X1 U11664 ( .A1(n9225), .A2(n9224), .ZN(n9226) );
  NAND2_X1 U11665 ( .A1(n7420), .A2(n9226), .ZN(n9230) );
  NAND2_X1 U11666 ( .A1(n11337), .A2(n9369), .ZN(n9228) );
  NAND2_X1 U11667 ( .A1(n13120), .A2(n9167), .ZN(n9227) );
  AOI22_X1 U11668 ( .A1(n11337), .A2(n9167), .B1(n9369), .B2(n13120), .ZN(
        n9229) );
  NAND2_X1 U11669 ( .A1(n11360), .A2(n9167), .ZN(n9232) );
  NAND2_X1 U11670 ( .A1(n13119), .A2(n9369), .ZN(n9231) );
  AOI22_X1 U11671 ( .A1(n11360), .A2(n9369), .B1(n9167), .B2(n13119), .ZN(
        n9233) );
  NAND2_X1 U11672 ( .A1(n11420), .A2(n9369), .ZN(n9235) );
  NAND2_X1 U11673 ( .A1(n13118), .A2(n9167), .ZN(n9234) );
  NAND2_X1 U11674 ( .A1(n9235), .A2(n9234), .ZN(n9236) );
  NAND2_X1 U11675 ( .A1(n11420), .A2(n9167), .ZN(n9238) );
  OAI21_X1 U11676 ( .B1(n9167), .B2(n7760), .A(n9238), .ZN(n9239) );
  NAND2_X1 U11677 ( .A1(n9240), .A2(n9239), .ZN(n9257) );
  AND2_X1 U11678 ( .A1(n13114), .A2(n9167), .ZN(n9241) );
  AOI21_X1 U11679 ( .B1(n13500), .B2(n9369), .A(n9241), .ZN(n9270) );
  NAND2_X1 U11680 ( .A1(n13500), .A2(n9167), .ZN(n9243) );
  NAND2_X1 U11681 ( .A1(n13114), .A2(n9369), .ZN(n9242) );
  NAND2_X1 U11682 ( .A1(n9243), .A2(n9242), .ZN(n9268) );
  NAND2_X1 U11683 ( .A1(n9270), .A2(n9268), .ZN(n9248) );
  AND2_X1 U11684 ( .A1(n13115), .A2(n9167), .ZN(n9244) );
  AOI21_X1 U11685 ( .B1(n13505), .B2(n9177), .A(n9244), .ZN(n9265) );
  NAND2_X1 U11686 ( .A1(n13505), .A2(n9167), .ZN(n9246) );
  NAND2_X1 U11687 ( .A1(n13115), .A2(n9369), .ZN(n9245) );
  NAND2_X1 U11688 ( .A1(n9246), .A2(n9245), .ZN(n9264) );
  NAND2_X1 U11689 ( .A1(n9265), .A2(n9264), .ZN(n9247) );
  NAND2_X1 U11690 ( .A1(n9248), .A2(n9247), .ZN(n9277) );
  AND2_X1 U11691 ( .A1(n13116), .A2(n9167), .ZN(n9249) );
  AOI21_X1 U11692 ( .B1(n11610), .B2(n9369), .A(n9249), .ZN(n9276) );
  NAND2_X1 U11693 ( .A1(n11610), .A2(n9167), .ZN(n9251) );
  NAND2_X1 U11694 ( .A1(n13116), .A2(n9369), .ZN(n9250) );
  NAND2_X1 U11695 ( .A1(n9251), .A2(n9250), .ZN(n9275) );
  AND2_X1 U11696 ( .A1(n9276), .A2(n9275), .ZN(n9252) );
  NOR2_X1 U11697 ( .A1(n9277), .A2(n9252), .ZN(n9259) );
  AND2_X1 U11698 ( .A1(n13117), .A2(n9167), .ZN(n9253) );
  AOI21_X1 U11699 ( .B1(n11490), .B2(n9369), .A(n9253), .ZN(n9261) );
  NAND2_X1 U11700 ( .A1(n11490), .A2(n9167), .ZN(n9255) );
  NAND2_X1 U11701 ( .A1(n13117), .A2(n9369), .ZN(n9254) );
  NAND2_X1 U11702 ( .A1(n9255), .A2(n9254), .ZN(n9260) );
  NAND2_X1 U11703 ( .A1(n9261), .A2(n9260), .ZN(n9256) );
  NAND3_X1 U11704 ( .A1(n9258), .A2(n9257), .A3(n7417), .ZN(n9283) );
  INV_X1 U11705 ( .A(n9259), .ZN(n9281) );
  INV_X1 U11706 ( .A(n9260), .ZN(n9263) );
  INV_X1 U11707 ( .A(n9261), .ZN(n9262) );
  NAND2_X1 U11708 ( .A1(n9263), .A2(n9262), .ZN(n9280) );
  INV_X1 U11709 ( .A(n9264), .ZN(n9267) );
  INV_X1 U11710 ( .A(n9265), .ZN(n9266) );
  NAND2_X1 U11711 ( .A1(n9267), .A2(n9266), .ZN(n9269) );
  INV_X1 U11712 ( .A(n13500), .ZN(n13061) );
  NAND3_X1 U11713 ( .A1(n9269), .A2(n13061), .A3(n13407), .ZN(n9274) );
  INV_X1 U11714 ( .A(n9268), .ZN(n9273) );
  INV_X1 U11715 ( .A(n9269), .ZN(n9272) );
  INV_X1 U11716 ( .A(n9270), .ZN(n9271) );
  AOI22_X1 U11717 ( .A1(n9274), .A2(n9273), .B1(n9272), .B2(n9271), .ZN(n9279)
         );
  OR3_X1 U11718 ( .A1(n9277), .A2(n9276), .A3(n9275), .ZN(n9278) );
  OAI211_X1 U11719 ( .C1(n9281), .C2(n9280), .A(n9279), .B(n9278), .ZN(n9282)
         );
  AND2_X1 U11720 ( .A1(n13113), .A2(n9177), .ZN(n9284) );
  AOI21_X1 U11721 ( .B1(n13375), .B2(n9167), .A(n9284), .ZN(n9288) );
  NAND2_X1 U11722 ( .A1(n13375), .A2(n9369), .ZN(n9286) );
  NAND2_X1 U11723 ( .A1(n13113), .A2(n9167), .ZN(n9285) );
  NAND2_X1 U11724 ( .A1(n9286), .A2(n9285), .ZN(n9287) );
  NAND2_X1 U11725 ( .A1(n13360), .A2(n9369), .ZN(n9290) );
  NAND2_X1 U11726 ( .A1(n13112), .A2(n9167), .ZN(n9289) );
  NAND2_X1 U11727 ( .A1(n9290), .A2(n9289), .ZN(n9292) );
  AOI22_X1 U11728 ( .A1(n13360), .A2(n9167), .B1(n9369), .B2(n13112), .ZN(
        n9291) );
  NAND2_X1 U11729 ( .A1(n13337), .A2(n9167), .ZN(n9295) );
  NAND2_X1 U11730 ( .A1(n13310), .A2(n9369), .ZN(n9294) );
  NAND2_X1 U11731 ( .A1(n9295), .A2(n9294), .ZN(n9297) );
  AOI22_X1 U11732 ( .A1(n13337), .A2(n9369), .B1(n9167), .B2(n13310), .ZN(
        n9296) );
  AOI21_X1 U11733 ( .B1(n9298), .B2(n9297), .A(n9296), .ZN(n9299) );
  NAND2_X1 U11734 ( .A1(n13319), .A2(n9177), .ZN(n9301) );
  NAND2_X1 U11735 ( .A1(n13111), .A2(n9167), .ZN(n9300) );
  AOI22_X1 U11736 ( .A1(n13319), .A2(n9167), .B1(n9369), .B2(n13111), .ZN(
        n9302) );
  NAND2_X1 U11737 ( .A1(n13299), .A2(n9167), .ZN(n9304) );
  NAND2_X1 U11738 ( .A1(n13313), .A2(n9369), .ZN(n9303) );
  NAND2_X1 U11739 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  OR2_X1 U11740 ( .A1(n9306), .A2(n9305), .ZN(n9311) );
  NAND2_X1 U11741 ( .A1(n9306), .A2(n9305), .ZN(n9309) );
  INV_X1 U11742 ( .A(n13313), .ZN(n13039) );
  NAND2_X1 U11743 ( .A1(n13299), .A2(n9177), .ZN(n9307) );
  OAI21_X1 U11744 ( .B1(n13039), .B2(n9369), .A(n9307), .ZN(n9308) );
  NAND2_X1 U11745 ( .A1(n9309), .A2(n9308), .ZN(n9310) );
  NAND2_X1 U11746 ( .A1(n9311), .A2(n9310), .ZN(n9316) );
  NAND2_X1 U11747 ( .A1(n13466), .A2(n9369), .ZN(n9313) );
  NAND2_X1 U11748 ( .A1(n13110), .A2(n9167), .ZN(n9312) );
  NAND2_X1 U11749 ( .A1(n9313), .A2(n9312), .ZN(n9315) );
  AOI22_X1 U11750 ( .A1(n13466), .A2(n9167), .B1(n9369), .B2(n13110), .ZN(
        n9314) );
  NAND2_X1 U11751 ( .A1(n13267), .A2(n9167), .ZN(n9318) );
  NAND2_X1 U11752 ( .A1(n13109), .A2(n9369), .ZN(n9317) );
  NAND2_X1 U11753 ( .A1(n9318), .A2(n9317), .ZN(n9320) );
  AOI22_X1 U11754 ( .A1(n13267), .A2(n9369), .B1(n9167), .B2(n13109), .ZN(
        n9319) );
  AOI21_X1 U11755 ( .B1(n9321), .B2(n9320), .A(n9319), .ZN(n9323) );
  AND2_X1 U11756 ( .A1(n13108), .A2(n9167), .ZN(n9324) );
  NAND2_X1 U11757 ( .A1(n13246), .A2(n9167), .ZN(n9325) );
  OAI21_X1 U11758 ( .B1(n9167), .B2(n13258), .A(n9325), .ZN(n9326) );
  AND2_X1 U11759 ( .A1(n13107), .A2(n9369), .ZN(n9328) );
  AOI21_X1 U11760 ( .B1(n13229), .B2(n9167), .A(n9328), .ZN(n9334) );
  INV_X1 U11761 ( .A(n9334), .ZN(n9329) );
  NAND2_X1 U11762 ( .A1(n9333), .A2(n9329), .ZN(n9332) );
  NAND2_X1 U11763 ( .A1(n13229), .A2(n9177), .ZN(n9330) );
  OAI21_X1 U11764 ( .B1(n13243), .B2(n9369), .A(n9330), .ZN(n9331) );
  NAND2_X1 U11765 ( .A1(n9332), .A2(n9331), .ZN(n9337) );
  INV_X1 U11766 ( .A(n9333), .ZN(n9335) );
  NAND2_X1 U11767 ( .A1(n9335), .A2(n9334), .ZN(n9336) );
  NAND2_X1 U11768 ( .A1(n13444), .A2(n9369), .ZN(n9339) );
  NAND2_X1 U11769 ( .A1(n13106), .A2(n9167), .ZN(n9338) );
  NAND2_X1 U11770 ( .A1(n9339), .A2(n9338), .ZN(n9371) );
  NAND2_X1 U11771 ( .A1(n9341), .A2(n9340), .ZN(n9344) );
  NAND2_X1 U11772 ( .A1(n9342), .A2(n12976), .ZN(n9343) );
  NAND2_X1 U11773 ( .A1(n9344), .A2(n9343), .ZN(n9355) );
  MUX2_X1 U11774 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n9812), .Z(n9345) );
  NAND2_X1 U11775 ( .A1(n9345), .A2(SI_30_), .ZN(n9347) );
  OAI21_X1 U11776 ( .B1(SI_30_), .B2(n9345), .A(n9347), .ZN(n9354) );
  MUX2_X1 U11777 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n9812), .Z(n9348) );
  XNOR2_X1 U11778 ( .A(n9348), .B(SI_31_), .ZN(n9349) );
  OR2_X1 U11779 ( .A1(n6410), .A2(n13553), .ZN(n9350) );
  INV_X1 U11780 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13430) );
  NAND2_X1 U11781 ( .A1(n7875), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U11782 ( .A1(n9351), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9352) );
  OAI211_X1 U11783 ( .C1(n7577), .C2(n13430), .A(n9353), .B(n9352), .ZN(n13183) );
  NAND2_X1 U11784 ( .A1(n9355), .A2(n9354), .ZN(n9356) );
  NAND2_X1 U11785 ( .A1(n12245), .A2(n6389), .ZN(n9359) );
  OR2_X1 U11786 ( .A1(n6410), .A2(n12246), .ZN(n9358) );
  AND2_X1 U11787 ( .A1(n13183), .A2(n9369), .ZN(n9386) );
  OAI21_X1 U11788 ( .B1(n9386), .B2(n9360), .A(n13103), .ZN(n9361) );
  AND2_X1 U11789 ( .A1(n13103), .A2(n9167), .ZN(n9362) );
  OAI22_X1 U11790 ( .A1(n9364), .A2(n9369), .B1(n9167), .B2(n9363), .ZN(n9373)
         );
  NAND2_X1 U11791 ( .A1(n13199), .A2(n9369), .ZN(n9366) );
  NAND2_X1 U11792 ( .A1(n13105), .A2(n9167), .ZN(n9365) );
  NAND2_X1 U11793 ( .A1(n9366), .A2(n9365), .ZN(n9374) );
  AND2_X1 U11794 ( .A1(n13105), .A2(n9369), .ZN(n9367) );
  AOI21_X1 U11795 ( .B1(n13199), .B2(n9167), .A(n9367), .ZN(n9375) );
  NOR2_X1 U11796 ( .A1(n9374), .A2(n9375), .ZN(n9368) );
  AOI22_X1 U11797 ( .A1(n13444), .A2(n9167), .B1(n9369), .B2(n13106), .ZN(
        n9370) );
  INV_X1 U11798 ( .A(n9372), .ZN(n9377) );
  INV_X1 U11799 ( .A(n9373), .ZN(n9376) );
  AOI22_X1 U11800 ( .A1(n9377), .A2(n9376), .B1(n9375), .B2(n9374), .ZN(n9380)
         );
  INV_X1 U11801 ( .A(n13183), .ZN(n9378) );
  OAI21_X1 U11802 ( .B1(n13513), .B2(n9378), .A(n9385), .ZN(n9387) );
  AOI21_X1 U11803 ( .B1(n9380), .B2(n9387), .A(n9379), .ZN(n9384) );
  INV_X1 U11804 ( .A(n9387), .ZN(n9420) );
  XNOR2_X1 U11805 ( .A(n6950), .B(n13103), .ZN(n9418) );
  XNOR2_X1 U11806 ( .A(n13360), .B(n13333), .ZN(n13348) );
  OR2_X1 U11807 ( .A1(n13131), .A2(n10243), .ZN(n9391) );
  NAND2_X1 U11808 ( .A1(n10231), .A2(n9391), .ZN(n10255) );
  NAND4_X1 U11809 ( .A1(n9394), .A2(n9393), .A3(n9392), .A4(n10255), .ZN(n9395) );
  NOR3_X1 U11810 ( .A1(n9395), .A2(n10446), .A3(n10366), .ZN(n9397) );
  OR4_X1 U11811 ( .A1(n11234), .A2(n9400), .A3(n10829), .A4(n9399), .ZN(n9403)
         );
  NAND2_X1 U11812 ( .A1(n9402), .A2(n9401), .ZN(n11412) );
  XNOR2_X1 U11813 ( .A(n11360), .B(n11225), .ZN(n11349) );
  OR4_X1 U11814 ( .A1(n9403), .A2(n11412), .A3(n11349), .A4(n10935), .ZN(n9404) );
  NOR2_X1 U11815 ( .A1(n9405), .A2(n9404), .ZN(n9407) );
  NAND4_X1 U11816 ( .A1(n9408), .A2(n9407), .A3(n9406), .A4(n13401), .ZN(n9409) );
  NOR4_X1 U11817 ( .A1(n13331), .A2(n13348), .A3(n9410), .A4(n9409), .ZN(n9411) );
  NAND4_X1 U11818 ( .A1(n7329), .A2(n9411), .A3(n13293), .A4(n13307), .ZN(
        n9412) );
  NOR2_X1 U11819 ( .A1(n13256), .A2(n9412), .ZN(n9414) );
  AND4_X1 U11820 ( .A1(n9415), .A2(n13227), .A3(n9414), .A4(n9413), .ZN(n9417)
         );
  NAND4_X1 U11821 ( .A1(n9418), .A2(n9417), .A3(n9416), .A4(n13206), .ZN(n9419) );
  NOR2_X1 U11822 ( .A1(n9420), .A2(n9419), .ZN(n9421) );
  XNOR2_X1 U11823 ( .A(n9421), .B(n9423), .ZN(n9422) );
  NAND2_X1 U11824 ( .A1(n9423), .A2(n9428), .ZN(n9425) );
  OAI21_X1 U11825 ( .B1(n9425), .B2(n11059), .A(n9424), .ZN(n9426) );
  NAND2_X1 U11826 ( .A1(n9427), .A2(n9426), .ZN(n9433) );
  NAND2_X1 U11827 ( .A1(n11405), .A2(n9428), .ZN(n9429) );
  OAI211_X1 U11828 ( .C1(n9500), .C2(n9436), .A(n9429), .B(n9627), .ZN(n9430)
         );
  OR2_X1 U11829 ( .A1(n9863), .A2(P2_U3088), .ZN(n11585) );
  INV_X1 U11830 ( .A(n14835), .ZN(n14837) );
  NOR4_X1 U11831 ( .A1(n14837), .A2(n13404), .A3(n13564), .A4(n9627), .ZN(
        n9438) );
  OAI21_X1 U11832 ( .B1(n11585), .B2(n9436), .A(P2_B_REG_SCAN_IN), .ZN(n9437)
         );
  OR2_X1 U11833 ( .A1(n9438), .A2(n9437), .ZN(n9439) );
  NAND2_X1 U11834 ( .A1(n9440), .A2(n10286), .ZN(n9441) );
  OR2_X1 U11835 ( .A1(n9442), .A2(n9441), .ZN(n9444) );
  NAND2_X1 U11836 ( .A1(n9445), .A2(n11024), .ZN(n9449) );
  NAND2_X1 U11837 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  NAND2_X1 U11838 ( .A1(n9449), .A2(n9448), .ZN(n9454) );
  NAND2_X1 U11839 ( .A1(n9451), .A2(n9450), .ZN(n10626) );
  NAND2_X1 U11840 ( .A1(n10626), .A2(n10629), .ZN(n9452) );
  NAND2_X1 U11841 ( .A1(n12966), .A2(n9452), .ZN(n9453) );
  OAI21_X1 U11842 ( .B1(n12966), .B2(n9454), .A(n9453), .ZN(n9455) );
  INV_X1 U11843 ( .A(n9455), .ZN(n9456) );
  NOR2_X1 U11844 ( .A1(n12494), .A2(n12899), .ZN(n9461) );
  INV_X1 U11845 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9459) );
  NOR2_X1 U11846 ( .A1(n9461), .A2(n9460), .ZN(n9462) );
  INV_X1 U11847 ( .A(n9863), .ZN(n9463) );
  NOR2_X1 U11848 ( .A1(n9464), .A2(n9463), .ZN(n9866) );
  INV_X1 U11849 ( .A(n9696), .ZN(n9473) );
  NOR2_X1 U11850 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .ZN(n9469) );
  NAND4_X1 U11851 ( .A1(n9469), .A2(n9468), .A3(n9467), .A4(n9466), .ZN(n9472)
         );
  NAND4_X1 U11852 ( .A1(n9856), .A2(n9470), .A3(n9849), .A4(n9839), .ZN(n9471)
         );
  INV_X1 U11853 ( .A(n9495), .ZN(n9480) );
  NAND2_X1 U11854 ( .A1(n9480), .A2(n9479), .ZN(n9491) );
  NOR2_X1 U11855 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9485) );
  NAND4_X1 U11856 ( .A1(n9485), .A2(n9484), .A3(n9483), .A4(n9482), .ZN(n9487)
         );
  NAND2_X1 U11857 ( .A1(n6445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9489) );
  MUX2_X1 U11858 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9489), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9490) );
  NAND2_X1 U11859 ( .A1(n9490), .A2(n9690), .ZN(n14240) );
  OAI21_X1 U11860 ( .B1(n9491), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9492) );
  MUX2_X1 U11861 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9492), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9493) );
  NAND2_X1 U11862 ( .A1(n9495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9496) );
  OR2_X1 U11863 ( .A1(n10014), .A2(n9498), .ZN(n9499) );
  AND2_X1 U11864 ( .A1(n10235), .A2(n9499), .ZN(n10009) );
  NAND2_X1 U11865 ( .A1(n10014), .A2(n13026), .ZN(n9502) );
  NAND2_X1 U11866 ( .A1(n10009), .A2(n9502), .ZN(n10152) );
  NAND2_X1 U11867 ( .A1(n13129), .A2(n9498), .ZN(n9505) );
  XNOR2_X1 U11868 ( .A(n9505), .B(n9503), .ZN(n10153) );
  NAND2_X1 U11869 ( .A1(n10152), .A2(n10153), .ZN(n10151) );
  INV_X1 U11870 ( .A(n9503), .ZN(n9504) );
  NAND2_X1 U11871 ( .A1(n9505), .A2(n9504), .ZN(n9506) );
  NAND2_X1 U11872 ( .A1(n10151), .A2(n9506), .ZN(n10191) );
  NAND2_X1 U11873 ( .A1(n9166), .A2(n9498), .ZN(n9508) );
  NAND2_X1 U11874 ( .A1(n9508), .A2(n9507), .ZN(n9510) );
  NAND2_X1 U11875 ( .A1(n10191), .A2(n10192), .ZN(n10190) );
  NAND2_X1 U11876 ( .A1(n13128), .A2(n9498), .ZN(n9511) );
  XNOR2_X1 U11877 ( .A(n6398), .B(n9588), .ZN(n9512) );
  XNOR2_X1 U11878 ( .A(n9511), .B(n9512), .ZN(n13004) );
  XNOR2_X1 U11879 ( .A(n10471), .B(n9588), .ZN(n9514) );
  NAND2_X1 U11880 ( .A1(n13127), .A2(n9498), .ZN(n9513) );
  NAND2_X1 U11881 ( .A1(n9514), .A2(n9513), .ZN(n9516) );
  OR2_X1 U11882 ( .A1(n9514), .A2(n9513), .ZN(n9515) );
  NAND2_X1 U11883 ( .A1(n9516), .A2(n9515), .ZN(n10374) );
  XNOR2_X1 U11884 ( .A(n10623), .B(n9588), .ZN(n9517) );
  NAND2_X1 U11885 ( .A1(n13126), .A2(n9498), .ZN(n9518) );
  NAND2_X1 U11886 ( .A1(n9517), .A2(n9518), .ZN(n9522) );
  INV_X1 U11887 ( .A(n9517), .ZN(n9520) );
  INV_X1 U11888 ( .A(n9518), .ZN(n9519) );
  NAND2_X1 U11889 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  AND2_X1 U11890 ( .A1(n9522), .A2(n9521), .ZN(n10572) );
  XNOR2_X1 U11891 ( .A(n10698), .B(n9588), .ZN(n9523) );
  NAND2_X1 U11892 ( .A1(n13125), .A2(n9498), .ZN(n9524) );
  XNOR2_X1 U11893 ( .A(n9523), .B(n9524), .ZN(n10607) );
  INV_X1 U11894 ( .A(n9523), .ZN(n9526) );
  INV_X1 U11895 ( .A(n9524), .ZN(n9525) );
  NAND2_X1 U11896 ( .A1(n9526), .A2(n9525), .ZN(n9527) );
  XNOR2_X1 U11897 ( .A(n10766), .B(n6712), .ZN(n9530) );
  NAND2_X1 U11898 ( .A1(n13124), .A2(n9498), .ZN(n9528) );
  XNOR2_X1 U11899 ( .A(n9530), .B(n9528), .ZN(n10761) );
  INV_X1 U11900 ( .A(n9528), .ZN(n9529) );
  XNOR2_X1 U11901 ( .A(n10853), .B(n9588), .ZN(n9531) );
  NAND2_X1 U11902 ( .A1(n13123), .A2(n9498), .ZN(n9532) );
  NAND2_X1 U11903 ( .A1(n9531), .A2(n9532), .ZN(n9536) );
  INV_X1 U11904 ( .A(n9531), .ZN(n9534) );
  INV_X1 U11905 ( .A(n9532), .ZN(n9533) );
  NAND2_X1 U11906 ( .A1(n9534), .A2(n9533), .ZN(n9535) );
  NAND2_X1 U11907 ( .A1(n9536), .A2(n9535), .ZN(n10749) );
  NAND2_X1 U11908 ( .A1(n10747), .A2(n9536), .ZN(n10908) );
  XNOR2_X1 U11909 ( .A(n11003), .B(n9588), .ZN(n9537) );
  NAND2_X1 U11910 ( .A1(n13122), .A2(n9498), .ZN(n9538) );
  NAND2_X1 U11911 ( .A1(n9537), .A2(n9538), .ZN(n9542) );
  INV_X1 U11912 ( .A(n9537), .ZN(n9540) );
  INV_X1 U11913 ( .A(n9538), .ZN(n9539) );
  NAND2_X1 U11914 ( .A1(n9540), .A2(n9539), .ZN(n9541) );
  AND2_X1 U11915 ( .A1(n9542), .A2(n9541), .ZN(n10909) );
  NAND2_X1 U11916 ( .A1(n10908), .A2(n10909), .ZN(n10907) );
  NAND2_X1 U11917 ( .A1(n10907), .A2(n9542), .ZN(n10919) );
  INV_X1 U11918 ( .A(n10919), .ZN(n9548) );
  XNOR2_X1 U11919 ( .A(n10945), .B(n9588), .ZN(n9543) );
  NAND2_X1 U11920 ( .A1(n13121), .A2(n9498), .ZN(n9544) );
  XNOR2_X1 U11921 ( .A(n9543), .B(n9544), .ZN(n10918) );
  INV_X1 U11922 ( .A(n10918), .ZN(n9547) );
  INV_X1 U11923 ( .A(n9543), .ZN(n9546) );
  INV_X1 U11924 ( .A(n9544), .ZN(n9545) );
  XNOR2_X1 U11925 ( .A(n11337), .B(n9588), .ZN(n9549) );
  NAND2_X1 U11926 ( .A1(n13120), .A2(n9498), .ZN(n9550) );
  NAND2_X1 U11927 ( .A1(n9549), .A2(n9550), .ZN(n9554) );
  INV_X1 U11928 ( .A(n9549), .ZN(n9552) );
  INV_X1 U11929 ( .A(n9550), .ZN(n9551) );
  NAND2_X1 U11930 ( .A1(n9552), .A2(n9551), .ZN(n9553) );
  AND2_X1 U11931 ( .A1(n9554), .A2(n9553), .ZN(n11222) );
  NAND2_X1 U11932 ( .A1(n11223), .A2(n11222), .ZN(n11221) );
  XNOR2_X1 U11933 ( .A(n11360), .B(n9588), .ZN(n9555) );
  NAND2_X1 U11934 ( .A1(n13119), .A2(n9498), .ZN(n9556) );
  NAND2_X1 U11935 ( .A1(n9555), .A2(n9556), .ZN(n9560) );
  INV_X1 U11936 ( .A(n9555), .ZN(n9558) );
  INV_X1 U11937 ( .A(n9556), .ZN(n9557) );
  NAND2_X1 U11938 ( .A1(n9558), .A2(n9557), .ZN(n9559) );
  AND2_X1 U11939 ( .A1(n9560), .A2(n9559), .ZN(n11342) );
  XNOR2_X1 U11940 ( .A(n11420), .B(n9588), .ZN(n9561) );
  NAND2_X1 U11941 ( .A1(n13118), .A2(n9498), .ZN(n9562) );
  XNOR2_X1 U11942 ( .A(n9561), .B(n9562), .ZN(n11363) );
  INV_X1 U11943 ( .A(n9561), .ZN(n9564) );
  INV_X1 U11944 ( .A(n9562), .ZN(n9563) );
  XNOR2_X1 U11945 ( .A(n11490), .B(n9588), .ZN(n9565) );
  NAND2_X1 U11946 ( .A1(n13117), .A2(n9498), .ZN(n9566) );
  NAND2_X1 U11947 ( .A1(n9565), .A2(n9566), .ZN(n9570) );
  INV_X1 U11948 ( .A(n9565), .ZN(n9568) );
  INV_X1 U11949 ( .A(n9566), .ZN(n9567) );
  NAND2_X1 U11950 ( .A1(n9568), .A2(n9567), .ZN(n9569) );
  AND2_X1 U11951 ( .A1(n9570), .A2(n9569), .ZN(n11559) );
  XNOR2_X1 U11952 ( .A(n11610), .B(n6712), .ZN(n9572) );
  AND2_X1 U11953 ( .A1(n13116), .A2(n13394), .ZN(n11602) );
  INV_X1 U11954 ( .A(n9571), .ZN(n9573) );
  XNOR2_X1 U11955 ( .A(n13505), .B(n9588), .ZN(n9575) );
  NAND2_X1 U11956 ( .A1(n13115), .A2(n9498), .ZN(n9576) );
  NAND2_X1 U11957 ( .A1(n9575), .A2(n9576), .ZN(n9581) );
  INV_X1 U11958 ( .A(n9575), .ZN(n9578) );
  INV_X1 U11959 ( .A(n9576), .ZN(n9577) );
  NAND2_X1 U11960 ( .A1(n9578), .A2(n9577), .ZN(n9579) );
  NAND2_X1 U11961 ( .A1(n9581), .A2(n9579), .ZN(n13047) );
  INV_X1 U11962 ( .A(n13047), .ZN(n9580) );
  NAND2_X1 U11963 ( .A1(n13044), .A2(n9581), .ZN(n13053) );
  XNOR2_X1 U11964 ( .A(n13500), .B(n9588), .ZN(n9582) );
  NAND2_X1 U11965 ( .A1(n13114), .A2(n9498), .ZN(n9583) );
  NAND2_X1 U11966 ( .A1(n9582), .A2(n9583), .ZN(n9587) );
  INV_X1 U11967 ( .A(n9582), .ZN(n9585) );
  INV_X1 U11968 ( .A(n9583), .ZN(n9584) );
  NAND2_X1 U11969 ( .A1(n9585), .A2(n9584), .ZN(n9586) );
  AND2_X1 U11970 ( .A1(n9587), .A2(n9586), .ZN(n13054) );
  NAND2_X1 U11971 ( .A1(n13052), .A2(n9587), .ZN(n13082) );
  XNOR2_X1 U11972 ( .A(n13375), .B(n9588), .ZN(n9589) );
  NAND2_X1 U11973 ( .A1(n13113), .A2(n9498), .ZN(n9590) );
  XNOR2_X1 U11974 ( .A(n9589), .B(n9590), .ZN(n13081) );
  INV_X1 U11975 ( .A(n9589), .ZN(n9592) );
  INV_X1 U11976 ( .A(n9590), .ZN(n9591) );
  NAND2_X1 U11977 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  OAI21_X2 U11978 ( .B1(n13082), .B2(n13081), .A(n9593), .ZN(n13017) );
  XNOR2_X1 U11979 ( .A(n13360), .B(n6712), .ZN(n9597) );
  INV_X1 U11980 ( .A(n9597), .ZN(n9595) );
  AND2_X1 U11981 ( .A1(n13112), .A2(n13394), .ZN(n9596) );
  INV_X1 U11982 ( .A(n9596), .ZN(n9594) );
  NAND2_X1 U11983 ( .A1(n9595), .A2(n9594), .ZN(n13013) );
  AND2_X1 U11984 ( .A1(n9597), .A2(n9596), .ZN(n13014) );
  XNOR2_X1 U11985 ( .A(n13337), .B(n6712), .ZN(n9598) );
  NAND2_X1 U11986 ( .A1(n13310), .A2(n9498), .ZN(n9599) );
  XNOR2_X1 U11987 ( .A(n9598), .B(n9599), .ZN(n13063) );
  INV_X1 U11988 ( .A(n9598), .ZN(n9600) );
  NAND2_X1 U11989 ( .A1(n9600), .A2(n9599), .ZN(n9601) );
  XNOR2_X1 U11990 ( .A(n13319), .B(n6712), .ZN(n9602) );
  AND2_X1 U11991 ( .A1(n13111), .A2(n13394), .ZN(n9603) );
  NAND2_X1 U11992 ( .A1(n9602), .A2(n9603), .ZN(n9607) );
  INV_X1 U11993 ( .A(n9602), .ZN(n9605) );
  INV_X1 U11994 ( .A(n9603), .ZN(n9604) );
  NAND2_X1 U11995 ( .A1(n9605), .A2(n9604), .ZN(n9606) );
  NAND2_X1 U11996 ( .A1(n9607), .A2(n9606), .ZN(n13035) );
  INV_X1 U11997 ( .A(n9611), .ZN(n9609) );
  XNOR2_X1 U11998 ( .A(n13299), .B(n6712), .ZN(n9610) );
  NAND2_X1 U11999 ( .A1(n9609), .A2(n9608), .ZN(n13071) );
  AND2_X1 U12000 ( .A1(n13313), .A2(n13394), .ZN(n13073) );
  NAND2_X1 U12001 ( .A1(n13071), .A2(n13073), .ZN(n9612) );
  NAND2_X1 U12002 ( .A1(n9611), .A2(n9610), .ZN(n13070) );
  XNOR2_X1 U12003 ( .A(n13466), .B(n6712), .ZN(n9613) );
  NOR2_X1 U12004 ( .A1(n7922), .A2(n13420), .ZN(n12998) );
  XNOR2_X1 U12005 ( .A(n13267), .B(n6712), .ZN(n9615) );
  AND2_X1 U12006 ( .A1(n13109), .A2(n13394), .ZN(n9614) );
  NAND2_X1 U12007 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  OAI21_X1 U12008 ( .B1(n9615), .B2(n9614), .A(n9616), .ZN(n9642) );
  INV_X1 U12009 ( .A(n9616), .ZN(n9617) );
  NOR2_X1 U12010 ( .A1(n9640), .A2(n9617), .ZN(n9625) );
  XNOR2_X1 U12011 ( .A(n13246), .B(n6712), .ZN(n9619) );
  AND2_X1 U12012 ( .A1(n13108), .A2(n13394), .ZN(n9618) );
  NAND2_X1 U12013 ( .A1(n9619), .A2(n9618), .ZN(n11947) );
  OAI21_X1 U12014 ( .B1(n9619), .B2(n9618), .A(n11947), .ZN(n9624) );
  OR2_X1 U12015 ( .A1(n14834), .A2(n14837), .ZN(n9620) );
  OR2_X1 U12016 ( .A1(n9631), .A2(n9620), .ZN(n9628) );
  INV_X1 U12017 ( .A(n9628), .ZN(n9623) );
  INV_X1 U12018 ( .A(n9864), .ZN(n9621) );
  AND2_X1 U12019 ( .A1(n14849), .A2(n9621), .ZN(n9622) );
  AOI211_X1 U12020 ( .C1(n9625), .C2(n9624), .A(n13088), .B(n11949), .ZN(n9639) );
  OAI21_X2 U12021 ( .B1(n9628), .B2(n9626), .A(n13412), .ZN(n13086) );
  NOR2_X1 U12022 ( .A1(n13526), .A2(n13102), .ZN(n9638) );
  NOR2_X2 U12023 ( .A1(n9628), .A2(n9627), .ZN(n13056) );
  NAND2_X1 U12024 ( .A1(n13056), .A2(n13311), .ZN(n13095) );
  INV_X1 U12025 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9629) );
  OAI22_X1 U12026 ( .A1(n13095), .A2(n13242), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9629), .ZN(n9637) );
  INV_X1 U12027 ( .A(n13408), .ZN(n13312) );
  NAND2_X1 U12028 ( .A1(n13056), .A2(n13312), .ZN(n13097) );
  OAI21_X1 U12029 ( .B1(n9631), .B2(n14834), .A(n9630), .ZN(n9635) );
  AND2_X1 U12030 ( .A1(n9633), .A2(n9632), .ZN(n9634) );
  NAND2_X1 U12031 ( .A1(n9635), .A2(n9634), .ZN(n10006) );
  OAI22_X1 U12032 ( .A1(n13097), .A2(n13243), .B1(n13096), .B2(n13247), .ZN(
        n9636) );
  OR4_X1 U12033 ( .A1(n9639), .A2(n9638), .A3(n9637), .A4(n9636), .ZN(P2_U3197) );
  AOI211_X1 U12034 ( .C1(n9642), .C2(n9641), .A(n13088), .B(n9640), .ZN(n9647)
         );
  NOR2_X1 U12035 ( .A1(n13461), .A2(n13102), .ZN(n9646) );
  OAI22_X1 U12036 ( .A1(n13095), .A2(n7922), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9643), .ZN(n9645) );
  OAI22_X1 U12037 ( .A1(n13097), .A2(n13258), .B1(n13096), .B2(n13264), .ZN(
        n9644) );
  OR4_X1 U12038 ( .A1(n9647), .A2(n9646), .A3(n9645), .A4(n9644), .ZN(P2_U3201) );
  NAND3_X1 U12039 ( .A1(n6402), .A2(n12905), .A3(n8973), .ZN(n9648) );
  AND2_X1 U12040 ( .A1(n9650), .A2(n14861), .ZN(n9657) );
  NOR2_X1 U12041 ( .A1(n12392), .A2(P3_U3151), .ZN(n14864) );
  INV_X1 U12042 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n9651) );
  NOR2_X1 U12043 ( .A1(n14864), .A2(n9651), .ZN(n9656) );
  NOR2_X1 U12044 ( .A1(n12395), .A2(n12908), .ZN(n9655) );
  OAI22_X1 U12045 ( .A1(n9653), .A2(n12390), .B1(n12378), .B2(n9652), .ZN(
        n9654) );
  OR4_X1 U12046 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(P3_U3162) );
  OAI21_X1 U12047 ( .B1(n9660), .B2(n9659), .A(n9658), .ZN(n9661) );
  AND2_X1 U12048 ( .A1(n9661), .A2(n14861), .ZN(n9666) );
  INV_X1 U12049 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n9662) );
  NOR2_X1 U12050 ( .A1(n14864), .A2(n9662), .ZN(n9665) );
  NOR2_X1 U12051 ( .A1(n12395), .A2(n15077), .ZN(n9664) );
  INV_X1 U12052 ( .A(n15082), .ZN(n15045) );
  OAI22_X1 U12053 ( .A1(n6694), .A2(n12390), .B1(n12378), .B2(n15045), .ZN(
        n9663) );
  OR4_X1 U12054 ( .A1(n9666), .A2(n9665), .A3(n9664), .A4(n9663), .ZN(P3_U3177) );
  AOI21_X1 U12055 ( .B1(n9702), .B2(n9704), .A(n9668), .ZN(n9671) );
  INV_X1 U12056 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9668) );
  AOI21_X2 U12057 ( .B1(n9671), .B2(P1_IR_REG_20__SCAN_IN), .A(n9670), .ZN(
        n9777) );
  AND2_X4 U12058 ( .A1(n9701), .A2(n9673), .ZN(n11929) );
  NAND2_X1 U12059 ( .A1(n6441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9674) );
  NAND2_X1 U12060 ( .A1(n12154), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9687) );
  OR2_X1 U12061 ( .A1(n9744), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9686) );
  NAND2_X4 U12062 ( .A1(n14233), .A2(n9682), .ZN(n12167) );
  INV_X1 U12063 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10021) );
  OR2_X1 U12064 ( .A1(n12167), .A2(n10021), .ZN(n9685) );
  INV_X1 U12065 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10048) );
  OR2_X1 U12066 ( .A1(n9745), .A2(n10048), .ZN(n9684) );
  INV_X1 U12067 ( .A(n13731), .ZN(n12006) );
  NAND2_X1 U12068 ( .A1(n9690), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9691) );
  NAND2_X1 U12069 ( .A1(n9694), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9695) );
  MUX2_X1 U12070 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9695), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9698) );
  NAND2_X1 U12071 ( .A1(n9698), .A2(n9697), .ZN(n13771) );
  NAND2_X1 U12072 ( .A1(n9826), .A2(n11085), .ZN(n9700) );
  OR2_X1 U12073 ( .A1(n12160), .A2(n9848), .ZN(n9699) );
  OAI211_X1 U12074 ( .C1(n11835), .C2(n13771), .A(n9700), .B(n9699), .ZN(
        n10885) );
  OAI22_X1 U12075 ( .A1(n9756), .A2(n12006), .B1(n14623), .B2(n9728), .ZN(
        n10773) );
  INV_X1 U12076 ( .A(n9702), .ZN(n9703) );
  NAND2_X1 U12077 ( .A1(n9703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9705) );
  XNOR2_X1 U12078 ( .A(n9706), .B(n11652), .ZN(n10772) );
  XOR2_X1 U12079 ( .A(n10773), .B(n10772), .Z(n9780) );
  INV_X1 U12080 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13735) );
  OR2_X1 U12081 ( .A1(n9721), .A2(n13735), .ZN(n9710) );
  INV_X1 U12082 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10044) );
  OR2_X1 U12083 ( .A1(n9745), .A2(n10044), .ZN(n9709) );
  INV_X1 U12084 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9707) );
  OR2_X1 U12085 ( .A1(n9845), .A2(n11849), .ZN(n9714) );
  INV_X1 U12086 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U12087 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9712) );
  XNOR2_X1 U12088 ( .A(n9713), .B(n9712), .ZN(n13738) );
  NOR2_X1 U12089 ( .A1(n9728), .A2(n6591), .ZN(n9715) );
  AOI21_X1 U12090 ( .B1(n11928), .B2(n13734), .A(n9715), .ZN(n9719) );
  INV_X1 U12091 ( .A(n9719), .ZN(n9716) );
  NAND2_X1 U12092 ( .A1(n9717), .A2(n9716), .ZN(n9720) );
  NAND2_X1 U12093 ( .A1(n9719), .A2(n9718), .ZN(n9743) );
  INV_X1 U12094 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10863) );
  INV_X1 U12095 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9722) );
  OR2_X1 U12096 ( .A1(n12167), .A2(n9722), .ZN(n9726) );
  INV_X4 U12097 ( .A(n9745), .ZN(n12164) );
  NAND2_X1 U12098 ( .A1(n12164), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9725) );
  INV_X1 U12099 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9723) );
  OR2_X1 U12100 ( .A1(n11178), .A2(n9723), .ZN(n9724) );
  INV_X1 U12101 ( .A(n11139), .ZN(n10358) );
  NAND2_X1 U12102 ( .A1(n9828), .A2(SI_0_), .ZN(n9730) );
  NAND2_X1 U12103 ( .A1(n9730), .A2(n9729), .ZN(n9732) );
  NAND2_X1 U12104 ( .A1(n9732), .A2(n9731), .ZN(n14252) );
  MUX2_X1 U12105 ( .A(n6927), .B(n14252), .S(n11835), .Z(n11138) );
  INV_X1 U12106 ( .A(n11138), .ZN(n10411) );
  INV_X1 U12107 ( .A(n9701), .ZN(n9734) );
  AOI22_X1 U12108 ( .A1(n11746), .A2(n10411), .B1(n9734), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9733) );
  NAND2_X1 U12109 ( .A1(n11746), .A2(n11139), .ZN(n9736) );
  NAND2_X1 U12110 ( .A1(n9734), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9735) );
  OAI211_X1 U12111 ( .C1(n9737), .C2(n11138), .A(n9736), .B(n9735), .ZN(n10268) );
  INV_X1 U12112 ( .A(n10268), .ZN(n9739) );
  NAND2_X1 U12113 ( .A1(n9739), .A2(n12232), .ZN(n9740) );
  INV_X1 U12114 ( .A(n10357), .ZN(n9741) );
  NAND2_X1 U12115 ( .A1(n9742), .A2(n9741), .ZN(n10355) );
  NAND2_X1 U12116 ( .A1(n10355), .A2(n9743), .ZN(n10390) );
  NAND2_X1 U12117 ( .A1(n11548), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9750) );
  INV_X1 U12118 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13751) );
  OR2_X1 U12119 ( .A1(n9744), .A2(n13751), .ZN(n9749) );
  INV_X1 U12120 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10043) );
  OR2_X1 U12121 ( .A1(n11923), .A2(n10043), .ZN(n9748) );
  INV_X1 U12122 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9746) );
  OR2_X1 U12123 ( .A1(n11178), .A2(n9746), .ZN(n9747) );
  INV_X1 U12124 ( .A(n13733), .ZN(n10882) );
  OR2_X1 U12125 ( .A1(n9751), .A2(n9668), .ZN(n9752) );
  XNOR2_X1 U12126 ( .A(n9752), .B(n12625), .ZN(n13759) );
  OR2_X1 U12127 ( .A1(n11835), .A2(n13759), .ZN(n9754) );
  INV_X1 U12128 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9830) );
  OR2_X1 U12129 ( .A1(n12160), .A2(n9830), .ZN(n9753) );
  INV_X1 U12130 ( .A(n14589), .ZN(n14616) );
  OAI22_X1 U12131 ( .A1(n10882), .A2(n9728), .B1(n9737), .B2(n14616), .ZN(
        n9755) );
  XNOR2_X1 U12132 ( .A(n9755), .B(n11652), .ZN(n9757) );
  OAI22_X1 U12133 ( .A1(n9756), .A2(n10882), .B1(n14616), .B2(n9728), .ZN(
        n9758) );
  XNOR2_X1 U12134 ( .A(n9757), .B(n9758), .ZN(n10391) );
  NAND2_X1 U12135 ( .A1(n10390), .A2(n10391), .ZN(n10389) );
  INV_X1 U12136 ( .A(n9757), .ZN(n9759) );
  NOR2_X1 U12137 ( .A1(n9765), .A2(n9761), .ZN(n9762) );
  MUX2_X1 U12138 ( .A(n9762), .B(n9761), .S(n9760), .Z(n9763) );
  INV_X1 U12139 ( .A(n9763), .ZN(n9764) );
  NAND2_X1 U12140 ( .A1(n9764), .A2(n9775), .ZN(n10405) );
  INV_X1 U12141 ( .A(n9765), .ZN(n14242) );
  NAND2_X1 U12142 ( .A1(n14242), .A2(n14240), .ZN(n10082) );
  NOR4_X1 U12143 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n9774) );
  NOR4_X1 U12144 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9773) );
  OR4_X1 U12145 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9771) );
  NOR4_X1 U12146 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9769) );
  NOR4_X1 U12147 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9768) );
  NOR4_X1 U12148 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9767) );
  NOR4_X1 U12149 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9766) );
  NAND4_X1 U12150 ( .A1(n9769), .A2(n9768), .A3(n9767), .A4(n9766), .ZN(n9770)
         );
  NOR4_X1 U12151 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9771), .A4(n9770), .ZN(n9772) );
  NAND3_X1 U12152 ( .A1(n9774), .A2(n9773), .A3(n9772), .ZN(n10402) );
  INV_X1 U12153 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n12670) );
  NOR2_X1 U12154 ( .A1(n10402), .A2(n12670), .ZN(n9776) );
  OAI21_X1 U12155 ( .B1(n10405), .B2(n9776), .A(n10404), .ZN(n10415) );
  OR2_X1 U12156 ( .A1(n10858), .A2(n10415), .ZN(n9796) );
  NOR2_X1 U12157 ( .A1(n9796), .A2(n9946), .ZN(n9785) );
  INV_X1 U12158 ( .A(n9785), .ZN(n9778) );
  INV_X1 U12159 ( .A(n11982), .ZN(n10409) );
  INV_X1 U12160 ( .A(n11979), .ZN(n9793) );
  NAND2_X1 U12161 ( .A1(n11977), .A2(n12226), .ZN(n9781) );
  AOI211_X1 U12162 ( .C1(n9780), .C2(n9779), .A(n13705), .B(n10775), .ZN(n9801) );
  NAND2_X1 U12163 ( .A1(n9796), .A2(n10399), .ZN(n10270) );
  AOI21_X1 U12164 ( .B1(n9781), .B2(n9793), .A(n9937), .ZN(n9782) );
  NAND2_X1 U12165 ( .A1(n9701), .A2(n9782), .ZN(n9797) );
  INV_X1 U12166 ( .A(n9797), .ZN(n9783) );
  NAND2_X1 U12167 ( .A1(n10270), .A2(n9783), .ZN(n9784) );
  MUX2_X1 U12168 ( .A(n13714), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n9800) );
  NOR2_X1 U12169 ( .A1(n11977), .A2(n11966), .ZN(n14557) );
  NAND2_X1 U12170 ( .A1(n9785), .A2(n14557), .ZN(n9786) );
  NAND2_X1 U12171 ( .A1(n12154), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9790) );
  INV_X1 U12172 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10024) );
  OR2_X1 U12173 ( .A1(n12167), .A2(n10024), .ZN(n9789) );
  NAND2_X1 U12174 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10781) );
  OAI21_X1 U12175 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n10781), .ZN(n11127) );
  OR2_X1 U12176 ( .A1(n9744), .A2(n11127), .ZN(n9788) );
  INV_X2 U12177 ( .A(n12164), .ZN(n11923) );
  INV_X1 U12178 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11129) );
  INV_X1 U12179 ( .A(n13691), .ZN(n14098) );
  OR2_X1 U12180 ( .A1(n12011), .A2(n14098), .ZN(n9795) );
  NAND2_X1 U12181 ( .A1(n13733), .A2(n14100), .ZN(n9794) );
  AND2_X1 U12182 ( .A1(n9795), .A2(n9794), .ZN(n14621) );
  INV_X1 U12183 ( .A(n9796), .ZN(n9798) );
  OR2_X1 U12184 ( .A1(n9797), .A2(P1_U3086), .ZN(n12222) );
  INV_X1 U12185 ( .A(n12222), .ZN(n10859) );
  OAI22_X1 U12186 ( .A1(n13718), .A2(n14623), .B1(n14621), .B2(n13712), .ZN(
        n9799) );
  OR3_X1 U12187 ( .A1(n9801), .A2(n9800), .A3(n9799), .ZN(P1_U3218) );
  OAI21_X1 U12188 ( .B1(n9803), .B2(P3_STATE_REG_SCAN_IN), .A(n9802), .ZN(
        P3_U3295) );
  INV_X1 U12189 ( .A(SI_3_), .ZN(n9804) );
  NAND2_X1 U12190 ( .A1(n11832), .A2(P3_U3151), .ZN(n12992) );
  OAI222_X1 U12191 ( .A1(n7120), .A2(P3_U3151), .B1(n14277), .B2(n9805), .C1(
        n9804), .C2(n12992), .ZN(P3_U3292) );
  INV_X1 U12192 ( .A(SI_2_), .ZN(n9806) );
  OAI222_X1 U12193 ( .A1(n10329), .A2(P3_U3151), .B1(n14277), .B2(n9807), .C1(
        n9806), .C2(n12992), .ZN(P3_U3293) );
  INV_X1 U12194 ( .A(SI_5_), .ZN(n9808) );
  OAI222_X1 U12195 ( .A1(n6844), .A2(P3_U3151), .B1(n14277), .B2(n9809), .C1(
        n9808), .C2(n12992), .ZN(P3_U3290) );
  INV_X1 U12196 ( .A(n10498), .ZN(n10492) );
  INV_X1 U12197 ( .A(SI_4_), .ZN(n9810) );
  OAI222_X1 U12198 ( .A1(n10492), .A2(P3_U3151), .B1(n14277), .B2(n9811), .C1(
        n9810), .C2(n12992), .ZN(P3_U3291) );
  NAND2_X1 U12199 ( .A1(n9828), .A2(P2_U3088), .ZN(n13561) );
  INV_X1 U12200 ( .A(n13561), .ZN(n11583) );
  INV_X1 U12201 ( .A(n11583), .ZN(n13573) );
  NOR2_X1 U12202 ( .A1(n9812), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13557) );
  INV_X2 U12203 ( .A(n13557), .ZN(n13575) );
  OAI222_X1 U12204 ( .A1(n13573), .A2(n12631), .B1(n13575), .B2(n9845), .C1(
        n9929), .C2(P2_U3088), .ZN(P2_U3326) );
  INV_X1 U12205 ( .A(n9813), .ZN(n9815) );
  OAI222_X1 U12206 ( .A1(n14277), .A2(n9815), .B1(n12992), .B2(n9814), .C1(
        n12442), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U12207 ( .A(n12992), .ZN(n14287) );
  INV_X1 U12208 ( .A(n9816), .ZN(n9817) );
  OAI222_X1 U12209 ( .A1(P3_U3151), .A2(n10525), .B1(n14275), .B2(n9818), .C1(
        n14277), .C2(n9817), .ZN(P3_U3289) );
  INV_X1 U12210 ( .A(n9819), .ZN(n9820) );
  INV_X1 U12211 ( .A(SI_7_), .ZN(n9822) );
  OAI222_X1 U12212 ( .A1(n10644), .A2(P3_U3151), .B1(n14277), .B2(n9823), .C1(
        n9822), .C2(n14275), .ZN(P3_U3288) );
  INV_X1 U12213 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9824) );
  INV_X1 U12214 ( .A(n10776), .ZN(n9837) );
  INV_X1 U12215 ( .A(n9897), .ZN(n10080) );
  OAI222_X1 U12216 ( .A1(n13561), .A2(n9824), .B1(n13575), .B2(n9837), .C1(
        n10080), .C2(P2_U3088), .ZN(P2_U3323) );
  OAI222_X1 U12217 ( .A1(n13561), .A2(n9825), .B1(n13575), .B2(n9829), .C1(
        n13136), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U12218 ( .A(n9826), .ZN(n9847) );
  OAI222_X1 U12219 ( .A1(n13561), .A2(n9827), .B1(n13575), .B2(n9847), .C1(
        n13154), .C2(P2_U3088), .ZN(P2_U3324) );
  AND2_X1 U12220 ( .A1(n9812), .A2(P1_U3086), .ZN(n14225) );
  INV_X2 U12221 ( .A(n14225), .ZN(n14244) );
  OAI222_X1 U12222 ( .A1(n14245), .A2(n9830), .B1(n14244), .B2(n9829), .C1(
        P1_U3086), .C2(n13759), .ZN(P1_U3353) );
  INV_X1 U12223 ( .A(n10803), .ZN(n9833) );
  INV_X1 U12224 ( .A(n9915), .ZN(n9907) );
  OAI222_X1 U12225 ( .A1(n13561), .A2(n9831), .B1(n13575), .B2(n9833), .C1(
        n9907), .C2(P2_U3088), .ZN(P2_U3322) );
  NOR2_X1 U12226 ( .A1(n9697), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9840) );
  OR2_X1 U12227 ( .A1(n9840), .A2(n9668), .ZN(n9832) );
  XNOR2_X1 U12228 ( .A(n9832), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10804) );
  INV_X1 U12229 ( .A(n10804), .ZN(n10149) );
  OAI222_X1 U12230 ( .A1(n14245), .A2(n9834), .B1(n14244), .B2(n9833), .C1(
        P1_U3086), .C2(n10149), .ZN(P1_U3350) );
  INV_X1 U12231 ( .A(n14245), .ZN(n11586) );
  NAND2_X1 U12232 ( .A1(n9697), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9835) );
  XNOR2_X1 U12233 ( .A(n9835), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13790) );
  AOI22_X1 U12234 ( .A1(n11586), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n13790), 
        .B2(P1_STATE_REG_SCAN_IN), .ZN(n9836) );
  OAI21_X1 U12235 ( .B1(n9837), .B2(n14244), .A(n9836), .ZN(P1_U3351) );
  INV_X1 U12236 ( .A(n10951), .ZN(n9843) );
  INV_X1 U12237 ( .A(n9960), .ZN(n9924) );
  OAI222_X1 U12238 ( .A1(n13561), .A2(n9838), .B1(n13575), .B2(n9843), .C1(
        n9924), .C2(P2_U3088), .ZN(P2_U3321) );
  AND2_X1 U12239 ( .A1(n9840), .A2(n9839), .ZN(n9850) );
  OR2_X1 U12240 ( .A1(n9850), .A2(n9668), .ZN(n9841) );
  XNOR2_X1 U12241 ( .A(n9841), .B(P1_IR_REG_6__SCAN_IN), .ZN(n13807) );
  INV_X1 U12242 ( .A(n13807), .ZN(n9842) );
  OAI222_X1 U12243 ( .A1(n14245), .A2(n9844), .B1(n14244), .B2(n9843), .C1(
        P1_U3086), .C2(n9842), .ZN(P1_U3349) );
  OAI222_X1 U12244 ( .A1(n14245), .A2(n9846), .B1(n14244), .B2(n9845), .C1(
        P1_U3086), .C2(n13738), .ZN(P1_U3354) );
  OAI222_X1 U12245 ( .A1(n14245), .A2(n9848), .B1(n14244), .B2(n9847), .C1(
        P1_U3086), .C2(n13771), .ZN(P1_U3352) );
  INV_X1 U12246 ( .A(n10962), .ZN(n9854) );
  NAND2_X1 U12247 ( .A1(n9850), .A2(n9849), .ZN(n9855) );
  NAND2_X1 U12248 ( .A1(n9855), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9851) );
  XNOR2_X1 U12249 ( .A(n9851), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10963) );
  INV_X1 U12250 ( .A(n10963), .ZN(n10182) );
  OAI222_X1 U12251 ( .A1(n14245), .A2(n9852), .B1(n14244), .B2(n9854), .C1(
        P1_U3086), .C2(n10182), .ZN(P1_U3348) );
  INV_X1 U12252 ( .A(n13171), .ZN(n9853) );
  OAI222_X1 U12253 ( .A1(n13573), .A2(n6669), .B1(n13575), .B2(n9854), .C1(
        n9853), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U12254 ( .A(n11081), .ZN(n9861) );
  NAND2_X1 U12255 ( .A1(n9858), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9857) );
  MUX2_X1 U12256 ( .A(n9857), .B(P1_IR_REG_31__SCAN_IN), .S(n9856), .Z(n9859)
         );
  NAND2_X1 U12257 ( .A1(n9859), .A2(n9940), .ZN(n10203) );
  OAI222_X1 U12258 ( .A1(n14245), .A2(n9860), .B1(n14244), .B2(n9861), .C1(
        P1_U3086), .C2(n10203), .ZN(P1_U3347) );
  INV_X1 U12259 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9862) );
  INV_X1 U12260 ( .A(n9981), .ZN(n9972) );
  OAI222_X1 U12261 ( .A1(n13573), .A2(n9862), .B1(n13575), .B2(n9861), .C1(
        n9972), .C2(P2_U3088), .ZN(P2_U3319) );
  NAND2_X1 U12262 ( .A1(n9864), .A2(n9863), .ZN(n9865) );
  AND2_X1 U12263 ( .A1(n7589), .A2(n9865), .ZN(n9867) );
  AND2_X1 U12264 ( .A1(n9869), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9868) );
  OR2_X1 U12265 ( .A1(n9869), .A2(P2_U3088), .ZN(n13558) );
  INV_X1 U12266 ( .A(n13558), .ZN(n9870) );
  NAND2_X1 U12267 ( .A1(n9900), .A2(n13564), .ZN(n14822) );
  INV_X1 U12268 ( .A(n14822), .ZN(n14779) );
  MUX2_X1 U12269 ( .A(n9871), .B(P2_REG1_REG_1__SCAN_IN), .S(n9929), .Z(n9926)
         );
  AND2_X1 U12270 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9872) );
  NAND2_X1 U12271 ( .A1(n9926), .A2(n9872), .ZN(n13133) );
  OR2_X1 U12272 ( .A1(n9929), .A2(n9871), .ZN(n13132) );
  NAND2_X1 U12273 ( .A1(n13133), .A2(n13132), .ZN(n9875) );
  INV_X1 U12274 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9873) );
  MUX2_X1 U12275 ( .A(n9873), .B(P2_REG1_REG_2__SCAN_IN), .S(n13136), .Z(n9874) );
  NAND2_X1 U12276 ( .A1(n9875), .A2(n9874), .ZN(n13150) );
  INV_X1 U12277 ( .A(n13136), .ZN(n13141) );
  NAND2_X1 U12278 ( .A1(n13141), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U12279 ( .A1(n13150), .A2(n13149), .ZN(n9878) );
  INV_X1 U12280 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9876) );
  MUX2_X1 U12281 ( .A(n9876), .B(P2_REG1_REG_3__SCAN_IN), .S(n13154), .Z(n9877) );
  NAND2_X1 U12282 ( .A1(n9878), .A2(n9877), .ZN(n13153) );
  INV_X1 U12283 ( .A(n13154), .ZN(n13148) );
  NAND2_X1 U12284 ( .A1(n13148), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9879) );
  NAND2_X1 U12285 ( .A1(n13153), .A2(n9879), .ZN(n10074) );
  MUX2_X1 U12286 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9880), .S(n9897), .Z(n10073) );
  NAND2_X1 U12287 ( .A1(n10074), .A2(n10073), .ZN(n10072) );
  NAND2_X1 U12288 ( .A1(n9897), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U12289 ( .A1(n10072), .A2(n9885), .ZN(n9883) );
  MUX2_X1 U12290 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9881), .S(n9915), .Z(n9882)
         );
  NAND2_X1 U12291 ( .A1(n9883), .A2(n9882), .ZN(n9913) );
  MUX2_X1 U12292 ( .A(n9881), .B(P2_REG1_REG_5__SCAN_IN), .S(n9915), .Z(n9884)
         );
  NAND3_X1 U12293 ( .A1(n10072), .A2(n9885), .A3(n9884), .ZN(n9886) );
  NAND3_X1 U12294 ( .A1(n14779), .A2(n9913), .A3(n9886), .ZN(n9906) );
  NOR2_X1 U12295 ( .A1(n9887), .A2(P2_U3088), .ZN(n14773) );
  NAND2_X1 U12296 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10577) );
  MUX2_X1 U12297 ( .A(n9888), .B(P2_REG2_REG_2__SCAN_IN), .S(n13136), .Z(n9893) );
  INV_X1 U12298 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9889) );
  MUX2_X1 U12299 ( .A(n9889), .B(P2_REG2_REG_1__SCAN_IN), .S(n9929), .Z(n9891)
         );
  AND2_X1 U12300 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9890) );
  NAND2_X1 U12301 ( .A1(n9891), .A2(n9890), .ZN(n13138) );
  OR2_X1 U12302 ( .A1(n9929), .A2(n9889), .ZN(n13137) );
  NAND2_X1 U12303 ( .A1(n13138), .A2(n13137), .ZN(n9892) );
  NAND2_X1 U12304 ( .A1(n9893), .A2(n9892), .ZN(n13156) );
  NAND2_X1 U12305 ( .A1(n13141), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U12306 ( .A1(n13156), .A2(n13155), .ZN(n9895) );
  MUX2_X1 U12307 ( .A(n10462), .B(P2_REG2_REG_3__SCAN_IN), .S(n13154), .Z(
        n9894) );
  NAND2_X1 U12308 ( .A1(n9895), .A2(n9894), .ZN(n13159) );
  NAND2_X1 U12309 ( .A1(n13148), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U12310 ( .A1(n13159), .A2(n9896), .ZN(n10071) );
  MUX2_X1 U12311 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10451), .S(n9897), .Z(
        n10070) );
  NAND2_X1 U12312 ( .A1(n10071), .A2(n10070), .ZN(n10069) );
  NAND2_X1 U12313 ( .A1(n9897), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U12314 ( .A1(n10069), .A2(n9898), .ZN(n9902) );
  MUX2_X1 U12315 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10599), .S(n9915), .Z(n9901) );
  INV_X1 U12316 ( .A(n13564), .ZN(n9899) );
  AND2_X1 U12317 ( .A1(n9900), .A2(n9899), .ZN(n14776) );
  NAND2_X1 U12318 ( .A1(n9902), .A2(n9901), .ZN(n9917) );
  OAI211_X1 U12319 ( .C1(n9902), .C2(n9901), .A(n14776), .B(n9917), .ZN(n9903)
         );
  NAND2_X1 U12320 ( .A1(n10577), .A2(n9903), .ZN(n9904) );
  AOI21_X1 U12321 ( .B1(n14773), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9904), .ZN(
        n9905) );
  OAI211_X1 U12322 ( .C1(n14807), .C2(n9907), .A(n9906), .B(n9905), .ZN(
        P2_U3219) );
  NAND2_X1 U12323 ( .A1(n9915), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9912) );
  NAND2_X1 U12324 ( .A1(n9913), .A2(n9912), .ZN(n9910) );
  MUX2_X1 U12325 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9908), .S(n9960), .Z(n9909)
         );
  NAND2_X1 U12326 ( .A1(n9910), .A2(n9909), .ZN(n13174) );
  MUX2_X1 U12327 ( .A(n9908), .B(P2_REG1_REG_6__SCAN_IN), .S(n9960), .Z(n9911)
         );
  NAND3_X1 U12328 ( .A1(n9913), .A2(n9912), .A3(n9911), .ZN(n9914) );
  NAND3_X1 U12329 ( .A1(n14779), .A2(n13174), .A3(n9914), .ZN(n9923) );
  NAND2_X1 U12330 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10613) );
  NAND2_X1 U12331 ( .A1(n9915), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U12332 ( .A1(n9917), .A2(n9916), .ZN(n9919) );
  MUX2_X1 U12333 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10670), .S(n9960), .Z(n9918) );
  NAND2_X1 U12334 ( .A1(n9919), .A2(n9918), .ZN(n13168) );
  OAI211_X1 U12335 ( .C1(n9919), .C2(n9918), .A(n14776), .B(n13168), .ZN(n9920) );
  NAND2_X1 U12336 ( .A1(n10613), .A2(n9920), .ZN(n9921) );
  AOI21_X1 U12337 ( .B1(n14773), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9921), .ZN(
        n9922) );
  OAI211_X1 U12338 ( .C1(n14807), .C2(n9924), .A(n9923), .B(n9922), .ZN(
        P2_U3220) );
  INV_X1 U12339 ( .A(n13133), .ZN(n9936) );
  INV_X1 U12340 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U12341 ( .A1(n14822), .A2(n9925), .ZN(n14710) );
  AOI22_X1 U12342 ( .A1(n14710), .A2(P2_IR_REG_0__SCAN_IN), .B1(n14779), .B2(
        n9926), .ZN(n9935) );
  INV_X1 U12343 ( .A(n9929), .ZN(n9928) );
  INV_X1 U12344 ( .A(n14807), .ZN(n14819) );
  OAI22_X1 U12345 ( .A1(n14827), .A2(n6785), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10536), .ZN(n9927) );
  AOI21_X1 U12346 ( .B1(n9928), .B2(n14819), .A(n9927), .ZN(n9934) );
  MUX2_X1 U12347 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9889), .S(n9929), .Z(n9930)
         );
  OAI21_X1 U12348 ( .B1(n7568), .B2(n9931), .A(n9930), .ZN(n9932) );
  NAND3_X1 U12349 ( .A1(n14776), .A2(n13138), .A3(n9932), .ZN(n9933) );
  OAI211_X1 U12350 ( .C1(n9936), .C2(n9935), .A(n9934), .B(n9933), .ZN(
        P2_U3215) );
  NAND2_X1 U12351 ( .A1(n9937), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12225) );
  NAND2_X1 U12352 ( .A1(n9946), .A2(n12225), .ZN(n9997) );
  OAI21_X1 U12353 ( .B1(n11979), .B2(n9937), .A(n11835), .ZN(n9995) );
  NAND2_X1 U12354 ( .A1(n9997), .A2(n9995), .ZN(n14544) );
  INV_X1 U12355 ( .A(n14544), .ZN(n13776) );
  NOR2_X1 U12356 ( .A1(n13776), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12357 ( .A(n11086), .ZN(n9944) );
  NAND2_X1 U12358 ( .A1(n9940), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9938) );
  MUX2_X1 U12359 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9938), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n9939) );
  INV_X1 U12360 ( .A(n9939), .ZN(n9941) );
  NOR2_X1 U12361 ( .A1(n9941), .A2(n10104), .ZN(n11087) );
  INV_X1 U12362 ( .A(n11087), .ZN(n9942) );
  OAI222_X1 U12363 ( .A1(n14245), .A2(n9943), .B1(n14244), .B2(n9944), .C1(
        P1_U3086), .C2(n9942), .ZN(P1_U3346) );
  INV_X1 U12364 ( .A(n9984), .ZN(n14727) );
  OAI222_X1 U12365 ( .A1(n13573), .A2(n9945), .B1(n13575), .B2(n9944), .C1(
        n14727), .C2(P2_U3088), .ZN(P2_U3318) );
  INV_X1 U12366 ( .A(n9946), .ZN(n9947) );
  INV_X1 U12367 ( .A(n10404), .ZN(n9949) );
  AOI22_X1 U12368 ( .A1(n14603), .A2(n12670), .B1(n9949), .B2(n9948), .ZN(
        P1_U3445) );
  INV_X1 U12369 ( .A(n11164), .ZN(n9993) );
  OR2_X1 U12370 ( .A1(n10104), .A2(n9668), .ZN(n9950) );
  XNOR2_X1 U12371 ( .A(n9950), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U12372 ( .A1(n11165), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n11586), .ZN(n9951) );
  OAI21_X1 U12373 ( .B1(n9993), .B2(n14244), .A(n9951), .ZN(P1_U3345) );
  NAND2_X1 U12374 ( .A1(n9960), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13167) );
  NAND2_X1 U12375 ( .A1(n13168), .A2(n13167), .ZN(n9953) );
  MUX2_X1 U12376 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10711), .S(n13171), .Z(
        n9952) );
  NAND2_X1 U12377 ( .A1(n9953), .A2(n9952), .ZN(n13170) );
  NAND2_X1 U12378 ( .A1(n13171), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U12379 ( .A1(n13170), .A2(n9958), .ZN(n9956) );
  MUX2_X1 U12380 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9954), .S(n9981), .Z(n9955)
         );
  NAND2_X1 U12381 ( .A1(n9956), .A2(n9955), .ZN(n9983) );
  MUX2_X1 U12382 ( .A(n9954), .B(P2_REG2_REG_8__SCAN_IN), .S(n9981), .Z(n9957)
         );
  NAND3_X1 U12383 ( .A1(n13170), .A2(n9958), .A3(n9957), .ZN(n9959) );
  NAND3_X1 U12384 ( .A1(n14776), .A2(n9983), .A3(n9959), .ZN(n9971) );
  NAND2_X1 U12385 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10751) );
  NAND2_X1 U12386 ( .A1(n9960), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U12387 ( .A1(n13174), .A2(n13173), .ZN(n9963) );
  MUX2_X1 U12388 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9961), .S(n13171), .Z(n9962) );
  NAND2_X1 U12389 ( .A1(n9963), .A2(n9962), .ZN(n13176) );
  NAND2_X1 U12390 ( .A1(n13171), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U12391 ( .A1(n13176), .A2(n9964), .ZN(n9967) );
  MUX2_X1 U12392 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9965), .S(n9981), .Z(n9966)
         );
  NAND2_X1 U12393 ( .A1(n9967), .A2(n9966), .ZN(n9975) );
  OAI211_X1 U12394 ( .C1(n9967), .C2(n9966), .A(n14779), .B(n9975), .ZN(n9968)
         );
  NAND2_X1 U12395 ( .A1(n10751), .A2(n9968), .ZN(n9969) );
  AOI21_X1 U12396 ( .B1(n14773), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9969), .ZN(
        n9970) );
  OAI211_X1 U12397 ( .C1(n14807), .C2(n9972), .A(n9971), .B(n9970), .ZN(
        P2_U3222) );
  NAND2_X1 U12398 ( .A1(P1_U4016), .A2(n11139), .ZN(n9973) );
  OAI21_X1 U12399 ( .B1(P1_U4016), .B2(n8086), .A(n9973), .ZN(P1_U3560) );
  INV_X1 U12400 ( .A(n10090), .ZN(n9992) );
  NAND2_X1 U12401 ( .A1(n9981), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U12402 ( .A1(n9975), .A2(n9974), .ZN(n14716) );
  MUX2_X1 U12403 ( .A(n9976), .B(P2_REG1_REG_9__SCAN_IN), .S(n9984), .Z(n14715) );
  OR2_X1 U12404 ( .A1(n14716), .A2(n14715), .ZN(n14718) );
  NAND2_X1 U12405 ( .A1(n14727), .A2(n9976), .ZN(n9977) );
  AND2_X1 U12406 ( .A1(n14718), .A2(n9977), .ZN(n9980) );
  MUX2_X1 U12407 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9978), .S(n10090), .Z(
        n9979) );
  NAND2_X1 U12408 ( .A1(n9980), .A2(n9979), .ZN(n10096) );
  OAI211_X1 U12409 ( .C1(n9980), .C2(n9979), .A(n10096), .B(n14779), .ZN(n9991) );
  NAND2_X1 U12410 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10920)
         );
  NAND2_X1 U12411 ( .A1(n9981), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U12412 ( .A1(n9983), .A2(n9982), .ZN(n14721) );
  MUX2_X1 U12413 ( .A(n10835), .B(P2_REG2_REG_9__SCAN_IN), .S(n9984), .Z(
        n14720) );
  OR2_X1 U12414 ( .A1(n14721), .A2(n14720), .ZN(n14723) );
  NAND2_X1 U12415 ( .A1(n14727), .A2(n10835), .ZN(n9985) );
  AND2_X1 U12416 ( .A1(n14723), .A2(n9985), .ZN(n9987) );
  MUX2_X1 U12417 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10942), .S(n10090), .Z(
        n9986) );
  NAND2_X1 U12418 ( .A1(n9987), .A2(n9986), .ZN(n10085) );
  OAI211_X1 U12419 ( .C1(n9987), .C2(n9986), .A(n14776), .B(n10085), .ZN(n9988) );
  NAND2_X1 U12420 ( .A1(n10920), .A2(n9988), .ZN(n9989) );
  AOI21_X1 U12421 ( .B1(n14773), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9989), .ZN(
        n9990) );
  OAI211_X1 U12422 ( .C1(n14807), .C2(n9992), .A(n9991), .B(n9990), .ZN(
        P2_U3224) );
  INV_X1 U12423 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9994) );
  OAI222_X1 U12424 ( .A1(n13573), .A2(n9994), .B1(n13575), .B2(n9993), .C1(
        n9992), .C2(P2_U3088), .ZN(P2_U3317) );
  INV_X1 U12425 ( .A(n9995), .ZN(n9996) );
  NAND2_X1 U12426 ( .A1(n9997), .A2(n9996), .ZN(n10037) );
  NOR2_X1 U12427 ( .A1(n6394), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9998) );
  OR2_X1 U12428 ( .A1(n9998), .A2(n6415), .ZN(n13748) );
  INV_X1 U12429 ( .A(n13748), .ZN(n10000) );
  NAND2_X1 U12430 ( .A1(n6394), .A2(n9722), .ZN(n9999) );
  NAND2_X1 U12431 ( .A1(n10000), .A2(n9999), .ZN(n10001) );
  MUX2_X1 U12432 ( .A(n10001), .B(n10000), .S(P1_IR_REG_0__SCAN_IN), .Z(n10002) );
  OAI22_X1 U12433 ( .A1(n10037), .A2(n10002), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10863), .ZN(n10003) );
  AOI21_X1 U12434 ( .B1(n13776), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n10003), .ZN(
        n10005) );
  INV_X1 U12435 ( .A(n6394), .ZN(n13745) );
  NAND3_X1 U12436 ( .A1(n13841), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9722), .ZN(
        n10004) );
  NAND2_X1 U12437 ( .A1(n10005), .A2(n10004), .ZN(P1_U3243) );
  NOR2_X1 U12438 ( .A1(n10006), .A2(P2_U3088), .ZN(n10197) );
  INV_X1 U12439 ( .A(n10197), .ZN(n10008) );
  INV_X1 U12440 ( .A(n13097), .ZN(n10007) );
  AOI22_X1 U12441 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n10008), .B1(n10007), 
        .B2(n13129), .ZN(n10013) );
  INV_X1 U12442 ( .A(n10009), .ZN(n10011) );
  NOR3_X1 U12443 ( .A1(n7987), .A2(n10243), .A3(n13420), .ZN(n10010) );
  OAI21_X1 U12444 ( .B1(n10011), .B2(n10010), .A(n13093), .ZN(n10012) );
  OAI211_X1 U12445 ( .C1(n13102), .C2(n10014), .A(n10013), .B(n10012), .ZN(
        P2_U3204) );
  INV_X1 U12446 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10015) );
  MUX2_X1 U12447 ( .A(n10015), .B(P1_REG1_REG_2__SCAN_IN), .S(n13759), .Z(
        n10020) );
  INV_X1 U12448 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10016) );
  MUX2_X1 U12449 ( .A(n10016), .B(P1_REG1_REG_1__SCAN_IN), .S(n13738), .Z(
        n10018) );
  AND2_X1 U12450 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10017) );
  NAND2_X1 U12451 ( .A1(n10018), .A2(n10017), .ZN(n13761) );
  OR2_X1 U12452 ( .A1(n13738), .A2(n10016), .ZN(n13760) );
  NAND2_X1 U12453 ( .A1(n13761), .A2(n13760), .ZN(n10019) );
  NAND2_X1 U12454 ( .A1(n10020), .A2(n10019), .ZN(n13768) );
  INV_X1 U12455 ( .A(n13759), .ZN(n13754) );
  NAND2_X1 U12456 ( .A1(n13754), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13767) );
  NAND2_X1 U12457 ( .A1(n13768), .A2(n13767), .ZN(n10023) );
  MUX2_X1 U12458 ( .A(n10021), .B(P1_REG1_REG_3__SCAN_IN), .S(n13771), .Z(
        n10022) );
  NAND2_X1 U12459 ( .A1(n10023), .A2(n10022), .ZN(n13787) );
  INV_X1 U12460 ( .A(n13771), .ZN(n13777) );
  NAND2_X1 U12461 ( .A1(n13777), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13786) );
  NAND2_X1 U12462 ( .A1(n13787), .A2(n13786), .ZN(n10026) );
  MUX2_X1 U12463 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10024), .S(n13790), .Z(
        n10025) );
  NAND2_X1 U12464 ( .A1(n10026), .A2(n10025), .ZN(n13789) );
  NAND2_X1 U12465 ( .A1(n13790), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10027) );
  AND2_X1 U12466 ( .A1(n13789), .A2(n10027), .ZN(n10139) );
  INV_X1 U12467 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14698) );
  MUX2_X1 U12468 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n14698), .S(n10804), .Z(
        n10140) );
  NAND2_X1 U12469 ( .A1(n10139), .A2(n10140), .ZN(n10138) );
  NAND2_X1 U12470 ( .A1(n10149), .A2(n14698), .ZN(n10028) );
  NAND2_X1 U12471 ( .A1(n10138), .A2(n10028), .ZN(n13803) );
  INV_X1 U12472 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14700) );
  MUX2_X1 U12473 ( .A(n14700), .B(P1_REG1_REG_6__SCAN_IN), .S(n13807), .Z(
        n10029) );
  OR2_X1 U12474 ( .A1(n13803), .A2(n10029), .ZN(n13804) );
  NAND2_X1 U12475 ( .A1(n13807), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10030) );
  NAND2_X1 U12476 ( .A1(n13804), .A2(n10030), .ZN(n10174) );
  INV_X1 U12477 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10966) );
  MUX2_X1 U12478 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10966), .S(n10963), .Z(
        n10173) );
  NAND2_X1 U12479 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  NAND2_X1 U12480 ( .A1(n10963), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U12481 ( .A1(n10172), .A2(n10031), .ZN(n10200) );
  INV_X1 U12482 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10979) );
  MUX2_X1 U12483 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10979), .S(n10203), .Z(
        n10201) );
  OR2_X1 U12484 ( .A1(n10200), .A2(n10201), .ZN(n10198) );
  NAND2_X1 U12485 ( .A1(n10203), .A2(n10979), .ZN(n10034) );
  NAND2_X1 U12486 ( .A1(n10198), .A2(n10034), .ZN(n10032) );
  INV_X1 U12487 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14704) );
  MUX2_X1 U12488 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14704), .S(n11087), .Z(
        n10033) );
  NAND2_X1 U12489 ( .A1(n10032), .A2(n10033), .ZN(n10157) );
  INV_X1 U12490 ( .A(n10033), .ZN(n10035) );
  NAND3_X1 U12491 ( .A1(n10198), .A2(n10035), .A3(n10034), .ZN(n10036) );
  AND2_X1 U12492 ( .A1(n10157), .A2(n10036), .ZN(n10068) );
  INV_X1 U12493 ( .A(n10037), .ZN(n10042) );
  AND2_X1 U12494 ( .A1(n10042), .A2(n6415), .ZN(n14536) );
  NAND2_X1 U12495 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10038) );
  OAI21_X1 U12496 ( .B1(n14544), .B2(n10039), .A(n10038), .ZN(n10040) );
  AOI21_X1 U12497 ( .B1(n11087), .B2(n14536), .A(n10040), .ZN(n10067) );
  NOR2_X1 U12498 ( .A1(n6415), .A2(n6394), .ZN(n10041) );
  MUX2_X1 U12499 ( .A(n10043), .B(P1_REG2_REG_2__SCAN_IN), .S(n13759), .Z(
        n10047) );
  MUX2_X1 U12500 ( .A(n10044), .B(P1_REG2_REG_1__SCAN_IN), .S(n13738), .Z(
        n13741) );
  AND2_X1 U12501 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10045) );
  NAND2_X1 U12502 ( .A1(n13741), .A2(n10045), .ZN(n13756) );
  OR2_X1 U12503 ( .A1(n13738), .A2(n10044), .ZN(n13755) );
  NAND2_X1 U12504 ( .A1(n13756), .A2(n13755), .ZN(n10046) );
  NAND2_X1 U12505 ( .A1(n10047), .A2(n10046), .ZN(n13773) );
  NAND2_X1 U12506 ( .A1(n13754), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13772) );
  NAND2_X1 U12507 ( .A1(n13773), .A2(n13772), .ZN(n10050) );
  MUX2_X1 U12508 ( .A(n10048), .B(P1_REG2_REG_3__SCAN_IN), .S(n13771), .Z(
        n10049) );
  NAND2_X1 U12509 ( .A1(n10050), .A2(n10049), .ZN(n13793) );
  NAND2_X1 U12510 ( .A1(n13777), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13792) );
  NAND2_X1 U12511 ( .A1(n13793), .A2(n13792), .ZN(n10052) );
  MUX2_X1 U12512 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11129), .S(n13790), .Z(
        n10051) );
  NAND2_X1 U12513 ( .A1(n10052), .A2(n10051), .ZN(n13795) );
  NAND2_X1 U12514 ( .A1(n13790), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10142) );
  NAND2_X1 U12515 ( .A1(n13795), .A2(n10142), .ZN(n10054) );
  INV_X1 U12516 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10895) );
  MUX2_X1 U12517 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10895), .S(n10804), .Z(
        n10053) );
  NAND2_X1 U12518 ( .A1(n10054), .A2(n10053), .ZN(n13810) );
  NAND2_X1 U12519 ( .A1(n10804), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n13809) );
  NAND2_X1 U12520 ( .A1(n13810), .A2(n13809), .ZN(n10056) );
  INV_X1 U12521 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10817) );
  MUX2_X1 U12522 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10817), .S(n13807), .Z(
        n10055) );
  NAND2_X1 U12523 ( .A1(n10056), .A2(n10055), .ZN(n13812) );
  NAND2_X1 U12524 ( .A1(n13807), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10178) );
  NAND2_X1 U12525 ( .A1(n13812), .A2(n10178), .ZN(n10058) );
  INV_X1 U12526 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10970) );
  MUX2_X1 U12527 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10970), .S(n10963), .Z(
        n10057) );
  NAND2_X1 U12528 ( .A1(n10058), .A2(n10057), .ZN(n10206) );
  NAND2_X1 U12529 ( .A1(n10963), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10205) );
  NAND2_X1 U12530 ( .A1(n10206), .A2(n10205), .ZN(n10060) );
  INV_X1 U12531 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10983) );
  MUX2_X1 U12532 ( .A(n10983), .B(P1_REG2_REG_8__SCAN_IN), .S(n10203), .Z(
        n10059) );
  NAND2_X1 U12533 ( .A1(n10060), .A2(n10059), .ZN(n10208) );
  INV_X1 U12534 ( .A(n10203), .ZN(n11082) );
  NAND2_X1 U12535 ( .A1(n11082), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U12536 ( .A1(n10208), .A2(n10063), .ZN(n10062) );
  INV_X1 U12537 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11115) );
  MUX2_X1 U12538 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11115), .S(n11087), .Z(
        n10061) );
  NAND2_X1 U12539 ( .A1(n10062), .A2(n10061), .ZN(n10165) );
  MUX2_X1 U12540 ( .A(n11115), .B(P1_REG2_REG_9__SCAN_IN), .S(n11087), .Z(
        n10064) );
  NAND3_X1 U12541 ( .A1(n10064), .A2(n10208), .A3(n10063), .ZN(n10065) );
  NAND3_X1 U12542 ( .A1(n13846), .A2(n10165), .A3(n10065), .ZN(n10066) );
  OAI211_X1 U12543 ( .C1(n10068), .C2(n14533), .A(n10067), .B(n10066), .ZN(
        P1_U3252) );
  OAI211_X1 U12544 ( .C1(n10071), .C2(n10070), .A(n14776), .B(n10069), .ZN(
        n10076) );
  OAI211_X1 U12545 ( .C1(n10074), .C2(n10073), .A(n14779), .B(n10072), .ZN(
        n10075) );
  NAND2_X1 U12546 ( .A1(n10076), .A2(n10075), .ZN(n10078) );
  NAND2_X1 U12547 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10380) );
  INV_X1 U12548 ( .A(n10380), .ZN(n10077) );
  AOI211_X1 U12549 ( .C1(n14773), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n10078), .B(
        n10077), .ZN(n10079) );
  OAI21_X1 U12550 ( .B1(n10080), .B2(n14807), .A(n10079), .ZN(P2_U3218) );
  INV_X1 U12551 ( .A(n14603), .ZN(n14602) );
  OAI22_X1 U12552 ( .A1(n14602), .A2(P1_D_REG_1__SCAN_IN), .B1(n10082), .B2(
        n10081), .ZN(n10083) );
  INV_X1 U12553 ( .A(n10083), .ZN(P1_U3446) );
  NAND2_X1 U12554 ( .A1(n10090), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U12555 ( .A1(n10085), .A2(n10084), .ZN(n10088) );
  MUX2_X1 U12556 ( .A(n11241), .B(P2_REG2_REG_11__SCAN_IN), .S(n11384), .Z(
        n10087) );
  INV_X1 U12557 ( .A(n14739), .ZN(n10086) );
  AOI21_X1 U12558 ( .B1(n10088), .B2(n10087), .A(n10086), .ZN(n10100) );
  AND2_X1 U12559 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11227) );
  INV_X1 U12560 ( .A(n11384), .ZN(n10101) );
  NOR2_X1 U12561 ( .A1(n14807), .A2(n10101), .ZN(n10089) );
  AOI211_X1 U12562 ( .C1(n14773), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11227), 
        .B(n10089), .ZN(n10099) );
  NAND2_X1 U12563 ( .A1(n10090), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U12564 ( .A1(n10096), .A2(n10095), .ZN(n10093) );
  MUX2_X1 U12565 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10091), .S(n11384), .Z(
        n10092) );
  NAND2_X1 U12566 ( .A1(n10093), .A2(n10092), .ZN(n11386) );
  MUX2_X1 U12567 ( .A(n10091), .B(P2_REG1_REG_11__SCAN_IN), .S(n11384), .Z(
        n10094) );
  NAND3_X1 U12568 ( .A1(n10096), .A2(n10095), .A3(n10094), .ZN(n10097) );
  NAND3_X1 U12569 ( .A1(n11386), .A2(n14779), .A3(n10097), .ZN(n10098) );
  OAI211_X1 U12570 ( .C1(n10100), .C2(n14816), .A(n10099), .B(n10098), .ZN(
        P2_U3225) );
  INV_X1 U12571 ( .A(n11171), .ZN(n10106) );
  OAI222_X1 U12572 ( .A1(n13573), .A2(n10102), .B1(n13575), .B2(n10106), .C1(
        n10101), .C2(P2_U3088), .ZN(P2_U3316) );
  INV_X1 U12573 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10103) );
  NAND2_X1 U12574 ( .A1(n10104), .A2(n10103), .ZN(n10183) );
  NAND2_X1 U12575 ( .A1(n10183), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10105) );
  XNOR2_X1 U12576 ( .A(n10105), .B(P1_IR_REG_11__SCAN_IN), .ZN(n13822) );
  INV_X1 U12577 ( .A(n13822), .ZN(n10221) );
  OAI222_X1 U12578 ( .A1(n14245), .A2(n10107), .B1(n14244), .B2(n10106), .C1(
        P1_U3086), .C2(n10221), .ZN(P1_U3344) );
  CLKBUF_X1 U12579 ( .A(n10111), .Z(n10135) );
  INV_X1 U12580 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10110) );
  NOR2_X1 U12581 ( .A1(n10135), .A2(n10110), .ZN(P3_U3256) );
  INV_X1 U12582 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10112) );
  NOR2_X1 U12583 ( .A1(n10135), .A2(n10112), .ZN(P3_U3258) );
  INV_X1 U12584 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10113) );
  NOR2_X1 U12585 ( .A1(n10135), .A2(n10113), .ZN(P3_U3257) );
  INV_X1 U12586 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10114) );
  NOR2_X1 U12587 ( .A1(n10135), .A2(n10114), .ZN(P3_U3254) );
  INV_X1 U12588 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10115) );
  NOR2_X1 U12589 ( .A1(n10135), .A2(n10115), .ZN(P3_U3259) );
  INV_X1 U12590 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10116) );
  NOR2_X1 U12591 ( .A1(n10111), .A2(n10116), .ZN(P3_U3262) );
  INV_X1 U12592 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10117) );
  NOR2_X1 U12593 ( .A1(n10135), .A2(n10117), .ZN(P3_U3263) );
  INV_X1 U12594 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10118) );
  NOR2_X1 U12595 ( .A1(n10135), .A2(n10118), .ZN(P3_U3247) );
  INV_X1 U12596 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10119) );
  NOR2_X1 U12597 ( .A1(n10135), .A2(n10119), .ZN(P3_U3251) );
  INV_X1 U12598 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10120) );
  NOR2_X1 U12599 ( .A1(n10111), .A2(n10120), .ZN(P3_U3260) );
  INV_X1 U12600 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10121) );
  NOR2_X1 U12601 ( .A1(n10135), .A2(n10121), .ZN(P3_U3253) );
  INV_X1 U12602 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10122) );
  NOR2_X1 U12603 ( .A1(n10111), .A2(n10122), .ZN(P3_U3237) );
  INV_X1 U12604 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U12605 ( .A1(n10135), .A2(n10123), .ZN(P3_U3255) );
  INV_X1 U12606 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10124) );
  NOR2_X1 U12607 ( .A1(n10111), .A2(n10124), .ZN(P3_U3239) );
  INV_X1 U12608 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U12609 ( .A1(n10111), .A2(n10125), .ZN(P3_U3240) );
  INV_X1 U12610 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10126) );
  NOR2_X1 U12611 ( .A1(n10111), .A2(n10126), .ZN(P3_U3241) );
  INV_X1 U12612 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10127) );
  NOR2_X1 U12613 ( .A1(n10111), .A2(n10127), .ZN(P3_U3242) );
  INV_X1 U12614 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U12615 ( .A1(n10111), .A2(n10128), .ZN(P3_U3243) );
  INV_X1 U12616 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10129) );
  NOR2_X1 U12617 ( .A1(n10135), .A2(n10129), .ZN(P3_U3261) );
  INV_X1 U12618 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U12619 ( .A1(n10111), .A2(n10130), .ZN(P3_U3245) );
  INV_X1 U12620 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n12661) );
  NOR2_X1 U12621 ( .A1(n10135), .A2(n12661), .ZN(P3_U3246) );
  INV_X1 U12622 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10131) );
  NOR2_X1 U12623 ( .A1(n10111), .A2(n10131), .ZN(P3_U3244) );
  INV_X1 U12624 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10132) );
  NOR2_X1 U12625 ( .A1(n10135), .A2(n10132), .ZN(P3_U3248) );
  INV_X1 U12626 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10133) );
  NOR2_X1 U12627 ( .A1(n10135), .A2(n10133), .ZN(P3_U3249) );
  INV_X1 U12628 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10134) );
  NOR2_X1 U12629 ( .A1(n10111), .A2(n10134), .ZN(P3_U3236) );
  INV_X1 U12630 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n12671) );
  NOR2_X1 U12631 ( .A1(n10135), .A2(n12671), .ZN(P3_U3234) );
  INV_X1 U12632 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n12644) );
  NOR2_X1 U12633 ( .A1(n10135), .A2(n12644), .ZN(P3_U3252) );
  INV_X1 U12634 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n12688) );
  NOR2_X1 U12635 ( .A1(n10135), .A2(n12688), .ZN(P3_U3250) );
  INV_X1 U12636 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10136) );
  NOR2_X1 U12637 ( .A1(n10135), .A2(n10136), .ZN(P3_U3235) );
  INV_X1 U12638 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10137) );
  NOR2_X1 U12639 ( .A1(n10135), .A2(n10137), .ZN(P3_U3238) );
  INV_X1 U12640 ( .A(n14536), .ZN(n11456) );
  OAI21_X1 U12641 ( .B1(n10140), .B2(n10139), .A(n10138), .ZN(n10145) );
  MUX2_X1 U12642 ( .A(n10895), .B(P1_REG2_REG_5__SCAN_IN), .S(n10804), .Z(
        n10141) );
  NAND3_X1 U12643 ( .A1(n13795), .A2(n10142), .A3(n10141), .ZN(n10143) );
  AND3_X1 U12644 ( .A1(n13846), .A2(n13810), .A3(n10143), .ZN(n10144) );
  AOI21_X1 U12645 ( .B1(n13841), .B2(n10145), .A(n10144), .ZN(n10148) );
  AND2_X1 U12646 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10146) );
  AOI21_X1 U12647 ( .B1(n13776), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10146), .ZN(
        n10147) );
  OAI211_X1 U12648 ( .C1(n10149), .C2(n11456), .A(n10148), .B(n10147), .ZN(
        P1_U3248) );
  AOI22_X1 U12649 ( .A1(n13311), .A2(n13131), .B1(n9166), .B2(n13312), .ZN(
        n10236) );
  INV_X1 U12650 ( .A(n10236), .ZN(n10150) );
  AOI22_X1 U12651 ( .A1(n13056), .A2(n10150), .B1(n13086), .B2(n10238), .ZN(
        n10156) );
  OAI21_X1 U12652 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(n10154) );
  NAND2_X1 U12653 ( .A1(n10154), .A2(n13093), .ZN(n10155) );
  OAI211_X1 U12654 ( .C1(n10197), .C2(n10536), .A(n10156), .B(n10155), .ZN(
        P2_U3194) );
  OAI21_X1 U12655 ( .B1(n11087), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10157), .ZN(
        n10159) );
  INV_X1 U12656 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14707) );
  MUX2_X1 U12657 ( .A(n14707), .B(P1_REG1_REG_10__SCAN_IN), .S(n11165), .Z(
        n10158) );
  NOR2_X1 U12658 ( .A1(n10159), .A2(n10158), .ZN(n10220) );
  AOI211_X1 U12659 ( .C1(n10159), .C2(n10158), .A(n14533), .B(n10220), .ZN(
        n10171) );
  INV_X1 U12660 ( .A(n11165), .ZN(n10169) );
  INV_X1 U12661 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10160) );
  NOR2_X1 U12662 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10160), .ZN(n13593) );
  AOI21_X1 U12663 ( .B1(n13776), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n13593), 
        .ZN(n10168) );
  NAND2_X1 U12664 ( .A1(n11087), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U12665 ( .A1(n10165), .A2(n10164), .ZN(n10162) );
  INV_X1 U12666 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11215) );
  MUX2_X1 U12667 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11215), .S(n11165), .Z(
        n10161) );
  NAND2_X1 U12668 ( .A1(n10162), .A2(n10161), .ZN(n13826) );
  MUX2_X1 U12669 ( .A(n11215), .B(P1_REG2_REG_10__SCAN_IN), .S(n11165), .Z(
        n10163) );
  NAND3_X1 U12670 ( .A1(n10165), .A2(n10164), .A3(n10163), .ZN(n10166) );
  NAND3_X1 U12671 ( .A1(n13846), .A2(n13826), .A3(n10166), .ZN(n10167) );
  OAI211_X1 U12672 ( .C1(n11456), .C2(n10169), .A(n10168), .B(n10167), .ZN(
        n10170) );
  OR2_X1 U12673 ( .A1(n10171), .A2(n10170), .ZN(P1_U3253) );
  NAND2_X1 U12674 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10990) );
  OAI211_X1 U12675 ( .C1(n10174), .C2(n10173), .A(n13841), .B(n10172), .ZN(
        n10175) );
  NAND2_X1 U12676 ( .A1(n10990), .A2(n10175), .ZN(n10176) );
  AOI21_X1 U12677 ( .B1(n13776), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10176), .ZN(
        n10181) );
  MUX2_X1 U12678 ( .A(n10970), .B(P1_REG2_REG_7__SCAN_IN), .S(n10963), .Z(
        n10177) );
  NAND3_X1 U12679 ( .A1(n13812), .A2(n10178), .A3(n10177), .ZN(n10179) );
  NAND3_X1 U12680 ( .A1(n13846), .A2(n10206), .A3(n10179), .ZN(n10180) );
  OAI211_X1 U12681 ( .C1(n11456), .C2(n10182), .A(n10181), .B(n10180), .ZN(
        P1_U3250) );
  INV_X1 U12682 ( .A(n11277), .ZN(n10188) );
  NAND2_X1 U12683 ( .A1(n10184), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10213) );
  XNOR2_X1 U12684 ( .A(n10213), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11278) );
  INV_X1 U12685 ( .A(n11278), .ZN(n10278) );
  OAI222_X1 U12686 ( .A1(n14244), .A2(n10188), .B1(n10278), .B2(P1_U3086), 
        .C1(n6711), .C2(n14245), .ZN(P1_U3343) );
  INV_X1 U12687 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n12674) );
  NAND2_X1 U12688 ( .A1(n11027), .A2(P3_U3897), .ZN(n10185) );
  OAI21_X1 U12689 ( .B1(P3_U3897), .B2(n12674), .A(n10185), .ZN(P3_U3497) );
  INV_X1 U12690 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n12715) );
  NAND2_X1 U12691 ( .A1(n11052), .A2(P3_U3897), .ZN(n10186) );
  OAI21_X1 U12692 ( .B1(P3_U3897), .B2(n12715), .A(n10186), .ZN(P3_U3496) );
  INV_X1 U12693 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n12706) );
  NAND2_X1 U12694 ( .A1(n11461), .A2(P3_U3897), .ZN(n10187) );
  OAI21_X1 U12695 ( .B1(P3_U3897), .B2(n12706), .A(n10187), .ZN(P3_U3501) );
  INV_X1 U12696 ( .A(n14742), .ZN(n11388) );
  OAI222_X1 U12697 ( .A1(n13573), .A2(n10189), .B1(n13575), .B2(n10188), .C1(
        P2_U3088), .C2(n11388), .ZN(P2_U3315) );
  OAI21_X1 U12698 ( .B1(n10192), .B2(n10191), .A(n10190), .ZN(n10193) );
  NAND2_X1 U12699 ( .A1(n10193), .A2(n13093), .ZN(n10196) );
  AOI22_X1 U12700 ( .A1(n13311), .A2(n13129), .B1(n13128), .B2(n13312), .ZN(
        n10264) );
  INV_X1 U12701 ( .A(n10264), .ZN(n10194) );
  AOI22_X1 U12702 ( .A1(n13056), .A2(n10194), .B1(n13086), .B2(n10266), .ZN(
        n10195) );
  OAI211_X1 U12703 ( .C1(n10197), .C2(n10545), .A(n10196), .B(n10195), .ZN(
        P2_U3209) );
  INV_X1 U12704 ( .A(n10198), .ZN(n10199) );
  AOI21_X1 U12705 ( .B1(n10201), .B2(n10200), .A(n10199), .ZN(n10211) );
  NOR2_X1 U12706 ( .A1(n10980), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11260) );
  NOR2_X1 U12707 ( .A1(n11456), .A2(n10203), .ZN(n10202) );
  AOI211_X1 U12708 ( .C1(n13776), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11260), .B(
        n10202), .ZN(n10210) );
  MUX2_X1 U12709 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10983), .S(n10203), .Z(
        n10204) );
  NAND3_X1 U12710 ( .A1(n10206), .A2(n10205), .A3(n10204), .ZN(n10207) );
  NAND3_X1 U12711 ( .A1(n13846), .A2(n10208), .A3(n10207), .ZN(n10209) );
  OAI211_X1 U12712 ( .C1(n10211), .C2(n14533), .A(n10210), .B(n10209), .ZN(
        P1_U3251) );
  INV_X1 U12713 ( .A(n11284), .ZN(n10250) );
  INV_X1 U12714 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10212) );
  NAND2_X1 U12715 ( .A1(n10213), .A2(n10212), .ZN(n10214) );
  NAND2_X1 U12716 ( .A1(n10214), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10421) );
  INV_X1 U12717 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10420) );
  XNOR2_X1 U12718 ( .A(n10421), .B(n10420), .ZN(n11286) );
  OAI222_X1 U12719 ( .A1(n14244), .A2(n10250), .B1(n11286), .B2(P1_U3086), 
        .C1(n11285), .C2(n14245), .ZN(P1_U3342) );
  INV_X1 U12720 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11189) );
  MUX2_X1 U12721 ( .A(n11189), .B(P1_REG2_REG_12__SCAN_IN), .S(n11278), .Z(
        n10219) );
  NAND2_X1 U12722 ( .A1(n11165), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n13825) );
  NAND2_X1 U12723 ( .A1(n13826), .A2(n13825), .ZN(n10216) );
  MUX2_X1 U12724 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n13823), .S(n13822), .Z(
        n10215) );
  NAND2_X1 U12725 ( .A1(n10216), .A2(n10215), .ZN(n13828) );
  NAND2_X1 U12726 ( .A1(n13822), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U12727 ( .A1(n13828), .A2(n10217), .ZN(n10218) );
  NOR2_X1 U12728 ( .A1(n10218), .A2(n10219), .ZN(n10277) );
  AOI21_X1 U12729 ( .B1(n10219), .B2(n10218), .A(n10277), .ZN(n10229) );
  INV_X1 U12730 ( .A(n13846), .ZN(n14539) );
  AOI21_X1 U12731 ( .B1(n11165), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10220), 
        .ZN(n13817) );
  INV_X1 U12732 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14503) );
  MUX2_X1 U12733 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14503), .S(n13822), .Z(
        n13818) );
  NAND2_X1 U12734 ( .A1(n13817), .A2(n13818), .ZN(n13816) );
  NAND2_X1 U12735 ( .A1(n10221), .A2(n14503), .ZN(n10222) );
  INV_X1 U12736 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11186) );
  MUX2_X1 U12737 ( .A(n11186), .B(P1_REG1_REG_12__SCAN_IN), .S(n11278), .Z(
        n10223) );
  AOI21_X1 U12738 ( .B1(n13816), .B2(n10222), .A(n10223), .ZN(n10274) );
  AND3_X1 U12739 ( .A1(n13816), .A2(n10223), .A3(n10222), .ZN(n10224) );
  OAI21_X1 U12740 ( .B1(n10274), .B2(n10224), .A(n13841), .ZN(n10228) );
  NOR2_X1 U12741 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11671), .ZN(n10226) );
  NOR2_X1 U12742 ( .A1(n11456), .A2(n10278), .ZN(n10225) );
  AOI211_X1 U12743 ( .C1(n13776), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n10226), 
        .B(n10225), .ZN(n10227) );
  OAI211_X1 U12744 ( .C1(n10229), .C2(n14539), .A(n10228), .B(n10227), .ZN(
        P1_U3255) );
  INV_X1 U12745 ( .A(n10260), .ZN(n10232) );
  AOI211_X1 U12746 ( .C1(n10243), .C2(n10238), .A(n13394), .B(n10232), .ZN(
        n10539) );
  INV_X1 U12747 ( .A(n10233), .ZN(n10234) );
  OAI21_X1 U12748 ( .B1(n10237), .B2(n13405), .A(n10236), .ZN(n10535) );
  AOI211_X1 U12749 ( .C1(n14440), .C2(n10534), .A(n10539), .B(n10535), .ZN(
        n10557) );
  AOI22_X1 U12750 ( .A1(n11336), .A2(n10238), .B1(n8929), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10239) );
  OAI21_X1 U12751 ( .B1(n10557), .B2(n8929), .A(n10239), .ZN(P2_U3500) );
  INV_X1 U12752 ( .A(n10240), .ZN(n10241) );
  NAND2_X1 U12753 ( .A1(n13356), .A2(n10241), .ZN(n13367) );
  NAND2_X1 U12754 ( .A1(n10243), .A2(n10242), .ZN(n10252) );
  AOI21_X1 U12755 ( .B1(n13405), .B2(n13355), .A(n10255), .ZN(n10244) );
  AOI21_X1 U12756 ( .B1(n13312), .B2(n13129), .A(n10244), .ZN(n10253) );
  OAI21_X1 U12757 ( .B1(n10245), .B2(n10252), .A(n10253), .ZN(n10248) );
  OAI22_X1 U12758 ( .A1(n13427), .A2(n7568), .B1(n10246), .B2(n13412), .ZN(
        n10247) );
  AOI21_X1 U12759 ( .B1(n10248), .B2(n13356), .A(n10247), .ZN(n10249) );
  OAI21_X1 U12760 ( .B1(n10255), .B2(n13367), .A(n10249), .ZN(P2_U3265) );
  INV_X1 U12761 ( .A(n11389), .ZN(n14749) );
  OAI222_X1 U12762 ( .A1(n13573), .A2(n10251), .B1(n13575), .B2(n10250), .C1(
        P2_U3088), .C2(n14749), .ZN(P2_U3314) );
  INV_X1 U12763 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10257) );
  OAI211_X1 U12764 ( .C1(n10255), .C2(n10254), .A(n10253), .B(n10252), .ZN(
        n13509) );
  NAND2_X1 U12765 ( .A1(n13509), .A2(n14854), .ZN(n10256) );
  OAI21_X1 U12766 ( .B1(n14457), .B2(n10257), .A(n10256), .ZN(P2_U3430) );
  OAI21_X1 U12767 ( .B1(n10259), .B2(n10263), .A(n10258), .ZN(n10543) );
  AOI21_X1 U12768 ( .B1(n10260), .B2(n10266), .A(n13394), .ZN(n10261) );
  AND2_X1 U12769 ( .A1(n10261), .A2(n10365), .ZN(n10548) );
  XNOR2_X1 U12770 ( .A(n10263), .B(n10262), .ZN(n10265) );
  OAI21_X1 U12771 ( .B1(n10265), .B2(n13405), .A(n10264), .ZN(n10544) );
  AOI211_X1 U12772 ( .C1(n14440), .C2(n10543), .A(n10548), .B(n10544), .ZN(
        n10569) );
  AOI22_X1 U12773 ( .A1(n11336), .A2(n10266), .B1(n8929), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10267) );
  OAI21_X1 U12774 ( .B1(n10569), .B2(n8929), .A(n10267), .ZN(P2_U3501) );
  XOR2_X1 U12775 ( .A(n10269), .B(n10268), .Z(n13747) );
  NAND2_X1 U12776 ( .A1(n10270), .A2(n10859), .ZN(n10393) );
  INV_X1 U12777 ( .A(n10393), .ZN(n10271) );
  CLKBUF_X1 U12778 ( .A(n13691), .Z(n13854) );
  NAND2_X1 U12779 ( .A1(n13734), .A2(n13854), .ZN(n10864) );
  OAI22_X1 U12780 ( .A1(n10271), .A2(n10863), .B1(n13712), .B2(n10864), .ZN(
        n10272) );
  AOI21_X1 U12781 ( .B1(n14470), .B2(n13747), .A(n10272), .ZN(n10273) );
  OAI21_X1 U12782 ( .B1(n13718), .B2(n11138), .A(n10273), .ZN(P1_U3232) );
  AOI21_X1 U12783 ( .B1(n11186), .B2(n10278), .A(n10274), .ZN(n10276) );
  INV_X1 U12784 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11290) );
  MUX2_X1 U12785 ( .A(n11290), .B(P1_REG1_REG_13__SCAN_IN), .S(n11286), .Z(
        n10275) );
  NAND2_X1 U12786 ( .A1(n10276), .A2(n10275), .ZN(n10431) );
  OAI211_X1 U12787 ( .C1(n10276), .C2(n10275), .A(n13841), .B(n10431), .ZN(
        n10284) );
  NAND2_X1 U12788 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13664)
         );
  AOI21_X1 U12789 ( .B1(n11189), .B2(n10278), .A(n10277), .ZN(n10280) );
  INV_X1 U12790 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11293) );
  MUX2_X1 U12791 ( .A(n11293), .B(P1_REG2_REG_13__SCAN_IN), .S(n11286), .Z(
        n10279) );
  NAND2_X1 U12792 ( .A1(n10279), .A2(n10280), .ZN(n10436) );
  OAI211_X1 U12793 ( .C1(n10280), .C2(n10279), .A(n10436), .B(n13846), .ZN(
        n10281) );
  NAND2_X1 U12794 ( .A1(n13664), .A2(n10281), .ZN(n10282) );
  AOI21_X1 U12795 ( .B1(n13776), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10282), 
        .ZN(n10283) );
  OAI211_X1 U12796 ( .C1(n11456), .C2(n11286), .A(n10284), .B(n10283), .ZN(
        P1_U3256) );
  MUX2_X1 U12797 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12449), .Z(n10312) );
  INV_X1 U12798 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n12667) );
  INV_X1 U12799 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10428) );
  MUX2_X1 U12800 ( .A(n12667), .B(n10428), .S(n12449), .Z(n14867) );
  XOR2_X1 U12801 ( .A(n10313), .B(n14866), .Z(n10310) );
  INV_X1 U12802 ( .A(n10311), .ZN(n10308) );
  INV_X1 U12803 ( .A(n10286), .ZN(n10287) );
  NAND2_X1 U12804 ( .A1(n10287), .A2(n11248), .ZN(n10299) );
  OR2_X1 U12805 ( .A1(n10288), .A2(n9450), .ZN(n10289) );
  AND2_X1 U12806 ( .A1(n6413), .A2(n10289), .ZN(n10297) );
  AND2_X1 U12807 ( .A1(n10299), .A2(n10297), .ZN(n10300) );
  MUX2_X1 U12808 ( .A(n10300), .B(P3_U3897), .S(n10291), .Z(n14865) );
  INV_X1 U12809 ( .A(n10292), .ZN(n10293) );
  INV_X1 U12810 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15111) );
  AND2_X1 U12811 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n8190), .ZN(n10295) );
  INV_X1 U12812 ( .A(n10327), .ZN(n10294) );
  OAI21_X1 U12813 ( .B1(n10311), .B2(n10295), .A(n10294), .ZN(n10296) );
  NOR2_X1 U12814 ( .A1(n10296), .A2(n15111), .ZN(n10328) );
  AOI21_X1 U12815 ( .B1(n15111), .B2(n10296), .A(n10328), .ZN(n10306) );
  INV_X1 U12816 ( .A(n10297), .ZN(n10298) );
  AOI22_X1 U12817 ( .A1(n14984), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10305) );
  NAND2_X1 U12818 ( .A1(n10300), .A2(n12449), .ZN(n14877) );
  INV_X1 U12819 ( .A(n14877), .ZN(n14989) );
  NAND2_X1 U12820 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n8190), .ZN(n10301) );
  NAND2_X1 U12821 ( .A1(n10302), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10319) );
  OAI21_X1 U12822 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n10302), .A(n10319), .ZN(
        n10303) );
  NAND2_X1 U12823 ( .A1(n14989), .A2(n10303), .ZN(n10304) );
  OAI211_X1 U12824 ( .C1(n14997), .C2(n10306), .A(n10305), .B(n10304), .ZN(
        n10307) );
  AOI21_X1 U12825 ( .B1(n10308), .B2(n14865), .A(n10307), .ZN(n10309) );
  OAI21_X1 U12826 ( .B1(n14952), .B2(n10310), .A(n10309), .ZN(P3_U3183) );
  MUX2_X1 U12827 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12449), .Z(n10486) );
  XNOR2_X1 U12828 ( .A(n10486), .B(n10498), .ZN(n10488) );
  MUX2_X1 U12829 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12449), .Z(n10314) );
  XNOR2_X1 U12830 ( .A(n10314), .B(n10351), .ZN(n10340) );
  INV_X1 U12831 ( .A(n10314), .ZN(n10315) );
  MUX2_X1 U12832 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12449), .Z(n10316) );
  XOR2_X1 U12833 ( .A(n10330), .B(n10316), .Z(n10474) );
  XOR2_X1 U12834 ( .A(n10488), .B(n10489), .Z(n10338) );
  INV_X1 U12835 ( .A(n14984), .ZN(n14886) );
  MUX2_X1 U12836 ( .A(n15147), .B(P3_REG1_REG_4__SCAN_IN), .S(n10498), .Z(
        n10323) );
  INV_X1 U12837 ( .A(n10317), .ZN(n10318) );
  NAND2_X1 U12838 ( .A1(n10319), .A2(n10318), .ZN(n10345) );
  XNOR2_X1 U12839 ( .A(n10351), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U12840 ( .A1(n10345), .A2(n10344), .B1(P3_REG1_REG_2__SCAN_IN), 
        .B2(n10329), .ZN(n10320) );
  XNOR2_X1 U12841 ( .A(n10320), .B(n10330), .ZN(n10477) );
  INV_X1 U12842 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10321) );
  OAI22_X1 U12843 ( .A1(n10477), .A2(n10321), .B1(n10330), .B2(n10320), .ZN(
        n10322) );
  NAND2_X1 U12844 ( .A1(n10322), .A2(n10323), .ZN(n10497) );
  OAI21_X1 U12845 ( .B1(n10323), .B2(n10322), .A(n10497), .ZN(n10324) );
  NAND2_X1 U12846 ( .A1(n14989), .A2(n10324), .ZN(n10326) );
  AND2_X1 U12847 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10795) );
  INV_X1 U12848 ( .A(n10795), .ZN(n10325) );
  OAI211_X1 U12849 ( .C1(n14886), .C2(n8825), .A(n10326), .B(n10325), .ZN(
        n10336) );
  NOR2_X1 U12850 ( .A1(n10328), .A2(n10327), .ZN(n10342) );
  XNOR2_X1 U12851 ( .A(n10329), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10343) );
  NOR2_X1 U12852 ( .A1(n10342), .A2(n10343), .ZN(n10341) );
  INV_X1 U12853 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10331) );
  XNOR2_X1 U12854 ( .A(n10498), .B(n10331), .ZN(n10332) );
  INV_X1 U12855 ( .A(n10491), .ZN(n10334) );
  NAND3_X1 U12856 ( .A1(n10475), .A2(n10332), .A3(n6440), .ZN(n10333) );
  AOI21_X1 U12857 ( .B1(n10334), .B2(n10333), .A(n14997), .ZN(n10335) );
  AOI211_X1 U12858 ( .C1(n14865), .C2(n10498), .A(n10336), .B(n10335), .ZN(
        n10337) );
  OAI21_X1 U12859 ( .B1(n10338), .B2(n14952), .A(n10337), .ZN(P3_U3186) );
  XOR2_X1 U12860 ( .A(n10339), .B(n10340), .Z(n10353) );
  AOI21_X1 U12861 ( .B1(n10343), .B2(n10342), .A(n10341), .ZN(n10349) );
  AOI22_X1 U12862 ( .A1(n14984), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10348) );
  XNOR2_X1 U12863 ( .A(n10345), .B(n10344), .ZN(n10346) );
  NAND2_X1 U12864 ( .A1(n14989), .A2(n10346), .ZN(n10347) );
  OAI211_X1 U12865 ( .C1(n14997), .C2(n10349), .A(n10348), .B(n10347), .ZN(
        n10350) );
  AOI21_X1 U12866 ( .B1(n10351), .B2(n14865), .A(n10350), .ZN(n10352) );
  OAI21_X1 U12867 ( .B1(n10353), .B2(n14952), .A(n10352), .ZN(P3_U3184) );
  INV_X1 U12868 ( .A(n10355), .ZN(n10356) );
  AOI21_X1 U12869 ( .B1(n10354), .B2(n10357), .A(n10356), .ZN(n10362) );
  NAND2_X1 U12870 ( .A1(n13733), .A2(n13854), .ZN(n11140) );
  OAI21_X1 U12871 ( .B1(n10358), .B2(n13903), .A(n11140), .ZN(n10359) );
  AOI22_X1 U12872 ( .A1(n14472), .A2(n10359), .B1(n10393), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10361) );
  NAND2_X1 U12873 ( .A1(n14475), .A2(n11992), .ZN(n10360) );
  OAI211_X1 U12874 ( .C1(n10362), .C2(n13705), .A(n10361), .B(n10360), .ZN(
        P1_U3222) );
  OAI21_X1 U12875 ( .B1(n10364), .B2(n10366), .A(n10363), .ZN(n10459) );
  AOI211_X1 U12876 ( .C1(n6399), .C2(n10365), .A(n13394), .B(n10452), .ZN(
        n10464) );
  XNOR2_X1 U12877 ( .A(n10367), .B(n10366), .ZN(n10370) );
  NAND2_X1 U12878 ( .A1(n13127), .A2(n13312), .ZN(n10369) );
  NAND2_X1 U12879 ( .A1(n9166), .A2(n13311), .ZN(n10368) );
  AND2_X1 U12880 ( .A1(n10369), .A2(n10368), .ZN(n13006) );
  OAI21_X1 U12881 ( .B1(n10370), .B2(n13405), .A(n13006), .ZN(n10460) );
  AOI211_X1 U12882 ( .C1(n14440), .C2(n10459), .A(n10464), .B(n10460), .ZN(
        n10566) );
  AOI22_X1 U12883 ( .A1(n11336), .A2(n6399), .B1(n8929), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10371) );
  OAI21_X1 U12884 ( .B1(n10566), .B2(n8929), .A(n10371), .ZN(P2_U3502) );
  INV_X1 U12885 ( .A(n10372), .ZN(n10373) );
  AOI21_X1 U12886 ( .B1(n10375), .B2(n10374), .A(n10373), .ZN(n10383) );
  NAND2_X1 U12887 ( .A1(n13126), .A2(n13312), .ZN(n10377) );
  NAND2_X1 U12888 ( .A1(n13128), .A2(n13311), .ZN(n10376) );
  AND2_X1 U12889 ( .A1(n10377), .A2(n10376), .ZN(n10448) );
  INV_X1 U12890 ( .A(n10448), .ZN(n10378) );
  NAND2_X1 U12891 ( .A1(n13056), .A2(n10378), .ZN(n10379) );
  OAI211_X1 U12892 ( .C1(n13096), .C2(n10454), .A(n10380), .B(n10379), .ZN(
        n10381) );
  AOI21_X1 U12893 ( .B1(n10471), .B2(n13086), .A(n10381), .ZN(n10382) );
  OAI21_X1 U12894 ( .B1(n10383), .B2(n13088), .A(n10382), .ZN(P2_U3202) );
  INV_X1 U12895 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U12896 ( .A1(n12581), .A2(P3_U3897), .ZN(n10384) );
  OAI21_X1 U12897 ( .B1(P3_U3897), .B2(n12668), .A(n10384), .ZN(P3_U3513) );
  INV_X1 U12898 ( .A(n11686), .ZN(n10425) );
  INV_X1 U12899 ( .A(n10385), .ZN(n10386) );
  NAND2_X1 U12900 ( .A1(n10386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10387) );
  MUX2_X1 U12901 ( .A(n10387), .B(P1_IR_REG_31__SCAN_IN), .S(n12612), .Z(
        n10388) );
  NAND2_X1 U12902 ( .A1(n10388), .A2(n9667), .ZN(n11012) );
  OAI222_X1 U12903 ( .A1(n14244), .A2(n10425), .B1(n11012), .B2(P1_U3086), 
        .C1(n12704), .C2(n14245), .ZN(P1_U3339) );
  OAI21_X1 U12904 ( .B1(n10391), .B2(n10390), .A(n10389), .ZN(n10392) );
  NAND2_X1 U12905 ( .A1(n10392), .A2(n14470), .ZN(n10395) );
  OAI22_X1 U12906 ( .A1(n12006), .A2(n14098), .B1(n10881), .B2(n13903), .ZN(
        n14583) );
  AOI22_X1 U12907 ( .A1(n14472), .A2(n14583), .B1(n10393), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10394) );
  OAI211_X1 U12908 ( .C1(n13718), .C2(n14616), .A(n10395), .B(n10394), .ZN(
        P1_U3237) );
  INV_X1 U12909 ( .A(n10396), .ZN(n10398) );
  OAI22_X1 U12910 ( .A1(n14361), .A2(P3_U3151), .B1(SI_17_), .B2(n14275), .ZN(
        n10397) );
  AOI21_X1 U12911 ( .B1(n10398), .B2(n14288), .A(n10397), .ZN(P3_U3278) );
  INV_X1 U12912 ( .A(n10399), .ZN(n10400) );
  NOR2_X1 U12913 ( .A1(n12222), .A2(n10400), .ZN(n10401) );
  AND2_X1 U12914 ( .A1(n10858), .A2(n10401), .ZN(n10417) );
  INV_X1 U12915 ( .A(n10405), .ZN(n10403) );
  NAND2_X1 U12916 ( .A1(n10403), .A2(n10402), .ZN(n10407) );
  OAI21_X1 U12917 ( .B1(n10405), .B2(P1_D_REG_0__SCAN_IN), .A(n10404), .ZN(
        n10406) );
  AND2_X1 U12918 ( .A1(n11985), .A2(n11971), .ZN(n10408) );
  NAND2_X1 U12919 ( .A1(n14561), .A2(n12226), .ZN(n14568) );
  NAND2_X1 U12920 ( .A1(n11970), .A2(n11977), .ZN(n14656) );
  NAND2_X1 U12921 ( .A1(n9777), .A2(n10409), .ZN(n11969) );
  NAND2_X1 U12922 ( .A1(n14250), .A2(n14559), .ZN(n10410) );
  NAND2_X2 U12923 ( .A1(n11969), .A2(n10410), .ZN(n14625) );
  OAI21_X1 U12924 ( .B1(n11139), .B2(n10411), .A(n11134), .ZN(n12184) );
  INV_X1 U12925 ( .A(n12184), .ZN(n10412) );
  OAI21_X1 U12926 ( .B1(n14683), .B2(n14625), .A(n10412), .ZN(n10413) );
  OAI211_X1 U12927 ( .C1(n11138), .C2(n11966), .A(n10413), .B(n10864), .ZN(
        n10418) );
  NAND2_X1 U12928 ( .A1(n14693), .A2(n10418), .ZN(n10414) );
  OAI21_X1 U12929 ( .B1(n14693), .B2(n9723), .A(n10414), .ZN(P1_U3459) );
  INV_X1 U12930 ( .A(n10415), .ZN(n10416) );
  NAND2_X1 U12931 ( .A1(n14709), .A2(n10418), .ZN(n10419) );
  OAI21_X1 U12932 ( .B1(n14709), .B2(n9722), .A(n10419), .ZN(P1_U3528) );
  INV_X1 U12933 ( .A(n11516), .ZN(n10442) );
  NAND2_X1 U12934 ( .A1(n10421), .A2(n10420), .ZN(n10422) );
  NAND2_X1 U12935 ( .A1(n10422), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10423) );
  XNOR2_X1 U12936 ( .A(n10423), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11517) );
  INV_X1 U12937 ( .A(n11517), .ZN(n10733) );
  OAI222_X1 U12938 ( .A1(n14244), .A2(n10442), .B1(n10733), .B2(P1_U3086), 
        .C1(n6630), .C2(n14245), .ZN(P1_U3341) );
  INV_X1 U12939 ( .A(n11383), .ZN(n14793) );
  OAI222_X1 U12940 ( .A1(P2_U3088), .A2(n14793), .B1(n13575), .B2(n10425), 
        .C1(n10424), .C2(n13573), .ZN(P2_U3311) );
  OR3_X1 U12941 ( .A1(n14858), .A2(n14410), .A3(n10426), .ZN(n10427) );
  OAI21_X1 U12942 ( .B1(n6694), .B2(n15046), .A(n10427), .ZN(n10633) );
  NOR2_X1 U12943 ( .A1(n15159), .A2(n10428), .ZN(n10429) );
  AOI21_X1 U12944 ( .B1(n15159), .B2(n10633), .A(n10429), .ZN(n10430) );
  OAI21_X1 U12945 ( .B1(n10588), .B2(n12899), .A(n10430), .ZN(P3_U3459) );
  INV_X1 U12946 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U12947 ( .A1(n11517), .A2(n14488), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10733), .ZN(n10433) );
  OAI21_X1 U12948 ( .B1(n11286), .B2(n11290), .A(n10431), .ZN(n10432) );
  NOR2_X1 U12949 ( .A1(n10433), .A2(n10432), .ZN(n10727) );
  AOI21_X1 U12950 ( .B1(n10433), .B2(n10432), .A(n10727), .ZN(n10441) );
  NAND2_X1 U12951 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14464)
         );
  OAI21_X1 U12952 ( .B1(n14544), .B2(n10434), .A(n14464), .ZN(n10435) );
  AOI21_X1 U12953 ( .B1(n11517), .B2(n14536), .A(n10435), .ZN(n10440) );
  INV_X1 U12954 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14105) );
  MUX2_X1 U12955 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14105), .S(n11517), .Z(
        n10438) );
  OAI21_X1 U12956 ( .B1(n11286), .B2(n11293), .A(n10436), .ZN(n10437) );
  NAND2_X1 U12957 ( .A1(n10438), .A2(n10437), .ZN(n10732) );
  OAI211_X1 U12958 ( .C1(n10438), .C2(n10437), .A(n13846), .B(n10732), .ZN(
        n10439) );
  OAI211_X1 U12959 ( .C1(n10441), .C2(n14533), .A(n10440), .B(n10439), .ZN(
        P1_U3257) );
  OAI222_X1 U12960 ( .A1(n13573), .A2(n10443), .B1(n13575), .B2(n10442), .C1(
        P2_U3088), .C2(n14772), .ZN(P2_U3313) );
  OAI21_X1 U12961 ( .B1(n10445), .B2(n10446), .A(n10444), .ZN(n10470) );
  INV_X1 U12962 ( .A(n10470), .ZN(n10458) );
  XNOR2_X1 U12963 ( .A(n10447), .B(n10446), .ZN(n10449) );
  OAI21_X1 U12964 ( .B1(n10449), .B2(n13405), .A(n10448), .ZN(n10468) );
  INV_X1 U12965 ( .A(n10468), .ZN(n10450) );
  MUX2_X1 U12966 ( .A(n10451), .B(n10450), .S(n13427), .Z(n10457) );
  OR2_X1 U12967 ( .A1(n10452), .A2(n10559), .ZN(n10453) );
  AND3_X1 U12968 ( .A1(n10601), .A2(n13420), .A3(n10453), .ZN(n10469) );
  OAI22_X1 U12969 ( .A1(n13376), .A2(n10559), .B1(n10454), .B2(n13412), .ZN(
        n10455) );
  AOI21_X1 U12970 ( .B1(n10469), .B2(n13422), .A(n10455), .ZN(n10456) );
  OAI211_X1 U12971 ( .C1(n13425), .C2(n10458), .A(n10457), .B(n10456), .ZN(
        P2_U3261) );
  INV_X1 U12972 ( .A(n10459), .ZN(n10467) );
  INV_X1 U12973 ( .A(n10460), .ZN(n10461) );
  MUX2_X1 U12974 ( .A(n10462), .B(n10461), .S(n13427), .Z(n10466) );
  OAI22_X1 U12975 ( .A1(n13376), .A2(n10563), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13412), .ZN(n10463) );
  AOI21_X1 U12976 ( .B1(n10464), .B2(n13422), .A(n10463), .ZN(n10465) );
  OAI211_X1 U12977 ( .C1(n10467), .C2(n13425), .A(n10466), .B(n10465), .ZN(
        P2_U3262) );
  AOI211_X1 U12978 ( .C1(n14440), .C2(n10470), .A(n10469), .B(n10468), .ZN(
        n10562) );
  AOI22_X1 U12979 ( .A1(n11336), .A2(n10471), .B1(n8929), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n10472) );
  OAI21_X1 U12980 ( .B1(n10562), .B2(n8929), .A(n10472), .ZN(P2_U3503) );
  XOR2_X1 U12981 ( .A(n10473), .B(n10474), .Z(n10485) );
  OAI21_X1 U12982 ( .B1(n10476), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10475), .ZN(
        n10483) );
  XOR2_X1 U12983 ( .A(P3_REG1_REG_3__SCAN_IN), .B(n10477), .Z(n10478) );
  NAND2_X1 U12984 ( .A1(n14989), .A2(n10478), .ZN(n10479) );
  NAND2_X1 U12985 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n10682) );
  OAI211_X1 U12986 ( .C1(n10480), .C2(n14886), .A(n10479), .B(n10682), .ZN(
        n10482) );
  NOR2_X1 U12987 ( .A1(n14987), .A2(n7120), .ZN(n10481) );
  AOI211_X1 U12988 ( .C1(n14385), .C2(n10483), .A(n10482), .B(n10481), .ZN(
        n10484) );
  OAI21_X1 U12989 ( .B1(n10485), .B2(n14952), .A(n10484), .ZN(P3_U3185) );
  INV_X1 U12990 ( .A(n10486), .ZN(n10487) );
  MUX2_X1 U12991 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12449), .Z(n10490) );
  XOR2_X1 U12992 ( .A(n10499), .B(n10490), .Z(n14873) );
  MUX2_X1 U12993 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12449), .Z(n10515) );
  XNOR2_X1 U12994 ( .A(n10515), .B(n10520), .ZN(n10517) );
  XNOR2_X1 U12995 ( .A(n10518), .B(n10517), .ZN(n10513) );
  INV_X1 U12996 ( .A(n14952), .ZN(n14991) );
  INV_X1 U12997 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15037) );
  NAND2_X1 U12998 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10525), .ZN(n10494) );
  OAI21_X1 U12999 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10525), .A(n10494), .ZN(
        n10495) );
  AOI21_X1 U13000 ( .B1(n10496), .B2(n10495), .A(n10524), .ZN(n10511) );
  INV_X1 U13001 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15151) );
  AOI22_X1 U13002 ( .A1(n10520), .A2(n15151), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n10525), .ZN(n10504) );
  INV_X1 U13003 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15147) );
  OAI21_X1 U13004 ( .B1(n10498), .B2(n15147), .A(n10497), .ZN(n10500) );
  NAND2_X1 U13005 ( .A1(n10500), .A2(n6844), .ZN(n10502) );
  XNOR2_X1 U13006 ( .A(n10500), .B(n10499), .ZN(n14875) );
  NAND2_X1 U13007 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14875), .ZN(n10501) );
  NAND2_X1 U13008 ( .A1(n10502), .A2(n10501), .ZN(n10503) );
  NAND2_X1 U13009 ( .A1(n10504), .A2(n10503), .ZN(n10519) );
  OAI21_X1 U13010 ( .B1(n10504), .B2(n10503), .A(n10519), .ZN(n10505) );
  INV_X1 U13011 ( .A(n10505), .ZN(n10507) );
  AND2_X1 U13012 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10931) );
  AOI21_X1 U13013 ( .B1(n14984), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10931), .ZN(
        n10506) );
  OAI21_X1 U13014 ( .B1(n14877), .B2(n10507), .A(n10506), .ZN(n10508) );
  INV_X1 U13015 ( .A(n10508), .ZN(n10510) );
  NAND2_X1 U13016 ( .A1(n14865), .A2(n10520), .ZN(n10509) );
  OAI211_X1 U13017 ( .C1(n14997), .C2(n10511), .A(n10510), .B(n10509), .ZN(
        n10512) );
  AOI21_X1 U13018 ( .B1(n10513), .B2(n14991), .A(n10512), .ZN(n10514) );
  INV_X1 U13019 ( .A(n10514), .ZN(P3_U3188) );
  MUX2_X1 U13020 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12449), .Z(n10645) );
  XNOR2_X1 U13021 ( .A(n10645), .B(n10644), .ZN(n10646) );
  INV_X1 U13022 ( .A(n10515), .ZN(n10516) );
  AOI22_X1 U13023 ( .A1(n10518), .A2(n10517), .B1(n10520), .B2(n10516), .ZN(
        n10647) );
  XOR2_X1 U13024 ( .A(n10647), .B(n10646), .Z(n10533) );
  OAI21_X1 U13025 ( .B1(n10520), .B2(n15151), .A(n10519), .ZN(n10639) );
  OAI21_X1 U13026 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10521), .A(n10640), .ZN(
        n10531) );
  INV_X1 U13027 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10522) );
  NOR2_X1 U13028 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10522), .ZN(n11040) );
  AOI21_X1 U13029 ( .B1(n14984), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11040), .ZN(
        n10523) );
  OAI21_X1 U13030 ( .B1(n14987), .B2(n10644), .A(n10523), .ZN(n10530) );
  INV_X1 U13031 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10526) );
  AOI21_X1 U13032 ( .B1(n10527), .B2(n10526), .A(n10653), .ZN(n10528) );
  NOR2_X1 U13033 ( .A1(n10528), .A2(n14997), .ZN(n10529) );
  AOI211_X1 U13034 ( .C1(n14989), .C2(n10531), .A(n10530), .B(n10529), .ZN(
        n10532) );
  OAI21_X1 U13035 ( .B1(n10533), .B2(n14952), .A(n10532), .ZN(P3_U3189) );
  INV_X1 U13036 ( .A(n10534), .ZN(n10542) );
  NAND2_X1 U13037 ( .A1(n10535), .A2(n13427), .ZN(n10541) );
  OAI22_X1 U13038 ( .A1(n13427), .A2(n9889), .B1(n10536), .B2(n13412), .ZN(
        n10538) );
  NOR2_X1 U13039 ( .A1(n13376), .A2(n10554), .ZN(n10537) );
  AOI211_X1 U13040 ( .C1(n10539), .C2(n13422), .A(n10538), .B(n10537), .ZN(
        n10540) );
  OAI211_X1 U13041 ( .C1(n13425), .C2(n10542), .A(n10541), .B(n10540), .ZN(
        P2_U3264) );
  INV_X1 U13042 ( .A(n10543), .ZN(n10551) );
  NAND2_X1 U13043 ( .A1(n10544), .A2(n13356), .ZN(n10550) );
  OAI22_X1 U13044 ( .A1(n13427), .A2(n9888), .B1(n10545), .B2(n13412), .ZN(
        n10547) );
  NOR2_X1 U13045 ( .A1(n13376), .A2(n7605), .ZN(n10546) );
  AOI211_X1 U13046 ( .C1(n10548), .C2(n13422), .A(n10547), .B(n10546), .ZN(
        n10549) );
  OAI211_X1 U13047 ( .C1(n10551), .C2(n13425), .A(n10550), .B(n10549), .ZN(
        P2_U3263) );
  INV_X1 U13048 ( .A(n11742), .ZN(n10590) );
  NAND2_X1 U13049 ( .A1(n9667), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10552) );
  MUX2_X1 U13050 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10552), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n10553) );
  AND2_X1 U13051 ( .A1(n10553), .A2(n10687), .ZN(n11743) );
  INV_X1 U13052 ( .A(n11743), .ZN(n11448) );
  OAI222_X1 U13053 ( .A1(n14244), .A2(n10590), .B1(n11448), .B2(P1_U3086), 
        .C1(n6632), .C2(n14245), .ZN(P1_U3338) );
  OAI22_X1 U13054 ( .A1(n13548), .A2(n10554), .B1(n14854), .B2(n7575), .ZN(
        n10555) );
  INV_X1 U13055 ( .A(n10555), .ZN(n10556) );
  OAI21_X1 U13056 ( .B1(n10557), .B2(n14450), .A(n10556), .ZN(P2_U3433) );
  INV_X1 U13057 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10558) );
  OAI22_X1 U13058 ( .A1(n13548), .A2(n10559), .B1(n14854), .B2(n10558), .ZN(
        n10560) );
  INV_X1 U13059 ( .A(n10560), .ZN(n10561) );
  OAI21_X1 U13060 ( .B1(n10562), .B2(n14450), .A(n10561), .ZN(P2_U3442) );
  OAI22_X1 U13061 ( .A1(n13548), .A2(n10563), .B1(n14854), .B2(n7607), .ZN(
        n10564) );
  INV_X1 U13062 ( .A(n10564), .ZN(n10565) );
  OAI21_X1 U13063 ( .B1(n10566), .B2(n14450), .A(n10565), .ZN(P2_U3439) );
  OAI22_X1 U13064 ( .A1(n13548), .A2(n7605), .B1(n14854), .B2(n7600), .ZN(
        n10567) );
  INV_X1 U13065 ( .A(n10567), .ZN(n10568) );
  OAI21_X1 U13066 ( .B1(n10569), .B2(n14450), .A(n10568), .ZN(P2_U3436) );
  OAI21_X1 U13067 ( .B1(n10572), .B2(n10571), .A(n10570), .ZN(n10580) );
  NOR2_X1 U13068 ( .A1(n13102), .A2(n6760), .ZN(n10579) );
  NAND2_X1 U13069 ( .A1(n13125), .A2(n13312), .ZN(n10574) );
  NAND2_X1 U13070 ( .A1(n13127), .A2(n13311), .ZN(n10573) );
  AND2_X1 U13071 ( .A1(n10574), .A2(n10573), .ZN(n10596) );
  INV_X1 U13072 ( .A(n10596), .ZN(n10575) );
  NAND2_X1 U13073 ( .A1(n13056), .A2(n10575), .ZN(n10576) );
  OAI211_X1 U13074 ( .C1(n13096), .C2(n10602), .A(n10577), .B(n10576), .ZN(
        n10578) );
  AOI211_X1 U13075 ( .C1(n10580), .C2(n13093), .A(n10579), .B(n10578), .ZN(
        n10581) );
  INV_X1 U13076 ( .A(n10581), .ZN(P2_U3199) );
  INV_X1 U13077 ( .A(n11520), .ZN(n10591) );
  NAND2_X1 U13078 ( .A1(n10583), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10584) );
  XNOR2_X1 U13079 ( .A(n10584), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14535) );
  INV_X1 U13080 ( .A(n14535), .ZN(n10734) );
  OAI222_X1 U13081 ( .A1(n14244), .A2(n10591), .B1(n10734), .B2(P1_U3086), 
        .C1(n6650), .C2(n14245), .ZN(P1_U3340) );
  NOR2_X1 U13082 ( .A1(n15143), .A2(n10585), .ZN(n10586) );
  AOI21_X1 U13083 ( .B1(n15143), .B2(n10633), .A(n10586), .ZN(n10587) );
  OAI21_X1 U13084 ( .B1(n10588), .B2(n12965), .A(n10587), .ZN(P3_U3390) );
  INV_X1 U13085 ( .A(n11382), .ZN(n14806) );
  OAI222_X1 U13086 ( .A1(P2_U3088), .A2(n14806), .B1(n13575), .B2(n10590), 
        .C1(n10589), .C2(n13573), .ZN(P2_U3310) );
  INV_X1 U13087 ( .A(n14774), .ZN(n11394) );
  OAI222_X1 U13088 ( .A1(P2_U3088), .A2(n11394), .B1(n13575), .B2(n10591), 
        .C1(n12681), .C2(n13573), .ZN(P2_U3312) );
  OAI21_X1 U13089 ( .B1(n10593), .B2(n10594), .A(n10592), .ZN(n10619) );
  INV_X1 U13090 ( .A(n10619), .ZN(n10606) );
  XNOR2_X1 U13091 ( .A(n10595), .B(n10594), .ZN(n10597) );
  OAI21_X1 U13092 ( .B1(n10597), .B2(n13405), .A(n10596), .ZN(n10617) );
  INV_X1 U13093 ( .A(n10617), .ZN(n10598) );
  MUX2_X1 U13094 ( .A(n10599), .B(n10598), .S(n13427), .Z(n10605) );
  INV_X1 U13095 ( .A(n10671), .ZN(n10600) );
  AOI211_X1 U13096 ( .C1(n10623), .C2(n10601), .A(n13394), .B(n10600), .ZN(
        n10618) );
  OAI22_X1 U13097 ( .A1(n13376), .A2(n6760), .B1(n13412), .B2(n10602), .ZN(
        n10603) );
  AOI21_X1 U13098 ( .B1(n10618), .B2(n13422), .A(n10603), .ZN(n10604) );
  OAI211_X1 U13099 ( .C1(n13425), .C2(n10606), .A(n10605), .B(n10604), .ZN(
        P2_U3260) );
  XNOR2_X1 U13100 ( .A(n10608), .B(n10607), .ZN(n10616) );
  NAND2_X1 U13101 ( .A1(n13124), .A2(n13312), .ZN(n10610) );
  NAND2_X1 U13102 ( .A1(n13126), .A2(n13311), .ZN(n10609) );
  AND2_X1 U13103 ( .A1(n10610), .A2(n10609), .ZN(n10667) );
  INV_X1 U13104 ( .A(n10667), .ZN(n10611) );
  NAND2_X1 U13105 ( .A1(n13056), .A2(n10611), .ZN(n10612) );
  OAI211_X1 U13106 ( .C1(n13096), .C2(n10672), .A(n10613), .B(n10612), .ZN(
        n10614) );
  AOI21_X1 U13107 ( .B1(n10698), .B2(n13086), .A(n10614), .ZN(n10615) );
  OAI21_X1 U13108 ( .B1(n10616), .B2(n13088), .A(n10615), .ZN(P2_U3211) );
  AOI211_X1 U13109 ( .C1(n14440), .C2(n10619), .A(n10618), .B(n10617), .ZN(
        n10625) );
  AOI22_X1 U13110 ( .A1(n11336), .A2(n10623), .B1(n8929), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10620) );
  OAI21_X1 U13111 ( .B1(n10625), .B2(n8929), .A(n10620), .ZN(P2_U3504) );
  INV_X1 U13112 ( .A(n13548), .ZN(n11002) );
  INV_X1 U13113 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10621) );
  NOR2_X1 U13114 ( .A1(n14854), .A2(n10621), .ZN(n10622) );
  AOI21_X1 U13115 ( .B1(n11002), .B2(n10623), .A(n10622), .ZN(n10624) );
  OAI21_X1 U13116 ( .B1(n10625), .B2(n14450), .A(n10624), .ZN(P2_U3445) );
  INV_X1 U13117 ( .A(n10626), .ZN(n10627) );
  XNOR2_X1 U13118 ( .A(n12966), .B(n10627), .ZN(n10628) );
  NAND3_X1 U13119 ( .A1(n10630), .A2(n10629), .A3(n10628), .ZN(n10632) );
  INV_X1 U13120 ( .A(n15101), .ZN(n15079) );
  OR2_X1 U13121 ( .A1(n10632), .A2(n15079), .ZN(n11047) );
  INV_X1 U13122 ( .A(n12826), .ZN(n15003) );
  NAND2_X1 U13123 ( .A1(n15003), .A2(n6906), .ZN(n10635) );
  AOI22_X1 U13124 ( .A1(n10633), .A2(n15109), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15103), .ZN(n10634) );
  OAI211_X1 U13125 ( .C1(n12667), .C2(n15109), .A(n10635), .B(n10634), .ZN(
        P3_U3233) );
  INV_X1 U13126 ( .A(n10636), .ZN(n10638) );
  OAI222_X1 U13127 ( .A1(n14277), .A2(n10638), .B1(n12992), .B2(n10637), .C1(
        n12477), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U13128 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15155) );
  MUX2_X1 U13129 ( .A(n15155), .B(P3_REG1_REG_8__SCAN_IN), .S(n12442), .Z(
        n10643) );
  NAND2_X1 U13130 ( .A1(n10644), .A2(n10639), .ZN(n10641) );
  AND2_X1 U13131 ( .A1(n10641), .A2(n10640), .ZN(n10642) );
  AOI21_X1 U13132 ( .B1(n10643), .B2(n10642), .A(n12413), .ZN(n10662) );
  OAI22_X1 U13133 ( .A1(n10647), .A2(n10646), .B1(n10645), .B2(n10644), .ZN(
        n10649) );
  MUX2_X1 U13134 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12449), .Z(n12443) );
  XOR2_X1 U13135 ( .A(n12442), .B(n12443), .Z(n10648) );
  NAND2_X1 U13136 ( .A1(n10649), .A2(n10648), .ZN(n12444) );
  OAI21_X1 U13137 ( .B1(n10649), .B2(n10648), .A(n12444), .ZN(n10650) );
  NAND2_X1 U13138 ( .A1(n10650), .A2(n14991), .ZN(n10661) );
  INV_X1 U13139 ( .A(n12442), .ZN(n12414) );
  NAND2_X1 U13140 ( .A1(n12442), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n12427) );
  OR2_X1 U13141 ( .A1(n12442), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10654) );
  NAND2_X1 U13142 ( .A1(n12427), .A2(n10654), .ZN(n10655) );
  AOI21_X1 U13143 ( .B1(n10656), .B2(n10655), .A(n6567), .ZN(n10658) );
  AND2_X1 U13144 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11269) );
  AOI21_X1 U13145 ( .B1(n14984), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11269), .ZN(
        n10657) );
  OAI21_X1 U13146 ( .B1(n14997), .B2(n10658), .A(n10657), .ZN(n10659) );
  AOI21_X1 U13147 ( .B1(n12414), .B2(n14865), .A(n10659), .ZN(n10660) );
  OAI211_X1 U13148 ( .C1(n10662), .C2(n14877), .A(n10661), .B(n10660), .ZN(
        P3_U3190) );
  OAI21_X1 U13149 ( .B1(n10664), .B2(n10665), .A(n10663), .ZN(n10694) );
  INV_X1 U13150 ( .A(n10694), .ZN(n10677) );
  XNOR2_X1 U13151 ( .A(n10666), .B(n10665), .ZN(n10668) );
  OAI21_X1 U13152 ( .B1(n10668), .B2(n13405), .A(n10667), .ZN(n10692) );
  INV_X1 U13153 ( .A(n10692), .ZN(n10669) );
  MUX2_X1 U13154 ( .A(n10670), .B(n10669), .S(n13427), .Z(n10676) );
  AOI211_X1 U13155 ( .C1(n10698), .C2(n10671), .A(n13394), .B(n10712), .ZN(
        n10693) );
  INV_X1 U13156 ( .A(n10698), .ZN(n10673) );
  OAI22_X1 U13157 ( .A1(n13376), .A2(n10673), .B1(n10672), .B2(n13412), .ZN(
        n10674) );
  AOI21_X1 U13158 ( .B1(n10693), .B2(n13422), .A(n10674), .ZN(n10675) );
  OAI211_X1 U13159 ( .C1(n13425), .C2(n10677), .A(n10676), .B(n10675), .ZN(
        P2_U3259) );
  OAI211_X1 U13160 ( .C1(n10680), .C2(n10679), .A(n10678), .B(n14861), .ZN(
        n10686) );
  INV_X1 U13161 ( .A(n12390), .ZN(n12375) );
  AOI22_X1 U13162 ( .A1(n14859), .A2(n10681), .B1(n12375), .B2(n15061), .ZN(
        n10683) );
  OAI211_X1 U13163 ( .C1(n15029), .C2(n12378), .A(n10683), .B(n10682), .ZN(
        n10684) );
  AOI21_X1 U13164 ( .B1(n8203), .B2(n12392), .A(n10684), .ZN(n10685) );
  NAND2_X1 U13165 ( .A1(n10686), .A2(n10685), .ZN(P3_U3158) );
  NAND2_X1 U13166 ( .A1(n10687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10688) );
  XNOR2_X1 U13167 ( .A(n10688), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13837) );
  INV_X1 U13168 ( .A(n13837), .ZN(n11455) );
  OAI222_X1 U13169 ( .A1(n14244), .A2(n11753), .B1(n11455), .B2(P1_U3086), 
        .C1(n6707), .C2(n14245), .ZN(P1_U3337) );
  OAI222_X1 U13170 ( .A1(P3_U3151), .A2(n10691), .B1(n12992), .B2(n10690), 
        .C1(n14277), .C2(n10689), .ZN(P3_U3276) );
  AOI211_X1 U13171 ( .C1(n14440), .C2(n10694), .A(n10693), .B(n10692), .ZN(
        n10700) );
  AOI22_X1 U13172 ( .A1(n11336), .A2(n10698), .B1(n8929), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10695) );
  OAI21_X1 U13173 ( .B1(n10700), .B2(n8929), .A(n10695), .ZN(P2_U3505) );
  INV_X1 U13174 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10696) );
  NOR2_X1 U13175 ( .A1(n14854), .A2(n10696), .ZN(n10697) );
  AOI21_X1 U13176 ( .B1(n11002), .B2(n10698), .A(n10697), .ZN(n10699) );
  OAI21_X1 U13177 ( .B1(n10700), .B2(n14450), .A(n10699), .ZN(P2_U3448) );
  INV_X1 U13178 ( .A(n14818), .ZN(n10702) );
  OAI222_X1 U13179 ( .A1(P2_U3088), .A2(n10702), .B1(n13575), .B2(n11753), 
        .C1(n10701), .C2(n13573), .ZN(P2_U3309) );
  OAI21_X1 U13180 ( .B1(n10704), .B2(n10705), .A(n10703), .ZN(n10720) );
  INV_X1 U13181 ( .A(n10720), .ZN(n10717) );
  XNOR2_X1 U13182 ( .A(n10706), .B(n10705), .ZN(n10709) );
  NAND2_X1 U13183 ( .A1(n13123), .A2(n13312), .ZN(n10708) );
  NAND2_X1 U13184 ( .A1(n13125), .A2(n13311), .ZN(n10707) );
  AND2_X1 U13185 ( .A1(n10708), .A2(n10707), .ZN(n10757) );
  OAI21_X1 U13186 ( .B1(n10709), .B2(n13405), .A(n10757), .ZN(n10718) );
  INV_X1 U13187 ( .A(n10718), .ZN(n10710) );
  MUX2_X1 U13188 ( .A(n10711), .B(n10710), .S(n13427), .Z(n10716) );
  INV_X1 U13189 ( .A(n10712), .ZN(n10713) );
  AOI211_X1 U13190 ( .C1(n10766), .C2(n10713), .A(n13394), .B(n10849), .ZN(
        n10719) );
  OAI22_X1 U13191 ( .A1(n10723), .A2(n13376), .B1(n13412), .B2(n10760), .ZN(
        n10714) );
  AOI21_X1 U13192 ( .B1(n10719), .B2(n13422), .A(n10714), .ZN(n10715) );
  OAI211_X1 U13193 ( .C1(n10717), .C2(n13425), .A(n10716), .B(n10715), .ZN(
        P2_U3258) );
  AOI211_X1 U13194 ( .C1(n14440), .C2(n10720), .A(n10719), .B(n10718), .ZN(
        n10726) );
  AOI22_X1 U13195 ( .A1(n11336), .A2(n10766), .B1(n8929), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10721) );
  OAI21_X1 U13196 ( .B1(n10726), .B2(n8929), .A(n10721), .ZN(P2_U3506) );
  INV_X1 U13197 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10722) );
  OAI22_X1 U13198 ( .A1(n13548), .A2(n10723), .B1(n14854), .B2(n10722), .ZN(
        n10724) );
  INV_X1 U13199 ( .A(n10724), .ZN(n10725) );
  OAI21_X1 U13200 ( .B1(n10726), .B2(n14450), .A(n10725), .ZN(P2_U3451) );
  AOI21_X1 U13201 ( .B1(n10733), .B2(n14488), .A(n10727), .ZN(n10728) );
  NOR2_X1 U13202 ( .A1(n14535), .A2(n10728), .ZN(n10729) );
  XNOR2_X1 U13203 ( .A(n10728), .B(n14535), .ZN(n14532) );
  NOR2_X1 U13204 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14532), .ZN(n14531) );
  NOR2_X1 U13205 ( .A1(n10729), .A2(n14531), .ZN(n11013) );
  XNOR2_X1 U13206 ( .A(n11012), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11014) );
  XNOR2_X1 U13207 ( .A(n11013), .B(n11014), .ZN(n10743) );
  NAND2_X1 U13208 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13631)
         );
  INV_X1 U13209 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U13210 ( .A1(n11012), .A2(n11549), .ZN(n10730) );
  OAI21_X1 U13211 ( .B1(n11012), .B2(n11549), .A(n10730), .ZN(n10731) );
  INV_X1 U13212 ( .A(n10731), .ZN(n10738) );
  OAI21_X1 U13213 ( .B1(n14105), .B2(n10733), .A(n10732), .ZN(n10735) );
  NOR2_X1 U13214 ( .A1(n14535), .A2(n10735), .ZN(n10736) );
  XOR2_X1 U13215 ( .A(n10735), .B(n10734), .Z(n14530) );
  NOR2_X1 U13216 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14530), .ZN(n14529) );
  NOR2_X1 U13217 ( .A1(n10736), .A2(n14529), .ZN(n10737) );
  NAND2_X1 U13218 ( .A1(n10737), .A2(n10738), .ZN(n11010) );
  OAI211_X1 U13219 ( .C1(n10738), .C2(n10737), .A(n13846), .B(n11010), .ZN(
        n10739) );
  NAND2_X1 U13220 ( .A1(n13631), .A2(n10739), .ZN(n10741) );
  NOR2_X1 U13221 ( .A1(n11456), .A2(n11012), .ZN(n10740) );
  AOI211_X1 U13222 ( .C1(n13776), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n10741), 
        .B(n10740), .ZN(n10742) );
  OAI21_X1 U13223 ( .B1(n10743), .B2(n14533), .A(n10742), .ZN(P1_U3259) );
  INV_X1 U13224 ( .A(n11772), .ZN(n12227) );
  OAI222_X1 U13225 ( .A1(n11405), .A2(P2_U3088), .B1(n13575), .B2(n12227), 
        .C1(n10744), .C2(n13573), .ZN(P2_U3308) );
  NAND2_X1 U13226 ( .A1(n12399), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10745) );
  OAI21_X1 U13227 ( .B1(n10746), .B2(n12399), .A(n10745), .ZN(P3_U3521) );
  INV_X1 U13228 ( .A(n10747), .ZN(n10748) );
  AOI21_X1 U13229 ( .B1(n10750), .B2(n10749), .A(n10748), .ZN(n10756) );
  OAI21_X1 U13230 ( .B1(n13095), .B2(n10752), .A(n10751), .ZN(n10754) );
  OAI22_X1 U13231 ( .A1(n13097), .A2(n10937), .B1(n13096), .B2(n10854), .ZN(
        n10753) );
  AOI211_X1 U13232 ( .C1(n10853), .C2(n13086), .A(n10754), .B(n10753), .ZN(
        n10755) );
  OAI21_X1 U13233 ( .B1(n10756), .B2(n13088), .A(n10755), .ZN(P2_U3193) );
  NAND2_X1 U13234 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13163) );
  INV_X1 U13235 ( .A(n10757), .ZN(n10758) );
  NAND2_X1 U13236 ( .A1(n13056), .A2(n10758), .ZN(n10759) );
  OAI211_X1 U13237 ( .C1(n13096), .C2(n10760), .A(n13163), .B(n10759), .ZN(
        n10765) );
  XNOR2_X1 U13238 ( .A(n10762), .B(n10761), .ZN(n10763) );
  NOR2_X1 U13239 ( .A1(n10763), .A2(n13088), .ZN(n10764) );
  AOI211_X1 U13240 ( .C1(n10766), .C2(n13086), .A(n10765), .B(n10764), .ZN(
        n10767) );
  INV_X1 U13241 ( .A(n10767), .ZN(P2_U3185) );
  INV_X1 U13242 ( .A(n10768), .ZN(n10769) );
  OAI222_X1 U13243 ( .A1(P3_U3151), .A2(n10771), .B1(n12992), .B2(n10770), 
        .C1(n14277), .C2(n10769), .ZN(P3_U3275) );
  INV_X1 U13244 ( .A(n10772), .ZN(n10774) );
  NAND2_X1 U13245 ( .A1(n10776), .A2(n11085), .ZN(n10778) );
  INV_X2 U13246 ( .A(n12160), .ZN(n11774) );
  AOI22_X1 U13247 ( .A1(n11774), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11773), 
        .B2(n13790), .ZN(n10777) );
  OAI22_X1 U13248 ( .A1(n9756), .A2(n12011), .B1(n14634), .B2(n9728), .ZN(
        n10800) );
  OAI22_X1 U13249 ( .A1(n12011), .A2(n9728), .B1(n9737), .B2(n14634), .ZN(
        n10779) );
  XOR2_X1 U13250 ( .A(n12232), .B(n10779), .Z(n10801) );
  XOR2_X1 U13251 ( .A(n10802), .B(n10801), .Z(n10780) );
  NAND2_X1 U13252 ( .A1(n10780), .A2(n14470), .ZN(n10791) );
  NAND2_X1 U13253 ( .A1(n13731), .A2(n14100), .ZN(n10788) );
  NAND2_X1 U13254 ( .A1(n12154), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10786) );
  OR2_X1 U13255 ( .A1(n12167), .A2(n14698), .ZN(n10785) );
  AND2_X1 U13256 ( .A1(n10781), .A2(n10824), .ZN(n10782) );
  NOR2_X1 U13257 ( .A1(n10781), .A2(n10824), .ZN(n10815) );
  OR2_X1 U13258 ( .A1(n10782), .A2(n10815), .ZN(n10877) );
  OR2_X1 U13259 ( .A1(n9744), .A2(n10877), .ZN(n10784) );
  NAND2_X1 U13260 ( .A1(n13730), .A2(n13691), .ZN(n10787) );
  AND2_X1 U13261 ( .A1(n10788), .A2(n10787), .ZN(n14632) );
  NAND2_X1 U13262 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13782) );
  OAI21_X1 U13263 ( .B1(n13712), .B2(n14632), .A(n13782), .ZN(n10789) );
  AOI21_X1 U13264 ( .B1(n7265), .B2(n14475), .A(n10789), .ZN(n10790) );
  OAI211_X1 U13265 ( .C1(n14479), .C2(n11127), .A(n10791), .B(n10790), .ZN(
        P1_U3230) );
  AOI21_X1 U13266 ( .B1(n10793), .B2(n10792), .A(n6571), .ZN(n10799) );
  INV_X1 U13267 ( .A(n12378), .ZN(n14860) );
  OAI22_X1 U13268 ( .A1(n12395), .A2(n15039), .B1(n12390), .B2(n15045), .ZN(
        n10794) );
  AOI211_X1 U13269 ( .C1(n14860), .C2(n11052), .A(n10795), .B(n10794), .ZN(
        n10798) );
  NAND2_X1 U13270 ( .A1(n12392), .A2(n10796), .ZN(n10797) );
  OAI211_X1 U13271 ( .C1(n10799), .C2(n12382), .A(n10798), .B(n10797), .ZN(
        P3_U3170) );
  NAND2_X1 U13272 ( .A1(n10803), .A2(n11085), .ZN(n10806) );
  AOI22_X1 U13273 ( .A1(n11774), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11773), 
        .B2(n10804), .ZN(n10805) );
  NAND2_X1 U13274 ( .A1(n10806), .A2(n10805), .ZN(n14641) );
  AOI22_X1 U13275 ( .A1(n11928), .A2(n13730), .B1(n11863), .B2(n14641), .ZN(
        n10811) );
  NAND2_X1 U13276 ( .A1(n14641), .A2(n11929), .ZN(n10808) );
  NAND2_X1 U13277 ( .A1(n11863), .A2(n13730), .ZN(n10807) );
  NAND2_X1 U13278 ( .A1(n10808), .A2(n10807), .ZN(n10809) );
  XNOR2_X1 U13279 ( .A(n10809), .B(n11652), .ZN(n10810) );
  OR2_X1 U13280 ( .A1(n10811), .A2(n10810), .ZN(n10948) );
  INV_X1 U13281 ( .A(n10948), .ZN(n10812) );
  AND2_X1 U13282 ( .A1(n10811), .A2(n10810), .ZN(n10949) );
  NOR2_X1 U13283 ( .A1(n10812), .A2(n10949), .ZN(n10813) );
  XNOR2_X1 U13284 ( .A(n10950), .B(n10813), .ZN(n10814) );
  NAND2_X1 U13285 ( .A1(n10814), .A2(n14470), .ZN(n10827) );
  OR2_X1 U13286 ( .A1(n12011), .A2(n13903), .ZN(n10823) );
  NAND2_X1 U13287 ( .A1(n12154), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10821) );
  OR2_X1 U13288 ( .A1(n12167), .A2(n14700), .ZN(n10820) );
  NAND2_X1 U13289 ( .A1(n10815), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10968) );
  OR2_X1 U13290 ( .A1(n10815), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10816) );
  NAND2_X1 U13291 ( .A1(n10968), .A2(n10816), .ZN(n14572) );
  OR2_X1 U13292 ( .A1(n9744), .A2(n14572), .ZN(n10819) );
  OR2_X1 U13293 ( .A1(n11923), .A2(n10817), .ZN(n10818) );
  NAND4_X1 U13294 ( .A1(n10821), .A2(n10820), .A3(n10819), .A4(n10818), .ZN(
        n13729) );
  NAND2_X1 U13295 ( .A1(n13729), .A2(n13691), .ZN(n10822) );
  AND2_X1 U13296 ( .A1(n10823), .A2(n10822), .ZN(n10892) );
  OAI22_X1 U13297 ( .A1(n13712), .A2(n10892), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10824), .ZN(n10825) );
  AOI21_X1 U13298 ( .B1(n14641), .B2(n14475), .A(n10825), .ZN(n10826) );
  OAI211_X1 U13299 ( .C1(n14479), .C2(n10877), .A(n10827), .B(n10826), .ZN(
        P1_U3227) );
  XNOR2_X1 U13300 ( .A(n10828), .B(n10829), .ZN(n10995) );
  XNOR2_X1 U13301 ( .A(n10830), .B(n10829), .ZN(n10833) );
  OAI22_X1 U13302 ( .A1(n10831), .A2(n13404), .B1(n10912), .B2(n13408), .ZN(
        n10832) );
  AOI21_X1 U13303 ( .B1(n10833), .B2(n13352), .A(n10832), .ZN(n10834) );
  OAI21_X1 U13304 ( .B1(n10995), .B2(n13355), .A(n10834), .ZN(n10996) );
  NAND2_X1 U13305 ( .A1(n10996), .A2(n13427), .ZN(n10839) );
  AOI211_X1 U13306 ( .C1(n11003), .C2(n10850), .A(n13394), .B(n6945), .ZN(
        n10997) );
  INV_X1 U13307 ( .A(n11003), .ZN(n10917) );
  NOR2_X1 U13308 ( .A1(n10917), .A2(n13376), .ZN(n10837) );
  OAI22_X1 U13309 ( .A1(n13427), .A2(n10835), .B1(n10911), .B2(n13412), .ZN(
        n10836) );
  AOI211_X1 U13310 ( .C1(n10997), .C2(n13422), .A(n10837), .B(n10836), .ZN(
        n10838) );
  OAI211_X1 U13311 ( .C1(n10995), .C2(n13367), .A(n10839), .B(n10838), .ZN(
        P2_U3256) );
  NAND2_X1 U13312 ( .A1(n10840), .A2(n10843), .ZN(n10841) );
  NAND2_X1 U13313 ( .A1(n10842), .A2(n10841), .ZN(n14839) );
  XNOR2_X1 U13314 ( .A(n10844), .B(n10843), .ZN(n10847) );
  OR2_X1 U13315 ( .A1(n14839), .A2(n13355), .ZN(n10846) );
  AOI22_X1 U13316 ( .A1(n13311), .A2(n13124), .B1(n13122), .B2(n13312), .ZN(
        n10845) );
  OAI211_X1 U13317 ( .C1(n13405), .C2(n10847), .A(n10846), .B(n10845), .ZN(
        n14843) );
  MUX2_X1 U13318 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n14843), .S(n13427), .Z(
        n10848) );
  INV_X1 U13319 ( .A(n10848), .ZN(n10857) );
  INV_X1 U13320 ( .A(n10849), .ZN(n10852) );
  INV_X1 U13321 ( .A(n10850), .ZN(n10851) );
  AOI211_X1 U13322 ( .C1(n10853), .C2(n10852), .A(n13394), .B(n10851), .ZN(
        n14840) );
  OAI22_X1 U13323 ( .A1(n14842), .A2(n13376), .B1(n10854), .B2(n13412), .ZN(
        n10855) );
  AOI21_X1 U13324 ( .B1(n14840), .B2(n13422), .A(n10855), .ZN(n10856) );
  OAI211_X1 U13325 ( .C1(n14839), .C2(n13367), .A(n10857), .B(n10856), .ZN(
        P2_U3257) );
  INV_X1 U13326 ( .A(n10858), .ZN(n10861) );
  NAND3_X1 U13327 ( .A1(n10861), .A2(n10860), .A3(n10859), .ZN(n13907) );
  AOI21_X1 U13328 ( .B1(n14595), .B2(n10862), .A(n14585), .ZN(n10868) );
  INV_X2 U13329 ( .A(n14562), .ZN(n14599) );
  OAI22_X1 U13330 ( .A1(n14599), .A2(n10864), .B1(n10863), .B2(n14555), .ZN(
        n10866) );
  AOI21_X1 U13331 ( .B1(n13930), .B2(n14092), .A(n12184), .ZN(n10865) );
  AOI211_X1 U13332 ( .C1(n14599), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10866), .B(
        n10865), .ZN(n10867) );
  OAI21_X1 U13333 ( .B1(n10868), .B2(n11138), .A(n10867), .ZN(P1_U3293) );
  NAND2_X1 U13334 ( .A1(n13734), .A2(n11992), .ZN(n10869) );
  INV_X1 U13335 ( .A(n14582), .ZN(n14587) );
  NAND2_X1 U13336 ( .A1(n14588), .A2(n14587), .ZN(n10871) );
  NAND2_X1 U13337 ( .A1(n10882), .A2(n14616), .ZN(n12001) );
  INV_X1 U13338 ( .A(n12003), .ZN(n12187) );
  NAND2_X1 U13339 ( .A1(n11149), .A2(n12187), .ZN(n10872) );
  NAND2_X1 U13340 ( .A1(n12006), .A2(n14623), .ZN(n12007) );
  NAND2_X1 U13341 ( .A1(n12011), .A2(n14634), .ZN(n10873) );
  INV_X1 U13342 ( .A(n13730), .ZN(n10874) );
  NAND2_X1 U13343 ( .A1(n14641), .A2(n10874), .ZN(n11068) );
  NAND2_X1 U13344 ( .A1(n11068), .A2(n10875), .ZN(n12188) );
  INV_X1 U13345 ( .A(n12188), .ZN(n10891) );
  XNOR2_X1 U13346 ( .A(n11060), .B(n10891), .ZN(n14645) );
  NOR2_X2 U13347 ( .A1(n14590), .A2(n14589), .ZN(n14594) );
  NAND2_X1 U13348 ( .A1(n14594), .A2(n14623), .ZN(n11157) );
  AOI21_X1 U13349 ( .B1(n11125), .B2(n14641), .A(n14575), .ZN(n10876) );
  AND2_X1 U13350 ( .A1(n10876), .A2(n14576), .ZN(n14643) );
  INV_X1 U13351 ( .A(n14641), .ZN(n10878) );
  OAI22_X1 U13352 ( .A1(n14088), .A2(n10878), .B1(n14555), .B2(n10877), .ZN(
        n10879) );
  AOI21_X1 U13353 ( .B1(n14595), .B2(n14643), .A(n10879), .ZN(n10897) );
  NOR2_X1 U13354 ( .A1(n11139), .A2(n11138), .ZN(n11989) );
  NAND2_X1 U13355 ( .A1(n13734), .A2(n6591), .ZN(n10880) );
  NAND2_X1 U13356 ( .A1(n11989), .A2(n10880), .ZN(n11988) );
  NAND2_X1 U13357 ( .A1(n10881), .A2(n11992), .ZN(n11986) );
  NAND2_X1 U13358 ( .A1(n11988), .A2(n11986), .ZN(n14581) );
  NAND2_X1 U13359 ( .A1(n14581), .A2(n14582), .ZN(n10884) );
  NAND2_X1 U13360 ( .A1(n10882), .A2(n14589), .ZN(n10883) );
  NAND2_X1 U13361 ( .A1(n10884), .A2(n10883), .ZN(n11150) );
  NAND2_X1 U13362 ( .A1(n11150), .A2(n12003), .ZN(n11152) );
  NAND2_X1 U13363 ( .A1(n12006), .A2(n10885), .ZN(n10886) );
  NAND2_X1 U13364 ( .A1(n11152), .A2(n10886), .ZN(n11123) );
  INV_X1 U13365 ( .A(n12186), .ZN(n10887) );
  NAND2_X1 U13366 ( .A1(n11123), .A2(n10887), .ZN(n10889) );
  NAND2_X1 U13367 ( .A1(n7265), .A2(n12011), .ZN(n10888) );
  OAI21_X1 U13368 ( .B1(n10891), .B2(n10890), .A(n11069), .ZN(n10894) );
  INV_X1 U13369 ( .A(n10892), .ZN(n10893) );
  AOI21_X1 U13370 ( .B1(n10894), .B2(n14625), .A(n10893), .ZN(n14648) );
  MUX2_X1 U13371 ( .A(n10895), .B(n14648), .S(n14562), .Z(n10896) );
  OAI211_X1 U13372 ( .C1(n14645), .C2(n14092), .A(n10897), .B(n10896), .ZN(
        P1_U3288) );
  XOR2_X1 U13373 ( .A(n10899), .B(n10898), .Z(n10904) );
  INV_X1 U13374 ( .A(n11027), .ZN(n15028) );
  AOI22_X1 U13375 ( .A1(n14859), .A2(n10900), .B1(n12375), .B2(n15060), .ZN(
        n10901) );
  NAND2_X1 U13376 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n14884) );
  OAI211_X1 U13377 ( .C1(n15028), .C2(n12378), .A(n10901), .B(n14884), .ZN(
        n10902) );
  AOI21_X1 U13378 ( .B1(n15035), .B2(n12392), .A(n10902), .ZN(n10903) );
  OAI21_X1 U13379 ( .B1(n10904), .B2(n12382), .A(n10903), .ZN(P3_U3167) );
  INV_X1 U13380 ( .A(n10905), .ZN(n10906) );
  OAI222_X1 U13381 ( .A1(n11024), .A2(P3_U3151), .B1(n14277), .B2(n10906), 
        .C1(n12626), .C2(n12992), .ZN(P3_U3274) );
  OAI21_X1 U13382 ( .B1(n10909), .B2(n10908), .A(n10907), .ZN(n10910) );
  NAND2_X1 U13383 ( .A1(n10910), .A2(n13093), .ZN(n10916) );
  INV_X1 U13384 ( .A(n13095), .ZN(n11564) );
  NAND2_X1 U13385 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14729) );
  INV_X1 U13386 ( .A(n14729), .ZN(n10914) );
  OAI22_X1 U13387 ( .A1(n13097), .A2(n10912), .B1(n13096), .B2(n10911), .ZN(
        n10913) );
  AOI211_X1 U13388 ( .C1(n11564), .C2(n13123), .A(n10914), .B(n10913), .ZN(
        n10915) );
  OAI211_X1 U13389 ( .C1(n10917), .C2(n13102), .A(n10916), .B(n10915), .ZN(
        P2_U3203) );
  XNOR2_X1 U13390 ( .A(n10919), .B(n10918), .ZN(n10924) );
  OAI21_X1 U13391 ( .B1(n13095), .B2(n10937), .A(n10920), .ZN(n10922) );
  OAI22_X1 U13392 ( .A1(n13097), .A2(n11351), .B1(n13096), .B2(n10941), .ZN(
        n10921) );
  AOI211_X1 U13393 ( .C1(n10945), .C2(n13086), .A(n10922), .B(n10921), .ZN(
        n10923) );
  OAI21_X1 U13394 ( .B1(n10924), .B2(n13088), .A(n10923), .ZN(P2_U3189) );
  INV_X1 U13395 ( .A(n10925), .ZN(n11046) );
  OAI211_X1 U13396 ( .C1(n10928), .C2(n10927), .A(n10926), .B(n14861), .ZN(
        n10933) );
  OAI22_X1 U13397 ( .A1(n12395), .A2(n10929), .B1(n12390), .B2(n15047), .ZN(
        n10930) );
  AOI211_X1 U13398 ( .C1(n14860), .C2(n12410), .A(n10931), .B(n10930), .ZN(
        n10932) );
  OAI211_X1 U13399 ( .C1(n11046), .C2(n11503), .A(n10933), .B(n10932), .ZN(
        P3_U3179) );
  XNOR2_X1 U13400 ( .A(n10934), .B(n10935), .ZN(n14847) );
  XNOR2_X1 U13401 ( .A(n10936), .B(n10935), .ZN(n10939) );
  OAI22_X1 U13402 ( .A1(n10937), .A2(n13404), .B1(n11351), .B2(n13408), .ZN(
        n10938) );
  AOI21_X1 U13403 ( .B1(n10939), .B2(n13352), .A(n10938), .ZN(n10940) );
  OAI21_X1 U13404 ( .B1(n14847), .B2(n13355), .A(n10940), .ZN(n14850) );
  NAND2_X1 U13405 ( .A1(n14850), .A2(n13356), .ZN(n10947) );
  INV_X1 U13406 ( .A(n13376), .ZN(n13416) );
  OAI22_X1 U13407 ( .A1(n13427), .A2(n10942), .B1(n10941), .B2(n13412), .ZN(
        n10944) );
  OAI211_X1 U13408 ( .C1(n6945), .C2(n6944), .A(n13420), .B(n11239), .ZN(
        n14848) );
  NOR2_X1 U13409 ( .A1(n14848), .A2(n13269), .ZN(n10943) );
  AOI211_X1 U13410 ( .C1(n13416), .C2(n10945), .A(n10944), .B(n10943), .ZN(
        n10946) );
  OAI211_X1 U13411 ( .C1(n14847), .C2(n13367), .A(n10947), .B(n10946), .ZN(
        P2_U3255) );
  NAND2_X1 U13412 ( .A1(n10951), .A2(n11085), .ZN(n10953) );
  AOI22_X1 U13413 ( .A1(n11774), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11773), 
        .B2(n13807), .ZN(n10952) );
  NAND2_X1 U13414 ( .A1(n10953), .A2(n10952), .ZN(n14651) );
  AOI22_X1 U13415 ( .A1(n11863), .A2(n14651), .B1(n11928), .B2(n13729), .ZN(
        n10958) );
  NAND2_X1 U13416 ( .A1(n14651), .A2(n11929), .ZN(n10955) );
  NAND2_X1 U13417 ( .A1(n11863), .A2(n13729), .ZN(n10954) );
  NAND2_X1 U13418 ( .A1(n10955), .A2(n10954), .ZN(n10956) );
  XNOR2_X1 U13419 ( .A(n10956), .B(n11652), .ZN(n10957) );
  XOR2_X1 U13420 ( .A(n10958), .B(n10957), .Z(n13689) );
  NAND2_X1 U13421 ( .A1(n13690), .A2(n13689), .ZN(n13688) );
  INV_X1 U13422 ( .A(n10957), .ZN(n10960) );
  INV_X1 U13423 ( .A(n10958), .ZN(n10959) );
  NAND2_X1 U13424 ( .A1(n10960), .A2(n10959), .ZN(n10961) );
  NAND2_X1 U13425 ( .A1(n10962), .A2(n11085), .ZN(n10965) );
  AOI22_X1 U13426 ( .A1(n11774), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11773), 
        .B2(n10963), .ZN(n10964) );
  NAND2_X1 U13427 ( .A1(n10965), .A2(n10964), .ZN(n12034) );
  NAND2_X1 U13428 ( .A1(n12154), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10974) );
  OR2_X1 U13429 ( .A1(n12167), .A2(n10966), .ZN(n10973) );
  NAND2_X1 U13430 ( .A1(n10968), .A2(n10967), .ZN(n10969) );
  NAND2_X1 U13431 ( .A1(n10981), .A2(n10969), .ZN(n11065) );
  OR2_X1 U13432 ( .A1(n9744), .A2(n11065), .ZN(n10972) );
  OR2_X1 U13433 ( .A1(n11923), .A2(n10970), .ZN(n10971) );
  NAND4_X1 U13434 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n13728) );
  AOI22_X1 U13435 ( .A1(n12034), .A2(n11929), .B1(n11863), .B2(n13728), .ZN(
        n10975) );
  XNOR2_X1 U13436 ( .A(n10975), .B(n12232), .ZN(n11252) );
  INV_X1 U13437 ( .A(n13728), .ZN(n11259) );
  NOR2_X1 U13438 ( .A1(n9756), .A2(n11259), .ZN(n10976) );
  AOI21_X1 U13439 ( .B1(n12034), .B2(n11863), .A(n10976), .ZN(n11253) );
  XNOR2_X1 U13440 ( .A(n11252), .B(n11253), .ZN(n10977) );
  NAND2_X1 U13441 ( .A1(n10978), .A2(n10977), .ZN(n11256) );
  OAI211_X1 U13442 ( .C1(n10978), .C2(n10977), .A(n11256), .B(n14470), .ZN(
        n10994) );
  NAND2_X1 U13443 ( .A1(n13729), .A2(n14100), .ZN(n10989) );
  NAND2_X1 U13444 ( .A1(n12154), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10987) );
  OR2_X1 U13445 ( .A1(n12167), .A2(n10979), .ZN(n10986) );
  NAND2_X1 U13446 ( .A1(n10981), .A2(n10980), .ZN(n10982) );
  NAND2_X1 U13447 ( .A1(n11090), .A2(n10982), .ZN(n14554) );
  OR2_X1 U13448 ( .A1(n9744), .A2(n14554), .ZN(n10985) );
  OR2_X1 U13449 ( .A1(n11923), .A2(n10983), .ZN(n10984) );
  NAND4_X1 U13450 ( .A1(n10987), .A2(n10986), .A3(n10985), .A4(n10984), .ZN(
        n13727) );
  NAND2_X1 U13451 ( .A1(n13727), .A2(n13854), .ZN(n10988) );
  AND2_X1 U13452 ( .A1(n10989), .A2(n10988), .ZN(n11072) );
  OAI21_X1 U13453 ( .B1(n13712), .B2(n11072), .A(n10990), .ZN(n10992) );
  NOR2_X1 U13454 ( .A1(n14479), .A2(n11065), .ZN(n10991) );
  AOI211_X1 U13455 ( .C1(n12034), .C2(n14475), .A(n10992), .B(n10991), .ZN(
        n10993) );
  NAND2_X1 U13456 ( .A1(n10994), .A2(n10993), .ZN(P1_U3213) );
  INV_X1 U13457 ( .A(n10995), .ZN(n10998) );
  AOI211_X1 U13458 ( .C1(n9151), .C2(n10998), .A(n10997), .B(n10996), .ZN(
        n11005) );
  AOI22_X1 U13459 ( .A1(n11003), .A2(n11336), .B1(n8929), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10999) );
  OAI21_X1 U13460 ( .B1(n11005), .B2(n8929), .A(n10999), .ZN(P2_U3508) );
  INV_X1 U13461 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11000) );
  NOR2_X1 U13462 ( .A1(n14854), .A2(n11000), .ZN(n11001) );
  AOI21_X1 U13463 ( .B1(n11003), .B2(n11002), .A(n11001), .ZN(n11004) );
  OAI21_X1 U13464 ( .B1(n11005), .B2(n14450), .A(n11004), .ZN(P2_U3457) );
  OAI222_X1 U13465 ( .A1(n14244), .A2(n11794), .B1(n11977), .B2(P1_U3086), 
        .C1(n7077), .C2(n14245), .ZN(P1_U3335) );
  INV_X1 U13466 ( .A(n11006), .ZN(n11009) );
  OAI22_X1 U13467 ( .A1(n11007), .A2(P3_U3151), .B1(SI_22_), .B2(n14275), .ZN(
        n11008) );
  AOI21_X1 U13468 ( .B1(n11009), .B2(n14288), .A(n11008), .ZN(P3_U3273) );
  OAI21_X1 U13469 ( .B1(n11549), .B2(n11012), .A(n11010), .ZN(n11443) );
  XNOR2_X1 U13470 ( .A(n11743), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n11441) );
  XNOR2_X1 U13471 ( .A(n11443), .B(n11441), .ZN(n11011) );
  NAND2_X1 U13472 ( .A1(n11011), .A2(n13846), .ZN(n11021) );
  NAND2_X1 U13473 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13643)
         );
  INV_X1 U13474 ( .A(n11012), .ZN(n11687) );
  AOI22_X1 U13475 ( .A1(n11687), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n11014), 
        .B2(n11013), .ZN(n11016) );
  XNOR2_X1 U13476 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n11743), .ZN(n11015) );
  AOI21_X1 U13477 ( .B1(n11016), .B2(n11015), .A(n14533), .ZN(n11017) );
  NAND2_X1 U13478 ( .A1(n11017), .A2(n11447), .ZN(n11018) );
  NAND2_X1 U13479 ( .A1(n13643), .A2(n11018), .ZN(n11019) );
  AOI21_X1 U13480 ( .B1(n13776), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11019), 
        .ZN(n11020) );
  OAI211_X1 U13481 ( .C1(n11456), .C2(n11448), .A(n11021), .B(n11020), .ZN(
        P1_U3260) );
  XNOR2_X1 U13482 ( .A(n11022), .B(n11023), .ZN(n15129) );
  OR2_X1 U13483 ( .A1(n15101), .A2(n11024), .ZN(n15106) );
  INV_X1 U13484 ( .A(n15106), .ZN(n15097) );
  INV_X1 U13485 ( .A(n12586), .ZN(n11033) );
  XNOR2_X1 U13486 ( .A(n11025), .B(n11026), .ZN(n11030) );
  INV_X1 U13487 ( .A(n15044), .ZN(n15084) );
  AOI22_X1 U13488 ( .A1(n15084), .A2(n11027), .B1(n12409), .B2(n15081), .ZN(
        n11028) );
  OAI21_X1 U13489 ( .B1(n15129), .B2(n15094), .A(n11028), .ZN(n11029) );
  AOI21_X1 U13490 ( .B1(n11030), .B2(n15089), .A(n11029), .ZN(n15130) );
  MUX2_X1 U13491 ( .A(n10526), .B(n15130), .S(n15109), .Z(n11032) );
  NOR2_X1 U13492 ( .A1(n11038), .A2(n15076), .ZN(n15132) );
  AOI22_X1 U13493 ( .A1(n15070), .A2(n15132), .B1(n15103), .B2(n11034), .ZN(
        n11031) );
  OAI211_X1 U13494 ( .C1(n15129), .C2(n11033), .A(n11032), .B(n11031), .ZN(
        P3_U3226) );
  INV_X1 U13495 ( .A(n11034), .ZN(n11043) );
  OAI211_X1 U13496 ( .C1(n11037), .C2(n11036), .A(n11035), .B(n14861), .ZN(
        n11042) );
  OAI22_X1 U13497 ( .A1(n12395), .A2(n11038), .B1(n12390), .B2(n15028), .ZN(
        n11039) );
  AOI211_X1 U13498 ( .C1(n14860), .C2(n12409), .A(n11040), .B(n11039), .ZN(
        n11041) );
  OAI211_X1 U13499 ( .C1(n11043), .C2(n11503), .A(n11042), .B(n11041), .ZN(
        P3_U3153) );
  XNOR2_X1 U13500 ( .A(n6408), .B(n11048), .ZN(n15128) );
  NAND2_X1 U13501 ( .A1(n11045), .A2(n14410), .ZN(n15125) );
  OAI22_X1 U13502 ( .A1(n11047), .A2(n15125), .B1(n11046), .B2(n15078), .ZN(
        n11057) );
  NAND2_X1 U13503 ( .A1(n11049), .A2(n11048), .ZN(n11050) );
  NAND3_X1 U13504 ( .A1(n11051), .A2(n15089), .A3(n11050), .ZN(n11055) );
  AOI22_X1 U13505 ( .A1(n15081), .A2(n12410), .B1(n11052), .B2(n15084), .ZN(
        n11054) );
  INV_X1 U13506 ( .A(n15094), .ZN(n15049) );
  NAND2_X1 U13507 ( .A1(n15128), .A2(n15049), .ZN(n11053) );
  NAND3_X1 U13508 ( .A1(n11055), .A2(n11054), .A3(n11053), .ZN(n15126) );
  MUX2_X1 U13509 ( .A(n15126), .B(P3_REG2_REG_6__SCAN_IN), .S(n15005), .Z(
        n11056) );
  AOI211_X1 U13510 ( .C1(n15128), .C2(n12586), .A(n11057), .B(n11056), .ZN(
        n11058) );
  INV_X1 U13511 ( .A(n11058), .ZN(P3_U3227) );
  OAI222_X1 U13512 ( .A1(P2_U3088), .A2(n11059), .B1(n13575), .B2(n11794), 
        .C1(n12660), .C2(n13573), .ZN(P2_U3307) );
  XNOR2_X1 U13513 ( .A(n14651), .B(n13729), .ZN(n14566) );
  INV_X1 U13514 ( .A(n14566), .ZN(n11061) );
  NAND2_X1 U13515 ( .A1(n14567), .A2(n11061), .ZN(n11063) );
  OR2_X1 U13516 ( .A1(n14651), .A2(n13729), .ZN(n11062) );
  XNOR2_X1 U13517 ( .A(n12034), .B(n13728), .ZN(n12189) );
  INV_X1 U13518 ( .A(n12189), .ZN(n11078) );
  XNOR2_X1 U13519 ( .A(n11079), .B(n11078), .ZN(n14659) );
  NAND2_X1 U13520 ( .A1(n11985), .A2(n14559), .ZN(n11981) );
  INV_X1 U13521 ( .A(n11981), .ZN(n11064) );
  AND2_X1 U13522 ( .A1(n14562), .A2(n11064), .ZN(n14577) );
  INV_X1 U13523 ( .A(n12034), .ZN(n14662) );
  NAND2_X1 U13524 ( .A1(n14574), .A2(n14662), .ZN(n14547) );
  OAI211_X1 U13525 ( .C1(n14574), .C2(n14662), .A(n14591), .B(n14547), .ZN(
        n14660) );
  INV_X1 U13526 ( .A(n14555), .ZN(n14586) );
  INV_X1 U13527 ( .A(n11065), .ZN(n11066) );
  AOI22_X1 U13528 ( .A1(n14585), .A2(n12034), .B1(n14586), .B2(n11066), .ZN(
        n11067) );
  OAI21_X1 U13529 ( .B1(n14109), .B2(n14660), .A(n11067), .ZN(n11076) );
  INV_X1 U13530 ( .A(n13729), .ZN(n11070) );
  NAND2_X1 U13531 ( .A1(n14651), .A2(n11070), .ZN(n11071) );
  NAND2_X1 U13532 ( .A1(n14564), .A2(n11071), .ZN(n11098) );
  XNOR2_X1 U13533 ( .A(n11098), .B(n11078), .ZN(n11074) );
  INV_X1 U13534 ( .A(n14568), .ZN(n14675) );
  NAND2_X1 U13535 ( .A1(n14659), .A2(n14675), .ZN(n11073) );
  OAI211_X1 U13536 ( .C1(n14635), .C2(n11074), .A(n11073), .B(n11072), .ZN(
        n14664) );
  MUX2_X1 U13537 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n14664), .S(n14562), .Z(
        n11075) );
  AOI211_X1 U13538 ( .C1(n14659), .C2(n14577), .A(n11076), .B(n11075), .ZN(
        n11077) );
  INV_X1 U13539 ( .A(n11077), .ZN(P1_U3286) );
  OR2_X1 U13540 ( .A1(n12034), .A2(n13728), .ZN(n11080) );
  NAND2_X1 U13541 ( .A1(n11081), .A2(n11085), .ZN(n11084) );
  AOI22_X1 U13542 ( .A1(n11774), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11773), 
        .B2(n11082), .ZN(n11083) );
  XNOR2_X1 U13543 ( .A(n14666), .B(n13727), .ZN(n12191) );
  NAND2_X1 U13544 ( .A1(n11086), .A2(n11085), .ZN(n11089) );
  AOI22_X1 U13545 ( .A1(n11087), .A2(n11773), .B1(n11774), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n11088) );
  NAND2_X1 U13546 ( .A1(n12154), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11096) );
  OR2_X1 U13547 ( .A1(n12167), .A2(n14704), .ZN(n11095) );
  INV_X1 U13548 ( .A(n11106), .ZN(n11092) );
  NAND2_X1 U13549 ( .A1(n11090), .A2(n11435), .ZN(n11091) );
  NAND2_X1 U13550 ( .A1(n11092), .A2(n11091), .ZN(n11434) );
  OR2_X1 U13551 ( .A1(n9744), .A2(n11434), .ZN(n11094) );
  OR2_X1 U13552 ( .A1(n11923), .A2(n11115), .ZN(n11093) );
  NAND4_X1 U13553 ( .A1(n11096), .A2(n11095), .A3(n11094), .A4(n11093), .ZN(
        n13726) );
  INV_X1 U13554 ( .A(n13726), .ZN(n11427) );
  XNOR2_X1 U13555 ( .A(n12046), .B(n11427), .ZN(n12193) );
  XNOR2_X1 U13556 ( .A(n11161), .B(n12193), .ZN(n14673) );
  INV_X1 U13557 ( .A(n14673), .ZN(n11122) );
  OR2_X1 U13558 ( .A1(n12034), .A2(n11259), .ZN(n11097) );
  NAND2_X1 U13559 ( .A1(n11098), .A2(n11097), .ZN(n11100) );
  NAND2_X1 U13560 ( .A1(n12034), .A2(n11259), .ZN(n11099) );
  INV_X1 U13561 ( .A(n13727), .ZN(n11101) );
  OR2_X1 U13562 ( .A1(n14666), .A2(n11101), .ZN(n11102) );
  NAND2_X1 U13563 ( .A1(n11103), .A2(n12193), .ZN(n11104) );
  NAND2_X1 U13564 ( .A1(n11206), .A2(n11104), .ZN(n11105) );
  NAND2_X1 U13565 ( .A1(n11105), .A2(n14625), .ZN(n11114) );
  NAND2_X1 U13566 ( .A1(n13727), .A2(n14100), .ZN(n11113) );
  NAND2_X1 U13567 ( .A1(n12154), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11111) );
  OR2_X1 U13568 ( .A1(n12167), .A2(n14707), .ZN(n11110) );
  NAND2_X1 U13569 ( .A1(n11106), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11175) );
  OR2_X1 U13570 ( .A1(n11106), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11107) );
  NAND2_X1 U13571 ( .A1(n11175), .A2(n11107), .ZN(n13596) );
  OR2_X1 U13572 ( .A1(n9744), .A2(n13596), .ZN(n11109) );
  OR2_X1 U13573 ( .A1(n11923), .A2(n11215), .ZN(n11108) );
  NAND4_X1 U13574 ( .A1(n11111), .A2(n11110), .A3(n11109), .A4(n11108), .ZN(
        n13725) );
  NAND2_X1 U13575 ( .A1(n13725), .A2(n13854), .ZN(n11112) );
  AND2_X1 U13576 ( .A1(n11113), .A2(n11112), .ZN(n11436) );
  NAND2_X1 U13577 ( .A1(n11114), .A2(n11436), .ZN(n14680) );
  NAND2_X1 U13578 ( .A1(n14680), .A2(n14562), .ZN(n11121) );
  OAI22_X1 U13579 ( .A1(n14562), .A2(n11115), .B1(n11434), .B2(n14555), .ZN(
        n11119) );
  NAND2_X1 U13580 ( .A1(n6438), .A2(n12046), .ZN(n11116) );
  NAND2_X1 U13581 ( .A1(n11116), .A2(n14591), .ZN(n11117) );
  OR2_X1 U13582 ( .A1(n11117), .A2(n11211), .ZN(n14677) );
  NOR2_X1 U13583 ( .A1(n14677), .A2(n14109), .ZN(n11118) );
  AOI211_X1 U13584 ( .C1(n14585), .C2(n12046), .A(n11119), .B(n11118), .ZN(
        n11120) );
  OAI211_X1 U13585 ( .C1(n14092), .C2(n11122), .A(n11121), .B(n11120), .ZN(
        P1_U3284) );
  XNOR2_X1 U13586 ( .A(n11123), .B(n12186), .ZN(n14636) );
  INV_X1 U13587 ( .A(n14092), .ZN(n14596) );
  XNOR2_X1 U13588 ( .A(n11124), .B(n12186), .ZN(n14639) );
  AOI21_X1 U13589 ( .B1(n11157), .B2(n7265), .A(n14575), .ZN(n11126) );
  NAND2_X1 U13590 ( .A1(n11126), .A2(n11125), .ZN(n14633) );
  NOR2_X1 U13591 ( .A1(n14555), .A2(n11127), .ZN(n11128) );
  AOI21_X1 U13592 ( .B1(n14585), .B2(n7265), .A(n11128), .ZN(n11131) );
  MUX2_X1 U13593 ( .A(n11129), .B(n14632), .S(n14562), .Z(n11130) );
  OAI211_X1 U13594 ( .C1(n14109), .C2(n14633), .A(n11131), .B(n11130), .ZN(
        n11132) );
  AOI21_X1 U13595 ( .B1(n14596), .B2(n14639), .A(n11132), .ZN(n11133) );
  OAI21_X1 U13596 ( .B1(n14636), .B2(n13930), .A(n11133), .ZN(P1_U3289) );
  INV_X1 U13597 ( .A(n11134), .ZN(n11135) );
  XNOR2_X1 U13598 ( .A(n12183), .B(n11135), .ZN(n14613) );
  NAND2_X1 U13599 ( .A1(n12183), .A2(n11139), .ZN(n11136) );
  NAND2_X1 U13600 ( .A1(n11136), .A2(n14625), .ZN(n11137) );
  NAND2_X1 U13601 ( .A1(n11137), .A2(n13903), .ZN(n14605) );
  OAI21_X1 U13602 ( .B1(n6591), .B2(n11138), .A(n14590), .ZN(n11145) );
  XNOR2_X1 U13603 ( .A(n11145), .B(n13734), .ZN(n14604) );
  NAND3_X1 U13604 ( .A1(n14063), .A2(n14605), .A3(n14604), .ZN(n11144) );
  NAND2_X1 U13605 ( .A1(n14605), .A2(n11139), .ZN(n11141) );
  NAND2_X1 U13606 ( .A1(n11141), .A2(n11140), .ZN(n14608) );
  NOR2_X1 U13607 ( .A1(n14555), .A2(n13735), .ZN(n11142) );
  AOI21_X1 U13608 ( .B1(n14562), .B2(n14608), .A(n11142), .ZN(n11143) );
  OAI211_X1 U13609 ( .C1(n10044), .C2(n14562), .A(n11144), .B(n11143), .ZN(
        n11147) );
  OR2_X1 U13610 ( .A1(n11145), .A2(n14575), .ZN(n14609) );
  OAI22_X1 U13611 ( .A1(n6591), .A2(n14088), .B1(n14109), .B2(n14609), .ZN(
        n11146) );
  AOI211_X1 U13612 ( .C1(n14613), .C2(n14596), .A(n11147), .B(n11146), .ZN(
        n11148) );
  INV_X1 U13613 ( .A(n11148), .ZN(P1_U3292) );
  XNOR2_X1 U13614 ( .A(n11149), .B(n12003), .ZN(n14628) );
  OR2_X1 U13615 ( .A1(n11150), .A2(n12003), .ZN(n11151) );
  NAND2_X1 U13616 ( .A1(n11152), .A2(n11151), .ZN(n14626) );
  INV_X1 U13617 ( .A(n14621), .ZN(n11153) );
  NAND2_X1 U13618 ( .A1(n14562), .A2(n11153), .ZN(n11156) );
  INV_X1 U13619 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11154) );
  NAND2_X1 U13620 ( .A1(n14586), .A2(n11154), .ZN(n11155) );
  OAI211_X1 U13621 ( .C1(n14562), .C2(n10048), .A(n11156), .B(n11155), .ZN(
        n11159) );
  OAI211_X1 U13622 ( .C1(n14594), .C2(n14623), .A(n11157), .B(n14591), .ZN(
        n14622) );
  OAI22_X1 U13623 ( .A1(n14623), .A2(n14088), .B1(n14109), .B2(n14622), .ZN(
        n11158) );
  AOI211_X1 U13624 ( .C1(n14063), .C2(n14626), .A(n11159), .B(n11158), .ZN(
        n11160) );
  OAI21_X1 U13625 ( .B1(n14092), .B2(n14628), .A(n11160), .ZN(P1_U3290) );
  OR2_X1 U13626 ( .A1(n12046), .A2(n13726), .ZN(n11162) );
  NAND2_X1 U13627 ( .A1(n11163), .A2(n11162), .ZN(n11203) );
  NAND2_X1 U13628 ( .A1(n11164), .A2(n11085), .ZN(n11167) );
  AOI22_X1 U13629 ( .A1(n11165), .A2(n11773), .B1(n11774), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n11166) );
  NAND2_X1 U13630 ( .A1(n11167), .A2(n11166), .ZN(n13595) );
  INV_X1 U13631 ( .A(n13725), .ZN(n11654) );
  OR2_X1 U13632 ( .A1(n13595), .A2(n11654), .ZN(n11184) );
  NAND2_X1 U13633 ( .A1(n13595), .A2(n11654), .ZN(n11168) );
  NAND2_X1 U13634 ( .A1(n11184), .A2(n11168), .ZN(n12194) );
  NAND2_X1 U13635 ( .A1(n11203), .A2(n12194), .ZN(n11170) );
  OR2_X1 U13636 ( .A1(n13595), .A2(n13725), .ZN(n11169) );
  NAND2_X1 U13637 ( .A1(n11171), .A2(n11085), .ZN(n11173) );
  AOI22_X1 U13638 ( .A1(n13822), .A2(n11773), .B1(n11774), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n11172) );
  NAND2_X1 U13639 ( .A1(n12164), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11182) );
  OR2_X1 U13640 ( .A1(n12167), .A2(n14503), .ZN(n11181) );
  NAND2_X1 U13641 ( .A1(n11175), .A2(n11174), .ZN(n11176) );
  NAND2_X1 U13642 ( .A1(n11187), .A2(n11176), .ZN(n14478) );
  OR2_X1 U13643 ( .A1(n9744), .A2(n14478), .ZN(n11180) );
  INV_X1 U13644 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11177) );
  OR2_X1 U13645 ( .A1(n11178), .A2(n11177), .ZN(n11179) );
  NAND4_X1 U13646 ( .A1(n11182), .A2(n11181), .A3(n11180), .A4(n11179), .ZN(
        n13724) );
  XNOR2_X1 U13647 ( .A(n14474), .B(n13724), .ZN(n12195) );
  INV_X1 U13648 ( .A(n12195), .ZN(n11273) );
  XNOR2_X1 U13649 ( .A(n11274), .B(n11273), .ZN(n14497) );
  INV_X1 U13650 ( .A(n14497), .ZN(n11202) );
  AND2_X1 U13651 ( .A1(n12046), .A2(n11427), .ZN(n11204) );
  NOR2_X1 U13652 ( .A1(n12194), .A2(n11204), .ZN(n11183) );
  NAND2_X1 U13653 ( .A1(n11208), .A2(n11184), .ZN(n11185) );
  NAND2_X1 U13654 ( .A1(n11185), .A2(n12195), .ZN(n11298) );
  OAI211_X1 U13655 ( .C1(n11185), .C2(n12195), .A(n11298), .B(n14625), .ZN(
        n11197) );
  NAND2_X1 U13656 ( .A1(n13725), .A2(n14100), .ZN(n11195) );
  NAND2_X1 U13657 ( .A1(n12154), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11193) );
  OR2_X1 U13658 ( .A1(n12167), .A2(n11186), .ZN(n11192) );
  AND2_X1 U13659 ( .A1(n11187), .A2(n11671), .ZN(n11188) );
  OR2_X1 U13660 ( .A1(n11188), .A2(n11291), .ZN(n11668) );
  OR2_X1 U13661 ( .A1(n9744), .A2(n11668), .ZN(n11191) );
  OR2_X1 U13662 ( .A1(n11923), .A2(n11189), .ZN(n11190) );
  NAND4_X1 U13663 ( .A1(n11193), .A2(n11192), .A3(n11191), .A4(n11190), .ZN(
        n13723) );
  NAND2_X1 U13664 ( .A1(n13723), .A2(n13691), .ZN(n11194) );
  NAND2_X1 U13665 ( .A1(n11195), .A2(n11194), .ZN(n14473) );
  INV_X1 U13666 ( .A(n14473), .ZN(n11196) );
  NAND2_X1 U13667 ( .A1(n11197), .A2(n11196), .ZN(n14501) );
  INV_X1 U13668 ( .A(n13595), .ZN(n14687) );
  INV_X1 U13669 ( .A(n14474), .ZN(n14499) );
  NAND2_X1 U13670 ( .A1(n11212), .A2(n14499), .ZN(n14306) );
  OAI211_X1 U13671 ( .C1(n11212), .C2(n14499), .A(n14591), .B(n14306), .ZN(
        n14498) );
  OAI22_X1 U13672 ( .A1(n14562), .A2(n13823), .B1(n14478), .B2(n14555), .ZN(
        n11198) );
  AOI21_X1 U13673 ( .B1(n14474), .B2(n14585), .A(n11198), .ZN(n11199) );
  OAI21_X1 U13674 ( .B1(n14498), .B2(n14109), .A(n11199), .ZN(n11200) );
  AOI21_X1 U13675 ( .B1(n14501), .B2(n14562), .A(n11200), .ZN(n11201) );
  OAI21_X1 U13676 ( .B1(n14092), .B2(n11202), .A(n11201), .ZN(P1_U3282) );
  XNOR2_X1 U13677 ( .A(n11203), .B(n12194), .ZN(n14684) );
  INV_X1 U13678 ( .A(n14684), .ZN(n11220) );
  INV_X1 U13679 ( .A(n11204), .ZN(n11205) );
  NAND2_X1 U13680 ( .A1(n11206), .A2(n11205), .ZN(n11207) );
  NAND2_X1 U13681 ( .A1(n11207), .A2(n12194), .ZN(n11209) );
  NAND3_X1 U13682 ( .A1(n11209), .A2(n14625), .A3(n11208), .ZN(n11210) );
  NAND2_X1 U13683 ( .A1(n13726), .A2(n14100), .ZN(n13591) );
  NAND2_X1 U13684 ( .A1(n11210), .A2(n13591), .ZN(n14689) );
  OAI21_X1 U13685 ( .B1(n11211), .B2(n14687), .A(n14591), .ZN(n11213) );
  OR2_X1 U13686 ( .A1(n11213), .A2(n11212), .ZN(n11214) );
  NAND2_X1 U13687 ( .A1(n13724), .A2(n13691), .ZN(n13592) );
  AND2_X1 U13688 ( .A1(n11214), .A2(n13592), .ZN(n14685) );
  OAI22_X1 U13689 ( .A1(n14562), .A2(n11215), .B1(n13596), .B2(n14555), .ZN(
        n11216) );
  AOI21_X1 U13690 ( .B1(n14585), .B2(n13595), .A(n11216), .ZN(n11217) );
  OAI21_X1 U13691 ( .B1(n14685), .B2(n14109), .A(n11217), .ZN(n11218) );
  AOI21_X1 U13692 ( .B1(n14689), .B2(n14562), .A(n11218), .ZN(n11219) );
  OAI21_X1 U13693 ( .B1(n11220), .B2(n14092), .A(n11219), .ZN(P1_U3283) );
  OAI21_X1 U13694 ( .B1(n11223), .B2(n11222), .A(n11221), .ZN(n11224) );
  NAND2_X1 U13695 ( .A1(n11224), .A2(n13093), .ZN(n11229) );
  OAI22_X1 U13696 ( .A1(n13097), .A2(n11225), .B1(n13096), .B2(n11240), .ZN(
        n11226) );
  AOI211_X1 U13697 ( .C1(n11564), .C2(n13121), .A(n11227), .B(n11226), .ZN(
        n11228) );
  OAI211_X1 U13698 ( .C1(n11333), .C2(n13102), .A(n11229), .B(n11228), .ZN(
        P2_U3208) );
  XOR2_X1 U13699 ( .A(n11230), .B(n11234), .Z(n11331) );
  INV_X1 U13700 ( .A(n11331), .ZN(n11246) );
  INV_X1 U13701 ( .A(n11231), .ZN(n11232) );
  AOI21_X1 U13702 ( .B1(n11234), .B2(n11233), .A(n11232), .ZN(n11238) );
  INV_X1 U13703 ( .A(n13355), .ZN(n11235) );
  NAND2_X1 U13704 ( .A1(n11331), .A2(n11235), .ZN(n11237) );
  AOI22_X1 U13705 ( .A1(n13311), .A2(n13121), .B1(n13119), .B2(n13312), .ZN(
        n11236) );
  OAI211_X1 U13706 ( .C1(n13405), .C2(n11238), .A(n11237), .B(n11236), .ZN(
        n11329) );
  NAND2_X1 U13707 ( .A1(n11329), .A2(n13356), .ZN(n11245) );
  AOI211_X1 U13708 ( .C1(n11337), .C2(n11239), .A(n13394), .B(n11357), .ZN(
        n11330) );
  NOR2_X1 U13709 ( .A1(n11333), .A2(n13376), .ZN(n11243) );
  OAI22_X1 U13710 ( .A1(n13427), .A2(n11241), .B1(n11240), .B2(n13412), .ZN(
        n11242) );
  AOI211_X1 U13711 ( .C1(n11330), .C2(n13422), .A(n11243), .B(n11242), .ZN(
        n11244) );
  OAI211_X1 U13712 ( .C1(n11246), .C2(n13367), .A(n11245), .B(n11244), .ZN(
        P2_U3254) );
  NAND2_X1 U13713 ( .A1(n11247), .A2(n14288), .ZN(n11249) );
  OAI211_X1 U13714 ( .C1(n11250), .C2(n12992), .A(n11249), .B(n11248), .ZN(
        P3_U3272) );
  AOI22_X1 U13715 ( .A1(n14666), .A2(n11863), .B1(n11928), .B2(n13727), .ZN(
        n11426) );
  AOI22_X1 U13716 ( .A1(n14666), .A2(n11929), .B1(n11863), .B2(n13727), .ZN(
        n11251) );
  XNOR2_X1 U13717 ( .A(n11251), .B(n12232), .ZN(n11423) );
  XOR2_X1 U13718 ( .A(n11426), .B(n11423), .Z(n11258) );
  INV_X1 U13719 ( .A(n11253), .ZN(n11254) );
  AOI21_X1 U13720 ( .B1(n11258), .B2(n11257), .A(n11424), .ZN(n11264) );
  OAI22_X1 U13721 ( .A1(n11259), .A2(n13903), .B1(n11427), .B2(n14098), .ZN(
        n14551) );
  AOI21_X1 U13722 ( .B1(n14472), .B2(n14551), .A(n11260), .ZN(n11261) );
  OAI21_X1 U13723 ( .B1(n14554), .B2(n14479), .A(n11261), .ZN(n11262) );
  AOI21_X1 U13724 ( .B1(n14666), .B2(n14475), .A(n11262), .ZN(n11263) );
  OAI21_X1 U13725 ( .B1(n11264), .B2(n13705), .A(n11263), .ZN(P1_U3221) );
  INV_X1 U13726 ( .A(n11812), .ZN(n11327) );
  OAI222_X1 U13727 ( .A1(n14244), .A2(n11327), .B1(n11982), .B2(P1_U3086), 
        .C1(n11813), .C2(n14245), .ZN(P1_U3334) );
  INV_X1 U13728 ( .A(n15011), .ZN(n11272) );
  OAI211_X1 U13729 ( .C1(n11267), .C2(n11266), .A(n11265), .B(n14861), .ZN(
        n11271) );
  INV_X1 U13730 ( .A(n12410), .ZN(n15016) );
  OAI22_X1 U13731 ( .A1(n12395), .A2(n15010), .B1(n12390), .B2(n15016), .ZN(
        n11268) );
  AOI211_X1 U13732 ( .C1(n14860), .C2(n12408), .A(n11269), .B(n11268), .ZN(
        n11270) );
  OAI211_X1 U13733 ( .C1(n11272), .C2(n11503), .A(n11271), .B(n11270), .ZN(
        P3_U3161) );
  NAND2_X1 U13734 ( .A1(n11274), .A2(n11273), .ZN(n11276) );
  OR2_X1 U13735 ( .A1(n14474), .A2(n13724), .ZN(n11275) );
  NAND2_X1 U13736 ( .A1(n11276), .A2(n11275), .ZN(n14297) );
  NAND2_X1 U13737 ( .A1(n11277), .A2(n11085), .ZN(n11280) );
  AOI22_X1 U13738 ( .A1(n11278), .A2(n11773), .B1(n11774), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n11279) );
  XNOR2_X1 U13739 ( .A(n14304), .B(n13723), .ZN(n14299) );
  INV_X1 U13740 ( .A(n14299), .ZN(n11281) );
  NAND2_X1 U13741 ( .A1(n14297), .A2(n11281), .ZN(n11283) );
  OR2_X1 U13742 ( .A1(n14304), .A2(n13723), .ZN(n11282) );
  NAND2_X1 U13743 ( .A1(n11284), .A2(n11085), .ZN(n11289) );
  OAI22_X1 U13744 ( .A1(n11286), .A2(n11835), .B1(n12160), .B2(n11285), .ZN(
        n11287) );
  INV_X1 U13745 ( .A(n11287), .ZN(n11288) );
  NAND2_X1 U13746 ( .A1(n12154), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11297) );
  OR2_X1 U13747 ( .A1(n12167), .A2(n11290), .ZN(n11296) );
  OR2_X1 U13748 ( .A1(n11291), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11292) );
  NAND2_X1 U13749 ( .A1(n11303), .A2(n11292), .ZN(n13665) );
  OR2_X1 U13750 ( .A1(n9744), .A2(n13665), .ZN(n11295) );
  OR2_X1 U13751 ( .A1(n11923), .A2(n11293), .ZN(n11294) );
  NAND4_X1 U13752 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(
        n14101) );
  XNOR2_X1 U13753 ( .A(n12068), .B(n14101), .ZN(n12197) );
  XNOR2_X1 U13754 ( .A(n11535), .B(n12197), .ZN(n14489) );
  INV_X1 U13755 ( .A(n13724), .ZN(n11643) );
  OAI21_X1 U13756 ( .B1(n11643), .B2(n14474), .A(n11298), .ZN(n14300) );
  INV_X1 U13757 ( .A(n13723), .ZN(n11661) );
  OAI211_X1 U13758 ( .C1(n11300), .C2(n12197), .A(n14625), .B(n11515), .ZN(
        n11301) );
  INV_X1 U13759 ( .A(n11301), .ZN(n14494) );
  NAND2_X1 U13760 ( .A1(n12154), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11308) );
  OR2_X1 U13761 ( .A1(n12167), .A2(n14488), .ZN(n11307) );
  NAND2_X1 U13762 ( .A1(n11303), .A2(n11302), .ZN(n11304) );
  NAND2_X1 U13763 ( .A1(n11525), .A2(n11304), .ZN(n14466) );
  OR2_X1 U13764 ( .A1(n9744), .A2(n14466), .ZN(n11306) );
  OR2_X1 U13765 ( .A1(n11923), .A2(n14105), .ZN(n11305) );
  OR2_X1 U13766 ( .A1(n11723), .A2(n14098), .ZN(n11310) );
  NAND2_X1 U13767 ( .A1(n13723), .A2(n14100), .ZN(n11309) );
  NAND2_X1 U13768 ( .A1(n11310), .A2(n11309), .ZN(n14490) );
  OAI21_X1 U13769 ( .B1(n14494), .B2(n14490), .A(n14562), .ZN(n11314) );
  OAI22_X1 U13770 ( .A1(n14562), .A2(n11293), .B1(n13665), .B2(n14555), .ZN(
        n11312) );
  INV_X1 U13771 ( .A(n12068), .ZN(n14493) );
  INV_X1 U13772 ( .A(n11543), .ZN(n14106) );
  OAI211_X1 U13773 ( .C1(n14493), .C2(n6929), .A(n14591), .B(n14106), .ZN(
        n14492) );
  NOR2_X1 U13774 ( .A1(n14492), .A2(n14109), .ZN(n11311) );
  AOI211_X1 U13775 ( .C1(n14585), .C2(n12068), .A(n11312), .B(n11311), .ZN(
        n11313) );
  OAI211_X1 U13776 ( .C1(n14489), .C2(n14092), .A(n11314), .B(n11313), .ZN(
        P1_U3280) );
  XNOR2_X1 U13777 ( .A(n11315), .B(n11316), .ZN(n11321) );
  XNOR2_X1 U13778 ( .A(n11317), .B(n11316), .ZN(n11318) );
  NAND2_X1 U13779 ( .A1(n11318), .A2(n15089), .ZN(n11320) );
  AOI22_X1 U13780 ( .A1(n15084), .A2(n12409), .B1(n11461), .B2(n15081), .ZN(
        n11319) );
  OAI211_X1 U13781 ( .C1(n15094), .C2(n11321), .A(n11320), .B(n11319), .ZN(
        n15138) );
  INV_X1 U13782 ( .A(n15138), .ZN(n11325) );
  INV_X1 U13783 ( .A(n11321), .ZN(n15141) );
  NOR2_X1 U13784 ( .A1(n11463), .A2(n15076), .ZN(n15139) );
  AOI22_X1 U13785 ( .A1(n15070), .A2(n15139), .B1(n15103), .B2(n11466), .ZN(
        n11322) );
  OAI21_X1 U13786 ( .B1(n14890), .B2(n15109), .A(n11322), .ZN(n11323) );
  AOI21_X1 U13787 ( .B1(n15141), .B2(n12586), .A(n11323), .ZN(n11324) );
  OAI21_X1 U13788 ( .B1(n11325), .B2(n15005), .A(n11324), .ZN(P3_U3224) );
  OAI222_X1 U13789 ( .A1(P2_U3088), .A2(n11328), .B1(n13575), .B2(n11327), 
        .C1(n11326), .C2(n13573), .ZN(P2_U3306) );
  AOI211_X1 U13790 ( .C1(n11331), .C2(n9151), .A(n11330), .B(n11329), .ZN(
        n11339) );
  INV_X1 U13791 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11332) );
  OAI22_X1 U13792 ( .A1(n11333), .A2(n13548), .B1(n14457), .B2(n11332), .ZN(
        n11334) );
  INV_X1 U13793 ( .A(n11334), .ZN(n11335) );
  OAI21_X1 U13794 ( .B1(n11339), .B2(n14450), .A(n11335), .ZN(P2_U3463) );
  AOI22_X1 U13795 ( .A1(n11337), .A2(n11336), .B1(n8929), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11338) );
  OAI21_X1 U13796 ( .B1(n11339), .B2(n8929), .A(n11338), .ZN(P2_U3510) );
  OAI21_X1 U13797 ( .B1(n11342), .B2(n11341), .A(n11340), .ZN(n11343) );
  NAND2_X1 U13798 ( .A1(n11343), .A2(n13093), .ZN(n11347) );
  NAND2_X1 U13799 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14746)
         );
  INV_X1 U13800 ( .A(n14746), .ZN(n11345) );
  OAI22_X1 U13801 ( .A1(n13097), .A2(n7760), .B1(n13096), .B2(n11355), .ZN(
        n11344) );
  AOI211_X1 U13802 ( .C1(n11564), .C2(n13120), .A(n11345), .B(n11344), .ZN(
        n11346) );
  OAI211_X1 U13803 ( .C1(n14444), .C2(n13102), .A(n11347), .B(n11346), .ZN(
        P2_U3196) );
  XOR2_X1 U13804 ( .A(n11349), .B(n11348), .Z(n14442) );
  XOR2_X1 U13805 ( .A(n11350), .B(n11349), .Z(n11353) );
  OAI22_X1 U13806 ( .A1(n11351), .A2(n13404), .B1(n7760), .B2(n13408), .ZN(
        n11352) );
  AOI21_X1 U13807 ( .B1(n11353), .B2(n13352), .A(n11352), .ZN(n11354) );
  OAI21_X1 U13808 ( .B1(n14442), .B2(n13355), .A(n11354), .ZN(n14445) );
  NAND2_X1 U13809 ( .A1(n14445), .A2(n13356), .ZN(n11362) );
  OAI22_X1 U13810 ( .A1(n13427), .A2(n11356), .B1(n11355), .B2(n13412), .ZN(
        n11359) );
  OAI211_X1 U13811 ( .C1(n11357), .C2(n14444), .A(n11416), .B(n13420), .ZN(
        n14443) );
  NOR2_X1 U13812 ( .A1(n14443), .A2(n13269), .ZN(n11358) );
  AOI211_X1 U13813 ( .C1(n13416), .C2(n11360), .A(n11359), .B(n11358), .ZN(
        n11361) );
  OAI211_X1 U13814 ( .C1(n14442), .C2(n13367), .A(n11362), .B(n11361), .ZN(
        P2_U3253) );
  XNOR2_X1 U13815 ( .A(n11364), .B(n11363), .ZN(n11370) );
  NAND2_X1 U13816 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n14748)
         );
  NAND2_X1 U13817 ( .A1(n13117), .A2(n13312), .ZN(n11366) );
  NAND2_X1 U13818 ( .A1(n13119), .A2(n13311), .ZN(n11365) );
  NAND2_X1 U13819 ( .A1(n11366), .A2(n11365), .ZN(n11410) );
  NAND2_X1 U13820 ( .A1(n13056), .A2(n11410), .ZN(n11367) );
  OAI211_X1 U13821 ( .C1(n13096), .C2(n11414), .A(n14748), .B(n11367), .ZN(
        n11368) );
  AOI21_X1 U13822 ( .B1(n11420), .B2(n13086), .A(n11368), .ZN(n11369) );
  OAI21_X1 U13823 ( .B1(n11370), .B2(n13088), .A(n11369), .ZN(P2_U3206) );
  NAND2_X1 U13824 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n11382), .ZN(n11378) );
  AOI22_X1 U13825 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n11382), .B1(n14806), 
        .B2(n13392), .ZN(n14800) );
  AOI22_X1 U13826 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n11383), .B1(n14793), 
        .B2(n13414), .ZN(n14787) );
  OR2_X1 U13827 ( .A1(n11384), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n14737) );
  NAND2_X1 U13828 ( .A1(n14739), .A2(n14737), .ZN(n11371) );
  MUX2_X1 U13829 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11356), .S(n14742), .Z(
        n14736) );
  NAND2_X1 U13830 ( .A1(n11371), .A2(n14736), .ZN(n14741) );
  NAND2_X1 U13831 ( .A1(n11388), .A2(n11356), .ZN(n11372) );
  OR2_X1 U13832 ( .A1(n11389), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U13833 ( .A1(n11389), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11374) );
  AND2_X1 U13834 ( .A1(n11373), .A2(n11374), .ZN(n14755) );
  NAND2_X1 U13835 ( .A1(n14756), .A2(n14755), .ZN(n14754) );
  AND3_X1 U13836 ( .A1(n14754), .A2(n14772), .A3(n11374), .ZN(n14760) );
  AOI21_X1 U13837 ( .B1(n14754), .B2(n11374), .A(n14772), .ZN(n14761) );
  INV_X1 U13838 ( .A(n14761), .ZN(n11375) );
  OAI21_X1 U13839 ( .B1(n14760), .B2(n11485), .A(n11375), .ZN(n11376) );
  NAND2_X1 U13840 ( .A1(n14774), .A2(n11376), .ZN(n11377) );
  XOR2_X1 U13841 ( .A(n14774), .B(n11376), .Z(n14777) );
  NAND2_X1 U13842 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14777), .ZN(n14775) );
  NAND2_X1 U13843 ( .A1(n11377), .A2(n14775), .ZN(n14786) );
  NAND2_X1 U13844 ( .A1(n14787), .A2(n14786), .ZN(n14785) );
  OAI21_X1 U13845 ( .B1(n14793), .B2(n13414), .A(n14785), .ZN(n14799) );
  NAND2_X1 U13846 ( .A1(n14800), .A2(n14799), .ZN(n14798) );
  NAND2_X1 U13847 ( .A1(n11378), .A2(n14798), .ZN(n11379) );
  XNOR2_X1 U13848 ( .A(n14818), .B(n11379), .ZN(n14815) );
  NOR2_X1 U13849 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14815), .ZN(n14814) );
  NOR2_X1 U13850 ( .A1(n14818), .A2(n11379), .ZN(n11380) );
  NOR2_X1 U13851 ( .A1(n14814), .A2(n11380), .ZN(n11381) );
  XOR2_X1 U13852 ( .A(n11381), .B(P2_REG2_REG_19__SCAN_IN), .Z(n11404) );
  INV_X1 U13853 ( .A(n11404), .ZN(n11402) );
  AOI22_X1 U13854 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n11382), .B1(n14806), 
        .B2(n11397), .ZN(n14803) );
  AOI22_X1 U13855 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n11383), .B1(n14793), 
        .B2(n11396), .ZN(n14790) );
  MUX2_X1 U13856 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7773), .S(n14772), .Z(
        n14763) );
  INV_X1 U13857 ( .A(n14763), .ZN(n11391) );
  NAND2_X1 U13858 ( .A1(n11384), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U13859 ( .A1(n11386), .A2(n11385), .ZN(n14733) );
  MUX2_X1 U13860 ( .A(n11387), .B(P2_REG1_REG_12__SCAN_IN), .S(n14742), .Z(
        n14732) );
  NOR2_X1 U13861 ( .A1(n14733), .A2(n14732), .ZN(n14735) );
  AOI21_X1 U13862 ( .B1(n11387), .B2(n11388), .A(n14735), .ZN(n14753) );
  MUX2_X1 U13863 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n11390), .S(n11389), .Z(
        n14752) );
  NAND2_X1 U13864 ( .A1(n14753), .A2(n14752), .ZN(n14751) );
  OAI21_X1 U13865 ( .B1(n11390), .B2(n14749), .A(n14751), .ZN(n14764) );
  NAND2_X1 U13866 ( .A1(n11391), .A2(n14764), .ZN(n11392) );
  OAI21_X1 U13867 ( .B1(n14772), .B2(n7773), .A(n11392), .ZN(n11393) );
  NAND2_X1 U13868 ( .A1(n14774), .A2(n11393), .ZN(n11395) );
  XNOR2_X1 U13869 ( .A(n11394), .B(n11393), .ZN(n14780) );
  NAND2_X1 U13870 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14780), .ZN(n14778) );
  NAND2_X1 U13871 ( .A1(n11395), .A2(n14778), .ZN(n14789) );
  NAND2_X1 U13872 ( .A1(n14790), .A2(n14789), .ZN(n14788) );
  OAI21_X1 U13873 ( .B1(n14793), .B2(n11396), .A(n14788), .ZN(n14802) );
  NAND2_X1 U13874 ( .A1(n14803), .A2(n14802), .ZN(n14801) );
  OAI21_X1 U13875 ( .B1(n14806), .B2(n11397), .A(n14801), .ZN(n11398) );
  XOR2_X1 U13876 ( .A(n14818), .B(n11398), .Z(n14813) );
  NAND2_X1 U13877 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14813), .ZN(n14812) );
  NAND2_X1 U13878 ( .A1(n14818), .A2(n11398), .ZN(n11399) );
  NAND2_X1 U13879 ( .A1(n14812), .A2(n11399), .ZN(n11400) );
  XOR2_X1 U13880 ( .A(n11400), .B(P2_REG1_REG_19__SCAN_IN), .Z(n11403) );
  OAI21_X1 U13881 ( .B1(n11403), .B2(n14822), .A(n14807), .ZN(n11401) );
  AOI21_X1 U13882 ( .B1(n11402), .B2(n14776), .A(n11401), .ZN(n11407) );
  AOI22_X1 U13883 ( .A1(n11404), .A2(n14776), .B1(n14779), .B2(n11403), .ZN(
        n11406) );
  MUX2_X1 U13884 ( .A(n11407), .B(n11406), .S(n11405), .Z(n11408) );
  NAND2_X1 U13885 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13018)
         );
  OAI211_X1 U13886 ( .C1(n7424), .C2(n14827), .A(n11408), .B(n13018), .ZN(
        P2_U3233) );
  XOR2_X1 U13887 ( .A(n11409), .B(n11412), .Z(n11411) );
  AOI21_X1 U13888 ( .B1(n11411), .B2(n13352), .A(n11410), .ZN(n14437) );
  XOR2_X1 U13889 ( .A(n11413), .B(n11412), .Z(n14441) );
  NAND2_X1 U13890 ( .A1(n14441), .A2(n13373), .ZN(n11422) );
  OAI22_X1 U13891 ( .A1(n13427), .A2(n11415), .B1(n11414), .B2(n13412), .ZN(
        n11419) );
  INV_X1 U13892 ( .A(n11416), .ZN(n11417) );
  OAI211_X1 U13893 ( .C1(n11417), .C2(n14438), .A(n13420), .B(n11486), .ZN(
        n14436) );
  NOR2_X1 U13894 ( .A1(n14436), .A2(n13269), .ZN(n11418) );
  AOI211_X1 U13895 ( .C1(n13416), .C2(n11420), .A(n11419), .B(n11418), .ZN(
        n11421) );
  OAI211_X1 U13896 ( .C1(n13384), .C2(n14437), .A(n11422), .B(n11421), .ZN(
        P2_U3252) );
  INV_X1 U13897 ( .A(n12046), .ZN(n14678) );
  INV_X1 U13898 ( .A(n11423), .ZN(n11425) );
  NOR2_X1 U13899 ( .A1(n9756), .A2(n11427), .ZN(n11428) );
  AOI21_X1 U13900 ( .B1(n12046), .B2(n11863), .A(n11428), .ZN(n11648) );
  NAND2_X1 U13901 ( .A1(n12046), .A2(n11929), .ZN(n11430) );
  NAND2_X1 U13902 ( .A1(n11863), .A2(n13726), .ZN(n11429) );
  NAND2_X1 U13903 ( .A1(n11430), .A2(n11429), .ZN(n11431) );
  XNOR2_X1 U13904 ( .A(n11431), .B(n11652), .ZN(n11649) );
  XOR2_X1 U13905 ( .A(n11648), .B(n11649), .Z(n11432) );
  OAI211_X1 U13906 ( .C1(n11433), .C2(n11432), .A(n6671), .B(n14470), .ZN(
        n11440) );
  NOR2_X1 U13907 ( .A1(n14479), .A2(n11434), .ZN(n11438) );
  OAI22_X1 U13908 ( .A1(n13712), .A2(n11436), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11435), .ZN(n11437) );
  NOR2_X1 U13909 ( .A1(n11438), .A2(n11437), .ZN(n11439) );
  OAI211_X1 U13910 ( .C1(n14678), .C2(n13718), .A(n11440), .B(n11439), .ZN(
        P1_U3231) );
  NAND2_X1 U13911 ( .A1(n11743), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11445) );
  INV_X1 U13912 ( .A(n11441), .ZN(n11442) );
  NAND2_X1 U13913 ( .A1(n11443), .A2(n11442), .ZN(n11444) );
  NAND2_X1 U13914 ( .A1(n11445), .A2(n11444), .ZN(n13836) );
  XOR2_X1 U13915 ( .A(n13837), .B(n13836), .Z(n11446) );
  NAND2_X1 U13916 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11446), .ZN(n13838) );
  OAI211_X1 U13917 ( .C1(n11446), .C2(P1_REG2_REG_18__SCAN_IN), .A(n13846), 
        .B(n13838), .ZN(n11454) );
  NAND2_X1 U13918 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13683)
         );
  INV_X1 U13919 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11449) );
  OAI21_X1 U13920 ( .B1(n11449), .B2(n11448), .A(n11447), .ZN(n13832) );
  XNOR2_X1 U13921 ( .A(n13832), .B(n11455), .ZN(n11450) );
  NAND2_X1 U13922 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n11450), .ZN(n13834) );
  OAI211_X1 U13923 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11450), .A(n13841), 
        .B(n13834), .ZN(n11451) );
  NAND2_X1 U13924 ( .A1(n13683), .A2(n11451), .ZN(n11452) );
  AOI21_X1 U13925 ( .B1(n13776), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11452), 
        .ZN(n11453) );
  OAI211_X1 U13926 ( .C1(n11456), .C2(n11455), .A(n11454), .B(n11453), .ZN(
        P1_U3261) );
  INV_X1 U13927 ( .A(n11457), .ZN(n11458) );
  AOI21_X1 U13928 ( .B1(n11460), .B2(n11459), .A(n11458), .ZN(n11468) );
  INV_X1 U13929 ( .A(n11461), .ZN(n11617) );
  OAI22_X1 U13930 ( .A1(n12378), .A2(n11617), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14891), .ZN(n11465) );
  INV_X1 U13931 ( .A(n12409), .ZN(n11462) );
  OAI22_X1 U13932 ( .A1(n12395), .A2(n11463), .B1(n12390), .B2(n11462), .ZN(
        n11464) );
  AOI211_X1 U13933 ( .C1(n11466), .C2(n12392), .A(n11465), .B(n11464), .ZN(
        n11467) );
  OAI21_X1 U13934 ( .B1(n11468), .B2(n12382), .A(n11467), .ZN(P3_U3171) );
  INV_X1 U13935 ( .A(n11469), .ZN(n11472) );
  OAI222_X1 U13936 ( .A1(n13575), .A2(n11472), .B1(n11471), .B2(P2_U3088), 
        .C1(n11470), .C2(n13573), .ZN(P2_U3305) );
  OAI21_X1 U13937 ( .B1(n6565), .B2(n11473), .A(n6436), .ZN(n15000) );
  OAI211_X1 U13938 ( .C1(n11476), .C2(n11475), .A(n11474), .B(n15089), .ZN(
        n11478) );
  AOI22_X1 U13939 ( .A1(n15081), .A2(n12407), .B1(n12408), .B2(n15084), .ZN(
        n11477) );
  NAND2_X1 U13940 ( .A1(n11478), .A2(n11477), .ZN(n14999) );
  AOI21_X1 U13941 ( .B1(n15136), .B2(n15000), .A(n14999), .ZN(n11480) );
  MUX2_X1 U13942 ( .A(n8319), .B(n11480), .S(n15143), .Z(n11479) );
  OAI21_X1 U13943 ( .B1(n12965), .B2(n11499), .A(n11479), .ZN(P3_U3420) );
  INV_X1 U13944 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12417) );
  MUX2_X1 U13945 ( .A(n12417), .B(n11480), .S(n15159), .Z(n11481) );
  OAI21_X1 U13946 ( .B1(n12899), .B2(n11499), .A(n11481), .ZN(P3_U3469) );
  OAI21_X1 U13947 ( .B1(n11483), .B2(n6780), .A(n11482), .ZN(n11484) );
  AOI222_X1 U13948 ( .A1(n13352), .A2(n11484), .B1(n13116), .B2(n13312), .C1(
        n13118), .C2(n13311), .ZN(n14431) );
  OAI22_X1 U13949 ( .A1(n13427), .A2(n11485), .B1(n11561), .B2(n13412), .ZN(
        n11489) );
  INV_X1 U13950 ( .A(n11490), .ZN(n14432) );
  INV_X1 U13951 ( .A(n11486), .ZN(n11487) );
  OAI211_X1 U13952 ( .C1(n14432), .C2(n11487), .A(n13420), .B(n11595), .ZN(
        n14430) );
  NOR2_X1 U13953 ( .A1(n14430), .A2(n13269), .ZN(n11488) );
  AOI211_X1 U13954 ( .C1(n13416), .C2(n11490), .A(n11489), .B(n11488), .ZN(
        n11494) );
  AND2_X1 U13955 ( .A1(n11491), .A2(n6780), .ZN(n14429) );
  INV_X1 U13956 ( .A(n14429), .ZN(n11492) );
  NAND3_X1 U13957 ( .A1(n11492), .A2(n13373), .A3(n14434), .ZN(n11493) );
  OAI211_X1 U13958 ( .C1(n14431), .C2(n13384), .A(n11494), .B(n11493), .ZN(
        P2_U3251) );
  AOI21_X1 U13959 ( .B1(n11496), .B2(n11495), .A(n12382), .ZN(n11498) );
  NAND2_X1 U13960 ( .A1(n11498), .A2(n11497), .ZN(n11502) );
  AND2_X1 U13961 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n14912) );
  OAI22_X1 U13962 ( .A1(n12395), .A2(n11499), .B1(n12390), .B2(n15017), .ZN(
        n11500) );
  AOI211_X1 U13963 ( .C1(n14860), .C2(n12407), .A(n14912), .B(n11500), .ZN(
        n11501) );
  OAI211_X1 U13964 ( .C1(n15009), .C2(n11503), .A(n11502), .B(n11501), .ZN(
        P3_U3157) );
  XNOR2_X1 U13965 ( .A(n11504), .B(n11506), .ZN(n11505) );
  OAI222_X1 U13966 ( .A1(n15044), .A2(n11617), .B1(n15046), .B2(n12352), .C1(
        n15052), .C2(n11505), .ZN(n14414) );
  INV_X1 U13967 ( .A(n14414), .ZN(n11514) );
  NAND2_X1 U13968 ( .A1(n6436), .A2(n11508), .ZN(n11507) );
  MUX2_X1 U13969 ( .A(n11508), .B(n11507), .S(n11506), .Z(n11510) );
  NAND2_X1 U13970 ( .A1(n11510), .A2(n11509), .ZN(n14416) );
  NAND2_X1 U13971 ( .A1(n15094), .A2(n15106), .ZN(n15001) );
  NAND2_X1 U13972 ( .A1(n15109), .A2(n15001), .ZN(n12498) );
  AOI22_X1 U13973 ( .A1(n15005), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15103), 
        .B2(n11619), .ZN(n11511) );
  OAI21_X1 U13974 ( .B1(n14413), .B2(n12826), .A(n11511), .ZN(n11512) );
  AOI21_X1 U13975 ( .B1(n14416), .B2(n15020), .A(n11512), .ZN(n11513) );
  OAI21_X1 U13976 ( .B1(n11514), .B2(n15005), .A(n11513), .ZN(P3_U3222) );
  INV_X1 U13977 ( .A(n14101), .ZN(n11717) );
  NAND2_X1 U13978 ( .A1(n11516), .A2(n11085), .ZN(n11519) );
  AOI22_X1 U13979 ( .A1(n11517), .A2(n11773), .B1(n11774), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U13980 ( .A1(n14481), .A2(n11723), .ZN(n12072) );
  NAND2_X1 U13981 ( .A1(n11520), .A2(n11085), .ZN(n11522) );
  AOI22_X1 U13982 ( .A1(n11774), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11773), 
        .B2(n14535), .ZN(n11521) );
  NAND2_X2 U13983 ( .A1(n11522), .A2(n11521), .ZN(n11704) );
  INV_X1 U13984 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U13985 ( .A1(n11525), .A2(n11524), .ZN(n11526) );
  NAND2_X1 U13986 ( .A1(n11546), .A2(n11526), .ZN(n13711) );
  OR2_X1 U13987 ( .A1(n13711), .A2(n9744), .ZN(n11532) );
  NAND2_X1 U13988 ( .A1(n12154), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11531) );
  INV_X1 U13989 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11527) );
  OR2_X1 U13990 ( .A1(n12167), .A2(n11527), .ZN(n11530) );
  INV_X1 U13991 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11528) );
  OR2_X1 U13992 ( .A1(n11923), .A2(n11528), .ZN(n11529) );
  OR2_X2 U13993 ( .A1(n11704), .A2(n14099), .ZN(n12078) );
  NAND2_X1 U13994 ( .A1(n11704), .A2(n14099), .ZN(n12079) );
  NAND2_X1 U13995 ( .A1(n12078), .A2(n12079), .ZN(n12199) );
  NAND2_X1 U13996 ( .A1(n11533), .A2(n11541), .ZN(n11685) );
  OAI21_X1 U13997 ( .B1(n11533), .B2(n11541), .A(n11685), .ZN(n14207) );
  INV_X1 U13998 ( .A(n12197), .ZN(n11534) );
  NAND2_X1 U13999 ( .A1(n11535), .A2(n11534), .ZN(n11537) );
  OR2_X1 U14000 ( .A1(n12068), .A2(n14101), .ZN(n11536) );
  INV_X1 U14001 ( .A(n11723), .ZN(n13722) );
  NAND2_X1 U14002 ( .A1(n14481), .A2(n13722), .ZN(n11540) );
  OAI21_X1 U14003 ( .B1(n6557), .B2(n12199), .A(n11705), .ZN(n14205) );
  NAND2_X1 U14004 ( .A1(n11704), .A2(n14107), .ZN(n11544) );
  NAND2_X1 U14005 ( .A1(n11544), .A2(n14591), .ZN(n11545) );
  NOR2_X1 U14006 ( .A1(n11699), .A2(n11545), .ZN(n14204) );
  NAND2_X1 U14007 ( .A1(n14204), .A2(n14595), .ZN(n11554) );
  NAND2_X1 U14008 ( .A1(n11546), .A2(n12613), .ZN(n11547) );
  NAND2_X1 U14009 ( .A1(n11692), .A2(n11547), .ZN(n13630) );
  AOI22_X1 U14010 ( .A1(n11548), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n12154), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n11551) );
  OR2_X1 U14011 ( .A1(n11923), .A2(n11549), .ZN(n11550) );
  OAI211_X1 U14012 ( .C1(n13630), .C2(n9744), .A(n11551), .B(n11550), .ZN(
        n13880) );
  AOI22_X1 U14013 ( .A1(n13722), .A2(n14100), .B1(n13880), .B2(n13854), .ZN(
        n14201) );
  OAI22_X1 U14014 ( .A1(n14599), .A2(n14201), .B1(n13711), .B2(n14555), .ZN(
        n11552) );
  AOI21_X1 U14015 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14599), .A(n11552), 
        .ZN(n11553) );
  OAI211_X1 U14016 ( .C1(n14202), .C2(n14088), .A(n11554), .B(n11553), .ZN(
        n11555) );
  AOI21_X1 U14017 ( .B1(n14205), .B2(n14596), .A(n11555), .ZN(n11556) );
  OAI21_X1 U14018 ( .B1(n14207), .B2(n13930), .A(n11556), .ZN(P1_U3278) );
  OAI21_X1 U14019 ( .B1(n11559), .B2(n11558), .A(n11557), .ZN(n11560) );
  NAND2_X1 U14020 ( .A1(n11560), .A2(n13093), .ZN(n11566) );
  NAND2_X1 U14021 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14766)
         );
  INV_X1 U14022 ( .A(n14766), .ZN(n11563) );
  OAI22_X1 U14023 ( .A1(n13097), .A2(n13403), .B1(n13096), .B2(n11561), .ZN(
        n11562) );
  AOI211_X1 U14024 ( .C1(n11564), .C2(n13118), .A(n11563), .B(n11562), .ZN(
        n11565) );
  OAI211_X1 U14025 ( .C1(n14432), .C2(n13102), .A(n11566), .B(n11565), .ZN(
        P2_U3187) );
  OAI22_X1 U14026 ( .A1(n11567), .A2(P3_U3151), .B1(n12683), .B2(n12992), .ZN(
        n11568) );
  AOI21_X1 U14027 ( .B1(n11569), .B2(n14288), .A(n11568), .ZN(n11570) );
  INV_X1 U14028 ( .A(n11570), .ZN(P3_U3271) );
  NAND2_X1 U14029 ( .A1(n11571), .A2(n11576), .ZN(n11572) );
  NAND3_X1 U14030 ( .A1(n11573), .A2(n15089), .A3(n11572), .ZN(n11575) );
  AOI22_X1 U14031 ( .A1(n15084), .A2(n12406), .B1(n12404), .B2(n15081), .ZN(
        n11574) );
  AND2_X1 U14032 ( .A1(n11575), .A2(n11574), .ZN(n12896) );
  OR2_X1 U14033 ( .A1(n11577), .A2(n11576), .ZN(n11578) );
  NAND2_X1 U14034 ( .A1(n11579), .A2(n11578), .ZN(n12894) );
  AOI22_X1 U14035 ( .A1(n15005), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15103), 
        .B2(n12355), .ZN(n11580) );
  OAI21_X1 U14036 ( .B1(n12964), .B2(n12826), .A(n11580), .ZN(n11581) );
  AOI21_X1 U14037 ( .B1(n12894), .B2(n15020), .A(n11581), .ZN(n11582) );
  OAI21_X1 U14038 ( .B1(n12896), .B2(n15005), .A(n11582), .ZN(P3_U3220) );
  NAND2_X1 U14039 ( .A1(n11583), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11584) );
  OAI211_X1 U14040 ( .C1(n11850), .C2(n13575), .A(n11585), .B(n11584), .ZN(
        P2_U3304) );
  NAND2_X1 U14041 ( .A1(n11586), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11587) );
  OAI211_X1 U14042 ( .C1(n11850), .C2(n14244), .A(n12225), .B(n11587), .ZN(
        P1_U3332) );
  AOI21_X1 U14043 ( .B1(n11588), .B2(n7799), .A(n13405), .ZN(n11591) );
  OAI22_X1 U14044 ( .A1(n11605), .A2(n13404), .B1(n11607), .B2(n13408), .ZN(
        n11589) );
  AOI21_X1 U14045 ( .B1(n11591), .B2(n11590), .A(n11589), .ZN(n14424) );
  OAI21_X1 U14046 ( .B1(n11593), .B2(n7799), .A(n11592), .ZN(n14427) );
  NAND2_X1 U14047 ( .A1(n14427), .A2(n13373), .ZN(n11601) );
  OAI22_X1 U14048 ( .A1(n13427), .A2(n11594), .B1(n11606), .B2(n13412), .ZN(
        n11599) );
  INV_X1 U14049 ( .A(n11610), .ZN(n14425) );
  INV_X1 U14050 ( .A(n11595), .ZN(n11597) );
  INV_X1 U14051 ( .A(n13418), .ZN(n11596) );
  OAI211_X1 U14052 ( .C1(n14425), .C2(n11597), .A(n11596), .B(n13420), .ZN(
        n14423) );
  NOR2_X1 U14053 ( .A1(n14423), .A2(n13269), .ZN(n11598) );
  AOI211_X1 U14054 ( .C1(n13416), .C2(n11610), .A(n11599), .B(n11598), .ZN(
        n11600) );
  OAI211_X1 U14055 ( .C1(n13384), .C2(n14424), .A(n11601), .B(n11600), .ZN(
        P2_U3250) );
  XNOR2_X1 U14056 ( .A(n11603), .B(n11602), .ZN(n11612) );
  OAI22_X1 U14057 ( .A1(n13095), .A2(n11605), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11604), .ZN(n11609) );
  OAI22_X1 U14058 ( .A1(n13097), .A2(n11607), .B1(n13096), .B2(n11606), .ZN(
        n11608) );
  AOI211_X1 U14059 ( .C1(n11610), .C2(n13086), .A(n11609), .B(n11608), .ZN(
        n11611) );
  OAI21_X1 U14060 ( .B1(n11612), .B2(n13088), .A(n11611), .ZN(P2_U3213) );
  NAND2_X1 U14061 ( .A1(n11614), .A2(n11613), .ZN(n11615) );
  XNOR2_X1 U14062 ( .A(n11615), .B(n11680), .ZN(n11622) );
  INV_X1 U14063 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11616) );
  NOR2_X1 U14064 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11616), .ZN(n14929) );
  OAI22_X1 U14065 ( .A1(n12395), .A2(n14413), .B1(n12390), .B2(n11617), .ZN(
        n11618) );
  AOI211_X1 U14066 ( .C1(n14860), .C2(n12406), .A(n14929), .B(n11618), .ZN(
        n11621) );
  NAND2_X1 U14067 ( .A1(n12392), .A2(n11619), .ZN(n11620) );
  OAI211_X1 U14068 ( .C1(n11622), .C2(n12382), .A(n11621), .B(n11620), .ZN(
        P3_U3176) );
  OAI211_X1 U14069 ( .C1(n11625), .C2(n11624), .A(n11623), .B(n15089), .ZN(
        n11627) );
  AOI22_X1 U14070 ( .A1(n15081), .A2(n12403), .B1(n12405), .B2(n15084), .ZN(
        n11626) );
  AND2_X1 U14071 ( .A1(n11627), .A2(n11626), .ZN(n12891) );
  XNOR2_X1 U14072 ( .A(n11629), .B(n11628), .ZN(n12889) );
  INV_X1 U14073 ( .A(n11630), .ZN(n12960) );
  AOI22_X1 U14074 ( .A1(n15005), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15103), 
        .B2(n12275), .ZN(n11631) );
  OAI21_X1 U14075 ( .B1(n12960), .B2(n12826), .A(n11631), .ZN(n11632) );
  AOI21_X1 U14076 ( .B1(n12889), .B2(n15020), .A(n11632), .ZN(n11633) );
  OAI21_X1 U14077 ( .B1(n12891), .B2(n15005), .A(n11633), .ZN(P3_U3219) );
  XNOR2_X1 U14078 ( .A(n11634), .B(n12406), .ZN(n11635) );
  XNOR2_X1 U14079 ( .A(n11636), .B(n11635), .ZN(n11642) );
  NAND2_X1 U14080 ( .A1(n12392), .A2(n11637), .ZN(n11639) );
  AND2_X1 U14081 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n14947) );
  AOI21_X1 U14082 ( .B1(n14860), .B2(n12405), .A(n14947), .ZN(n11638) );
  OAI211_X1 U14083 ( .C1(n11680), .C2(n12390), .A(n11639), .B(n11638), .ZN(
        n11640) );
  AOI21_X1 U14084 ( .B1(n14401), .B2(n14859), .A(n11640), .ZN(n11641) );
  OAI21_X1 U14085 ( .B1(n11642), .B2(n12382), .A(n11641), .ZN(P3_U3164) );
  INV_X1 U14086 ( .A(n14304), .ZN(n14314) );
  NOR2_X1 U14087 ( .A1(n9756), .A2(n11643), .ZN(n11644) );
  AOI21_X1 U14088 ( .B1(n14474), .B2(n11863), .A(n11644), .ZN(n11660) );
  NAND2_X1 U14089 ( .A1(n14474), .A2(n11929), .ZN(n11646) );
  NAND2_X1 U14090 ( .A1(n11863), .A2(n13724), .ZN(n11645) );
  NAND2_X1 U14091 ( .A1(n11646), .A2(n11645), .ZN(n11647) );
  XNOR2_X1 U14092 ( .A(n11647), .B(n12232), .ZN(n11659) );
  OR2_X1 U14093 ( .A1(n11649), .A2(n11648), .ZN(n11650) );
  AOI22_X1 U14094 ( .A1(n13595), .A2(n11929), .B1(n11863), .B2(n13725), .ZN(
        n11653) );
  XNOR2_X1 U14095 ( .A(n11653), .B(n11652), .ZN(n11656) );
  NOR2_X1 U14096 ( .A1(n9756), .A2(n11654), .ZN(n11655) );
  AOI21_X1 U14097 ( .B1(n13595), .B2(n11863), .A(n11655), .ZN(n11657) );
  XNOR2_X1 U14098 ( .A(n11656), .B(n11657), .ZN(n13590) );
  INV_X1 U14099 ( .A(n11656), .ZN(n11658) );
  NOR2_X1 U14100 ( .A1(n11658), .A2(n11657), .ZN(n14468) );
  XNOR2_X1 U14101 ( .A(n11659), .B(n11660), .ZN(n14467) );
  NOR2_X1 U14102 ( .A1(n9756), .A2(n11661), .ZN(n11662) );
  AOI21_X1 U14103 ( .B1(n14304), .B2(n11863), .A(n11662), .ZN(n11712) );
  NAND2_X1 U14104 ( .A1(n14304), .A2(n11929), .ZN(n11664) );
  NAND2_X1 U14105 ( .A1(n11863), .A2(n13723), .ZN(n11663) );
  NAND2_X1 U14106 ( .A1(n11664), .A2(n11663), .ZN(n11665) );
  XNOR2_X1 U14107 ( .A(n11665), .B(n12232), .ZN(n11713) );
  XOR2_X1 U14108 ( .A(n11712), .B(n11713), .Z(n11666) );
  OAI211_X1 U14109 ( .C1(n11667), .C2(n11666), .A(n6609), .B(n14470), .ZN(
        n11674) );
  INV_X1 U14110 ( .A(n11668), .ZN(n14303) );
  NAND2_X1 U14111 ( .A1(n13724), .A2(n14100), .ZN(n11670) );
  NAND2_X1 U14112 ( .A1(n14101), .A2(n13691), .ZN(n11669) );
  AND2_X1 U14113 ( .A1(n11670), .A2(n11669), .ZN(n14302) );
  OAI22_X1 U14114 ( .A1(n13712), .A2(n14302), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11671), .ZN(n11672) );
  AOI21_X1 U14115 ( .B1(n14303), .B2(n13714), .A(n11672), .ZN(n11673) );
  OAI211_X1 U14116 ( .C1(n14314), .C2(n13718), .A(n11674), .B(n11673), .ZN(
        P1_U3224) );
  OAI21_X1 U14117 ( .B1(n11676), .B2(n11677), .A(n11675), .ZN(n14400) );
  XOR2_X1 U14118 ( .A(n11678), .B(n11677), .Z(n11679) );
  OAI222_X1 U14119 ( .A1(n15046), .A2(n12273), .B1(n15044), .B2(n11680), .C1(
        n11679), .C2(n15052), .ZN(n14399) );
  AOI21_X1 U14120 ( .B1(n15136), .B2(n14400), .A(n14399), .ZN(n11682) );
  MUX2_X1 U14121 ( .A(n8360), .B(n11682), .S(n15143), .Z(n11681) );
  OAI21_X1 U14122 ( .B1(n12965), .B2(n11684), .A(n11681), .ZN(P3_U3426) );
  INV_X1 U14123 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12420) );
  MUX2_X1 U14124 ( .A(n12420), .B(n11682), .S(n15159), .Z(n11683) );
  OAI21_X1 U14125 ( .B1(n12899), .B2(n11684), .A(n11683), .ZN(P3_U3471) );
  NAND2_X1 U14126 ( .A1(n11686), .A2(n11085), .ZN(n11689) );
  AOI22_X1 U14127 ( .A1(n11774), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11773), 
        .B2(n11687), .ZN(n11688) );
  XNOR2_X1 U14128 ( .A(n14197), .B(n13880), .ZN(n12200) );
  XNOR2_X1 U14129 ( .A(n13883), .B(n13882), .ZN(n11698) );
  INV_X1 U14130 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11696) );
  INV_X1 U14131 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11691) );
  NAND2_X1 U14132 ( .A1(n11692), .A2(n11691), .ZN(n11693) );
  NAND2_X1 U14133 ( .A1(n11757), .A2(n11693), .ZN(n13641) );
  OR2_X1 U14134 ( .A1(n13641), .A2(n9744), .ZN(n11695) );
  AOI22_X1 U14135 ( .A1(n11548), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n12154), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n11694) );
  OAI211_X1 U14136 ( .C1(n11923), .C2(n11696), .A(n11695), .B(n11694), .ZN(
        n13884) );
  INV_X1 U14137 ( .A(n14099), .ZN(n13721) );
  AOI22_X1 U14138 ( .A1(n13884), .A2(n13854), .B1(n13721), .B2(n14100), .ZN(
        n13632) );
  INV_X1 U14139 ( .A(n13632), .ZN(n11697) );
  AOI21_X1 U14140 ( .B1(n11698), .B2(n14625), .A(n11697), .ZN(n14199) );
  INV_X1 U14141 ( .A(n11699), .ZN(n11701) );
  INV_X1 U14142 ( .A(n14197), .ZN(n13881) );
  INV_X1 U14143 ( .A(n14084), .ZN(n11700) );
  AOI211_X1 U14144 ( .C1(n14197), .C2(n11701), .A(n14575), .B(n11700), .ZN(
        n14196) );
  INV_X1 U14145 ( .A(n13630), .ZN(n11702) );
  AOI22_X1 U14146 ( .A1(n14599), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11702), 
        .B2(n14586), .ZN(n11703) );
  OAI21_X1 U14147 ( .B1(n13881), .B2(n14088), .A(n11703), .ZN(n11707) );
  XNOR2_X1 U14148 ( .A(n13865), .B(n12200), .ZN(n14200) );
  NOR2_X1 U14149 ( .A1(n14200), .A2(n14092), .ZN(n11706) );
  AOI211_X1 U14150 ( .C1(n14196), .C2(n14595), .A(n11707), .B(n11706), .ZN(
        n11708) );
  OAI21_X1 U14151 ( .B1(n14599), .B2(n14199), .A(n11708), .ZN(P1_U3277) );
  INV_X1 U14152 ( .A(n12147), .ZN(n11945) );
  OAI222_X1 U14153 ( .A1(n14244), .A2(n11945), .B1(n11709), .B2(P1_U3086), 
        .C1(n12148), .C2(n14245), .ZN(P1_U3326) );
  NAND2_X1 U14154 ( .A1(n13562), .A2(n11085), .ZN(n11711) );
  OR2_X1 U14155 ( .A1(n12160), .A2(n7103), .ZN(n11710) );
  OR2_X1 U14156 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  AOI22_X1 U14157 ( .A1(n12068), .A2(n11929), .B1(n11863), .B2(n14101), .ZN(
        n11716) );
  XNOR2_X1 U14158 ( .A(n11716), .B(n12232), .ZN(n11727) );
  NOR2_X1 U14159 ( .A1(n9756), .A2(n11717), .ZN(n11718) );
  AOI21_X1 U14160 ( .B1(n12068), .B2(n11863), .A(n11718), .ZN(n11725) );
  XNOR2_X1 U14161 ( .A(n11727), .B(n11725), .ZN(n13662) );
  NAND2_X1 U14162 ( .A1(n14481), .A2(n11929), .ZN(n11720) );
  OR2_X1 U14163 ( .A1(n11723), .A2(n9728), .ZN(n11719) );
  NAND2_X1 U14164 ( .A1(n11720), .A2(n11719), .ZN(n11722) );
  XNOR2_X1 U14165 ( .A(n11722), .B(n11721), .ZN(n11731) );
  NOR2_X1 U14166 ( .A1(n9756), .A2(n11723), .ZN(n11724) );
  AOI21_X1 U14167 ( .B1(n14481), .B2(n11863), .A(n11724), .ZN(n11729) );
  XNOR2_X1 U14168 ( .A(n11731), .B(n11729), .ZN(n14461) );
  INV_X1 U14169 ( .A(n11725), .ZN(n11726) );
  NAND2_X1 U14170 ( .A1(n11727), .A2(n11726), .ZN(n14458) );
  INV_X1 U14171 ( .A(n11729), .ZN(n11730) );
  OAI22_X1 U14172 ( .A1(n14202), .A2(n9737), .B1(n14099), .B2(n9728), .ZN(
        n11732) );
  XOR2_X1 U14173 ( .A(n12232), .B(n11732), .Z(n11734) );
  XNOR2_X1 U14174 ( .A(n11733), .B(n11734), .ZN(n13710) );
  OAI22_X1 U14175 ( .A1(n14202), .A2(n9728), .B1(n14099), .B2(n9756), .ZN(
        n13709) );
  INV_X1 U14176 ( .A(n11733), .ZN(n11735) );
  NAND2_X1 U14177 ( .A1(n11735), .A2(n11734), .ZN(n11736) );
  AOI22_X1 U14178 ( .A1(n14197), .A2(n11863), .B1(n11928), .B2(n13880), .ZN(
        n11739) );
  AOI22_X1 U14179 ( .A1(n14197), .A2(n11929), .B1(n11863), .B2(n13880), .ZN(
        n11737) );
  XNOR2_X1 U14180 ( .A(n11737), .B(n12232), .ZN(n11738) );
  XOR2_X1 U14181 ( .A(n11739), .B(n11738), .Z(n13629) );
  INV_X1 U14182 ( .A(n11738), .ZN(n11740) );
  NAND2_X1 U14183 ( .A1(n11740), .A2(n11739), .ZN(n11741) );
  NAND2_X1 U14184 ( .A1(n11742), .A2(n11085), .ZN(n11745) );
  AOI22_X1 U14185 ( .A1(n11774), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11773), 
        .B2(n11743), .ZN(n11744) );
  AOI22_X1 U14186 ( .A1(n14192), .A2(n11863), .B1(n11928), .B2(n13884), .ZN(
        n11750) );
  NAND2_X1 U14187 ( .A1(n14192), .A2(n11929), .ZN(n11748) );
  NAND2_X1 U14188 ( .A1(n13884), .A2(n11863), .ZN(n11747) );
  NAND2_X1 U14189 ( .A1(n11748), .A2(n11747), .ZN(n11749) );
  XNOR2_X1 U14190 ( .A(n11749), .B(n12232), .ZN(n11751) );
  XOR2_X1 U14191 ( .A(n11750), .B(n11751), .Z(n13639) );
  NAND2_X1 U14192 ( .A1(n11751), .A2(n11750), .ZN(n11752) );
  OR2_X1 U14193 ( .A1(n11753), .A2(n6647), .ZN(n11755) );
  AOI22_X1 U14194 ( .A1(n11774), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11773), 
        .B2(n13837), .ZN(n11754) );
  INV_X1 U14195 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11756) );
  NAND2_X1 U14196 ( .A1(n11757), .A2(n11756), .ZN(n11758) );
  NAND2_X1 U14197 ( .A1(n11778), .A2(n11758), .ZN(n14072) );
  OR2_X1 U14198 ( .A1(n14072), .A2(n9744), .ZN(n11765) );
  INV_X1 U14199 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U14200 ( .A1(n12154), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11761) );
  INV_X1 U14201 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n11759) );
  OR2_X1 U14202 ( .A1(n11923), .A2(n11759), .ZN(n11760) );
  OAI211_X1 U14203 ( .C1(n12167), .C2(n11762), .A(n11761), .B(n11760), .ZN(
        n11763) );
  INV_X1 U14204 ( .A(n11763), .ZN(n11764) );
  NAND2_X1 U14205 ( .A1(n11765), .A2(n11764), .ZN(n13886) );
  AOI22_X1 U14206 ( .A1(n14187), .A2(n11863), .B1(n11928), .B2(n13886), .ZN(
        n11769) );
  NAND2_X1 U14207 ( .A1(n14187), .A2(n11929), .ZN(n11767) );
  NAND2_X1 U14208 ( .A1(n13886), .A2(n11863), .ZN(n11766) );
  NAND2_X1 U14209 ( .A1(n11767), .A2(n11766), .ZN(n11768) );
  XNOR2_X1 U14210 ( .A(n11768), .B(n12232), .ZN(n11770) );
  XOR2_X1 U14211 ( .A(n11769), .B(n11770), .Z(n13679) );
  NAND2_X1 U14212 ( .A1(n11770), .A2(n11769), .ZN(n11771) );
  NAND2_X1 U14213 ( .A1(n11772), .A2(n11085), .ZN(n11776) );
  AOI22_X1 U14214 ( .A1(n11774), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14559), 
        .B2(n11773), .ZN(n11775) );
  NAND2_X1 U14215 ( .A1(n14060), .A2(n11929), .ZN(n11787) );
  INV_X1 U14216 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11777) );
  NAND2_X1 U14217 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  AND2_X1 U14218 ( .A1(n11798), .A2(n11779), .ZN(n14055) );
  NAND2_X1 U14219 ( .A1(n14055), .A2(n11933), .ZN(n11785) );
  INV_X1 U14220 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n11782) );
  NAND2_X1 U14221 ( .A1(n12154), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11781) );
  NAND2_X1 U14222 ( .A1(n12164), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11780) );
  OAI211_X1 U14223 ( .C1(n12167), .C2(n11782), .A(n11781), .B(n11780), .ZN(
        n11783) );
  INV_X1 U14224 ( .A(n11783), .ZN(n11784) );
  NAND2_X1 U14225 ( .A1(n13887), .A2(n11863), .ZN(n11786) );
  NAND2_X1 U14226 ( .A1(n11787), .A2(n11786), .ZN(n11788) );
  XNOR2_X1 U14227 ( .A(n11788), .B(n12232), .ZN(n11792) );
  NOR2_X1 U14228 ( .A1(n13682), .A2(n9756), .ZN(n11789) );
  AOI21_X1 U14229 ( .B1(n14060), .B2(n11863), .A(n11789), .ZN(n11791) );
  XNOR2_X1 U14230 ( .A(n11792), .B(n11791), .ZN(n13601) );
  INV_X1 U14231 ( .A(n13601), .ZN(n11790) );
  OR2_X1 U14232 ( .A1(n11792), .A2(n11791), .ZN(n11793) );
  OR2_X1 U14233 ( .A1(n11794), .A2(n6647), .ZN(n11796) );
  OR2_X1 U14234 ( .A1(n12160), .A2(n7077), .ZN(n11795) );
  INV_X1 U14235 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13658) );
  NAND2_X1 U14236 ( .A1(n11798), .A2(n13658), .ZN(n11799) );
  AND2_X1 U14237 ( .A1(n11818), .A2(n11799), .ZN(n14038) );
  NAND2_X1 U14238 ( .A1(n14038), .A2(n11933), .ZN(n11805) );
  INV_X1 U14239 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n11802) );
  NAND2_X1 U14240 ( .A1(n12154), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U14241 ( .A1(n12164), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11800) );
  OAI211_X1 U14242 ( .C1(n12167), .C2(n11802), .A(n11801), .B(n11800), .ZN(
        n11803) );
  INV_X1 U14243 ( .A(n11803), .ZN(n11804) );
  NAND2_X1 U14244 ( .A1(n11805), .A2(n11804), .ZN(n13888) );
  AOI22_X1 U14245 ( .A1(n14175), .A2(n11929), .B1(n11863), .B2(n13888), .ZN(
        n11806) );
  XNOR2_X1 U14246 ( .A(n11806), .B(n12232), .ZN(n11810) );
  AND2_X1 U14247 ( .A1(n13888), .A2(n11928), .ZN(n11807) );
  AOI21_X1 U14248 ( .B1(n14175), .B2(n11863), .A(n11807), .ZN(n11808) );
  XNOR2_X1 U14249 ( .A(n11810), .B(n11808), .ZN(n13656) );
  INV_X1 U14250 ( .A(n11808), .ZN(n11809) );
  NAND2_X1 U14251 ( .A1(n11810), .A2(n11809), .ZN(n11811) );
  NAND2_X1 U14252 ( .A1(n11812), .A2(n11085), .ZN(n11815) );
  OR2_X1 U14253 ( .A1(n12160), .A2(n11813), .ZN(n11814) );
  INV_X1 U14254 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n11817) );
  NAND2_X1 U14255 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  NAND2_X1 U14256 ( .A1(n11836), .A2(n11819), .ZN(n14024) );
  OR2_X1 U14257 ( .A1(n14024), .A2(n9744), .ZN(n11825) );
  INV_X1 U14258 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n11822) );
  NAND2_X1 U14259 ( .A1(n12154), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11821) );
  NAND2_X1 U14260 ( .A1(n12164), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11820) );
  OAI211_X1 U14261 ( .C1(n12167), .C2(n11822), .A(n11821), .B(n11820), .ZN(
        n11823) );
  INV_X1 U14262 ( .A(n11823), .ZN(n11824) );
  AOI22_X1 U14263 ( .A1(n14170), .A2(n11863), .B1(n11928), .B2(n13874), .ZN(
        n11829) );
  AOI22_X1 U14264 ( .A1(n14170), .A2(n11929), .B1(n11863), .B2(n13874), .ZN(
        n11826) );
  XNOR2_X1 U14265 ( .A(n11826), .B(n12232), .ZN(n11828) );
  XOR2_X1 U14266 ( .A(n11829), .B(n11828), .Z(n13612) );
  INV_X1 U14267 ( .A(n11828), .ZN(n11830) );
  NAND2_X1 U14268 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  INV_X1 U14269 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U14270 ( .A1(n11836), .A2(n13675), .ZN(n11837) );
  AND2_X1 U14271 ( .A1(n11856), .A2(n11837), .ZN(n14005) );
  NAND2_X1 U14272 ( .A1(n14005), .A2(n11933), .ZN(n11843) );
  INV_X1 U14273 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11840) );
  NAND2_X1 U14274 ( .A1(n12154), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11839) );
  NAND2_X1 U14275 ( .A1(n12164), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11838) );
  OAI211_X1 U14276 ( .C1(n12167), .C2(n11840), .A(n11839), .B(n11838), .ZN(
        n11841) );
  INV_X1 U14277 ( .A(n11841), .ZN(n11842) );
  OAI22_X1 U14278 ( .A1(n14007), .A2(n9737), .B1(n13875), .B2(n9728), .ZN(
        n11844) );
  XNOR2_X1 U14279 ( .A(n11844), .B(n12232), .ZN(n11845) );
  OAI22_X1 U14280 ( .A1(n14007), .A2(n9728), .B1(n13875), .B2(n9756), .ZN(
        n11846) );
  XNOR2_X1 U14281 ( .A(n11845), .B(n11846), .ZN(n13672) );
  NAND2_X1 U14282 ( .A1(n13671), .A2(n13672), .ZN(n13670) );
  INV_X1 U14283 ( .A(n11845), .ZN(n11847) );
  OR2_X1 U14284 ( .A1(n11847), .A2(n11846), .ZN(n11848) );
  OR2_X1 U14285 ( .A1(n12160), .A2(n11851), .ZN(n11852) );
  INV_X1 U14286 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n11855) );
  NAND2_X1 U14287 ( .A1(n11856), .A2(n11855), .ZN(n11857) );
  NAND2_X1 U14288 ( .A1(n11872), .A2(n11857), .ZN(n13992) );
  INV_X1 U14289 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U14290 ( .A1(n12154), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11859) );
  NAND2_X1 U14291 ( .A1(n11548), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11858) );
  OAI211_X1 U14292 ( .C1(n12685), .C2(n11923), .A(n11859), .B(n11858), .ZN(
        n11860) );
  INV_X1 U14293 ( .A(n11860), .ZN(n11861) );
  AOI22_X1 U14294 ( .A1(n14159), .A2(n11863), .B1(n11928), .B2(n13876), .ZN(
        n11867) );
  NAND2_X1 U14295 ( .A1(n14159), .A2(n11929), .ZN(n11865) );
  NAND2_X1 U14296 ( .A1(n13876), .A2(n11863), .ZN(n11864) );
  NAND2_X1 U14297 ( .A1(n11865), .A2(n11864), .ZN(n11866) );
  XNOR2_X1 U14298 ( .A(n11866), .B(n12232), .ZN(n11868) );
  XOR2_X1 U14299 ( .A(n11867), .B(n11868), .Z(n13579) );
  NAND2_X1 U14300 ( .A1(n11868), .A2(n11867), .ZN(n11869) );
  OR2_X1 U14301 ( .A1(n12160), .A2(n14246), .ZN(n11870) );
  INV_X1 U14302 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13650) );
  NAND2_X1 U14303 ( .A1(n11872), .A2(n13650), .ZN(n11873) );
  AND2_X1 U14304 ( .A1(n11887), .A2(n11873), .ZN(n13982) );
  NAND2_X1 U14305 ( .A1(n13982), .A2(n11933), .ZN(n11878) );
  INV_X1 U14306 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n12653) );
  NAND2_X1 U14307 ( .A1(n12154), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U14308 ( .A1(n11548), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11874) );
  OAI211_X1 U14309 ( .C1(n12653), .C2(n11923), .A(n11875), .B(n11874), .ZN(
        n11876) );
  INV_X1 U14310 ( .A(n11876), .ZN(n11877) );
  AOI22_X1 U14311 ( .A1(n13983), .A2(n11863), .B1(n11928), .B2(n13893), .ZN(
        n11882) );
  NAND2_X1 U14312 ( .A1(n13983), .A2(n11929), .ZN(n11880) );
  NAND2_X1 U14313 ( .A1(n13893), .A2(n11863), .ZN(n11879) );
  NAND2_X1 U14314 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  XNOR2_X1 U14315 ( .A(n11881), .B(n12232), .ZN(n11883) );
  XOR2_X1 U14316 ( .A(n11882), .B(n11883), .Z(n13648) );
  OR2_X1 U14317 ( .A1(n12160), .A2(n6685), .ZN(n11884) );
  INV_X1 U14318 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11886) );
  NAND2_X1 U14319 ( .A1(n11887), .A2(n11886), .ZN(n11888) );
  NAND2_X1 U14320 ( .A1(n13965), .A2(n11933), .ZN(n11894) );
  INV_X1 U14321 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U14322 ( .A1(n12154), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11890) );
  NAND2_X1 U14323 ( .A1(n12164), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11889) );
  OAI211_X1 U14324 ( .C1(n12167), .C2(n11891), .A(n11890), .B(n11889), .ZN(
        n11892) );
  INV_X1 U14325 ( .A(n11892), .ZN(n11893) );
  AOI22_X1 U14326 ( .A1(n13969), .A2(n11863), .B1(n11928), .B2(n13894), .ZN(
        n11898) );
  NAND2_X1 U14327 ( .A1(n13969), .A2(n11929), .ZN(n11896) );
  NAND2_X1 U14328 ( .A1(n13894), .A2(n11863), .ZN(n11895) );
  NAND2_X1 U14329 ( .A1(n11896), .A2(n11895), .ZN(n11897) );
  XNOR2_X1 U14330 ( .A(n11897), .B(n12232), .ZN(n11899) );
  XOR2_X1 U14331 ( .A(n11898), .B(n11899), .Z(n13620) );
  NAND2_X1 U14332 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  NAND2_X1 U14333 ( .A1(n13565), .A2(n11085), .ZN(n11902) );
  OR2_X1 U14334 ( .A1(n12160), .A2(n6709), .ZN(n11901) );
  NAND2_X2 U14335 ( .A1(n11902), .A2(n11901), .ZN(n14142) );
  INV_X1 U14336 ( .A(n11905), .ZN(n11903) );
  NAND2_X1 U14337 ( .A1(n11903), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11919) );
  INV_X1 U14338 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11904) );
  NAND2_X1 U14339 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  NAND2_X1 U14340 ( .A1(n11919), .A2(n11906), .ZN(n13949) );
  OR2_X1 U14341 ( .A1(n13949), .A2(n9744), .ZN(n11912) );
  INV_X1 U14342 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n11909) );
  NAND2_X1 U14343 ( .A1(n12154), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11908) );
  NAND2_X1 U14344 ( .A1(n12164), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11907) );
  OAI211_X1 U14345 ( .C1(n12167), .C2(n11909), .A(n11908), .B(n11907), .ZN(
        n11910) );
  INV_X1 U14346 ( .A(n11910), .ZN(n11911) );
  AOI22_X1 U14347 ( .A1(n14142), .A2(n11863), .B1(n11928), .B2(n13720), .ZN(
        n11916) );
  NAND2_X1 U14348 ( .A1(n14142), .A2(n11929), .ZN(n11914) );
  NAND2_X1 U14349 ( .A1(n13720), .A2(n11863), .ZN(n11913) );
  NAND2_X1 U14350 ( .A1(n11914), .A2(n11913), .ZN(n11915) );
  XNOR2_X1 U14351 ( .A(n11915), .B(n12232), .ZN(n11917) );
  XOR2_X1 U14352 ( .A(n11916), .B(n11917), .Z(n13699) );
  NAND2_X1 U14353 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  INV_X1 U14354 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11940) );
  NAND2_X1 U14355 ( .A1(n11919), .A2(n11940), .ZN(n11920) );
  NAND2_X1 U14356 ( .A1(n13937), .A2(n11933), .ZN(n11927) );
  INV_X1 U14357 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U14358 ( .A1(n12154), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11922) );
  NAND2_X1 U14359 ( .A1(n11548), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11921) );
  OAI211_X1 U14360 ( .C1(n11924), .C2(n11923), .A(n11922), .B(n11921), .ZN(
        n11925) );
  INV_X1 U14361 ( .A(n11925), .ZN(n11926) );
  AOI22_X1 U14362 ( .A1(n6701), .A2(n11863), .B1(n11928), .B2(n13896), .ZN(
        n12229) );
  NAND2_X1 U14363 ( .A1(n14135), .A2(n11929), .ZN(n11931) );
  NAND2_X1 U14364 ( .A1(n13896), .A2(n11863), .ZN(n11930) );
  NAND2_X1 U14365 ( .A1(n11931), .A2(n11930), .ZN(n11932) );
  XNOR2_X1 U14366 ( .A(n11932), .B(n12232), .ZN(n12230) );
  XOR2_X1 U14367 ( .A(n12229), .B(n12230), .Z(n12231) );
  XNOR2_X1 U14368 ( .A(n13909), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n13923) );
  NAND2_X1 U14369 ( .A1(n13923), .A2(n11933), .ZN(n11939) );
  INV_X1 U14370 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n11936) );
  NAND2_X1 U14371 ( .A1(n12154), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11935) );
  NAND2_X1 U14372 ( .A1(n12164), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11934) );
  OAI211_X1 U14373 ( .C1(n12167), .C2(n11936), .A(n11935), .B(n11934), .ZN(
        n11937) );
  INV_X1 U14374 ( .A(n11937), .ZN(n11938) );
  OAI22_X1 U14375 ( .A1(n13904), .A2(n14098), .B1(n13895), .B2(n13903), .ZN(
        n13933) );
  INV_X1 U14376 ( .A(n13937), .ZN(n11941) );
  OAI22_X1 U14377 ( .A1(n11941), .A2(n14479), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11940), .ZN(n11942) );
  AOI21_X1 U14378 ( .B1(n13933), .B2(n14472), .A(n11942), .ZN(n11943) );
  OAI222_X1 U14379 ( .A1(P2_U3088), .A2(n11946), .B1(n13575), .B2(n11945), 
        .C1(n11944), .C2(n13573), .ZN(P2_U3298) );
  NAND2_X1 U14380 ( .A1(n13107), .A2(n9498), .ZN(n11950) );
  INV_X1 U14381 ( .A(n11950), .ZN(n11952) );
  XNOR2_X1 U14382 ( .A(n13229), .B(n6712), .ZN(n11951) );
  INV_X1 U14383 ( .A(n11947), .ZN(n11948) );
  XNOR2_X1 U14384 ( .A(n11951), .B(n11950), .ZN(n13091) );
  XNOR2_X1 U14385 ( .A(n13444), .B(n6712), .ZN(n11954) );
  AND2_X1 U14386 ( .A1(n13106), .A2(n13394), .ZN(n11953) );
  NAND2_X1 U14387 ( .A1(n11954), .A2(n11953), .ZN(n13023) );
  OAI21_X1 U14388 ( .B1(n11954), .B2(n11953), .A(n13023), .ZN(n11955) );
  OAI22_X1 U14389 ( .A1(n11957), .A2(n13408), .B1(n13243), .B2(n13404), .ZN(
        n13208) );
  AOI22_X1 U14390 ( .A1(n13208), .A2(n13056), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11958) );
  OAI21_X1 U14391 ( .B1(n13212), .B2(n13096), .A(n11958), .ZN(n11959) );
  INV_X1 U14392 ( .A(n11959), .ZN(n11960) );
  NAND2_X1 U14393 ( .A1(n14226), .A2(n11085), .ZN(n11965) );
  OR2_X1 U14394 ( .A1(n12160), .A2(n14231), .ZN(n11964) );
  NAND2_X1 U14395 ( .A1(n11971), .A2(n11982), .ZN(n11967) );
  OAI21_X1 U14396 ( .B1(n11971), .B2(n11970), .A(n9777), .ZN(n11972) );
  NOR2_X1 U14397 ( .A1(n13856), .A2(n12128), .ZN(n12212) );
  INV_X1 U14398 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n11975) );
  NAND2_X1 U14399 ( .A1(n12164), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11974) );
  NAND2_X1 U14400 ( .A1(n12154), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11973) );
  OAI211_X1 U14401 ( .C1(n12167), .C2(n11975), .A(n11974), .B(n11973), .ZN(
        n13855) );
  NAND2_X1 U14402 ( .A1(n11977), .A2(n11976), .ZN(n11978) );
  NAND2_X1 U14403 ( .A1(n11979), .A2(n11978), .ZN(n11980) );
  NAND2_X1 U14404 ( .A1(n11981), .A2(n11980), .ZN(n12219) );
  NAND2_X1 U14405 ( .A1(n9777), .A2(n11982), .ZN(n12216) );
  NAND2_X1 U14406 ( .A1(n12219), .A2(n12216), .ZN(n12208) );
  NAND2_X1 U14407 ( .A1(n13856), .A2(n12128), .ZN(n12210) );
  NOR2_X1 U14408 ( .A1(n12210), .A2(n13855), .ZN(n11983) );
  AOI211_X1 U14409 ( .C1(n12212), .C2(n13855), .A(n12208), .B(n11983), .ZN(
        n11984) );
  MUX2_X1 U14410 ( .A(n13896), .B(n14135), .S(n12173), .Z(n12139) );
  MUX2_X1 U14411 ( .A(n13880), .B(n14197), .S(n12173), .Z(n12084) );
  MUX2_X1 U14412 ( .A(n14101), .B(n12068), .S(n12173), .Z(n12070) );
  NAND2_X1 U14413 ( .A1(n12184), .A2(n11985), .ZN(n11987) );
  NAND2_X1 U14414 ( .A1(n11987), .A2(n11986), .ZN(n11996) );
  INV_X1 U14415 ( .A(n11988), .ZN(n11991) );
  NAND2_X1 U14416 ( .A1(n11989), .A2(n12037), .ZN(n11990) );
  OAI21_X1 U14417 ( .B1(n11991), .B2(n12037), .A(n11990), .ZN(n11995) );
  MUX2_X1 U14418 ( .A(n13734), .B(n11992), .S(n12037), .Z(n11993) );
  OAI22_X1 U14419 ( .A1(n11996), .A2(n11995), .B1(n11994), .B2(n11993), .ZN(
        n11999) );
  MUX2_X1 U14420 ( .A(n13733), .B(n14589), .S(n12037), .Z(n12000) );
  NAND2_X1 U14421 ( .A1(n13733), .A2(n14589), .ZN(n11997) );
  NAND2_X1 U14422 ( .A1(n12000), .A2(n11997), .ZN(n11998) );
  NAND2_X1 U14423 ( .A1(n11999), .A2(n11998), .ZN(n12005) );
  INV_X1 U14424 ( .A(n12000), .ZN(n12002) );
  NAND2_X1 U14425 ( .A1(n12002), .A2(n12001), .ZN(n12004) );
  NAND2_X1 U14426 ( .A1(n12005), .A2(n7419), .ZN(n12010) );
  MUX2_X1 U14427 ( .A(n14623), .B(n12006), .S(n12037), .Z(n12008) );
  NAND2_X1 U14428 ( .A1(n12008), .A2(n12007), .ZN(n12009) );
  MUX2_X1 U14429 ( .A(n14634), .B(n12011), .S(n12037), .Z(n12013) );
  OAI21_X1 U14430 ( .B1(n12014), .B2(n12013), .A(n12012), .ZN(n12016) );
  NAND2_X1 U14431 ( .A1(n12014), .A2(n12013), .ZN(n12015) );
  NAND2_X1 U14432 ( .A1(n12016), .A2(n12015), .ZN(n12019) );
  MUX2_X1 U14433 ( .A(n13730), .B(n14641), .S(n12173), .Z(n12020) );
  NAND2_X1 U14434 ( .A1(n12019), .A2(n12020), .ZN(n12018) );
  MUX2_X1 U14435 ( .A(n14641), .B(n13730), .S(n12173), .Z(n12017) );
  NAND2_X1 U14436 ( .A1(n12018), .A2(n12017), .ZN(n12024) );
  INV_X1 U14437 ( .A(n12019), .ZN(n12022) );
  INV_X1 U14438 ( .A(n12020), .ZN(n12021) );
  NAND2_X1 U14439 ( .A1(n12022), .A2(n12021), .ZN(n12023) );
  NAND2_X1 U14440 ( .A1(n12024), .A2(n12023), .ZN(n12027) );
  MUX2_X1 U14441 ( .A(n13729), .B(n14651), .S(n12033), .Z(n12028) );
  NAND2_X1 U14442 ( .A1(n12027), .A2(n12028), .ZN(n12026) );
  MUX2_X1 U14443 ( .A(n13729), .B(n14651), .S(n12173), .Z(n12025) );
  NAND2_X1 U14444 ( .A1(n12026), .A2(n12025), .ZN(n12032) );
  INV_X1 U14445 ( .A(n12027), .ZN(n12030) );
  INV_X1 U14446 ( .A(n12028), .ZN(n12029) );
  NAND2_X1 U14447 ( .A1(n12030), .A2(n12029), .ZN(n12031) );
  MUX2_X1 U14448 ( .A(n13728), .B(n12034), .S(n12173), .Z(n12036) );
  MUX2_X1 U14449 ( .A(n13728), .B(n12034), .S(n12033), .Z(n12035) );
  MUX2_X1 U14450 ( .A(n13727), .B(n14666), .S(n12128), .Z(n12041) );
  NAND2_X1 U14451 ( .A1(n12040), .A2(n12041), .ZN(n12039) );
  MUX2_X1 U14452 ( .A(n13727), .B(n14666), .S(n12173), .Z(n12038) );
  NAND2_X1 U14453 ( .A1(n12039), .A2(n12038), .ZN(n12045) );
  INV_X1 U14454 ( .A(n12040), .ZN(n12043) );
  INV_X1 U14455 ( .A(n12041), .ZN(n12042) );
  NAND2_X1 U14456 ( .A1(n12043), .A2(n12042), .ZN(n12044) );
  MUX2_X1 U14457 ( .A(n13726), .B(n12046), .S(n12173), .Z(n12048) );
  MUX2_X1 U14458 ( .A(n13726), .B(n12046), .S(n12128), .Z(n12047) );
  INV_X1 U14459 ( .A(n12048), .ZN(n12049) );
  MUX2_X1 U14460 ( .A(n13725), .B(n13595), .S(n12128), .Z(n12053) );
  NAND2_X1 U14461 ( .A1(n12052), .A2(n12053), .ZN(n12051) );
  MUX2_X1 U14462 ( .A(n13725), .B(n13595), .S(n12173), .Z(n12050) );
  NAND2_X1 U14463 ( .A1(n12051), .A2(n12050), .ZN(n12057) );
  INV_X1 U14464 ( .A(n12052), .ZN(n12055) );
  INV_X1 U14465 ( .A(n12053), .ZN(n12054) );
  NAND2_X1 U14466 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  MUX2_X1 U14467 ( .A(n13724), .B(n14474), .S(n12173), .Z(n12059) );
  MUX2_X1 U14468 ( .A(n13724), .B(n14474), .S(n12128), .Z(n12058) );
  MUX2_X1 U14469 ( .A(n13723), .B(n14304), .S(n12128), .Z(n12063) );
  NAND2_X1 U14470 ( .A1(n12062), .A2(n12063), .ZN(n12061) );
  MUX2_X1 U14471 ( .A(n13723), .B(n14304), .S(n12173), .Z(n12060) );
  NAND2_X1 U14472 ( .A1(n12061), .A2(n12060), .ZN(n12067) );
  INV_X1 U14473 ( .A(n12062), .ZN(n12065) );
  INV_X1 U14474 ( .A(n12063), .ZN(n12064) );
  NAND2_X1 U14475 ( .A1(n12065), .A2(n12064), .ZN(n12066) );
  MUX2_X1 U14476 ( .A(n14101), .B(n12068), .S(n12128), .Z(n12069) );
  NAND2_X1 U14477 ( .A1(n12071), .A2(n14112), .ZN(n12077) );
  AND2_X1 U14478 ( .A1(n12079), .A2(n12072), .ZN(n12075) );
  AND2_X1 U14479 ( .A1(n12078), .A2(n12073), .ZN(n12074) );
  MUX2_X1 U14480 ( .A(n12075), .B(n12074), .S(n12173), .Z(n12076) );
  NAND2_X1 U14481 ( .A1(n12077), .A2(n12076), .ZN(n12081) );
  MUX2_X1 U14482 ( .A(n12079), .B(n12078), .S(n12128), .Z(n12080) );
  MUX2_X1 U14483 ( .A(n13880), .B(n14197), .S(n12128), .Z(n12082) );
  XNOR2_X1 U14484 ( .A(n14187), .B(n12128), .ZN(n12091) );
  XNOR2_X1 U14485 ( .A(n13886), .B(n12173), .ZN(n12085) );
  NAND2_X1 U14486 ( .A1(n14192), .A2(n13884), .ZN(n13869) );
  MUX2_X1 U14487 ( .A(n13884), .B(n14192), .S(n12128), .Z(n12089) );
  AOI22_X1 U14488 ( .A1(n12091), .A2(n12085), .B1(n13869), .B2(n12089), .ZN(
        n12083) );
  XNOR2_X1 U14489 ( .A(n14060), .B(n13682), .ZN(n13873) );
  INV_X1 U14490 ( .A(n12089), .ZN(n12086) );
  OR2_X1 U14491 ( .A1(n14192), .A2(n13884), .ZN(n13867) );
  INV_X1 U14492 ( .A(n12085), .ZN(n12087) );
  AOI21_X1 U14493 ( .B1(n12086), .B2(n13867), .A(n12087), .ZN(n12090) );
  NAND2_X1 U14494 ( .A1(n13867), .A2(n12087), .ZN(n12088) );
  OAI22_X1 U14495 ( .A1(n12091), .A2(n12090), .B1(n12089), .B2(n12088), .ZN(
        n12092) );
  NOR2_X1 U14496 ( .A1(n13873), .A2(n12092), .ZN(n12093) );
  NAND2_X1 U14497 ( .A1(n12094), .A2(n12093), .ZN(n12098) );
  NAND2_X1 U14498 ( .A1(n13887), .A2(n12173), .ZN(n12096) );
  OR2_X1 U14499 ( .A1(n13887), .A2(n12173), .ZN(n12095) );
  MUX2_X1 U14500 ( .A(n12096), .B(n12095), .S(n14060), .Z(n12097) );
  MUX2_X1 U14501 ( .A(n13888), .B(n14175), .S(n12037), .Z(n12099) );
  INV_X1 U14502 ( .A(n12099), .ZN(n12101) );
  MUX2_X1 U14503 ( .A(n14175), .B(n13888), .S(n12173), .Z(n12100) );
  MUX2_X1 U14504 ( .A(n14170), .B(n13874), .S(n12037), .Z(n12104) );
  MUX2_X1 U14505 ( .A(n13874), .B(n14170), .S(n12037), .Z(n12102) );
  NAND2_X1 U14506 ( .A1(n12103), .A2(n12102), .ZN(n12106) );
  NAND2_X1 U14507 ( .A1(n6516), .A2(n7223), .ZN(n12105) );
  NAND2_X1 U14508 ( .A1(n12106), .A2(n12105), .ZN(n12110) );
  MUX2_X1 U14509 ( .A(n14007), .B(n13875), .S(n12128), .Z(n12107) );
  INV_X1 U14510 ( .A(n12107), .ZN(n12109) );
  MUX2_X1 U14511 ( .A(n14007), .B(n13875), .S(n12037), .Z(n12108) );
  MUX2_X1 U14512 ( .A(n13876), .B(n14159), .S(n12037), .Z(n12113) );
  MUX2_X1 U14513 ( .A(n13893), .B(n13983), .S(n12173), .Z(n12119) );
  NAND2_X1 U14514 ( .A1(n12118), .A2(n12119), .ZN(n12117) );
  MUX2_X1 U14515 ( .A(n13983), .B(n13893), .S(n12173), .Z(n12116) );
  NAND2_X1 U14516 ( .A1(n12117), .A2(n12116), .ZN(n12123) );
  INV_X1 U14517 ( .A(n12118), .ZN(n12121) );
  INV_X1 U14518 ( .A(n12119), .ZN(n12120) );
  NAND2_X1 U14519 ( .A1(n12121), .A2(n12120), .ZN(n12122) );
  NAND2_X1 U14520 ( .A1(n12123), .A2(n12122), .ZN(n12125) );
  MUX2_X1 U14521 ( .A(n13894), .B(n13969), .S(n12128), .Z(n12126) );
  MUX2_X1 U14522 ( .A(n13894), .B(n13969), .S(n12173), .Z(n12124) );
  INV_X1 U14523 ( .A(n12126), .ZN(n12127) );
  MUX2_X1 U14524 ( .A(n13720), .B(n14142), .S(n12173), .Z(n12131) );
  MUX2_X1 U14525 ( .A(n13720), .B(n14142), .S(n12128), .Z(n12129) );
  NAND2_X1 U14526 ( .A1(n12130), .A2(n12129), .ZN(n12133) );
  NAND2_X1 U14527 ( .A1(n12133), .A2(n12132), .ZN(n12134) );
  MUX2_X1 U14528 ( .A(n13896), .B(n6701), .S(n12128), .Z(n12135) );
  NAND2_X1 U14529 ( .A1(n12134), .A2(n12135), .ZN(n12138) );
  INV_X1 U14530 ( .A(n12134), .ZN(n12137) );
  INV_X1 U14531 ( .A(n12135), .ZN(n12136) );
  NAND2_X1 U14532 ( .A1(n14235), .A2(n11085), .ZN(n12141) );
  OR2_X1 U14533 ( .A1(n12160), .A2(n14236), .ZN(n12140) );
  MUX2_X1 U14534 ( .A(n13904), .B(n14130), .S(n12173), .Z(n12143) );
  MUX2_X1 U14535 ( .A(n13926), .B(n13897), .S(n12173), .Z(n12142) );
  NAND2_X1 U14536 ( .A1(n12146), .A2(n12145), .ZN(n12177) );
  NAND2_X1 U14537 ( .A1(n12147), .A2(n11085), .ZN(n12150) );
  OR2_X1 U14538 ( .A1(n12160), .A2(n12148), .ZN(n12149) );
  INV_X1 U14539 ( .A(n13909), .ZN(n12153) );
  INV_X1 U14540 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12151) );
  NOR2_X1 U14541 ( .A1(n9744), .A2(n12151), .ZN(n12152) );
  NAND2_X1 U14542 ( .A1(n12153), .A2(n12152), .ZN(n12159) );
  INV_X1 U14543 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n12620) );
  NAND2_X1 U14544 ( .A1(n12154), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12156) );
  NAND2_X1 U14545 ( .A1(n12164), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12155) );
  OAI211_X1 U14546 ( .C1(n12167), .C2(n12620), .A(n12156), .B(n12155), .ZN(
        n12157) );
  INV_X1 U14547 ( .A(n12157), .ZN(n12158) );
  NAND2_X1 U14548 ( .A1(n12159), .A2(n12158), .ZN(n13719) );
  MUX2_X1 U14549 ( .A(n14126), .B(n13719), .S(n12173), .Z(n12176) );
  NAND2_X1 U14550 ( .A1(n12245), .A2(n11085), .ZN(n12162) );
  OR2_X1 U14551 ( .A1(n12160), .A2(n14232), .ZN(n12161) );
  INV_X1 U14552 ( .A(n12163), .ZN(n12168) );
  INV_X1 U14553 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U14554 ( .A1(n12164), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U14555 ( .A1(n12154), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12165) );
  OAI211_X1 U14556 ( .C1(n12167), .C2(n12717), .A(n12166), .B(n12165), .ZN(
        n13905) );
  OAI21_X1 U14557 ( .B1(n12168), .B2(n13855), .A(n13905), .ZN(n12169) );
  INV_X1 U14558 ( .A(n12169), .ZN(n12170) );
  MUX2_X1 U14559 ( .A(n13859), .B(n12170), .S(n12173), .Z(n12178) );
  INV_X1 U14560 ( .A(n13855), .ZN(n12181) );
  OAI21_X1 U14561 ( .B1(n12173), .B2(n12181), .A(n12171), .ZN(n12172) );
  AOI22_X1 U14562 ( .A1(n13859), .A2(n12173), .B1(n13905), .B2(n12172), .ZN(
        n12179) );
  INV_X1 U14563 ( .A(n13719), .ZN(n12205) );
  INV_X1 U14564 ( .A(n14126), .ZN(n12174) );
  MUX2_X1 U14565 ( .A(n12205), .B(n12174), .S(n12037), .Z(n12175) );
  INV_X1 U14566 ( .A(n12179), .ZN(n12180) );
  INV_X1 U14567 ( .A(n13896), .ZN(n13879) );
  NAND2_X1 U14568 ( .A1(n13969), .A2(n13894), .ZN(n13878) );
  OR2_X1 U14569 ( .A1(n13969), .A2(n13894), .ZN(n12182) );
  XNOR2_X1 U14570 ( .A(n14007), .B(n13891), .ZN(n13890) );
  INV_X1 U14571 ( .A(n13888), .ZN(n13613) );
  XNOR2_X1 U14572 ( .A(n14175), .B(n13613), .ZN(n14041) );
  NAND2_X1 U14573 ( .A1(n14028), .A2(n13874), .ZN(n13889) );
  OAI21_X1 U14574 ( .B1(n14028), .B2(n13874), .A(n13889), .ZN(n14021) );
  NAND3_X1 U14575 ( .A1(n14582), .A2(n12184), .A3(n12183), .ZN(n12185) );
  NOR4_X1 U14576 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n12190) );
  NAND4_X1 U14577 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n14566), .ZN(
        n12192) );
  NOR3_X1 U14578 ( .A1(n12194), .A2(n12193), .A3(n12192), .ZN(n12196) );
  NAND4_X1 U14579 ( .A1(n12197), .A2(n12196), .A3(n14299), .A4(n12195), .ZN(
        n12198) );
  NOR4_X1 U14580 ( .A1(n14090), .A2(n12199), .A3(n11538), .A4(n12198), .ZN(
        n12201) );
  XNOR2_X1 U14581 ( .A(n14187), .B(n13886), .ZN(n13885) );
  NAND4_X1 U14582 ( .A1(n14050), .A2(n12201), .A3(n13885), .A4(n12200), .ZN(
        n12202) );
  NOR4_X1 U14583 ( .A1(n13890), .A2(n14041), .A3(n14021), .A4(n12202), .ZN(
        n12203) );
  NAND4_X1 U14584 ( .A1(n13961), .A2(n12203), .A3(n13973), .A4(n13997), .ZN(
        n12204) );
  XOR2_X1 U14585 ( .A(n12205), .B(n14126), .Z(n13898) );
  XNOR2_X1 U14586 ( .A(n13859), .B(n13905), .ZN(n12206) );
  INV_X1 U14587 ( .A(n13856), .ZN(n14118) );
  NOR3_X1 U14588 ( .A1(n14118), .A2(n13855), .A3(n12208), .ZN(n12211) );
  NOR3_X1 U14589 ( .A1(n12210), .A2(n13855), .A3(n12219), .ZN(n12209) );
  AOI21_X1 U14590 ( .B1(n12211), .B2(n12210), .A(n12209), .ZN(n12215) );
  XOR2_X1 U14591 ( .A(n12219), .B(n12212), .Z(n12213) );
  NAND3_X1 U14592 ( .A1(n12213), .A2(n14118), .A3(n13855), .ZN(n12214) );
  OAI211_X1 U14593 ( .C1(n12217), .C2(n12216), .A(n12215), .B(n12214), .ZN(
        n12218) );
  INV_X1 U14594 ( .A(n12218), .ZN(n12221) );
  INV_X1 U14595 ( .A(n12219), .ZN(n12220) );
  NOR3_X1 U14596 ( .A1(n12222), .A2(n6394), .A3(n13903), .ZN(n12224) );
  OAI21_X1 U14597 ( .B1(n12225), .B2(n14250), .A(P1_B_REG_SCAN_IN), .ZN(n12223) );
  OAI222_X1 U14598 ( .A1(n14245), .A2(n12228), .B1(n14244), .B2(n12227), .C1(
        P1_U3086), .C2(n12226), .ZN(P1_U3336) );
  OAI22_X1 U14599 ( .A1(n14130), .A2(n9728), .B1(n13904), .B2(n9756), .ZN(
        n12233) );
  XNOR2_X1 U14600 ( .A(n12233), .B(n12232), .ZN(n12235) );
  OAI22_X1 U14601 ( .A1(n14130), .A2(n9737), .B1(n13904), .B2(n9728), .ZN(
        n12234) );
  XNOR2_X1 U14602 ( .A(n12235), .B(n12234), .ZN(n12236) );
  NAND2_X1 U14603 ( .A1(n13896), .A2(n14100), .ZN(n12238) );
  NAND2_X1 U14604 ( .A1(n13719), .A2(n13854), .ZN(n12237) );
  AND2_X1 U14605 ( .A1(n12238), .A2(n12237), .ZN(n14128) );
  AOI22_X1 U14606 ( .A1(n13923), .A2(n13714), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12239) );
  OAI21_X1 U14607 ( .B1(n14128), .B2(n13712), .A(n12239), .ZN(n12240) );
  AOI21_X1 U14608 ( .B1(n13926), .B2(n14475), .A(n12240), .ZN(n12241) );
  OAI21_X1 U14609 ( .B1(n12242), .B2(n13705), .A(n12241), .ZN(P1_U3220) );
  INV_X1 U14610 ( .A(n12243), .ZN(n12244) );
  OAI222_X1 U14611 ( .A1(P3_U3151), .A2(n8152), .B1(n12992), .B2(n12658), .C1(
        n14277), .C2(n12244), .ZN(P3_U3265) );
  INV_X1 U14612 ( .A(n12245), .ZN(n14234) );
  OAI222_X1 U14613 ( .A1(P2_U3088), .A2(n12247), .B1(n13575), .B2(n14234), 
        .C1(n12246), .C2(n13573), .ZN(P2_U3297) );
  XNOR2_X1 U14614 ( .A(n12524), .B(n8764), .ZN(n12292) );
  XNOR2_X1 U14615 ( .A(n12292), .B(n12536), .ZN(n12294) );
  AOI22_X1 U14616 ( .A1(n12252), .A2(n12582), .B1(n12253), .B2(n12564), .ZN(
        n12251) );
  AND2_X1 U14617 ( .A1(n12251), .A2(n7411), .ZN(n12248) );
  NAND3_X1 U14618 ( .A1(n12251), .A2(n12743), .A3(n12250), .ZN(n12258) );
  INV_X1 U14619 ( .A(n12252), .ZN(n12256) );
  OAI21_X1 U14620 ( .B1(n12253), .B2(n12564), .A(n12582), .ZN(n12255) );
  NOR3_X1 U14621 ( .A1(n12253), .A2(n12564), .A3(n12582), .ZN(n12254) );
  AOI21_X1 U14622 ( .B1(n12256), .B2(n12255), .A(n12254), .ZN(n12257) );
  XNOR2_X1 U14623 ( .A(n12845), .B(n8764), .ZN(n12260) );
  XNOR2_X1 U14624 ( .A(n12260), .B(n12535), .ZN(n12315) );
  INV_X1 U14625 ( .A(n12260), .ZN(n12261) );
  AOI22_X1 U14626 ( .A1(n12314), .A2(n12315), .B1(n12535), .B2(n12261), .ZN(
        n12373) );
  XNOR2_X1 U14627 ( .A(n12838), .B(n6402), .ZN(n12262) );
  XNOR2_X1 U14628 ( .A(n12262), .B(n12550), .ZN(n12374) );
  OAI22_X1 U14629 ( .A1(n12373), .A2(n12374), .B1(n12262), .B2(n12550), .ZN(
        n12295) );
  XOR2_X1 U14630 ( .A(n12294), .B(n12295), .Z(n12268) );
  AOI22_X1 U14631 ( .A1(n12550), .A2(n12375), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12264) );
  NAND2_X1 U14632 ( .A1(n12525), .A2(n12392), .ZN(n12263) );
  OAI211_X1 U14633 ( .C1(n12265), .C2(n12378), .A(n12264), .B(n12263), .ZN(
        n12266) );
  AOI21_X1 U14634 ( .B1(n12524), .B2(n14859), .A(n12266), .ZN(n12267) );
  OAI21_X1 U14635 ( .B1(n12268), .B2(n12382), .A(n12267), .ZN(P3_U3154) );
  OAI211_X1 U14636 ( .C1(n12271), .C2(n12270), .A(n12269), .B(n14861), .ZN(
        n12277) );
  AND2_X1 U14637 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n14983) );
  AOI21_X1 U14638 ( .B1(n14860), .B2(n12403), .A(n14983), .ZN(n12272) );
  OAI21_X1 U14639 ( .B1(n12273), .B2(n12390), .A(n12272), .ZN(n12274) );
  AOI21_X1 U14640 ( .B1(n12275), .B2(n12392), .A(n12274), .ZN(n12276) );
  OAI211_X1 U14641 ( .C1(n12960), .C2(n12395), .A(n12277), .B(n12276), .ZN(
        P3_U3155) );
  XNOR2_X1 U14642 ( .A(n12278), .B(n12731), .ZN(n12284) );
  AOI22_X1 U14643 ( .A1(n12582), .A2(n14860), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12280) );
  NAND2_X1 U14644 ( .A1(n12392), .A2(n12587), .ZN(n12279) );
  OAI211_X1 U14645 ( .C1(n12743), .C2(n12390), .A(n12280), .B(n12279), .ZN(
        n12281) );
  AOI21_X1 U14646 ( .B1(n12282), .B2(n14859), .A(n12281), .ZN(n12283) );
  OAI21_X1 U14647 ( .B1(n12284), .B2(n12382), .A(n12283), .ZN(P3_U3156) );
  OAI211_X1 U14648 ( .C1(n12287), .C2(n12286), .A(n12285), .B(n14861), .ZN(
        n12291) );
  NAND2_X1 U14649 ( .A1(n12375), .A2(n12766), .ZN(n12288) );
  NAND2_X1 U14650 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12485)
         );
  OAI211_X1 U14651 ( .C1(n12742), .C2(n12378), .A(n12288), .B(n12485), .ZN(
        n12289) );
  AOI21_X1 U14652 ( .B1(n12773), .B2(n12392), .A(n12289), .ZN(n12290) );
  OAI211_X1 U14653 ( .C1(n12395), .C2(n12940), .A(n12291), .B(n12290), .ZN(
        P3_U3159) );
  INV_X1 U14654 ( .A(n12292), .ZN(n12293) );
  XNOR2_X1 U14655 ( .A(n12504), .B(n6401), .ZN(n12297) );
  XNOR2_X1 U14656 ( .A(n12298), .B(n12297), .ZN(n12304) );
  AOI22_X1 U14657 ( .A1(n12397), .A2(n12375), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12300) );
  NAND2_X1 U14658 ( .A1(n12506), .A2(n12392), .ZN(n12299) );
  OAI211_X1 U14659 ( .C1(n12301), .C2(n12378), .A(n12300), .B(n12299), .ZN(
        n12302) );
  AOI21_X1 U14660 ( .B1(n6688), .B2(n14859), .A(n12302), .ZN(n12303) );
  OAI21_X1 U14661 ( .B1(n12304), .B2(n12382), .A(n12303), .ZN(P3_U3160) );
  INV_X1 U14662 ( .A(n12305), .ZN(n12306) );
  AOI21_X1 U14663 ( .B1(n12308), .B2(n12307), .A(n12306), .ZN(n12313) );
  NAND2_X1 U14664 ( .A1(n12392), .A2(n12747), .ZN(n12310) );
  AOI22_X1 U14665 ( .A1(n12581), .A2(n14860), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12309) );
  OAI211_X1 U14666 ( .C1(n12742), .C2(n12390), .A(n12310), .B(n12309), .ZN(
        n12311) );
  AOI21_X1 U14667 ( .B1(n12746), .B2(n14859), .A(n12311), .ZN(n12312) );
  OAI21_X1 U14668 ( .B1(n12313), .B2(n12382), .A(n12312), .ZN(P3_U3163) );
  XOR2_X1 U14669 ( .A(n12315), .B(n12314), .Z(n12321) );
  AOI22_X1 U14670 ( .A1(n12582), .A2(n12375), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12317) );
  NAND2_X1 U14671 ( .A1(n12555), .A2(n12392), .ZN(n12316) );
  OAI211_X1 U14672 ( .C1(n12318), .C2(n12378), .A(n12317), .B(n12316), .ZN(
        n12319) );
  AOI21_X1 U14673 ( .B1(n12845), .B2(n14859), .A(n12319), .ZN(n12320) );
  OAI21_X1 U14674 ( .B1(n12321), .B2(n12382), .A(n12320), .ZN(P3_U3165) );
  OAI211_X1 U14675 ( .C1(n12325), .C2(n12324), .A(n12323), .B(n14861), .ZN(
        n12330) );
  NOR2_X1 U14676 ( .A1(n12326), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14347) );
  AOI21_X1 U14677 ( .B1(n14860), .B2(n12401), .A(n14347), .ZN(n12327) );
  OAI21_X1 U14678 ( .B1(n12807), .B2(n12390), .A(n12327), .ZN(n12328) );
  AOI21_X1 U14679 ( .B1(n12812), .B2(n12392), .A(n12328), .ZN(n12329) );
  OAI211_X1 U14680 ( .C1(n12952), .C2(n12395), .A(n12330), .B(n12329), .ZN(
        P3_U3166) );
  AOI21_X1 U14681 ( .B1(n12332), .B2(n12331), .A(n6559), .ZN(n12337) );
  NAND2_X1 U14682 ( .A1(n12392), .A2(n12796), .ZN(n12334) );
  AOI22_X1 U14683 ( .A1(n14860), .A2(n12766), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12333) );
  OAI211_X1 U14684 ( .C1(n12820), .C2(n12390), .A(n12334), .B(n12333), .ZN(
        n12335) );
  AOI21_X1 U14685 ( .B1(n12795), .B2(n14859), .A(n12335), .ZN(n12336) );
  OAI21_X1 U14686 ( .B1(n12337), .B2(n12382), .A(n12336), .ZN(P3_U3168) );
  OAI211_X1 U14687 ( .C1(n12341), .C2(n12340), .A(n12339), .B(n14861), .ZN(
        n12345) );
  AOI22_X1 U14688 ( .A1(n12398), .A2(n14860), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12342) );
  OAI21_X1 U14689 ( .B1(n12781), .B2(n12390), .A(n12342), .ZN(n12343) );
  AOI21_X1 U14690 ( .B1(n12758), .B2(n12392), .A(n12343), .ZN(n12344) );
  OAI211_X1 U14691 ( .C1(n12936), .C2(n12395), .A(n12345), .B(n12344), .ZN(
        P3_U3173) );
  NAND2_X1 U14692 ( .A1(n12347), .A2(n12346), .ZN(n12349) );
  XOR2_X1 U14693 ( .A(n12349), .B(n12348), .Z(n12357) );
  NOR2_X1 U14694 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12350), .ZN(n14965) );
  AOI21_X1 U14695 ( .B1(n14860), .B2(n12404), .A(n14965), .ZN(n12351) );
  OAI21_X1 U14696 ( .B1(n12352), .B2(n12390), .A(n12351), .ZN(n12354) );
  NOR2_X1 U14697 ( .A1(n12964), .A2(n12395), .ZN(n12353) );
  AOI211_X1 U14698 ( .C1(n12355), .C2(n12392), .A(n12354), .B(n12353), .ZN(
        n12356) );
  OAI21_X1 U14699 ( .B1(n12357), .B2(n12382), .A(n12356), .ZN(P3_U3174) );
  XNOR2_X1 U14700 ( .A(n12358), .B(n12581), .ZN(n12363) );
  AOI22_X1 U14701 ( .A1(n12564), .A2(n14860), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12360) );
  NAND2_X1 U14702 ( .A1(n12392), .A2(n12735), .ZN(n12359) );
  OAI211_X1 U14703 ( .C1(n12754), .C2(n12390), .A(n12360), .B(n12359), .ZN(
        n12361) );
  AOI21_X1 U14704 ( .B1(n12734), .B2(n14859), .A(n12361), .ZN(n12362) );
  OAI21_X1 U14705 ( .B1(n12363), .B2(n12382), .A(n12362), .ZN(P3_U3175) );
  AOI21_X1 U14706 ( .B1(n12366), .B2(n12365), .A(n12382), .ZN(n12368) );
  NAND2_X1 U14707 ( .A1(n12368), .A2(n12367), .ZN(n12372) );
  NAND2_X1 U14708 ( .A1(n12375), .A2(n12401), .ZN(n12369) );
  NAND2_X1 U14709 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14390)
         );
  OAI211_X1 U14710 ( .C1(n12781), .C2(n12378), .A(n12369), .B(n14390), .ZN(
        n12370) );
  AOI21_X1 U14711 ( .B1(n12784), .B2(n12392), .A(n12370), .ZN(n12371) );
  OAI211_X1 U14712 ( .C1(n12944), .C2(n12395), .A(n12372), .B(n12371), .ZN(
        P3_U3178) );
  XOR2_X1 U14713 ( .A(n12374), .B(n12373), .Z(n12383) );
  AOI22_X1 U14714 ( .A1(n12565), .A2(n12375), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12377) );
  NAND2_X1 U14715 ( .A1(n12540), .A2(n12392), .ZN(n12376) );
  OAI211_X1 U14716 ( .C1(n12536), .C2(n12378), .A(n12377), .B(n12376), .ZN(
        n12379) );
  AOI21_X1 U14717 ( .B1(n12380), .B2(n14859), .A(n12379), .ZN(n12381) );
  OAI21_X1 U14718 ( .B1(n12383), .B2(n12382), .A(n12381), .ZN(P3_U3180) );
  OAI211_X1 U14719 ( .C1(n12387), .C2(n12386), .A(n12385), .B(n14861), .ZN(
        n12394) );
  INV_X1 U14720 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n12388) );
  NOR2_X1 U14721 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12388), .ZN(n14329) );
  AOI21_X1 U14722 ( .B1(n14860), .B2(n12402), .A(n14329), .ZN(n12389) );
  OAI21_X1 U14723 ( .B1(n12819), .B2(n12390), .A(n12389), .ZN(n12391) );
  AOI21_X1 U14724 ( .B1(n12824), .B2(n12392), .A(n12391), .ZN(n12393) );
  OAI211_X1 U14725 ( .C1(n12956), .C2(n12395), .A(n12394), .B(n12393), .ZN(
        P3_U3181) );
  MUX2_X1 U14726 ( .A(n12396), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12399), .Z(
        P3_U3522) );
  MUX2_X1 U14727 ( .A(n12503), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12399), .Z(
        P3_U3520) );
  MUX2_X1 U14728 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12516), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14729 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12397), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14730 ( .A(n12550), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12399), .Z(
        P3_U3517) );
  MUX2_X1 U14731 ( .A(n12565), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12399), .Z(
        P3_U3516) );
  MUX2_X1 U14732 ( .A(n12582), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12399), .Z(
        P3_U3515) );
  MUX2_X1 U14733 ( .A(n12564), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12399), .Z(
        P3_U3514) );
  MUX2_X1 U14734 ( .A(n12398), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12399), .Z(
        P3_U3512) );
  MUX2_X1 U14735 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12767), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14736 ( .A(n12400), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12399), .Z(
        P3_U3510) );
  MUX2_X1 U14737 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12766), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14738 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12401), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14739 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12402), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14740 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12403), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14741 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12404), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14742 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12405), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14743 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12406), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14744 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12407), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14745 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12408), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14746 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12409), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14747 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12410), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14748 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n15060), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14749 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15082), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14750 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15061), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14751 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n15083), .S(P3_U3897), .Z(
        P3_U3492) );
  INV_X1 U14752 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12875) );
  AOI22_X1 U14753 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12477), .B1(n14376), 
        .B2(n12875), .ZN(n14379) );
  INV_X1 U14754 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12883) );
  AOI22_X1 U14755 ( .A1(n12471), .A2(n12883), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n14349), .ZN(n14346) );
  NAND2_X1 U14756 ( .A1(n14986), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12465) );
  INV_X1 U14757 ( .A(n14986), .ZN(n12411) );
  INV_X1 U14758 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U14759 ( .A1(n12411), .A2(n12892), .ZN(n12412) );
  AND2_X1 U14760 ( .A1(n12412), .A2(n12465), .ZN(n14982) );
  AOI22_X1 U14761 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n14949), .B1(n12433), 
        .B2(n12420), .ZN(n14946) );
  AOI22_X1 U14762 ( .A1(n12451), .A2(n12417), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n14914), .ZN(n14911) );
  NAND2_X1 U14763 ( .A1(n14896), .A2(n12415), .ZN(n12416) );
  XNOR2_X1 U14764 ( .A(n12446), .B(n12415), .ZN(n14901) );
  NAND2_X1 U14765 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14901), .ZN(n14900) );
  NAND2_X1 U14766 ( .A1(n12416), .A2(n14900), .ZN(n14910) );
  NAND2_X1 U14767 ( .A1(n14911), .A2(n14910), .ZN(n14909) );
  NAND2_X1 U14768 ( .A1(n14931), .A2(n12418), .ZN(n12419) );
  XNOR2_X1 U14769 ( .A(n12455), .B(n12418), .ZN(n14928) );
  NAND2_X1 U14770 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n14928), .ZN(n14927) );
  NAND2_X1 U14771 ( .A1(n12419), .A2(n14927), .ZN(n14945) );
  NAND2_X1 U14772 ( .A1(n14946), .A2(n14945), .ZN(n14944) );
  NAND2_X1 U14773 ( .A1(n14967), .A2(n12421), .ZN(n12422) );
  XNOR2_X1 U14774 ( .A(n12461), .B(n12421), .ZN(n14964) );
  NAND2_X1 U14775 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n14964), .ZN(n14963) );
  NAND2_X1 U14776 ( .A1(n12422), .A2(n14963), .ZN(n14981) );
  NAND2_X1 U14777 ( .A1(n14982), .A2(n14981), .ZN(n14980) );
  NAND2_X1 U14778 ( .A1(n12465), .A2(n14980), .ZN(n12423) );
  NAND2_X1 U14779 ( .A1(n14331), .A2(n12423), .ZN(n12424) );
  XNOR2_X1 U14780 ( .A(n12469), .B(n12423), .ZN(n14328) );
  NAND2_X1 U14781 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14328), .ZN(n14327) );
  NAND2_X1 U14782 ( .A1(n12424), .A2(n14327), .ZN(n14345) );
  NAND2_X1 U14783 ( .A1(n14346), .A2(n14345), .ZN(n14344) );
  OAI21_X1 U14784 ( .B1(n12471), .B2(n12883), .A(n14344), .ZN(n12425) );
  NAND2_X1 U14785 ( .A1(n12474), .A2(n12425), .ZN(n12426) );
  XNOR2_X1 U14786 ( .A(n14361), .B(n12425), .ZN(n14363) );
  NAND2_X1 U14787 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14363), .ZN(n14362) );
  NAND2_X1 U14788 ( .A1(n12426), .A2(n14362), .ZN(n14378) );
  NAND2_X1 U14789 ( .A1(n14379), .A2(n14378), .ZN(n14377) );
  NAND2_X1 U14790 ( .A1(n14986), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12466) );
  NOR2_X1 U14791 ( .A1(n12446), .A2(n12428), .ZN(n12429) );
  INV_X1 U14792 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14890) );
  XOR2_X1 U14793 ( .A(n14896), .B(n12428), .Z(n14889) );
  INV_X1 U14794 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U14795 ( .A1(n12451), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n12430), 
        .B2(n14914), .ZN(n14907) );
  INV_X1 U14796 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14926) );
  INV_X1 U14797 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U14798 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12433), .B1(n14949), 
        .B2(n12432), .ZN(n14942) );
  INV_X1 U14799 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14962) );
  OAI21_X1 U14800 ( .B1(n14986), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12466), 
        .ZN(n14978) );
  INV_X1 U14801 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14326) );
  INV_X1 U14802 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U14803 ( .A1(n12471), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12441), 
        .B2(n14349), .ZN(n14342) );
  NOR2_X1 U14804 ( .A1(n14361), .A2(n12435), .ZN(n12436) );
  INV_X1 U14805 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14370) );
  INV_X1 U14806 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U14807 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14376), .B1(n12477), 
        .B2(n12440), .ZN(n14386) );
  NOR2_X1 U14808 ( .A1(n14387), .A2(n14386), .ZN(n14388) );
  INV_X1 U14809 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12437) );
  MUX2_X1 U14810 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n12437), .S(n6403), .Z(
        n12481) );
  XNOR2_X1 U14811 ( .A(n12438), .B(n12481), .ZN(n12439) );
  MUX2_X1 U14812 ( .A(n12440), .B(n12875), .S(n12449), .Z(n14381) );
  MUX2_X1 U14813 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12449), .Z(n12475) );
  AND2_X1 U14814 ( .A1(n12475), .A2(n12474), .ZN(n12476) );
  MUX2_X1 U14815 ( .A(n12441), .B(n12883), .S(n12449), .Z(n12472) );
  NOR2_X1 U14816 ( .A1(n12472), .A2(n12471), .ZN(n14354) );
  INV_X1 U14817 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15157) );
  MUX2_X1 U14818 ( .A(n14890), .B(n15157), .S(n12449), .Z(n12447) );
  OR2_X1 U14819 ( .A1(n12447), .A2(n12446), .ZN(n14892) );
  OR2_X1 U14820 ( .A1(n12443), .A2(n12442), .ZN(n12445) );
  NAND2_X1 U14821 ( .A1(n12447), .A2(n12446), .ZN(n14893) );
  MUX2_X1 U14822 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12449), .Z(n12450) );
  XNOR2_X1 U14823 ( .A(n12450), .B(n12451), .ZN(n14918) );
  INV_X1 U14824 ( .A(n12450), .ZN(n12452) );
  NAND2_X1 U14825 ( .A1(n12452), .A2(n12451), .ZN(n12453) );
  NAND2_X1 U14826 ( .A1(n14917), .A2(n12453), .ZN(n14936) );
  MUX2_X1 U14827 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12449), .Z(n12454) );
  XNOR2_X1 U14828 ( .A(n12454), .B(n12455), .ZN(n14935) );
  INV_X1 U14829 ( .A(n12454), .ZN(n12456) );
  NAND2_X1 U14830 ( .A1(n12456), .A2(n12455), .ZN(n12457) );
  NAND2_X1 U14831 ( .A1(n14934), .A2(n12457), .ZN(n14954) );
  MUX2_X1 U14832 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12449), .Z(n12458) );
  XNOR2_X1 U14833 ( .A(n12458), .B(n14949), .ZN(n14953) );
  NAND2_X1 U14834 ( .A1(n12458), .A2(n14949), .ZN(n12459) );
  MUX2_X1 U14835 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12449), .Z(n12460) );
  XNOR2_X1 U14836 ( .A(n12460), .B(n12461), .ZN(n14971) );
  INV_X1 U14837 ( .A(n12460), .ZN(n12462) );
  NAND2_X1 U14838 ( .A1(n12462), .A2(n12461), .ZN(n12463) );
  INV_X1 U14839 ( .A(n14978), .ZN(n12464) );
  MUX2_X1 U14840 ( .A(n12464), .B(n14982), .S(n12449), .Z(n14993) );
  NAND2_X1 U14841 ( .A1(n14994), .A2(n14993), .ZN(n14992) );
  MUX2_X1 U14842 ( .A(n12466), .B(n12465), .S(n12449), .Z(n12467) );
  INV_X1 U14843 ( .A(n12468), .ZN(n12470) );
  XNOR2_X1 U14844 ( .A(n12468), .B(n14331), .ZN(n14335) );
  MUX2_X1 U14845 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12449), .Z(n14336) );
  NOR2_X1 U14846 ( .A1(n14335), .A2(n14336), .ZN(n14334) );
  NAND2_X1 U14847 ( .A1(n12472), .A2(n12471), .ZN(n14352) );
  OAI21_X1 U14848 ( .B1(n14354), .B2(n14357), .A(n14352), .ZN(n14366) );
  INV_X1 U14849 ( .A(n12476), .ZN(n12473) );
  OAI21_X1 U14850 ( .B1(n12475), .B2(n12474), .A(n12473), .ZN(n14365) );
  NOR2_X1 U14851 ( .A1(n12476), .A2(n14364), .ZN(n12478) );
  NAND2_X1 U14852 ( .A1(n14381), .A2(n14382), .ZN(n14380) );
  NAND2_X1 U14853 ( .A1(n14376), .A2(n12478), .ZN(n12479) );
  NAND2_X1 U14854 ( .A1(n14380), .A2(n12479), .ZN(n12483) );
  MUX2_X1 U14855 ( .A(n6569), .B(n12481), .S(n12480), .Z(n12482) );
  XNOR2_X1 U14856 ( .A(n12483), .B(n12482), .ZN(n12484) );
  NOR2_X1 U14857 ( .A1(n14952), .A2(n12484), .ZN(n12487) );
  OAI21_X1 U14858 ( .B1(n14886), .B2(n12642), .A(n12485), .ZN(n12486) );
  INV_X1 U14859 ( .A(n12491), .ZN(n12499) );
  NAND2_X1 U14860 ( .A1(n12492), .A2(n15109), .ZN(n12497) );
  NOR2_X1 U14861 ( .A1(n12493), .A2(n15078), .ZN(n14395) );
  NOR2_X1 U14862 ( .A1(n12494), .A2(n12826), .ZN(n12495) );
  AOI211_X1 U14863 ( .C1(n15005), .C2(P3_REG2_REG_29__SCAN_IN), .A(n14395), 
        .B(n12495), .ZN(n12496) );
  OAI211_X1 U14864 ( .C1(n12499), .C2(n12498), .A(n12497), .B(n12496), .ZN(
        P3_U3204) );
  NOR2_X1 U14865 ( .A1(n12536), .A2(n15044), .ZN(n12502) );
  XNOR2_X1 U14866 ( .A(n12505), .B(n12504), .ZN(n12831) );
  INV_X1 U14867 ( .A(n6688), .ZN(n12508) );
  AOI22_X1 U14868 ( .A1(n12506), .A2(n15103), .B1(n15005), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12507) );
  OAI21_X1 U14869 ( .B1(n12508), .B2(n12826), .A(n12507), .ZN(n12509) );
  AOI21_X1 U14870 ( .B1(n12831), .B2(n15020), .A(n12509), .ZN(n12510) );
  OAI21_X1 U14871 ( .B1(n12833), .B2(n15005), .A(n12510), .ZN(P3_U3205) );
  AOI21_X1 U14872 ( .B1(n12512), .B2(n12530), .A(n12511), .ZN(n12515) );
  INV_X1 U14873 ( .A(n12513), .ZN(n12514) );
  AOI22_X1 U14874 ( .A1(n12516), .A2(n15081), .B1(n15084), .B2(n12550), .ZN(
        n12522) );
  OAI21_X1 U14875 ( .B1(n12519), .B2(n12518), .A(n12517), .ZN(n12520) );
  NAND2_X1 U14876 ( .A1(n12520), .A2(n15089), .ZN(n12521) );
  OAI211_X1 U14877 ( .C1(n12523), .C2(n15094), .A(n12522), .B(n12521), .ZN(
        n12834) );
  INV_X1 U14878 ( .A(n12834), .ZN(n12529) );
  INV_X1 U14879 ( .A(n12523), .ZN(n12835) );
  AOI22_X1 U14880 ( .A1(n12525), .A2(n15103), .B1(n15005), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12526) );
  OAI21_X1 U14881 ( .B1(n12915), .B2(n12826), .A(n12526), .ZN(n12527) );
  AOI21_X1 U14882 ( .B1(n12835), .B2(n12586), .A(n12527), .ZN(n12528) );
  OAI21_X1 U14883 ( .B1(n12529), .B2(n15005), .A(n12528), .ZN(P3_U3206) );
  OAI21_X1 U14884 ( .B1(n12531), .B2(n12533), .A(n12530), .ZN(n12840) );
  XNOR2_X1 U14885 ( .A(n12532), .B(n12533), .ZN(n12534) );
  NAND2_X1 U14886 ( .A1(n12534), .A2(n15089), .ZN(n12539) );
  OAI22_X1 U14887 ( .A1(n12536), .A2(n15046), .B1(n12535), .B2(n15044), .ZN(
        n12537) );
  INV_X1 U14888 ( .A(n12537), .ZN(n12538) );
  OAI211_X1 U14889 ( .C1(n12840), .C2(n15094), .A(n12539), .B(n12538), .ZN(
        n12842) );
  INV_X1 U14890 ( .A(n12842), .ZN(n12545) );
  INV_X1 U14891 ( .A(n12840), .ZN(n12543) );
  AOI22_X1 U14892 ( .A1(n12540), .A2(n15103), .B1(n15005), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12541) );
  OAI21_X1 U14893 ( .B1(n12838), .B2(n12826), .A(n12541), .ZN(n12542) );
  AOI21_X1 U14894 ( .B1(n12543), .B2(n12586), .A(n12542), .ZN(n12544) );
  OAI21_X1 U14895 ( .B1(n12545), .B2(n15005), .A(n12544), .ZN(P3_U3207) );
  XNOR2_X1 U14896 ( .A(n6409), .B(n12548), .ZN(n12554) );
  OAI211_X1 U14897 ( .C1(n12549), .C2(n12548), .A(n12547), .B(n15089), .ZN(
        n12552) );
  AOI22_X1 U14898 ( .A1(n15084), .A2(n12582), .B1(n12550), .B2(n15081), .ZN(
        n12551) );
  OAI211_X1 U14899 ( .C1(n15094), .C2(n12554), .A(n12552), .B(n12551), .ZN(
        n12553) );
  INV_X1 U14900 ( .A(n12553), .ZN(n12848) );
  INV_X1 U14901 ( .A(n12554), .ZN(n12846) );
  INV_X1 U14902 ( .A(n12845), .ZN(n12557) );
  AOI22_X1 U14903 ( .A1(n12555), .A2(n15103), .B1(n15005), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12556) );
  OAI21_X1 U14904 ( .B1(n12557), .B2(n12826), .A(n12556), .ZN(n12558) );
  AOI21_X1 U14905 ( .B1(n12846), .B2(n12586), .A(n12558), .ZN(n12559) );
  OAI21_X1 U14906 ( .B1(n12848), .B2(n15005), .A(n12559), .ZN(P3_U3208) );
  XNOR2_X1 U14907 ( .A(n12561), .B(n12560), .ZN(n12568) );
  AOI21_X1 U14908 ( .B1(n12563), .B2(n12562), .A(n8639), .ZN(n12569) );
  AOI22_X1 U14909 ( .A1(n12565), .A2(n15081), .B1(n15084), .B2(n12564), .ZN(
        n12566) );
  OAI21_X1 U14910 ( .B1(n12569), .B2(n15094), .A(n12566), .ZN(n12567) );
  AOI21_X1 U14911 ( .B1(n15089), .B2(n12568), .A(n12567), .ZN(n12852) );
  INV_X1 U14912 ( .A(n12569), .ZN(n12850) );
  AOI22_X1 U14913 ( .A1(n15005), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12570), 
        .B2(n15103), .ZN(n12571) );
  OAI21_X1 U14914 ( .B1(n6392), .B2(n12826), .A(n12571), .ZN(n12573) );
  AOI21_X1 U14915 ( .B1(n12850), .B2(n12586), .A(n12573), .ZN(n12574) );
  OAI21_X1 U14916 ( .B1(n12852), .B2(n15005), .A(n12574), .ZN(P3_U3209) );
  OR2_X1 U14917 ( .A1(n12575), .A2(n12578), .ZN(n12576) );
  NAND2_X1 U14918 ( .A1(n12577), .A2(n12576), .ZN(n12585) );
  XNOR2_X1 U14919 ( .A(n12579), .B(n12578), .ZN(n12580) );
  NAND2_X1 U14920 ( .A1(n12580), .A2(n15089), .ZN(n12584) );
  AOI22_X1 U14921 ( .A1(n12582), .A2(n15081), .B1(n15084), .B2(n12581), .ZN(
        n12583) );
  OAI211_X1 U14922 ( .C1(n15094), .C2(n12585), .A(n12584), .B(n12583), .ZN(
        n12853) );
  INV_X1 U14923 ( .A(n12585), .ZN(n12854) );
  NAND2_X1 U14924 ( .A1(n12854), .A2(n12586), .ZN(n12589) );
  AOI22_X1 U14925 ( .A1(n15005), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15103), 
        .B2(n12587), .ZN(n12588) );
  OAI211_X1 U14926 ( .C1(n12924), .C2(n12826), .A(n12589), .B(n12588), .ZN(
        n12590) );
  AOI21_X1 U14927 ( .B1(n12853), .B2(n15109), .A(n12590), .ZN(n12728) );
  INV_X1 U14928 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12879) );
  NAND4_X1 U14929 ( .A1(P3_REG0_REG_14__SCAN_IN), .A2(P3_REG1_REG_13__SCAN_IN), 
        .A3(n12879), .A4(n15155), .ZN(n12593) );
  NAND4_X1 U14930 ( .A1(SI_3_), .A2(P3_REG1_REG_6__SCAN_IN), .A3(
        P3_REG1_REG_4__SCAN_IN), .A4(P3_REG0_REG_3__SCAN_IN), .ZN(n12592) );
  NAND3_X1 U14931 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_REG2_REG_0__SCAN_IN), 
        .A3(n8170), .ZN(n12591) );
  NOR4_X1 U14932 ( .A1(P3_D_REG_13__SCAN_IN), .A2(n12593), .A3(n12592), .A4(
        n12591), .ZN(n12611) );
  INV_X1 U14933 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12712) );
  NAND4_X1 U14934 ( .A1(P3_DATAO_REG_5__SCAN_IN), .A2(P3_DATAO_REG_6__SCAN_IN), 
        .A3(n12712), .A4(n10863), .ZN(n12597) );
  NAND4_X1 U14935 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_REG1_REG_13__SCAN_IN), 
        .A3(P2_REG1_REG_1__SCAN_IN), .A4(P1_REG1_REG_29__SCAN_IN), .ZN(n12596)
         );
  NAND4_X1 U14936 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), 
        .A3(P1_REG2_REG_24__SCAN_IN), .A4(P1_REG1_REG_30__SCAN_IN), .ZN(n12595) );
  NAND4_X1 U14937 ( .A1(SI_24_), .A2(P2_DATAO_REG_28__SCAN_IN), .A3(
        P3_REG1_REG_30__SCAN_IN), .A4(P1_REG3_REG_16__SCAN_IN), .ZN(n12594) );
  NOR4_X1 U14938 ( .A1(n12597), .A2(n12596), .A3(n12595), .A4(n12594), .ZN(
        n12610) );
  NOR4_X1 U14939 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), 
        .A3(P1_D_REG_0__SCAN_IN), .A4(n12661), .ZN(n12609) );
  NOR4_X1 U14940 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        P1_DATAO_REG_1__SCAN_IN), .A4(P2_DATAO_REG_5__SCAN_IN), .ZN(n12601) );
  NAND4_X1 U14941 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(P3_ADDR_REG_19__SCAN_IN), .A3(P1_DATAO_REG_15__SCAN_IN), .A4(n12660), .ZN(n12599) );
  INV_X1 U14942 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12687) );
  NAND4_X1 U14943 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_REG2_REG_24__SCAN_IN), 
        .A3(n12656), .A4(n12687), .ZN(n12598) );
  NOR4_X1 U14944 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(n12599), .A3(n12598), .A4(
        P1_ADDR_REG_0__SCAN_IN), .ZN(n12600) );
  NAND4_X1 U14945 ( .A1(n12601), .A2(P1_DATAO_REG_8__SCAN_IN), .A3(n12600), 
        .A4(n12626), .ZN(n12607) );
  NOR4_X1 U14946 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(P3_DATAO_REG_22__SCAN_IN), 
        .A3(P3_DATAO_REG_10__SCAN_IN), .A4(P3_RD_REG_SCAN_IN), .ZN(n12605) );
  NOR4_X1 U14947 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_REG2_REG_1__SCAN_IN), 
        .A3(P1_D_REG_15__SCAN_IN), .A4(P1_REG2_REG_23__SCAN_IN), .ZN(n12604)
         );
  NOR4_X1 U14948 ( .A1(SI_30_), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_REG3_REG_4__SCAN_IN), .A4(P1_REG1_REG_12__SCAN_IN), .ZN(n12603) );
  NOR4_X1 U14949 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(P1_DATAO_REG_31__SCAN_IN), 
        .A3(P1_REG2_REG_27__SCAN_IN), .A4(P1_REG2_REG_13__SCAN_IN), .ZN(n12602) );
  NAND4_X1 U14950 ( .A1(n12605), .A2(n12604), .A3(n12603), .A4(n12602), .ZN(
        n12606) );
  NOR2_X1 U14951 ( .A1(n12607), .A2(n12606), .ZN(n12608) );
  NAND4_X1 U14952 ( .A1(n12611), .A2(n12610), .A3(n12609), .A4(n12608), .ZN(
        n12726) );
  XNOR2_X1 U14953 ( .A(n12612), .B(keyinput57), .ZN(n12619) );
  XNOR2_X1 U14954 ( .A(n12613), .B(keyinput10), .ZN(n12618) );
  XNOR2_X1 U14955 ( .A(n12614), .B(keyinput12), .ZN(n12617) );
  XNOR2_X1 U14956 ( .A(n12615), .B(keyinput30), .ZN(n12616) );
  NOR4_X1 U14957 ( .A1(n12619), .A2(n12618), .A3(n12617), .A4(n12616), .ZN(
        n12640) );
  XOR2_X1 U14958 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput1), .Z(n12624) );
  XOR2_X1 U14959 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput6), .Z(n12623) );
  XNOR2_X1 U14960 ( .A(n12957), .B(keyinput63), .ZN(n12622) );
  XNOR2_X1 U14961 ( .A(n12620), .B(keyinput11), .ZN(n12621) );
  NOR4_X1 U14962 ( .A1(n12624), .A2(n12623), .A3(n12622), .A4(n12621), .ZN(
        n12639) );
  XOR2_X1 U14963 ( .A(SI_3_), .B(keyinput24), .Z(n12630) );
  XOR2_X1 U14964 ( .A(P3_REG1_REG_13__SCAN_IN), .B(keyinput38), .Z(n12629) );
  XNOR2_X1 U14965 ( .A(n12625), .B(keyinput18), .ZN(n12628) );
  XNOR2_X1 U14966 ( .A(n12626), .B(keyinput27), .ZN(n12627) );
  NOR4_X1 U14967 ( .A1(n12630), .A2(n12629), .A3(n12628), .A4(n12627), .ZN(
        n12638) );
  XNOR2_X1 U14968 ( .A(n12631), .B(keyinput36), .ZN(n12636) );
  XNOR2_X1 U14969 ( .A(n12632), .B(keyinput41), .ZN(n12635) );
  XNOR2_X1 U14970 ( .A(keyinput28), .B(n13320), .ZN(n12634) );
  XNOR2_X1 U14971 ( .A(keyinput45), .B(n11186), .ZN(n12633) );
  NOR4_X1 U14972 ( .A1(n12636), .A2(n12635), .A3(n12634), .A4(n12633), .ZN(
        n12637) );
  NAND4_X1 U14973 ( .A1(n12640), .A2(n12639), .A3(n12638), .A4(n12637), .ZN(
        n12651) );
  AOI22_X1 U14974 ( .A1(n12642), .A2(keyinput20), .B1(keyinput16), .B2(n15155), 
        .ZN(n12641) );
  OAI221_X1 U14975 ( .B1(n12642), .B2(keyinput20), .C1(n15155), .C2(keyinput16), .A(n12641), .ZN(n12650) );
  AOI22_X1 U14976 ( .A1(n12644), .A2(keyinput49), .B1(keyinput54), .B2(n14412), 
        .ZN(n12643) );
  OAI221_X1 U14977 ( .B1(n12644), .B2(keyinput49), .C1(n14412), .C2(keyinput54), .A(n12643), .ZN(n12649) );
  XOR2_X1 U14978 ( .A(n11293), .B(keyinput31), .Z(n12647) );
  XNOR2_X1 U14979 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput55), .ZN(n12646)
         );
  XNOR2_X1 U14980 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput34), .ZN(n12645) );
  NAND3_X1 U14981 ( .A1(n12647), .A2(n12646), .A3(n12645), .ZN(n12648) );
  NOR4_X1 U14982 ( .A1(n12651), .A2(n12650), .A3(n12649), .A4(n12648), .ZN(
        n12698) );
  AOI22_X1 U14983 ( .A1(n12654), .A2(keyinput59), .B1(n12653), .B2(keyinput60), 
        .ZN(n12652) );
  OAI221_X1 U14984 ( .B1(n12654), .B2(keyinput59), .C1(n12653), .C2(keyinput60), .A(n12652), .ZN(n12665) );
  AOI22_X1 U14985 ( .A1(n9871), .A2(keyinput37), .B1(keyinput33), .B2(n12656), 
        .ZN(n12655) );
  OAI221_X1 U14986 ( .B1(n9871), .B2(keyinput37), .C1(n12656), .C2(keyinput33), 
        .A(n12655), .ZN(n12664) );
  INV_X1 U14987 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14830) );
  AOI22_X1 U14988 ( .A1(n12658), .A2(keyinput14), .B1(n14830), .B2(keyinput26), 
        .ZN(n12657) );
  OAI221_X1 U14989 ( .B1(n12658), .B2(keyinput14), .C1(n14830), .C2(keyinput26), .A(n12657), .ZN(n12663) );
  AOI22_X1 U14990 ( .A1(n12661), .A2(keyinput40), .B1(n12660), .B2(keyinput53), 
        .ZN(n12659) );
  OAI221_X1 U14991 ( .B1(n12661), .B2(keyinput40), .C1(n12660), .C2(keyinput53), .A(n12659), .ZN(n12662) );
  NOR4_X1 U14992 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12697) );
  AOI22_X1 U14993 ( .A1(n12668), .A2(keyinput43), .B1(n12667), .B2(keyinput21), 
        .ZN(n12666) );
  OAI221_X1 U14994 ( .B1(n12668), .B2(keyinput43), .C1(n12667), .C2(keyinput21), .A(n12666), .ZN(n12679) );
  AOI22_X1 U14995 ( .A1(n12671), .A2(keyinput0), .B1(keyinput2), .B2(n12670), 
        .ZN(n12669) );
  OAI221_X1 U14996 ( .B1(n12671), .B2(keyinput0), .C1(n12670), .C2(keyinput2), 
        .A(n12669), .ZN(n12678) );
  AOI22_X1 U14997 ( .A1(n10863), .A2(keyinput42), .B1(n9889), .B2(keyinput13), 
        .ZN(n12672) );
  OAI221_X1 U14998 ( .B1(n10863), .B2(keyinput42), .C1(n9889), .C2(keyinput13), 
        .A(n12672), .ZN(n12677) );
  INV_X1 U14999 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U15000 ( .A1(n12675), .A2(keyinput9), .B1(keyinput35), .B2(n12674), 
        .ZN(n12673) );
  OAI221_X1 U15001 ( .B1(n12675), .B2(keyinput9), .C1(n12674), .C2(keyinput35), 
        .A(n12673), .ZN(n12676) );
  NOR4_X1 U15002 ( .A1(n12679), .A2(n12678), .A3(n12677), .A4(n12676), .ZN(
        n12696) );
  AOI22_X1 U15003 ( .A1(n12681), .A2(keyinput17), .B1(keyinput50), .B2(n15147), 
        .ZN(n12680) );
  OAI221_X1 U15004 ( .B1(n12681), .B2(keyinput17), .C1(n15147), .C2(keyinput50), .A(n12680), .ZN(n12694) );
  AOI22_X1 U15005 ( .A1(n12683), .A2(keyinput8), .B1(keyinput46), .B2(n11390), 
        .ZN(n12682) );
  OAI221_X1 U15006 ( .B1(n12683), .B2(keyinput8), .C1(n11390), .C2(keyinput46), 
        .A(n12682), .ZN(n12693) );
  AOI22_X1 U15007 ( .A1(n8037), .A2(keyinput19), .B1(keyinput58), .B2(n12685), 
        .ZN(n12684) );
  OAI221_X1 U15008 ( .B1(n8037), .B2(keyinput19), .C1(n12685), .C2(keyinput58), 
        .A(n12684), .ZN(n12691) );
  AOI22_X1 U15009 ( .A1(n12687), .A2(keyinput32), .B1(keyinput52), .B2(n13553), 
        .ZN(n12686) );
  OAI221_X1 U15010 ( .B1(n12687), .B2(keyinput32), .C1(n13553), .C2(keyinput52), .A(n12686), .ZN(n12690) );
  XNOR2_X1 U15011 ( .A(n12688), .B(keyinput61), .ZN(n12689) );
  OR3_X1 U15012 ( .A1(n12691), .A2(n12690), .A3(n12689), .ZN(n12692) );
  NOR3_X1 U15013 ( .A1(n12694), .A2(n12693), .A3(n12692), .ZN(n12695) );
  AND4_X1 U15014 ( .A1(n12698), .A2(n12697), .A3(n12696), .A4(n12695), .ZN(
        n12724) );
  INV_X1 U15015 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U15016 ( .A1(n15151), .A2(keyinput3), .B1(n12700), .B2(keyinput22), 
        .ZN(n12699) );
  OAI221_X1 U15017 ( .B1(n15151), .B2(keyinput3), .C1(n12700), .C2(keyinput22), 
        .A(n12699), .ZN(n12710) );
  INV_X1 U15018 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15019 ( .A1(n12702), .A2(keyinput23), .B1(n12879), .B2(keyinput7), 
        .ZN(n12701) );
  OAI221_X1 U15020 ( .B1(n12702), .B2(keyinput23), .C1(n12879), .C2(keyinput7), 
        .A(n12701), .ZN(n12709) );
  INV_X1 U15021 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14601) );
  AOI22_X1 U15022 ( .A1(n14601), .A2(keyinput48), .B1(n12704), .B2(keyinput47), 
        .ZN(n12703) );
  OAI221_X1 U15023 ( .B1(n14601), .B2(keyinput48), .C1(n12704), .C2(keyinput47), .A(n12703), .ZN(n12708) );
  INV_X1 U15024 ( .A(P3_RD_REG_SCAN_IN), .ZN(n14256) );
  AOI22_X1 U15025 ( .A1(n12706), .A2(keyinput56), .B1(keyinput5), .B2(n14256), 
        .ZN(n12705) );
  OAI221_X1 U15026 ( .B1(n12706), .B2(keyinput56), .C1(n14256), .C2(keyinput5), 
        .A(n12705), .ZN(n12707) );
  NOR4_X1 U15027 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12723) );
  AOI22_X1 U15028 ( .A1(n12712), .A2(keyinput62), .B1(n14236), .B2(keyinput15), 
        .ZN(n12711) );
  OAI221_X1 U15029 ( .B1(n12712), .B2(keyinput62), .C1(n14236), .C2(keyinput15), .A(n12711), .ZN(n12721) );
  INV_X1 U15030 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14600) );
  AOI22_X1 U15031 ( .A1(n14600), .A2(keyinput25), .B1(n8204), .B2(keyinput39), 
        .ZN(n12713) );
  OAI221_X1 U15032 ( .B1(n14600), .B2(keyinput25), .C1(n8204), .C2(keyinput39), 
        .A(n12713), .ZN(n12720) );
  AOI22_X1 U15033 ( .A1(n8170), .A2(keyinput4), .B1(keyinput44), .B2(n12715), 
        .ZN(n12714) );
  OAI221_X1 U15034 ( .B1(n8170), .B2(keyinput4), .C1(n12715), .C2(keyinput44), 
        .A(n12714), .ZN(n12719) );
  AOI22_X1 U15035 ( .A1(n11924), .A2(keyinput51), .B1(keyinput29), .B2(n12717), 
        .ZN(n12716) );
  OAI221_X1 U15036 ( .B1(n11924), .B2(keyinput51), .C1(n12717), .C2(keyinput29), .A(n12716), .ZN(n12718) );
  NOR4_X1 U15037 ( .A1(n12721), .A2(n12720), .A3(n12719), .A4(n12718), .ZN(
        n12722) );
  NAND3_X1 U15038 ( .A1(n12724), .A2(n12723), .A3(n12722), .ZN(n12725) );
  XOR2_X1 U15039 ( .A(n12726), .B(n12725), .Z(n12727) );
  XNOR2_X1 U15040 ( .A(n12728), .B(n12727), .ZN(P3_U3210) );
  XNOR2_X1 U15041 ( .A(n12729), .B(n12732), .ZN(n12730) );
  OAI222_X1 U15042 ( .A1(n15046), .A2(n12731), .B1(n15044), .B2(n12754), .C1(
        n12730), .C2(n15052), .ZN(n12857) );
  INV_X1 U15043 ( .A(n12857), .ZN(n12739) );
  XNOR2_X1 U15044 ( .A(n12733), .B(n12732), .ZN(n12858) );
  INV_X1 U15045 ( .A(n12734), .ZN(n12928) );
  AOI22_X1 U15046 ( .A1(n15005), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15103), 
        .B2(n12735), .ZN(n12736) );
  OAI21_X1 U15047 ( .B1(n12928), .B2(n12826), .A(n12736), .ZN(n12737) );
  AOI21_X1 U15048 ( .B1(n12858), .B2(n15020), .A(n12737), .ZN(n12738) );
  OAI21_X1 U15049 ( .B1(n12739), .B2(n15005), .A(n12738), .ZN(P3_U3211) );
  XNOR2_X1 U15050 ( .A(n12740), .B(n12745), .ZN(n12741) );
  OAI222_X1 U15051 ( .A1(n15046), .A2(n12743), .B1(n15044), .B2(n12742), .C1(
        n15052), .C2(n12741), .ZN(n12861) );
  INV_X1 U15052 ( .A(n12861), .ZN(n12751) );
  XNOR2_X1 U15053 ( .A(n12744), .B(n12745), .ZN(n12862) );
  INV_X1 U15054 ( .A(n12746), .ZN(n12932) );
  AOI22_X1 U15055 ( .A1(n15005), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15103), 
        .B2(n12747), .ZN(n12748) );
  OAI21_X1 U15056 ( .B1(n12932), .B2(n12826), .A(n12748), .ZN(n12749) );
  AOI21_X1 U15057 ( .B1(n12862), .B2(n15020), .A(n12749), .ZN(n12750) );
  OAI21_X1 U15058 ( .B1(n12751), .B2(n15005), .A(n12750), .ZN(P3_U3212) );
  XNOR2_X1 U15059 ( .A(n12752), .B(n12757), .ZN(n12753) );
  OAI222_X1 U15060 ( .A1(n15046), .A2(n12754), .B1(n15044), .B2(n12781), .C1(
        n12753), .C2(n15052), .ZN(n12865) );
  INV_X1 U15061 ( .A(n12865), .ZN(n12762) );
  AOI21_X1 U15062 ( .B1(n12757), .B2(n12756), .A(n12755), .ZN(n12866) );
  AOI22_X1 U15063 ( .A1(n15005), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15103), 
        .B2(n12758), .ZN(n12759) );
  OAI21_X1 U15064 ( .B1(n12936), .B2(n12826), .A(n12759), .ZN(n12760) );
  AOI21_X1 U15065 ( .B1(n12866), .B2(n15020), .A(n12760), .ZN(n12761) );
  OAI21_X1 U15066 ( .B1(n12762), .B2(n15005), .A(n12761), .ZN(P3_U3213) );
  NAND2_X1 U15067 ( .A1(n12763), .A2(n15089), .ZN(n12770) );
  AOI21_X1 U15068 ( .B1(n12764), .B2(n12765), .A(n12771), .ZN(n12769) );
  AOI22_X1 U15069 ( .A1(n12767), .A2(n15081), .B1(n15084), .B2(n12766), .ZN(
        n12768) );
  OAI21_X1 U15070 ( .B1(n12770), .B2(n12769), .A(n12768), .ZN(n12869) );
  INV_X1 U15071 ( .A(n12869), .ZN(n12777) );
  XNOR2_X1 U15072 ( .A(n12772), .B(n12771), .ZN(n12870) );
  AOI22_X1 U15073 ( .A1(n15005), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15103), 
        .B2(n12773), .ZN(n12774) );
  OAI21_X1 U15074 ( .B1(n12940), .B2(n12826), .A(n12774), .ZN(n12775) );
  AOI21_X1 U15075 ( .B1(n12870), .B2(n15020), .A(n12775), .ZN(n12776) );
  OAI21_X1 U15076 ( .B1(n12777), .B2(n15005), .A(n12776), .ZN(P3_U3214) );
  INV_X1 U15077 ( .A(n12764), .ZN(n12778) );
  AOI21_X1 U15078 ( .B1(n12782), .B2(n12779), .A(n12778), .ZN(n12780) );
  OAI222_X1 U15079 ( .A1(n15046), .A2(n12781), .B1(n15044), .B2(n12808), .C1(
        n15052), .C2(n12780), .ZN(n12873) );
  INV_X1 U15080 ( .A(n12873), .ZN(n12788) );
  XNOR2_X1 U15081 ( .A(n12783), .B(n12782), .ZN(n12874) );
  AOI22_X1 U15082 ( .A1(n15005), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15103), 
        .B2(n12784), .ZN(n12785) );
  OAI21_X1 U15083 ( .B1(n12944), .B2(n12826), .A(n12785), .ZN(n12786) );
  AOI21_X1 U15084 ( .B1(n12874), .B2(n15020), .A(n12786), .ZN(n12787) );
  OAI21_X1 U15085 ( .B1(n12788), .B2(n15005), .A(n12787), .ZN(P3_U3215) );
  XNOR2_X1 U15086 ( .A(n12789), .B(n12790), .ZN(n12791) );
  OAI222_X1 U15087 ( .A1(n15046), .A2(n12792), .B1(n15044), .B2(n12820), .C1(
        n12791), .C2(n15052), .ZN(n12877) );
  INV_X1 U15088 ( .A(n12877), .ZN(n12800) );
  XNOR2_X1 U15089 ( .A(n12794), .B(n12793), .ZN(n12878) );
  INV_X1 U15090 ( .A(n12795), .ZN(n12948) );
  AOI22_X1 U15091 ( .A1(n15005), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15103), 
        .B2(n12796), .ZN(n12797) );
  OAI21_X1 U15092 ( .B1(n12948), .B2(n12826), .A(n12797), .ZN(n12798) );
  AOI21_X1 U15093 ( .B1(n12878), .B2(n15020), .A(n12798), .ZN(n12799) );
  OAI21_X1 U15094 ( .B1(n12800), .B2(n15005), .A(n12799), .ZN(P3_U3216) );
  NAND2_X1 U15095 ( .A1(n12817), .A2(n12801), .ZN(n12803) );
  NAND2_X1 U15096 ( .A1(n12803), .A2(n12802), .ZN(n12805) );
  XNOR2_X1 U15097 ( .A(n12805), .B(n12804), .ZN(n12806) );
  OAI222_X1 U15098 ( .A1(n15046), .A2(n12808), .B1(n15044), .B2(n12807), .C1(
        n12806), .C2(n15052), .ZN(n12881) );
  INV_X1 U15099 ( .A(n12881), .ZN(n12816) );
  OAI21_X1 U15100 ( .B1(n12811), .B2(n12810), .A(n12809), .ZN(n12882) );
  AOI22_X1 U15101 ( .A1(n15005), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15103), 
        .B2(n12812), .ZN(n12813) );
  OAI21_X1 U15102 ( .B1(n12952), .B2(n12826), .A(n12813), .ZN(n12814) );
  AOI21_X1 U15103 ( .B1(n12882), .B2(n15020), .A(n12814), .ZN(n12815) );
  OAI21_X1 U15104 ( .B1(n12816), .B2(n15005), .A(n12815), .ZN(P3_U3217) );
  XOR2_X1 U15105 ( .A(n12817), .B(n12822), .Z(n12818) );
  OAI222_X1 U15106 ( .A1(n15046), .A2(n12820), .B1(n15044), .B2(n12819), .C1(
        n12818), .C2(n15052), .ZN(n12885) );
  INV_X1 U15107 ( .A(n12885), .ZN(n12829) );
  OAI21_X1 U15108 ( .B1(n12823), .B2(n12822), .A(n12821), .ZN(n12886) );
  AOI22_X1 U15109 ( .A1(n15005), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12824), 
        .B2(n15103), .ZN(n12825) );
  OAI21_X1 U15110 ( .B1(n12956), .B2(n12826), .A(n12825), .ZN(n12827) );
  AOI21_X1 U15111 ( .B1(n12886), .B2(n15020), .A(n12827), .ZN(n12828) );
  OAI21_X1 U15112 ( .B1(n12829), .B2(n15005), .A(n12828), .ZN(P3_U3218) );
  AOI22_X1 U15113 ( .A1(n12831), .A2(n15136), .B1(n14410), .B2(n6688), .ZN(
        n12832) );
  INV_X1 U15114 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12836) );
  AOI21_X1 U15115 ( .B1(n15140), .B2(n12835), .A(n12834), .ZN(n12912) );
  MUX2_X1 U15116 ( .A(n12836), .B(n12912), .S(n15159), .Z(n12837) );
  INV_X1 U15117 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12843) );
  OAI22_X1 U15118 ( .A1(n12840), .A2(n12839), .B1(n12838), .B2(n15076), .ZN(
        n12841) );
  NOR2_X1 U15119 ( .A1(n12842), .A2(n12841), .ZN(n12916) );
  MUX2_X1 U15120 ( .A(n12843), .B(n12916), .S(n15159), .Z(n12844) );
  INV_X1 U15121 ( .A(n12844), .ZN(P3_U3485) );
  AOI22_X1 U15122 ( .A1(n12846), .A2(n15140), .B1(n14410), .B2(n12845), .ZN(
        n12847) );
  NAND2_X1 U15123 ( .A1(n12848), .A2(n12847), .ZN(n12919) );
  MUX2_X1 U15124 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12919), .S(n15159), .Z(
        P3_U3484) );
  AOI22_X1 U15125 ( .A1(n12850), .A2(n15140), .B1(n14410), .B2(n12849), .ZN(
        n12851) );
  NAND2_X1 U15126 ( .A1(n12852), .A2(n12851), .ZN(n12920) );
  MUX2_X1 U15127 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12920), .S(n15159), .Z(
        P3_U3483) );
  INV_X1 U15128 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12855) );
  AOI21_X1 U15129 ( .B1(n15140), .B2(n12854), .A(n12853), .ZN(n12921) );
  MUX2_X1 U15130 ( .A(n12855), .B(n12921), .S(n15159), .Z(n12856) );
  OAI21_X1 U15131 ( .B1(n12924), .B2(n12899), .A(n12856), .ZN(P3_U3482) );
  INV_X1 U15132 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12859) );
  AOI21_X1 U15133 ( .B1(n15136), .B2(n12858), .A(n12857), .ZN(n12925) );
  MUX2_X1 U15134 ( .A(n12859), .B(n12925), .S(n15159), .Z(n12860) );
  OAI21_X1 U15135 ( .B1(n12928), .B2(n12899), .A(n12860), .ZN(P3_U3481) );
  INV_X1 U15136 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12863) );
  AOI21_X1 U15137 ( .B1(n12862), .B2(n15136), .A(n12861), .ZN(n12929) );
  MUX2_X1 U15138 ( .A(n12863), .B(n12929), .S(n15159), .Z(n12864) );
  OAI21_X1 U15139 ( .B1(n12932), .B2(n12899), .A(n12864), .ZN(P3_U3480) );
  INV_X1 U15140 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12867) );
  AOI21_X1 U15141 ( .B1(n12866), .B2(n15136), .A(n12865), .ZN(n12933) );
  MUX2_X1 U15142 ( .A(n12867), .B(n12933), .S(n15159), .Z(n12868) );
  OAI21_X1 U15143 ( .B1(n12936), .B2(n12899), .A(n12868), .ZN(P3_U3479) );
  INV_X1 U15144 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12871) );
  AOI21_X1 U15145 ( .B1(n12870), .B2(n15136), .A(n12869), .ZN(n12937) );
  MUX2_X1 U15146 ( .A(n12871), .B(n12937), .S(n15159), .Z(n12872) );
  OAI21_X1 U15147 ( .B1(n12899), .B2(n12940), .A(n12872), .ZN(P3_U3478) );
  AOI21_X1 U15148 ( .B1(n12874), .B2(n15136), .A(n12873), .ZN(n12941) );
  MUX2_X1 U15149 ( .A(n12875), .B(n12941), .S(n15159), .Z(n12876) );
  OAI21_X1 U15150 ( .B1(n12944), .B2(n12899), .A(n12876), .ZN(P3_U3477) );
  AOI21_X1 U15151 ( .B1(n12878), .B2(n15136), .A(n12877), .ZN(n12945) );
  MUX2_X1 U15152 ( .A(n12879), .B(n12945), .S(n15159), .Z(n12880) );
  OAI21_X1 U15153 ( .B1(n12948), .B2(n12899), .A(n12880), .ZN(P3_U3476) );
  AOI21_X1 U15154 ( .B1(n15136), .B2(n12882), .A(n12881), .ZN(n12949) );
  MUX2_X1 U15155 ( .A(n12883), .B(n12949), .S(n15159), .Z(n12884) );
  OAI21_X1 U15156 ( .B1(n12952), .B2(n12899), .A(n12884), .ZN(P3_U3475) );
  INV_X1 U15157 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12887) );
  AOI21_X1 U15158 ( .B1(n15136), .B2(n12886), .A(n12885), .ZN(n12953) );
  MUX2_X1 U15159 ( .A(n12887), .B(n12953), .S(n15159), .Z(n12888) );
  OAI21_X1 U15160 ( .B1(n12956), .B2(n12899), .A(n12888), .ZN(P3_U3474) );
  NAND2_X1 U15161 ( .A1(n12889), .A2(n15136), .ZN(n12890) );
  AND2_X1 U15162 ( .A1(n12891), .A2(n12890), .ZN(n12958) );
  MUX2_X1 U15163 ( .A(n12958), .B(n12892), .S(n9457), .Z(n12893) );
  OAI21_X1 U15164 ( .B1(n12960), .B2(n12899), .A(n12893), .ZN(P3_U3473) );
  NAND2_X1 U15165 ( .A1(n12894), .A2(n15136), .ZN(n12895) );
  NAND2_X1 U15166 ( .A1(n12896), .A2(n12895), .ZN(n12961) );
  MUX2_X1 U15167 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n12961), .S(n15159), .Z(
        n12897) );
  INV_X1 U15168 ( .A(n12897), .ZN(n12898) );
  OAI21_X1 U15169 ( .B1(n12899), .B2(n12964), .A(n12898), .ZN(P3_U3472) );
  OAI21_X1 U15170 ( .B1(n8973), .B2(n12900), .A(n15088), .ZN(n12904) );
  NAND2_X1 U15171 ( .A1(n15061), .A2(n15081), .ZN(n12901) );
  NAND2_X1 U15172 ( .A1(n12902), .A2(n12901), .ZN(n12903) );
  AOI21_X1 U15173 ( .B1(n12904), .B2(n15089), .A(n12903), .ZN(n12907) );
  XNOR2_X1 U15174 ( .A(n8973), .B(n12905), .ZN(n15100) );
  NAND2_X1 U15175 ( .A1(n15100), .A2(n15049), .ZN(n12906) );
  AND2_X1 U15176 ( .A1(n12907), .A2(n12906), .ZN(n15105) );
  NOR2_X1 U15177 ( .A1(n12908), .A2(n15076), .ZN(n15102) );
  AOI21_X1 U15178 ( .B1(n15100), .B2(n15140), .A(n15102), .ZN(n12909) );
  AND2_X1 U15179 ( .A1(n15105), .A2(n12909), .ZN(n15112) );
  INV_X1 U15180 ( .A(n15112), .ZN(n12910) );
  MUX2_X1 U15181 ( .A(n12910), .B(P3_REG1_REG_1__SCAN_IN), .S(n9457), .Z(
        P3_U3460) );
  MUX2_X1 U15182 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n12911), .S(n15143), .Z(
        P3_U3455) );
  MUX2_X1 U15183 ( .A(n12913), .B(n12912), .S(n15143), .Z(n12914) );
  MUX2_X1 U15184 ( .A(n12917), .B(n12916), .S(n15143), .Z(n12918) );
  INV_X1 U15185 ( .A(n12918), .ZN(P3_U3453) );
  MUX2_X1 U15186 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12919), .S(n15143), .Z(
        P3_U3452) );
  MUX2_X1 U15187 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12920), .S(n15143), .Z(
        P3_U3451) );
  MUX2_X1 U15188 ( .A(n12922), .B(n12921), .S(n15143), .Z(n12923) );
  OAI21_X1 U15189 ( .B1(n12924), .B2(n12965), .A(n12923), .ZN(P3_U3450) );
  MUX2_X1 U15190 ( .A(n12926), .B(n12925), .S(n15143), .Z(n12927) );
  OAI21_X1 U15191 ( .B1(n12928), .B2(n12965), .A(n12927), .ZN(P3_U3449) );
  MUX2_X1 U15192 ( .A(n12930), .B(n12929), .S(n15143), .Z(n12931) );
  OAI21_X1 U15193 ( .B1(n12932), .B2(n12965), .A(n12931), .ZN(P3_U3448) );
  MUX2_X1 U15194 ( .A(n12934), .B(n12933), .S(n15143), .Z(n12935) );
  OAI21_X1 U15195 ( .B1(n12936), .B2(n12965), .A(n12935), .ZN(P3_U3447) );
  INV_X1 U15196 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12938) );
  MUX2_X1 U15197 ( .A(n12938), .B(n12937), .S(n15143), .Z(n12939) );
  OAI21_X1 U15198 ( .B1(n12965), .B2(n12940), .A(n12939), .ZN(P3_U3446) );
  MUX2_X1 U15199 ( .A(n12942), .B(n12941), .S(n15143), .Z(n12943) );
  OAI21_X1 U15200 ( .B1(n12944), .B2(n12965), .A(n12943), .ZN(P3_U3444) );
  MUX2_X1 U15201 ( .A(n12946), .B(n12945), .S(n15143), .Z(n12947) );
  OAI21_X1 U15202 ( .B1(n12948), .B2(n12965), .A(n12947), .ZN(P3_U3441) );
  MUX2_X1 U15203 ( .A(n12950), .B(n12949), .S(n15143), .Z(n12951) );
  OAI21_X1 U15204 ( .B1(n12952), .B2(n12965), .A(n12951), .ZN(P3_U3438) );
  MUX2_X1 U15205 ( .A(n12954), .B(n12953), .S(n15143), .Z(n12955) );
  OAI21_X1 U15206 ( .B1(n12956), .B2(n12965), .A(n12955), .ZN(P3_U3435) );
  MUX2_X1 U15207 ( .A(n12958), .B(n12957), .S(n15142), .Z(n12959) );
  OAI21_X1 U15208 ( .B1(n12960), .B2(n12965), .A(n12959), .ZN(P3_U3432) );
  MUX2_X1 U15209 ( .A(n12961), .B(P3_REG0_REG_13__SCAN_IN), .S(n15142), .Z(
        n12962) );
  INV_X1 U15210 ( .A(n12962), .ZN(n12963) );
  OAI21_X1 U15211 ( .B1(n12965), .B2(n12964), .A(n12963), .ZN(P3_U3429) );
  MUX2_X1 U15212 ( .A(P3_D_REG_1__SCAN_IN), .B(n12966), .S(n12967), .Z(
        P3_U3377) );
  MUX2_X1 U15213 ( .A(P3_D_REG_0__SCAN_IN), .B(n12968), .S(n12967), .Z(
        P3_U3376) );
  NAND3_X1 U15214 ( .A1(n12969), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n12973) );
  NAND2_X1 U15215 ( .A1(n12970), .A2(n14288), .ZN(n12972) );
  NAND2_X1 U15216 ( .A1(n14287), .A2(SI_31_), .ZN(n12971) );
  OAI211_X1 U15217 ( .C1(n12974), .C2(n12973), .A(n12972), .B(n12971), .ZN(
        P3_U3264) );
  NAND2_X1 U15218 ( .A1(n8153), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12975) );
  OAI21_X1 U15219 ( .B1(n14275), .B2(n12976), .A(n12975), .ZN(n12977) );
  AOI21_X1 U15220 ( .B1(n12978), .B2(n14288), .A(n12977), .ZN(n12979) );
  INV_X1 U15221 ( .A(n12979), .ZN(P3_U3266) );
  NAND2_X1 U15222 ( .A1(n12980), .A2(n14288), .ZN(n12982) );
  OAI211_X1 U15223 ( .C1(n12983), .C2(n12992), .A(n12982), .B(n12981), .ZN(
        P3_U3267) );
  INV_X1 U15224 ( .A(n12984), .ZN(n12985) );
  OAI222_X1 U15225 ( .A1(P3_U3151), .A2(n12449), .B1(n12992), .B2(n12986), 
        .C1(n14277), .C2(n12985), .ZN(P3_U3268) );
  INV_X1 U15226 ( .A(n12987), .ZN(n12988) );
  OAI222_X1 U15227 ( .A1(n12990), .A2(P3_U3151), .B1(n12992), .B2(n12989), 
        .C1(n14277), .C2(n12988), .ZN(P3_U3269) );
  INV_X1 U15228 ( .A(n12991), .ZN(n12996) );
  OAI222_X1 U15229 ( .A1(n14277), .A2(n12996), .B1(P3_U3151), .B2(n12994), 
        .C1(n12993), .C2(n12992), .ZN(P3_U3270) );
  XOR2_X1 U15230 ( .A(n12998), .B(n12997), .Z(n13002) );
  OAI22_X1 U15231 ( .A1(n13039), .A2(n13404), .B1(n13242), .B2(n13408), .ZN(
        n13284) );
  AOI22_X1 U15232 ( .A1(n13284), .A2(n13056), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12999) );
  OAI21_X1 U15233 ( .B1(n13286), .B2(n13096), .A(n12999), .ZN(n13000) );
  AOI21_X1 U15234 ( .B1(n13466), .B2(n13086), .A(n13000), .ZN(n13001) );
  OAI21_X1 U15235 ( .B1(n13002), .B2(n13088), .A(n13001), .ZN(P2_U3188) );
  XOR2_X1 U15236 ( .A(n13004), .B(n13003), .Z(n13005) );
  NAND2_X1 U15237 ( .A1(n13005), .A2(n13093), .ZN(n13012) );
  INV_X1 U15238 ( .A(n13006), .ZN(n13007) );
  AOI22_X1 U15239 ( .A1(n13056), .A2(n13007), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13011) );
  INV_X1 U15240 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n13146) );
  OR2_X1 U15241 ( .A1(n13096), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n13010) );
  NAND2_X1 U15242 ( .A1(n13086), .A2(n6399), .ZN(n13009) );
  NAND4_X1 U15243 ( .A1(n13012), .A2(n13011), .A3(n13010), .A4(n13009), .ZN(
        P2_U3190) );
  INV_X1 U15244 ( .A(n13013), .ZN(n13015) );
  NOR2_X1 U15245 ( .A1(n13015), .A2(n13014), .ZN(n13016) );
  XNOR2_X1 U15246 ( .A(n13017), .B(n13016), .ZN(n13022) );
  OAI21_X1 U15247 ( .B1(n13097), .B2(n13350), .A(n13018), .ZN(n13020) );
  OAI22_X1 U15248 ( .A1(n13095), .A2(n13349), .B1(n13096), .B2(n13361), .ZN(
        n13019) );
  AOI211_X1 U15249 ( .C1(n13360), .C2(n13086), .A(n13020), .B(n13019), .ZN(
        n13021) );
  OAI21_X1 U15250 ( .B1(n13022), .B2(n13088), .A(n13021), .ZN(P2_U3191) );
  INV_X1 U15251 ( .A(n13023), .ZN(n13024) );
  NAND2_X1 U15252 ( .A1(n13105), .A2(n9498), .ZN(n13025) );
  XOR2_X1 U15253 ( .A(n6712), .B(n13025), .Z(n13027) );
  XNOR2_X1 U15254 ( .A(n13199), .B(n13027), .ZN(n13028) );
  XNOR2_X1 U15255 ( .A(n13029), .B(n13028), .ZN(n13034) );
  AOI22_X1 U15256 ( .A1(n13030), .A2(n13056), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13031) );
  OAI21_X1 U15257 ( .B1(n13193), .B2(n13096), .A(n13031), .ZN(n13032) );
  AOI21_X1 U15258 ( .B1(n13199), .B2(n13086), .A(n13032), .ZN(n13033) );
  OAI21_X1 U15259 ( .B1(n13034), .B2(n13088), .A(n13033), .ZN(P2_U3192) );
  AOI21_X1 U15260 ( .B1(n13036), .B2(n13035), .A(n13088), .ZN(n13038) );
  NAND2_X1 U15261 ( .A1(n13038), .A2(n13037), .ZN(n13043) );
  NOR2_X1 U15262 ( .A1(n13095), .A2(n13350), .ZN(n13041) );
  OAI22_X1 U15263 ( .A1(n13039), .A2(n13097), .B1(n13321), .B2(n13096), .ZN(
        n13040) );
  AOI211_X1 U15264 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(P2_U3088), .A(n13041), 
        .B(n13040), .ZN(n13042) );
  OAI211_X1 U15265 ( .C1(n13536), .C2(n13102), .A(n13043), .B(n13042), .ZN(
        P2_U3195) );
  INV_X1 U15266 ( .A(n13044), .ZN(n13045) );
  AOI21_X1 U15267 ( .B1(n13047), .B2(n13046), .A(n13045), .ZN(n13051) );
  NAND2_X1 U15268 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14795)
         );
  OAI21_X1 U15269 ( .B1(n13095), .B2(n13403), .A(n14795), .ZN(n13049) );
  OAI22_X1 U15270 ( .A1(n13097), .A2(n13407), .B1(n13096), .B2(n13413), .ZN(
        n13048) );
  AOI211_X1 U15271 ( .C1(n13505), .C2(n13086), .A(n13049), .B(n13048), .ZN(
        n13050) );
  OAI21_X1 U15272 ( .B1(n13051), .B2(n13088), .A(n13050), .ZN(P2_U3198) );
  OAI21_X1 U15273 ( .B1(n13054), .B2(n13053), .A(n13052), .ZN(n13055) );
  NAND2_X1 U15274 ( .A1(n13055), .A2(n13093), .ZN(n13060) );
  INV_X1 U15275 ( .A(n13391), .ZN(n13058) );
  INV_X1 U15276 ( .A(n13096), .ZN(n13078) );
  INV_X1 U15277 ( .A(n13056), .ZN(n13083) );
  AOI22_X1 U15278 ( .A1(n13113), .A2(n13312), .B1(n13115), .B2(n13311), .ZN(
        n13386) );
  NAND2_X1 U15279 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14809)
         );
  OAI21_X1 U15280 ( .B1(n13083), .B2(n13386), .A(n14809), .ZN(n13057) );
  AOI21_X1 U15281 ( .B1(n13058), .B2(n13078), .A(n13057), .ZN(n13059) );
  OAI211_X1 U15282 ( .C1(n13061), .C2(n13102), .A(n13060), .B(n13059), .ZN(
        P2_U3200) );
  OAI21_X1 U15283 ( .B1(n6644), .B2(n13063), .A(n13062), .ZN(n13065) );
  NAND2_X1 U15284 ( .A1(n13065), .A2(n13093), .ZN(n13069) );
  NOR2_X1 U15285 ( .A1(n13095), .A2(n13333), .ZN(n13067) );
  OAI22_X1 U15286 ( .A1(n13334), .A2(n13097), .B1(n13338), .B2(n13096), .ZN(
        n13066) );
  AOI211_X1 U15287 ( .C1(P2_REG3_REG_20__SCAN_IN), .C2(P2_U3088), .A(n13067), 
        .B(n13066), .ZN(n13068) );
  OAI211_X1 U15288 ( .C1(n13540), .C2(n13102), .A(n13069), .B(n13068), .ZN(
        P2_U3205) );
  NAND2_X1 U15289 ( .A1(n13071), .A2(n13070), .ZN(n13072) );
  XOR2_X1 U15290 ( .A(n13073), .B(n13072), .Z(n13080) );
  AND2_X1 U15291 ( .A1(n13110), .A2(n13312), .ZN(n13074) );
  AOI21_X1 U15292 ( .B1(n13111), .B2(n13311), .A(n13074), .ZN(n13296) );
  INV_X1 U15293 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13075) );
  OAI22_X1 U15294 ( .A1(n13296), .A2(n13083), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13075), .ZN(n13077) );
  NOR2_X1 U15295 ( .A1(n13532), .A2(n13102), .ZN(n13076) );
  AOI211_X1 U15296 ( .C1(n13078), .C2(n13302), .A(n13077), .B(n13076), .ZN(
        n13079) );
  OAI21_X1 U15297 ( .B1(n13080), .B2(n13088), .A(n13079), .ZN(P2_U3207) );
  XNOR2_X1 U15298 ( .A(n13082), .B(n13081), .ZN(n13089) );
  NOR2_X1 U15299 ( .A1(n13096), .A2(n13377), .ZN(n13085) );
  AOI22_X1 U15300 ( .A1(n13112), .A2(n13312), .B1(n13311), .B2(n13114), .ZN(
        n13369) );
  NAND2_X1 U15301 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14825)
         );
  OAI21_X1 U15302 ( .B1(n13369), .B2(n13083), .A(n14825), .ZN(n13084) );
  AOI211_X1 U15303 ( .C1(n13375), .C2(n13086), .A(n13085), .B(n13084), .ZN(
        n13087) );
  OAI21_X1 U15304 ( .B1(n13089), .B2(n13088), .A(n13087), .ZN(P2_U3210) );
  OAI21_X1 U15305 ( .B1(n13092), .B2(n13091), .A(n13090), .ZN(n13094) );
  NAND2_X1 U15306 ( .A1(n13094), .A2(n13093), .ZN(n13101) );
  NOR2_X1 U15307 ( .A1(n13095), .A2(n13258), .ZN(n13099) );
  OAI22_X1 U15308 ( .A1(n13097), .A2(n13223), .B1(n13096), .B2(n13224), .ZN(
        n13098) );
  AOI211_X1 U15309 ( .C1(P2_REG3_REG_26__SCAN_IN), .C2(P2_U3088), .A(n13099), 
        .B(n13098), .ZN(n13100) );
  OAI211_X1 U15310 ( .C1(n13522), .C2(n13102), .A(n13101), .B(n13100), .ZN(
        P2_U3212) );
  MUX2_X1 U15311 ( .A(n13183), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13130), .Z(
        P2_U3562) );
  MUX2_X1 U15312 ( .A(n13103), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13130), .Z(
        P2_U3561) );
  MUX2_X1 U15313 ( .A(n13104), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13130), .Z(
        P2_U3560) );
  MUX2_X1 U15314 ( .A(n13105), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13130), .Z(
        P2_U3559) );
  MUX2_X1 U15315 ( .A(n13106), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13130), .Z(
        P2_U3558) );
  MUX2_X1 U15316 ( .A(n13107), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13130), .Z(
        P2_U3557) );
  MUX2_X1 U15317 ( .A(n13108), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13130), .Z(
        P2_U3556) );
  MUX2_X1 U15318 ( .A(n13109), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13130), .Z(
        P2_U3555) );
  MUX2_X1 U15319 ( .A(n13110), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13130), .Z(
        P2_U3554) );
  MUX2_X1 U15320 ( .A(n13313), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13130), .Z(
        P2_U3553) );
  MUX2_X1 U15321 ( .A(n13111), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13130), .Z(
        P2_U3552) );
  MUX2_X1 U15322 ( .A(n13310), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13130), .Z(
        P2_U3551) );
  INV_X2 U15323 ( .A(P2_U3947), .ZN(n13130) );
  MUX2_X1 U15324 ( .A(n13112), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13130), .Z(
        P2_U3550) );
  MUX2_X1 U15325 ( .A(n13113), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13130), .Z(
        P2_U3549) );
  MUX2_X1 U15326 ( .A(n13114), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13130), .Z(
        P2_U3548) );
  MUX2_X1 U15327 ( .A(n13115), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13130), .Z(
        P2_U3547) );
  MUX2_X1 U15328 ( .A(n13116), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13130), .Z(
        P2_U3546) );
  MUX2_X1 U15329 ( .A(n13117), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13130), .Z(
        P2_U3545) );
  MUX2_X1 U15330 ( .A(n13118), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13130), .Z(
        P2_U3544) );
  MUX2_X1 U15331 ( .A(n13119), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13130), .Z(
        P2_U3543) );
  MUX2_X1 U15332 ( .A(n13120), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13130), .Z(
        P2_U3542) );
  MUX2_X1 U15333 ( .A(n13121), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13130), .Z(
        P2_U3541) );
  MUX2_X1 U15334 ( .A(n13122), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13130), .Z(
        P2_U3540) );
  MUX2_X1 U15335 ( .A(n13123), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13130), .Z(
        P2_U3539) );
  MUX2_X1 U15336 ( .A(n13124), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13130), .Z(
        P2_U3538) );
  MUX2_X1 U15337 ( .A(n13125), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13130), .Z(
        P2_U3537) );
  MUX2_X1 U15338 ( .A(n13126), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13130), .Z(
        P2_U3536) );
  MUX2_X1 U15339 ( .A(n13127), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13130), .Z(
        P2_U3535) );
  MUX2_X1 U15340 ( .A(n13128), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13130), .Z(
        P2_U3534) );
  MUX2_X1 U15341 ( .A(n9166), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13130), .Z(
        P2_U3533) );
  MUX2_X1 U15342 ( .A(n13129), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13130), .Z(
        P2_U3532) );
  MUX2_X1 U15343 ( .A(n13131), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13130), .Z(
        P2_U3531) );
  MUX2_X1 U15344 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9873), .S(n13136), .Z(
        n13134) );
  NAND3_X1 U15345 ( .A1(n13134), .A2(n13133), .A3(n13132), .ZN(n13135) );
  NAND3_X1 U15346 ( .A1(n14779), .A2(n13150), .A3(n13135), .ZN(n13145) );
  AOI22_X1 U15347 ( .A1(n14773), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n13144) );
  MUX2_X1 U15348 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9888), .S(n13136), .Z(
        n13139) );
  NAND3_X1 U15349 ( .A1(n13139), .A2(n13138), .A3(n13137), .ZN(n13140) );
  NAND3_X1 U15350 ( .A1(n14776), .A2(n13156), .A3(n13140), .ZN(n13143) );
  NAND2_X1 U15351 ( .A1(n14819), .A2(n13141), .ZN(n13142) );
  NAND4_X1 U15352 ( .A1(n13145), .A2(n13144), .A3(n13143), .A4(n13142), .ZN(
        P2_U3216) );
  OAI22_X1 U15353 ( .A1(n14827), .A2(n15170), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13146), .ZN(n13147) );
  AOI21_X1 U15354 ( .B1(n13148), .B2(n14819), .A(n13147), .ZN(n13162) );
  MUX2_X1 U15355 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9876), .S(n13154), .Z(
        n13151) );
  NAND3_X1 U15356 ( .A1(n13151), .A2(n13150), .A3(n13149), .ZN(n13152) );
  NAND3_X1 U15357 ( .A1(n14779), .A2(n13153), .A3(n13152), .ZN(n13161) );
  MUX2_X1 U15358 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10462), .S(n13154), .Z(
        n13157) );
  NAND3_X1 U15359 ( .A1(n13157), .A2(n13156), .A3(n13155), .ZN(n13158) );
  NAND3_X1 U15360 ( .A1(n14776), .A2(n13159), .A3(n13158), .ZN(n13160) );
  NAND3_X1 U15361 ( .A1(n13162), .A2(n13161), .A3(n13160), .ZN(P2_U3217) );
  INV_X1 U15362 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n13164) );
  OAI21_X1 U15363 ( .B1(n14827), .B2(n13164), .A(n13163), .ZN(n13165) );
  AOI21_X1 U15364 ( .B1(n13171), .B2(n14819), .A(n13165), .ZN(n13179) );
  MUX2_X1 U15365 ( .A(n10711), .B(P2_REG2_REG_7__SCAN_IN), .S(n13171), .Z(
        n13166) );
  NAND3_X1 U15366 ( .A1(n13168), .A2(n13167), .A3(n13166), .ZN(n13169) );
  NAND3_X1 U15367 ( .A1(n14776), .A2(n13170), .A3(n13169), .ZN(n13178) );
  MUX2_X1 U15368 ( .A(n9961), .B(P2_REG1_REG_7__SCAN_IN), .S(n13171), .Z(
        n13172) );
  NAND3_X1 U15369 ( .A1(n13174), .A2(n13173), .A3(n13172), .ZN(n13175) );
  NAND3_X1 U15370 ( .A1(n14779), .A2(n13176), .A3(n13175), .ZN(n13177) );
  NAND3_X1 U15371 ( .A1(n13179), .A2(n13178), .A3(n13177), .ZN(P2_U3221) );
  XNOR2_X1 U15372 ( .A(n13180), .B(n13187), .ZN(n13181) );
  NAND2_X1 U15373 ( .A1(n13429), .A2(n13422), .ZN(n13186) );
  AND2_X1 U15374 ( .A1(n13183), .A2(n13182), .ZN(n13432) );
  INV_X1 U15375 ( .A(n13432), .ZN(n13184) );
  NOR2_X1 U15376 ( .A1(n13384), .A2(n13184), .ZN(n13190) );
  AOI21_X1 U15377 ( .B1(n13384), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13190), 
        .ZN(n13185) );
  OAI211_X1 U15378 ( .C1(n13513), .C2(n13376), .A(n13186), .B(n13185), .ZN(
        P2_U3234) );
  INV_X1 U15379 ( .A(n13187), .ZN(n13188) );
  NAND2_X1 U15380 ( .A1(n13433), .A2(n13422), .ZN(n13192) );
  AOI21_X1 U15381 ( .B1(n13384), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13190), 
        .ZN(n13191) );
  OAI211_X1 U15382 ( .C1(n13517), .C2(n13376), .A(n13192), .B(n13191), .ZN(
        P2_U3235) );
  INV_X1 U15383 ( .A(n13193), .ZN(n13195) );
  AOI21_X1 U15384 ( .B1(n13195), .B2(n13339), .A(n13194), .ZN(n13205) );
  INV_X1 U15385 ( .A(n13196), .ZN(n13203) );
  NOR2_X1 U15386 ( .A1(n13356), .A2(n13197), .ZN(n13198) );
  AOI21_X1 U15387 ( .B1(n13199), .B2(n13416), .A(n13198), .ZN(n13200) );
  OAI21_X1 U15388 ( .B1(n13201), .B2(n13269), .A(n13200), .ZN(n13202) );
  AOI21_X1 U15389 ( .B1(n13203), .B2(n13373), .A(n13202), .ZN(n13204) );
  OAI21_X1 U15390 ( .B1(n13384), .B2(n13205), .A(n13204), .ZN(P2_U3237) );
  XNOR2_X1 U15391 ( .A(n13207), .B(n13206), .ZN(n13209) );
  AOI21_X1 U15392 ( .B1(n13209), .B2(n13352), .A(n13208), .ZN(n13446) );
  OR2_X1 U15393 ( .A1(n13211), .A2(n13210), .ZN(n13442) );
  NAND3_X1 U15394 ( .A1(n13442), .A2(n13441), .A3(n13373), .ZN(n13220) );
  OAI22_X1 U15395 ( .A1(n13427), .A2(n13213), .B1(n13212), .B2(n13412), .ZN(
        n13214) );
  AOI21_X1 U15396 ( .B1(n13444), .B2(n13416), .A(n13214), .ZN(n13219) );
  OAI21_X1 U15397 ( .B1(n13232), .B2(n13215), .A(n13420), .ZN(n13217) );
  NOR2_X1 U15398 ( .A1(n13217), .A2(n13216), .ZN(n13443) );
  NAND2_X1 U15399 ( .A1(n13443), .A2(n13422), .ZN(n13218) );
  OAI21_X1 U15400 ( .B1(n13384), .B2(n13446), .A(n13221), .ZN(P2_U3238) );
  NAND2_X1 U15401 ( .A1(n13448), .A2(n13427), .ZN(n13236) );
  OAI22_X1 U15402 ( .A1(n13356), .A2(n13225), .B1(n13224), .B2(n13412), .ZN(
        n13226) );
  AOI21_X1 U15403 ( .B1(n13229), .B2(n13416), .A(n13226), .ZN(n13235) );
  XNOR2_X1 U15404 ( .A(n13228), .B(n13227), .ZN(n13450) );
  NAND2_X1 U15405 ( .A1(n13450), .A2(n13373), .ZN(n13234) );
  NAND2_X1 U15406 ( .A1(n13244), .A2(n13229), .ZN(n13230) );
  NAND2_X1 U15407 ( .A1(n13230), .A2(n13420), .ZN(n13231) );
  NOR2_X1 U15408 ( .A1(n13232), .A2(n13231), .ZN(n13449) );
  NAND2_X1 U15409 ( .A1(n13449), .A2(n13422), .ZN(n13233) );
  NAND4_X1 U15410 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        P2_U3239) );
  XNOR2_X1 U15411 ( .A(n13237), .B(n13239), .ZN(n13455) );
  INV_X1 U15412 ( .A(n13455), .ZN(n13253) );
  AOI21_X1 U15413 ( .B1(n13240), .B2(n13239), .A(n13238), .ZN(n13241) );
  OAI222_X1 U15414 ( .A1(n13408), .A2(n13243), .B1(n13404), .B2(n13242), .C1(
        n13405), .C2(n13241), .ZN(n13453) );
  NAND2_X1 U15415 ( .A1(n13453), .A2(n13427), .ZN(n13252) );
  INV_X1 U15416 ( .A(n13244), .ZN(n13245) );
  AOI211_X1 U15417 ( .C1(n13246), .C2(n13262), .A(n13394), .B(n13245), .ZN(
        n13454) );
  NOR2_X1 U15418 ( .A1(n13526), .A2(n13376), .ZN(n13250) );
  OAI22_X1 U15419 ( .A1(n13427), .A2(n13248), .B1(n13247), .B2(n13412), .ZN(
        n13249) );
  AOI211_X1 U15420 ( .C1(n13454), .C2(n13422), .A(n13250), .B(n13249), .ZN(
        n13251) );
  OAI211_X1 U15421 ( .C1(n13253), .C2(n13425), .A(n13252), .B(n13251), .ZN(
        P2_U3240) );
  AOI21_X1 U15422 ( .B1(n13256), .B2(n13255), .A(n13254), .ZN(n13257) );
  OAI222_X1 U15423 ( .A1(n13408), .A2(n13258), .B1(n13404), .B2(n7922), .C1(
        n13405), .C2(n13257), .ZN(n13464) );
  AND2_X1 U15424 ( .A1(n13260), .A2(n13259), .ZN(n13458) );
  NOR3_X1 U15425 ( .A1(n13459), .A2(n13458), .A3(n13425), .ZN(n13271) );
  INV_X1 U15426 ( .A(n13279), .ZN(n13261) );
  AOI21_X1 U15427 ( .B1(n13261), .B2(n13267), .A(n13394), .ZN(n13263) );
  NAND2_X1 U15428 ( .A1(n13263), .A2(n13262), .ZN(n13460) );
  OAI22_X1 U15429 ( .A1(n13427), .A2(n13265), .B1(n13264), .B2(n13412), .ZN(
        n13266) );
  AOI21_X1 U15430 ( .B1(n13267), .B2(n13416), .A(n13266), .ZN(n13268) );
  OAI21_X1 U15431 ( .B1(n13460), .B2(n13269), .A(n13268), .ZN(n13270) );
  AOI211_X1 U15432 ( .C1(n13464), .C2(n13356), .A(n13271), .B(n13270), .ZN(
        n13272) );
  INV_X1 U15433 ( .A(n13272), .ZN(P2_U3241) );
  OAI21_X1 U15434 ( .B1(n13275), .B2(n13274), .A(n13273), .ZN(n13276) );
  INV_X1 U15435 ( .A(n13276), .ZN(n13469) );
  NAND2_X1 U15436 ( .A1(n13466), .A2(n13301), .ZN(n13277) );
  NAND2_X1 U15437 ( .A1(n13277), .A2(n13420), .ZN(n13278) );
  NOR2_X1 U15438 ( .A1(n13279), .A2(n13278), .ZN(n13465) );
  OAI22_X1 U15439 ( .A1(n13281), .A2(n13376), .B1(n13427), .B2(n13280), .ZN(
        n13282) );
  AOI21_X1 U15440 ( .B1(n13465), .B2(n13422), .A(n13282), .ZN(n13289) );
  XNOR2_X1 U15441 ( .A(n13283), .B(n7329), .ZN(n13285) );
  AOI21_X1 U15442 ( .B1(n13285), .B2(n13352), .A(n13284), .ZN(n13468) );
  OAI21_X1 U15443 ( .B1(n13286), .B2(n13412), .A(n13468), .ZN(n13287) );
  NAND2_X1 U15444 ( .A1(n13287), .A2(n13427), .ZN(n13288) );
  OAI211_X1 U15445 ( .C1(n13469), .C2(n13425), .A(n13289), .B(n13288), .ZN(
        P2_U3242) );
  NAND2_X1 U15446 ( .A1(n13291), .A2(n13293), .ZN(n13292) );
  NAND2_X1 U15447 ( .A1(n13290), .A2(n13292), .ZN(n13473) );
  NOR2_X1 U15448 ( .A1(n6539), .A2(n13293), .ZN(n13295) );
  OR3_X1 U15449 ( .A1(n13295), .A2(n13294), .A3(n13405), .ZN(n13297) );
  NAND2_X1 U15450 ( .A1(n13297), .A2(n13296), .ZN(n13471) );
  INV_X1 U15451 ( .A(n13318), .ZN(n13298) );
  AOI21_X1 U15452 ( .B1(n13299), .B2(n13298), .A(n13394), .ZN(n13300) );
  AND2_X1 U15453 ( .A1(n13301), .A2(n13300), .ZN(n13470) );
  NAND2_X1 U15454 ( .A1(n13470), .A2(n13422), .ZN(n13304) );
  AOI22_X1 U15455 ( .A1(n13302), .A2(n13339), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n13384), .ZN(n13303) );
  OAI211_X1 U15456 ( .C1(n13532), .C2(n13376), .A(n13304), .B(n13303), .ZN(
        n13305) );
  AOI21_X1 U15457 ( .B1(n13471), .B2(n13356), .A(n13305), .ZN(n13306) );
  OAI21_X1 U15458 ( .B1(n13473), .B2(n13425), .A(n13306), .ZN(P2_U3243) );
  XNOR2_X1 U15459 ( .A(n13308), .B(n13307), .ZN(n13309) );
  NAND2_X1 U15460 ( .A1(n13309), .A2(n13352), .ZN(n13315) );
  AOI22_X1 U15461 ( .A1(n13313), .A2(n13312), .B1(n13311), .B2(n13310), .ZN(
        n13314) );
  NAND2_X1 U15462 ( .A1(n13315), .A2(n13314), .ZN(n13476) );
  INV_X1 U15463 ( .A(n13476), .ZN(n13326) );
  XNOR2_X1 U15464 ( .A(n13317), .B(n13316), .ZN(n13478) );
  NAND2_X1 U15465 ( .A1(n13478), .A2(n13373), .ZN(n13325) );
  AOI211_X1 U15466 ( .C1(n13319), .C2(n13335), .A(n13394), .B(n13318), .ZN(
        n13477) );
  NOR2_X1 U15467 ( .A1(n13536), .A2(n13376), .ZN(n13323) );
  OAI22_X1 U15468 ( .A1(n13321), .A2(n13412), .B1(n13320), .B2(n13356), .ZN(
        n13322) );
  AOI211_X1 U15469 ( .C1(n13477), .C2(n13422), .A(n13323), .B(n13322), .ZN(
        n13324) );
  OAI211_X1 U15470 ( .C1(n13384), .C2(n13326), .A(n13325), .B(n13324), .ZN(
        P2_U3244) );
  XOR2_X1 U15471 ( .A(n13331), .B(n13327), .Z(n13483) );
  INV_X1 U15472 ( .A(n13483), .ZN(n13345) );
  INV_X1 U15473 ( .A(n13328), .ZN(n13329) );
  AOI21_X1 U15474 ( .B1(n13331), .B2(n13330), .A(n13329), .ZN(n13332) );
  OAI222_X1 U15475 ( .A1(n13408), .A2(n13334), .B1(n13404), .B2(n13333), .C1(
        n13405), .C2(n13332), .ZN(n13481) );
  INV_X1 U15476 ( .A(n13335), .ZN(n13336) );
  AOI211_X1 U15477 ( .C1(n13337), .C2(n13357), .A(n13394), .B(n13336), .ZN(
        n13482) );
  NAND2_X1 U15478 ( .A1(n13482), .A2(n13422), .ZN(n13342) );
  INV_X1 U15479 ( .A(n13338), .ZN(n13340) );
  AOI22_X1 U15480 ( .A1(n13384), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13340), 
        .B2(n13339), .ZN(n13341) );
  OAI211_X1 U15481 ( .C1(n13540), .C2(n13376), .A(n13342), .B(n13341), .ZN(
        n13343) );
  AOI21_X1 U15482 ( .B1(n13481), .B2(n13356), .A(n13343), .ZN(n13344) );
  OAI21_X1 U15483 ( .B1(n13345), .B2(n13425), .A(n13344), .ZN(P2_U3245) );
  XOR2_X1 U15484 ( .A(n13348), .B(n13346), .Z(n13486) );
  XOR2_X1 U15485 ( .A(n13348), .B(n13347), .Z(n13353) );
  OAI22_X1 U15486 ( .A1(n13350), .A2(n13408), .B1(n13349), .B2(n13404), .ZN(
        n13351) );
  AOI21_X1 U15487 ( .B1(n13353), .B2(n13352), .A(n13351), .ZN(n13354) );
  OAI21_X1 U15488 ( .B1(n13486), .B2(n13355), .A(n13354), .ZN(n13487) );
  NAND2_X1 U15489 ( .A1(n13487), .A2(n13356), .ZN(n13366) );
  INV_X1 U15490 ( .A(n13357), .ZN(n13358) );
  AOI211_X1 U15491 ( .C1(n13360), .C2(n13359), .A(n13394), .B(n13358), .ZN(
        n13488) );
  NOR2_X1 U15492 ( .A1(n13544), .A2(n13376), .ZN(n13364) );
  OAI22_X1 U15493 ( .A1(n13427), .A2(n13362), .B1(n13361), .B2(n13412), .ZN(
        n13363) );
  AOI211_X1 U15494 ( .C1(n13488), .C2(n13422), .A(n13364), .B(n13363), .ZN(
        n13365) );
  OAI211_X1 U15495 ( .C1(n13486), .C2(n13367), .A(n13366), .B(n13365), .ZN(
        P2_U3246) );
  XNOR2_X1 U15496 ( .A(n13368), .B(n13371), .ZN(n13370) );
  OAI21_X1 U15497 ( .B1(n13370), .B2(n13405), .A(n13369), .ZN(n13492) );
  INV_X1 U15498 ( .A(n13492), .ZN(n13383) );
  XNOR2_X1 U15499 ( .A(n13372), .B(n13371), .ZN(n13494) );
  NAND2_X1 U15500 ( .A1(n13494), .A2(n13373), .ZN(n13382) );
  AOI211_X1 U15501 ( .C1(n13375), .C2(n13395), .A(n13394), .B(n13374), .ZN(
        n13493) );
  NOR2_X1 U15502 ( .A1(n6951), .A2(n13376), .ZN(n13380) );
  OAI22_X1 U15503 ( .A1(n13427), .A2(n13378), .B1(n13377), .B2(n13412), .ZN(
        n13379) );
  AOI211_X1 U15504 ( .C1(n13493), .C2(n13422), .A(n13380), .B(n13379), .ZN(
        n13381) );
  OAI211_X1 U15505 ( .C1(n13384), .C2(n13383), .A(n13382), .B(n13381), .ZN(
        P2_U3247) );
  XNOR2_X1 U15506 ( .A(n13385), .B(n13389), .ZN(n13387) );
  OAI21_X1 U15507 ( .B1(n13387), .B2(n13405), .A(n13386), .ZN(n13498) );
  OAI21_X1 U15508 ( .B1(n13390), .B2(n13389), .A(n13388), .ZN(n13502) );
  OAI22_X1 U15509 ( .A1(n13427), .A2(n13392), .B1(n13391), .B2(n13412), .ZN(
        n13393) );
  AOI21_X1 U15510 ( .B1(n13500), .B2(n13416), .A(n13393), .ZN(n13398) );
  AOI21_X1 U15511 ( .B1(n13421), .B2(n13500), .A(n13394), .ZN(n13396) );
  AND2_X1 U15512 ( .A1(n13396), .A2(n13395), .ZN(n13499) );
  NAND2_X1 U15513 ( .A1(n13499), .A2(n13422), .ZN(n13397) );
  OAI211_X1 U15514 ( .C1(n13502), .C2(n13425), .A(n13398), .B(n13397), .ZN(
        n13399) );
  AOI21_X1 U15515 ( .B1(n13427), .B2(n13498), .A(n13399), .ZN(n13400) );
  INV_X1 U15516 ( .A(n13400), .ZN(P2_U3248) );
  XNOR2_X1 U15517 ( .A(n13402), .B(n13401), .ZN(n13406) );
  OAI222_X1 U15518 ( .A1(n13408), .A2(n13407), .B1(n13406), .B2(n13405), .C1(
        n13404), .C2(n13403), .ZN(n13503) );
  OAI21_X1 U15519 ( .B1(n13411), .B2(n13410), .A(n13409), .ZN(n13508) );
  OAI22_X1 U15520 ( .A1(n13427), .A2(n13414), .B1(n13413), .B2(n13412), .ZN(
        n13415) );
  AOI21_X1 U15521 ( .B1(n13505), .B2(n13416), .A(n13415), .ZN(n13424) );
  OR2_X1 U15522 ( .A1(n13418), .A2(n13417), .ZN(n13419) );
  AND3_X1 U15523 ( .A1(n13421), .A2(n13420), .A3(n13419), .ZN(n13504) );
  NAND2_X1 U15524 ( .A1(n13504), .A2(n13422), .ZN(n13423) );
  OAI211_X1 U15525 ( .C1(n13508), .C2(n13425), .A(n13424), .B(n13423), .ZN(
        n13426) );
  AOI21_X1 U15526 ( .B1(n13427), .B2(n13503), .A(n13426), .ZN(n13428) );
  INV_X1 U15527 ( .A(n13428), .ZN(P2_U3249) );
  NOR2_X1 U15528 ( .A1(n13429), .A2(n13432), .ZN(n13510) );
  MUX2_X1 U15529 ( .A(n13430), .B(n13510), .S(n14857), .Z(n13431) );
  OAI21_X1 U15530 ( .B1(n13513), .B2(n13497), .A(n13431), .ZN(P2_U3530) );
  NOR2_X1 U15531 ( .A1(n13433), .A2(n13432), .ZN(n13514) );
  MUX2_X1 U15532 ( .A(n13434), .B(n13514), .S(n14857), .Z(n13435) );
  OAI21_X1 U15533 ( .B1(n13517), .B2(n13497), .A(n13435), .ZN(P2_U3529) );
  AOI21_X1 U15534 ( .B1(n13506), .B2(n13437), .A(n13436), .ZN(n13438) );
  MUX2_X1 U15535 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13518), .S(n14857), .Z(
        P2_U3528) );
  NAND3_X1 U15536 ( .A1(n13442), .A2(n13441), .A3(n14440), .ZN(n13447) );
  AOI21_X1 U15537 ( .B1(n13506), .B2(n13444), .A(n13443), .ZN(n13445) );
  NAND3_X1 U15538 ( .A1(n13447), .A2(n13446), .A3(n13445), .ZN(n13519) );
  MUX2_X1 U15539 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13519), .S(n14857), .Z(
        P2_U3526) );
  MUX2_X1 U15540 ( .A(n13451), .B(n13520), .S(n14857), .Z(n13452) );
  OAI21_X1 U15541 ( .B1(n13522), .B2(n13497), .A(n13452), .ZN(P2_U3525) );
  AOI211_X1 U15542 ( .C1(n14440), .C2(n13455), .A(n13454), .B(n13453), .ZN(
        n13523) );
  MUX2_X1 U15543 ( .A(n13456), .B(n13523), .S(n14857), .Z(n13457) );
  OAI21_X1 U15544 ( .B1(n13526), .B2(n13497), .A(n13457), .ZN(P2_U3524) );
  NOR3_X1 U15545 ( .A1(n13459), .A2(n13458), .A3(n14428), .ZN(n13463) );
  OAI21_X1 U15546 ( .B1(n13461), .B2(n14849), .A(n13460), .ZN(n13462) );
  MUX2_X1 U15547 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13527), .S(n14857), .Z(
        P2_U3523) );
  AOI21_X1 U15548 ( .B1(n13506), .B2(n13466), .A(n13465), .ZN(n13467) );
  OAI211_X1 U15549 ( .C1(n13469), .C2(n14428), .A(n13468), .B(n13467), .ZN(
        n13528) );
  MUX2_X1 U15550 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13528), .S(n14857), .Z(
        P2_U3522) );
  NOR2_X1 U15551 ( .A1(n13471), .A2(n13470), .ZN(n13472) );
  OAI21_X1 U15552 ( .B1(n13473), .B2(n14428), .A(n13472), .ZN(n13529) );
  MUX2_X1 U15553 ( .A(n13529), .B(P2_REG1_REG_22__SCAN_IN), .S(n8929), .Z(
        n13474) );
  INV_X1 U15554 ( .A(n13474), .ZN(n13475) );
  OAI21_X1 U15555 ( .B1(n13532), .B2(n13497), .A(n13475), .ZN(P2_U3521) );
  INV_X1 U15556 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13479) );
  AOI211_X1 U15557 ( .C1(n13478), .C2(n14440), .A(n13477), .B(n13476), .ZN(
        n13533) );
  MUX2_X1 U15558 ( .A(n13479), .B(n13533), .S(n14857), .Z(n13480) );
  OAI21_X1 U15559 ( .B1(n13536), .B2(n13497), .A(n13480), .ZN(P2_U3520) );
  INV_X1 U15560 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n13484) );
  AOI211_X1 U15561 ( .C1(n13483), .C2(n14440), .A(n13482), .B(n13481), .ZN(
        n13537) );
  MUX2_X1 U15562 ( .A(n13484), .B(n13537), .S(n14857), .Z(n13485) );
  OAI21_X1 U15563 ( .B1(n13540), .B2(n13497), .A(n13485), .ZN(P2_U3519) );
  INV_X1 U15564 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13490) );
  INV_X1 U15565 ( .A(n13486), .ZN(n13489) );
  AOI211_X1 U15566 ( .C1(n13489), .C2(n9151), .A(n13488), .B(n13487), .ZN(
        n13541) );
  MUX2_X1 U15567 ( .A(n13490), .B(n13541), .S(n14857), .Z(n13491) );
  OAI21_X1 U15568 ( .B1(n13544), .B2(n13497), .A(n13491), .ZN(P2_U3518) );
  AOI211_X1 U15569 ( .C1(n13494), .C2(n14440), .A(n13493), .B(n13492), .ZN(
        n13545) );
  MUX2_X1 U15570 ( .A(n13495), .B(n13545), .S(n14857), .Z(n13496) );
  OAI21_X1 U15571 ( .B1(n6951), .B2(n13497), .A(n13496), .ZN(P2_U3517) );
  AOI211_X1 U15572 ( .C1(n13506), .C2(n13500), .A(n13499), .B(n13498), .ZN(
        n13501) );
  OAI21_X1 U15573 ( .B1(n14428), .B2(n13502), .A(n13501), .ZN(n13549) );
  MUX2_X1 U15574 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13549), .S(n14857), .Z(
        P2_U3516) );
  AOI211_X1 U15575 ( .C1(n13506), .C2(n13505), .A(n13504), .B(n13503), .ZN(
        n13507) );
  OAI21_X1 U15576 ( .B1(n14428), .B2(n13508), .A(n13507), .ZN(n13550) );
  MUX2_X1 U15577 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13550), .S(n14857), .Z(
        P2_U3515) );
  MUX2_X1 U15578 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n13509), .S(n14857), .Z(
        P2_U3499) );
  INV_X1 U15579 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13511) );
  MUX2_X1 U15580 ( .A(n13511), .B(n13510), .S(n14457), .Z(n13512) );
  OAI21_X1 U15581 ( .B1(n13513), .B2(n13548), .A(n13512), .ZN(P2_U3498) );
  INV_X1 U15582 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13515) );
  MUX2_X1 U15583 ( .A(n13515), .B(n13514), .S(n14457), .Z(n13516) );
  OAI21_X1 U15584 ( .B1(n13517), .B2(n13548), .A(n13516), .ZN(P2_U3497) );
  MUX2_X1 U15585 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13518), .S(n14457), .Z(
        P2_U3496) );
  MUX2_X1 U15586 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13519), .S(n14457), .Z(
        P2_U3494) );
  INV_X1 U15587 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n13521) );
  INV_X1 U15588 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13524) );
  MUX2_X1 U15589 ( .A(n13524), .B(n13523), .S(n14457), .Z(n13525) );
  OAI21_X1 U15590 ( .B1(n13526), .B2(n13548), .A(n13525), .ZN(P2_U3492) );
  MUX2_X1 U15591 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13527), .S(n14457), .Z(
        P2_U3491) );
  MUX2_X1 U15592 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13528), .S(n14457), .Z(
        P2_U3490) );
  MUX2_X1 U15593 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13529), .S(n14457), .Z(
        n13530) );
  INV_X1 U15594 ( .A(n13530), .ZN(n13531) );
  OAI21_X1 U15595 ( .B1(n13532), .B2(n13548), .A(n13531), .ZN(P2_U3489) );
  INV_X1 U15596 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13534) );
  MUX2_X1 U15597 ( .A(n13534), .B(n13533), .S(n14854), .Z(n13535) );
  OAI21_X1 U15598 ( .B1(n13536), .B2(n13548), .A(n13535), .ZN(P2_U3488) );
  INV_X1 U15599 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n13538) );
  MUX2_X1 U15600 ( .A(n13538), .B(n13537), .S(n14854), .Z(n13539) );
  OAI21_X1 U15601 ( .B1(n13540), .B2(n13548), .A(n13539), .ZN(P2_U3487) );
  INV_X1 U15602 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13542) );
  MUX2_X1 U15603 ( .A(n13542), .B(n13541), .S(n14457), .Z(n13543) );
  OAI21_X1 U15604 ( .B1(n13544), .B2(n13548), .A(n13543), .ZN(P2_U3486) );
  INV_X1 U15605 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n13546) );
  MUX2_X1 U15606 ( .A(n13546), .B(n13545), .S(n14457), .Z(n13547) );
  OAI21_X1 U15607 ( .B1(n6951), .B2(n13548), .A(n13547), .ZN(P2_U3484) );
  MUX2_X1 U15608 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13549), .S(n14457), .Z(
        P2_U3481) );
  MUX2_X1 U15609 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13550), .S(n14457), .Z(
        P2_U3478) );
  NAND3_X1 U15610 ( .A1(n13552), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13554) );
  OAI22_X1 U15611 ( .A1(n13551), .A2(n13554), .B1(n13553), .B2(n13573), .ZN(
        n13555) );
  AOI21_X1 U15612 ( .B1(n14226), .B2(n13557), .A(n13555), .ZN(n13556) );
  INV_X1 U15613 ( .A(n13556), .ZN(P2_U3296) );
  NAND2_X1 U15614 ( .A1(n14235), .A2(n13557), .ZN(n13559) );
  OAI211_X1 U15615 ( .C1(n13561), .C2(n13560), .A(n13559), .B(n13558), .ZN(
        P2_U3299) );
  INV_X1 U15616 ( .A(n13562), .ZN(n14239) );
  OAI222_X1 U15617 ( .A1(n13564), .A2(P2_U3088), .B1(n13575), .B2(n14239), 
        .C1(n13563), .C2(n13573), .ZN(P2_U3300) );
  INV_X1 U15618 ( .A(n13565), .ZN(n14241) );
  OAI222_X1 U15619 ( .A1(P2_U3088), .A2(n13567), .B1(n13575), .B2(n14241), 
        .C1(n13566), .C2(n13573), .ZN(P2_U3301) );
  INV_X1 U15620 ( .A(n13568), .ZN(n14243) );
  OAI222_X1 U15621 ( .A1(n13570), .A2(P2_U3088), .B1(n13575), .B2(n14243), 
        .C1(n13569), .C2(n13573), .ZN(P2_U3302) );
  INV_X1 U15622 ( .A(n13571), .ZN(n13576) );
  INV_X1 U15623 ( .A(n13572), .ZN(n14249) );
  OAI222_X1 U15624 ( .A1(P2_U3088), .A2(n13576), .B1(n13575), .B2(n14249), 
        .C1(n13574), .C2(n13573), .ZN(P2_U3303) );
  INV_X1 U15625 ( .A(n13577), .ZN(n13578) );
  MUX2_X1 U15626 ( .A(n13578), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15627 ( .A(n13580), .B(n13579), .Z(n13586) );
  NAND2_X1 U15628 ( .A1(n13893), .A2(n13691), .ZN(n13582) );
  NAND2_X1 U15629 ( .A1(n13891), .A2(n14100), .ZN(n13581) );
  NAND2_X1 U15630 ( .A1(n13582), .A2(n13581), .ZN(n13990) );
  AOI22_X1 U15631 ( .A1(n13990), .A2(n14472), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13583) );
  OAI21_X1 U15632 ( .B1(n13992), .B2(n14479), .A(n13583), .ZN(n13584) );
  AOI21_X1 U15633 ( .B1(n14159), .B2(n14475), .A(n13584), .ZN(n13585) );
  OAI21_X1 U15634 ( .B1(n13586), .B2(n13705), .A(n13585), .ZN(P1_U3216) );
  INV_X1 U15635 ( .A(n13587), .ZN(n13588) );
  OAI211_X1 U15636 ( .C1(n13590), .C2(n13589), .A(n13588), .B(n14470), .ZN(
        n13600) );
  NAND2_X1 U15637 ( .A1(n13592), .A2(n13591), .ZN(n13594) );
  AOI21_X1 U15638 ( .B1(n14472), .B2(n13594), .A(n13593), .ZN(n13599) );
  NAND2_X1 U15639 ( .A1(n14475), .A2(n13595), .ZN(n13598) );
  OR2_X1 U15640 ( .A1(n14479), .A2(n13596), .ZN(n13597) );
  NAND4_X1 U15641 ( .A1(n13600), .A2(n13599), .A3(n13598), .A4(n13597), .ZN(
        P1_U3217) );
  INV_X1 U15642 ( .A(n14060), .ZN(n14181) );
  AOI21_X1 U15643 ( .B1(n13602), .B2(n13601), .A(n13705), .ZN(n13604) );
  NAND2_X1 U15644 ( .A1(n13604), .A2(n13603), .ZN(n13608) );
  AND2_X1 U15645 ( .A1(n13886), .A2(n14100), .ZN(n13605) );
  AOI21_X1 U15646 ( .B1(n13888), .B2(n13854), .A(n13605), .ZN(n14179) );
  NAND2_X1 U15647 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13849)
         );
  OAI21_X1 U15648 ( .B1(n14179), .B2(n13712), .A(n13849), .ZN(n13606) );
  AOI21_X1 U15649 ( .B1(n14055), .B2(n13714), .A(n13606), .ZN(n13607) );
  OAI211_X1 U15650 ( .C1(n14181), .C2(n13718), .A(n13608), .B(n13607), .ZN(
        P1_U3219) );
  INV_X1 U15651 ( .A(n13609), .ZN(n13610) );
  AOI21_X1 U15652 ( .B1(n13612), .B2(n13611), .A(n13610), .ZN(n13617) );
  OAI22_X1 U15653 ( .A1(n13875), .A2(n14098), .B1(n13613), .B2(n13903), .ZN(
        n14169) );
  AOI22_X1 U15654 ( .A1(n14169), .A2(n14472), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13614) );
  OAI21_X1 U15655 ( .B1(n14024), .B2(n14479), .A(n13614), .ZN(n13615) );
  AOI21_X1 U15656 ( .B1(n14170), .B2(n14475), .A(n13615), .ZN(n13616) );
  OAI21_X1 U15657 ( .B1(n13617), .B2(n13705), .A(n13616), .ZN(P1_U3223) );
  XOR2_X1 U15658 ( .A(n13620), .B(n13619), .Z(n13625) );
  AND2_X1 U15659 ( .A1(n13893), .A2(n14100), .ZN(n13621) );
  AOI21_X1 U15660 ( .B1(n13720), .B2(n13854), .A(n13621), .ZN(n14146) );
  AOI22_X1 U15661 ( .A1(n13965), .A2(n13714), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13622) );
  OAI21_X1 U15662 ( .B1(n14146), .B2(n13712), .A(n13622), .ZN(n13623) );
  AOI21_X1 U15663 ( .B1(n13969), .B2(n14475), .A(n13623), .ZN(n13624) );
  OAI21_X1 U15664 ( .B1(n13625), .B2(n13705), .A(n13624), .ZN(P1_U3225) );
  INV_X1 U15665 ( .A(n13627), .ZN(n13628) );
  AOI21_X1 U15666 ( .B1(n13629), .B2(n13626), .A(n13628), .ZN(n13636) );
  NOR2_X1 U15667 ( .A1(n14479), .A2(n13630), .ZN(n13634) );
  OAI21_X1 U15668 ( .B1(n13712), .B2(n13632), .A(n13631), .ZN(n13633) );
  AOI211_X1 U15669 ( .C1(n14197), .C2(n14475), .A(n13634), .B(n13633), .ZN(
        n13635) );
  OAI21_X1 U15670 ( .B1(n13636), .B2(n13705), .A(n13635), .ZN(P1_U3226) );
  INV_X1 U15671 ( .A(n14192), .ZN(n14089) );
  OAI21_X1 U15672 ( .B1(n13639), .B2(n13638), .A(n13637), .ZN(n13640) );
  NAND2_X1 U15673 ( .A1(n13640), .A2(n14470), .ZN(n13646) );
  INV_X1 U15674 ( .A(n13641), .ZN(n14086) );
  AND2_X1 U15675 ( .A1(n13880), .A2(n14100), .ZN(n13642) );
  AOI21_X1 U15676 ( .B1(n13886), .B2(n13691), .A(n13642), .ZN(n14081) );
  OAI21_X1 U15677 ( .B1(n13712), .B2(n14081), .A(n13643), .ZN(n13644) );
  AOI21_X1 U15678 ( .B1(n14086), .B2(n13714), .A(n13644), .ZN(n13645) );
  OAI211_X1 U15679 ( .C1(n14089), .C2(n13718), .A(n13646), .B(n13645), .ZN(
        P1_U3228) );
  XOR2_X1 U15680 ( .A(n13648), .B(n13647), .Z(n13654) );
  AND2_X1 U15681 ( .A1(n13876), .A2(n14100), .ZN(n13649) );
  AOI21_X1 U15682 ( .B1(n13894), .B2(n13691), .A(n13649), .ZN(n13975) );
  OAI22_X1 U15683 ( .A1(n13975), .A2(n13712), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13650), .ZN(n13652) );
  NOR2_X1 U15684 ( .A1(n14153), .A2(n13718), .ZN(n13651) );
  AOI211_X1 U15685 ( .C1(n13714), .C2(n13982), .A(n13652), .B(n13651), .ZN(
        n13653) );
  OAI21_X1 U15686 ( .B1(n13654), .B2(n13705), .A(n13653), .ZN(P1_U3229) );
  INV_X1 U15687 ( .A(n14175), .ZN(n14040) );
  OAI211_X1 U15688 ( .C1(n13657), .C2(n13656), .A(n13655), .B(n14470), .ZN(
        n13661) );
  AOI22_X1 U15689 ( .A1(n13874), .A2(n13854), .B1(n13887), .B2(n14100), .ZN(
        n14034) );
  OAI22_X1 U15690 ( .A1(n14034), .A2(n13712), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13658), .ZN(n13659) );
  AOI21_X1 U15691 ( .B1(n14038), .B2(n13714), .A(n13659), .ZN(n13660) );
  OAI211_X1 U15692 ( .C1(n14040), .C2(n13718), .A(n13661), .B(n13660), .ZN(
        P1_U3233) );
  OAI211_X1 U15693 ( .C1(n13663), .C2(n13662), .A(n14459), .B(n14470), .ZN(
        n13669) );
  INV_X1 U15694 ( .A(n13664), .ZN(n13667) );
  NOR2_X1 U15695 ( .A1(n14479), .A2(n13665), .ZN(n13666) );
  AOI211_X1 U15696 ( .C1(n14472), .C2(n14490), .A(n13667), .B(n13666), .ZN(
        n13668) );
  OAI211_X1 U15697 ( .C1(n14493), .C2(n13718), .A(n13669), .B(n13668), .ZN(
        P1_U3234) );
  OAI21_X1 U15698 ( .B1(n13672), .B2(n13671), .A(n13670), .ZN(n13673) );
  NAND2_X1 U15699 ( .A1(n13673), .A2(n14470), .ZN(n13678) );
  AND2_X1 U15700 ( .A1(n13874), .A2(n14100), .ZN(n13674) );
  AOI21_X1 U15701 ( .B1(n13876), .B2(n13691), .A(n13674), .ZN(n14011) );
  OAI22_X1 U15702 ( .A1(n14011), .A2(n13712), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13675), .ZN(n13676) );
  AOI21_X1 U15703 ( .B1(n14005), .B2(n13714), .A(n13676), .ZN(n13677) );
  OAI211_X1 U15704 ( .C1(n13718), .C2(n14007), .A(n13678), .B(n13677), .ZN(
        P1_U3235) );
  XOR2_X1 U15705 ( .A(n13680), .B(n13679), .Z(n13687) );
  INV_X1 U15706 ( .A(n13884), .ZN(n13681) );
  OAI22_X1 U15707 ( .A1(n13682), .A2(n14098), .B1(n13681), .B2(n13903), .ZN(
        n14067) );
  NAND2_X1 U15708 ( .A1(n14472), .A2(n14067), .ZN(n13684) );
  OAI211_X1 U15709 ( .C1(n14479), .C2(n14072), .A(n13684), .B(n13683), .ZN(
        n13685) );
  AOI21_X1 U15710 ( .B1(n14187), .B2(n14475), .A(n13685), .ZN(n13686) );
  OAI21_X1 U15711 ( .B1(n13687), .B2(n13705), .A(n13686), .ZN(P1_U3238) );
  OAI211_X1 U15712 ( .C1(n13690), .C2(n13689), .A(n13688), .B(n14470), .ZN(
        n13697) );
  NAND2_X1 U15713 ( .A1(n13730), .A2(n14100), .ZN(n13693) );
  NAND2_X1 U15714 ( .A1(n13728), .A2(n13691), .ZN(n13692) );
  NAND2_X1 U15715 ( .A1(n13693), .A2(n13692), .ZN(n14570) );
  AND2_X1 U15716 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n13802) );
  AOI21_X1 U15717 ( .B1(n14472), .B2(n14570), .A(n13802), .ZN(n13696) );
  NAND2_X1 U15718 ( .A1(n14475), .A2(n14651), .ZN(n13695) );
  OR2_X1 U15719 ( .A1(n14479), .A2(n14572), .ZN(n13694) );
  NAND4_X1 U15720 ( .A1(n13697), .A2(n13696), .A3(n13695), .A4(n13694), .ZN(
        P1_U3239) );
  XOR2_X1 U15721 ( .A(n13699), .B(n13698), .Z(n13706) );
  AND2_X1 U15722 ( .A1(n13894), .A2(n14100), .ZN(n13700) );
  AOI21_X1 U15723 ( .B1(n13896), .B2(n13854), .A(n13700), .ZN(n14139) );
  INV_X1 U15724 ( .A(n13949), .ZN(n13701) );
  AOI22_X1 U15725 ( .A1(n13701), .A2(n13714), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13702) );
  OAI21_X1 U15726 ( .B1(n14139), .B2(n13712), .A(n13702), .ZN(n13703) );
  AOI21_X1 U15727 ( .B1(n14142), .B2(n14475), .A(n13703), .ZN(n13704) );
  OAI21_X1 U15728 ( .B1(n13706), .B2(n13705), .A(n13704), .ZN(P1_U3240) );
  OAI211_X1 U15729 ( .C1(n13710), .C2(n13709), .A(n13708), .B(n14470), .ZN(
        n13717) );
  INV_X1 U15730 ( .A(n13711), .ZN(n13715) );
  NAND2_X1 U15731 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14542)
         );
  OAI21_X1 U15732 ( .B1(n13712), .B2(n14201), .A(n14542), .ZN(n13713) );
  AOI21_X1 U15733 ( .B1(n13715), .B2(n13714), .A(n13713), .ZN(n13716) );
  OAI211_X1 U15734 ( .C1(n14202), .C2(n13718), .A(n13717), .B(n13716), .ZN(
        P1_U3241) );
  MUX2_X1 U15735 ( .A(n13855), .B(P1_DATAO_REG_31__SCAN_IN), .S(n13732), .Z(
        P1_U3591) );
  MUX2_X1 U15736 ( .A(n13905), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13732), .Z(
        P1_U3590) );
  MUX2_X1 U15737 ( .A(n13719), .B(P1_DATAO_REG_29__SCAN_IN), .S(n13732), .Z(
        P1_U3589) );
  MUX2_X1 U15738 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13897), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15739 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13896), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15740 ( .A(n13720), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13732), .Z(
        P1_U3586) );
  MUX2_X1 U15741 ( .A(n13894), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13732), .Z(
        P1_U3585) );
  MUX2_X1 U15742 ( .A(n13893), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13732), .Z(
        P1_U3584) );
  MUX2_X1 U15743 ( .A(n13876), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13732), .Z(
        P1_U3583) );
  MUX2_X1 U15744 ( .A(n13891), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13732), .Z(
        P1_U3582) );
  MUX2_X1 U15745 ( .A(n13874), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13732), .Z(
        P1_U3581) );
  MUX2_X1 U15746 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13888), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15747 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13887), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15748 ( .A(n13886), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13732), .Z(
        P1_U3578) );
  MUX2_X1 U15749 ( .A(n13884), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13732), .Z(
        P1_U3577) );
  MUX2_X1 U15750 ( .A(n13880), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13732), .Z(
        P1_U3576) );
  MUX2_X1 U15751 ( .A(n13721), .B(P1_DATAO_REG_15__SCAN_IN), .S(n13732), .Z(
        P1_U3575) );
  MUX2_X1 U15752 ( .A(n13722), .B(P1_DATAO_REG_14__SCAN_IN), .S(n13732), .Z(
        P1_U3574) );
  MUX2_X1 U15753 ( .A(n14101), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13732), .Z(
        P1_U3573) );
  MUX2_X1 U15754 ( .A(n13723), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13732), .Z(
        P1_U3572) );
  MUX2_X1 U15755 ( .A(n13724), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13732), .Z(
        P1_U3571) );
  MUX2_X1 U15756 ( .A(n13725), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13732), .Z(
        P1_U3570) );
  MUX2_X1 U15757 ( .A(n13726), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13732), .Z(
        P1_U3569) );
  MUX2_X1 U15758 ( .A(n13727), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13732), .Z(
        P1_U3568) );
  MUX2_X1 U15759 ( .A(n13728), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13732), .Z(
        P1_U3567) );
  MUX2_X1 U15760 ( .A(n13729), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13732), .Z(
        P1_U3566) );
  MUX2_X1 U15761 ( .A(n13730), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13732), .Z(
        P1_U3565) );
  MUX2_X1 U15762 ( .A(n13731), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13732), .Z(
        P1_U3563) );
  MUX2_X1 U15763 ( .A(n13733), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13732), .Z(
        P1_U3562) );
  MUX2_X1 U15764 ( .A(n13734), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13732), .Z(
        P1_U3561) );
  INV_X1 U15765 ( .A(n13738), .ZN(n13737) );
  OAI22_X1 U15766 ( .A1(n14544), .A2(n8819), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13735), .ZN(n13736) );
  AOI21_X1 U15767 ( .B1(n13737), .B2(n14536), .A(n13736), .ZN(n13744) );
  MUX2_X1 U15768 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10016), .S(n13738), .Z(
        n13739) );
  OAI21_X1 U15769 ( .B1(n9722), .B2(n6927), .A(n13739), .ZN(n13740) );
  NAND3_X1 U15770 ( .A1(n13841), .A2(n13761), .A3(n13740), .ZN(n13743) );
  NAND2_X1 U15771 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13746) );
  OAI211_X1 U15772 ( .C1(n10045), .C2(n13741), .A(n13846), .B(n13756), .ZN(
        n13742) );
  NAND3_X1 U15773 ( .A1(n13744), .A2(n13743), .A3(n13742), .ZN(P1_U3244) );
  MUX2_X1 U15774 ( .A(n13747), .B(n13746), .S(n13745), .Z(n13750) );
  AOI21_X1 U15775 ( .B1(n6927), .B2(n13748), .A(n13732), .ZN(n13749) );
  OAI21_X1 U15776 ( .B1(n13750), .B2(n6415), .A(n13749), .ZN(n13799) );
  OAI22_X1 U15777 ( .A1(n14544), .A2(n13752), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13751), .ZN(n13753) );
  AOI21_X1 U15778 ( .B1(n13754), .B2(n14536), .A(n13753), .ZN(n13766) );
  MUX2_X1 U15779 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10043), .S(n13759), .Z(
        n13757) );
  NAND3_X1 U15780 ( .A1(n13757), .A2(n13756), .A3(n13755), .ZN(n13758) );
  NAND3_X1 U15781 ( .A1(n13846), .A2(n13773), .A3(n13758), .ZN(n13765) );
  MUX2_X1 U15782 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10015), .S(n13759), .Z(
        n13762) );
  NAND3_X1 U15783 ( .A1(n13762), .A2(n13761), .A3(n13760), .ZN(n13763) );
  NAND3_X1 U15784 ( .A1(n13841), .A2(n13768), .A3(n13763), .ZN(n13764) );
  NAND4_X1 U15785 ( .A1(n13799), .A2(n13766), .A3(n13765), .A4(n13764), .ZN(
        P1_U3245) );
  MUX2_X1 U15786 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10021), .S(n13771), .Z(
        n13769) );
  NAND3_X1 U15787 ( .A1(n13769), .A2(n13768), .A3(n13767), .ZN(n13770) );
  NAND3_X1 U15788 ( .A1(n13841), .A2(n13787), .A3(n13770), .ZN(n13781) );
  MUX2_X1 U15789 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10048), .S(n13771), .Z(
        n13774) );
  NAND3_X1 U15790 ( .A1(n13774), .A2(n13773), .A3(n13772), .ZN(n13775) );
  NAND3_X1 U15791 ( .A1(n13846), .A2(n13793), .A3(n13775), .ZN(n13780) );
  AOI22_X1 U15792 ( .A1(n13776), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n13779) );
  NAND2_X1 U15793 ( .A1(n14536), .A2(n13777), .ZN(n13778) );
  NAND4_X1 U15794 ( .A1(n13781), .A2(n13780), .A3(n13779), .A4(n13778), .ZN(
        P1_U3246) );
  INV_X1 U15795 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n13783) );
  OAI21_X1 U15796 ( .B1(n14544), .B2(n13783), .A(n13782), .ZN(n13784) );
  AOI21_X1 U15797 ( .B1(n13790), .B2(n14536), .A(n13784), .ZN(n13798) );
  MUX2_X1 U15798 ( .A(n10024), .B(P1_REG1_REG_4__SCAN_IN), .S(n13790), .Z(
        n13785) );
  NAND3_X1 U15799 ( .A1(n13787), .A2(n13786), .A3(n13785), .ZN(n13788) );
  NAND3_X1 U15800 ( .A1(n13841), .A2(n13789), .A3(n13788), .ZN(n13797) );
  MUX2_X1 U15801 ( .A(n11129), .B(P1_REG2_REG_4__SCAN_IN), .S(n13790), .Z(
        n13791) );
  NAND3_X1 U15802 ( .A1(n13793), .A2(n13792), .A3(n13791), .ZN(n13794) );
  NAND3_X1 U15803 ( .A1(n13846), .A2(n13795), .A3(n13794), .ZN(n13796) );
  NAND4_X1 U15804 ( .A1(n13799), .A2(n13798), .A3(n13797), .A4(n13796), .ZN(
        P1_U3247) );
  NOR2_X1 U15805 ( .A1(n14544), .A2(n13800), .ZN(n13801) );
  AOI211_X1 U15806 ( .C1(n14536), .C2(n13807), .A(n13802), .B(n13801), .ZN(
        n13815) );
  INV_X1 U15807 ( .A(n13803), .ZN(n13806) );
  MUX2_X1 U15808 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n14700), .S(n13807), .Z(
        n13805) );
  OAI211_X1 U15809 ( .C1(n13806), .C2(n13805), .A(n13841), .B(n13804), .ZN(
        n13814) );
  MUX2_X1 U15810 ( .A(n10817), .B(P1_REG2_REG_6__SCAN_IN), .S(n13807), .Z(
        n13808) );
  NAND3_X1 U15811 ( .A1(n13810), .A2(n13809), .A3(n13808), .ZN(n13811) );
  NAND3_X1 U15812 ( .A1(n13846), .A2(n13812), .A3(n13811), .ZN(n13813) );
  NAND3_X1 U15813 ( .A1(n13815), .A2(n13814), .A3(n13813), .ZN(P1_U3249) );
  OAI21_X1 U15814 ( .B1(n13818), .B2(n13817), .A(n13816), .ZN(n13819) );
  NAND2_X1 U15815 ( .A1(n13819), .A2(n13841), .ZN(n13831) );
  NAND2_X1 U15816 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14476)
         );
  OAI21_X1 U15817 ( .B1(n14544), .B2(n13820), .A(n14476), .ZN(n13821) );
  AOI21_X1 U15818 ( .B1(n13822), .B2(n14536), .A(n13821), .ZN(n13830) );
  INV_X1 U15819 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n13823) );
  MUX2_X1 U15820 ( .A(n13823), .B(P1_REG2_REG_11__SCAN_IN), .S(n13822), .Z(
        n13824) );
  NAND3_X1 U15821 ( .A1(n13826), .A2(n13825), .A3(n13824), .ZN(n13827) );
  NAND3_X1 U15822 ( .A1(n13846), .A2(n13828), .A3(n13827), .ZN(n13829) );
  NAND3_X1 U15823 ( .A1(n13831), .A2(n13830), .A3(n13829), .ZN(P1_U3254) );
  INV_X1 U15824 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13851) );
  NAND2_X1 U15825 ( .A1(n13837), .A2(n13832), .ZN(n13833) );
  NAND2_X1 U15826 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  XOR2_X1 U15827 ( .A(n13835), .B(P1_REG1_REG_19__SCAN_IN), .Z(n13843) );
  NAND2_X1 U15828 ( .A1(n13837), .A2(n13836), .ZN(n13839) );
  NAND2_X1 U15829 ( .A1(n13839), .A2(n13838), .ZN(n13840) );
  XOR2_X1 U15830 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13840), .Z(n13842) );
  AOI22_X1 U15831 ( .A1(n13843), .A2(n13841), .B1(n13846), .B2(n13842), .ZN(
        n13848) );
  INV_X1 U15832 ( .A(n13842), .ZN(n13845) );
  NOR2_X1 U15833 ( .A1(n13843), .A2(n14533), .ZN(n13844) );
  AOI211_X1 U15834 ( .C1(n13846), .C2(n13845), .A(n14536), .B(n13844), .ZN(
        n13847) );
  MUX2_X1 U15835 ( .A(n13848), .B(n13847), .S(n14559), .Z(n13850) );
  OAI211_X1 U15836 ( .C1(n13851), .C2(n14544), .A(n13850), .B(n13849), .ZN(
        P1_U3262) );
  NAND2_X1 U15837 ( .A1(n13935), .A2(n14130), .ZN(n13900) );
  XNOR2_X1 U15838 ( .A(n13860), .B(n13856), .ZN(n13852) );
  NAND2_X1 U15839 ( .A1(n13852), .A2(n14591), .ZN(n14117) );
  OR2_X1 U15840 ( .A1(n6394), .A2(n9761), .ZN(n13853) );
  AND2_X1 U15841 ( .A1(n13854), .A2(n13853), .ZN(n13906) );
  NAND2_X1 U15842 ( .A1(n13906), .A2(n13855), .ZN(n14119) );
  NOR2_X1 U15843 ( .A1(n14599), .A2(n14119), .ZN(n13863) );
  AOI21_X1 U15844 ( .B1(n14599), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13863), 
        .ZN(n13858) );
  NAND2_X1 U15845 ( .A1(n13856), .A2(n14585), .ZN(n13857) );
  OAI211_X1 U15846 ( .C1(n14117), .C2(n14109), .A(n13858), .B(n13857), .ZN(
        P1_U3263) );
  INV_X1 U15847 ( .A(n13860), .ZN(n13861) );
  NOR2_X1 U15848 ( .A1(n14121), .A2(n14088), .ZN(n13862) );
  AOI211_X1 U15849 ( .C1(n14599), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13863), 
        .B(n13862), .ZN(n13864) );
  OAI21_X1 U15850 ( .B1(n14109), .B2(n14120), .A(n13864), .ZN(P1_U3264) );
  OR2_X1 U15851 ( .A1(n14197), .A2(n13880), .ZN(n13866) );
  INV_X1 U15852 ( .A(n13867), .ZN(n13868) );
  AND2_X1 U15853 ( .A1(n14187), .A2(n13886), .ZN(n13871) );
  OR2_X1 U15854 ( .A1(n14187), .A2(n13886), .ZN(n13870) );
  NOR2_X1 U15855 ( .A1(n14060), .A2(n13887), .ZN(n13872) );
  INV_X1 U15856 ( .A(n14159), .ZN(n13995) );
  INV_X1 U15857 ( .A(n13876), .ZN(n13892) );
  NAND2_X1 U15858 ( .A1(n13995), .A2(n13892), .ZN(n13877) );
  INV_X1 U15859 ( .A(n13973), .ZN(n13979) );
  INV_X1 U15860 ( .A(n14142), .ZN(n13953) );
  INV_X1 U15861 ( .A(n13931), .ZN(n13942) );
  NAND2_X1 U15862 ( .A1(n13921), .A2(n13920), .ZN(n13919) );
  NAND2_X1 U15863 ( .A1(n14051), .A2(n14050), .ZN(n14049) );
  OAI21_X1 U15864 ( .B1(n13891), .B2(n14007), .A(n14008), .ZN(n13989) );
  INV_X1 U15865 ( .A(n13898), .ZN(n13899) );
  NAND2_X1 U15866 ( .A1(n14122), .A2(n14063), .ZN(n13917) );
  AOI21_X1 U15867 ( .B1(n13900), .B2(n14126), .A(n14575), .ZN(n13902) );
  OR2_X1 U15868 ( .A1(n13904), .A2(n13903), .ZN(n14124) );
  NAND2_X1 U15869 ( .A1(n14126), .A2(n14585), .ZN(n13914) );
  NAND2_X1 U15870 ( .A1(n14586), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13908) );
  NAND2_X1 U15871 ( .A1(n13906), .A2(n13905), .ZN(n14123) );
  OAI22_X1 U15872 ( .A1(n13909), .A2(n13908), .B1(n14123), .B2(n13907), .ZN(
        n13912) );
  INV_X1 U15873 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n13910) );
  NOR2_X1 U15874 ( .A1(n14562), .A2(n13910), .ZN(n13911) );
  NOR2_X1 U15875 ( .A1(n13912), .A2(n13911), .ZN(n13913) );
  OAI211_X1 U15876 ( .C1(n14599), .C2(n14124), .A(n13914), .B(n13913), .ZN(
        n13915) );
  AOI21_X1 U15877 ( .B1(n14125), .B2(n14595), .A(n13915), .ZN(n13916) );
  OAI211_X1 U15878 ( .C1(n14127), .C2(n14092), .A(n13917), .B(n13916), .ZN(
        P1_U3356) );
  XNOR2_X1 U15879 ( .A(n13918), .B(n13920), .ZN(n14133) );
  OAI21_X1 U15880 ( .B1(n13921), .B2(n13920), .A(n13919), .ZN(n13922) );
  INV_X1 U15881 ( .A(n13922), .ZN(n14132) );
  OAI211_X1 U15882 ( .C1(n13935), .C2(n14130), .A(n14591), .B(n13900), .ZN(
        n14129) );
  AOI22_X1 U15883 ( .A1(n13923), .A2(n14586), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n14599), .ZN(n13924) );
  OAI21_X1 U15884 ( .B1(n14128), .B2(n14599), .A(n13924), .ZN(n13925) );
  AOI21_X1 U15885 ( .B1(n13926), .B2(n14585), .A(n13925), .ZN(n13927) );
  OAI21_X1 U15886 ( .B1(n14129), .B2(n14109), .A(n13927), .ZN(n13928) );
  AOI21_X1 U15887 ( .B1(n14132), .B2(n14596), .A(n13928), .ZN(n13929) );
  OAI21_X1 U15888 ( .B1(n14133), .B2(n13930), .A(n13929), .ZN(P1_U3265) );
  XNOR2_X1 U15889 ( .A(n13932), .B(n13931), .ZN(n13934) );
  INV_X1 U15890 ( .A(n13951), .ZN(n13936) );
  AOI211_X1 U15891 ( .C1(n6701), .C2(n13936), .A(n14575), .B(n13935), .ZN(
        n14134) );
  AOI22_X1 U15892 ( .A1(n13937), .A2(n14586), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n14599), .ZN(n13938) );
  OAI21_X1 U15893 ( .B1(n13939), .B2(n14088), .A(n13938), .ZN(n13944) );
  AOI21_X1 U15894 ( .B1(n13942), .B2(n13941), .A(n13940), .ZN(n14138) );
  NOR2_X1 U15895 ( .A1(n14138), .A2(n14092), .ZN(n13943) );
  AOI211_X1 U15896 ( .C1(n14134), .C2(n14595), .A(n13944), .B(n13943), .ZN(
        n13945) );
  OAI21_X1 U15897 ( .B1(n14137), .B2(n14599), .A(n13945), .ZN(P1_U3266) );
  XNOR2_X1 U15898 ( .A(n6530), .B(n13946), .ZN(n14145) );
  XNOR2_X1 U15899 ( .A(n13947), .B(n13946), .ZN(n13948) );
  NAND2_X1 U15900 ( .A1(n13948), .A2(n14625), .ZN(n14144) );
  OAI211_X1 U15901 ( .C1(n14555), .C2(n13949), .A(n14144), .B(n14139), .ZN(
        n13950) );
  NAND2_X1 U15902 ( .A1(n13950), .A2(n14562), .ZN(n13956) );
  AOI211_X1 U15903 ( .C1(n14142), .C2(n13963), .A(n14575), .B(n13951), .ZN(
        n14140) );
  INV_X1 U15904 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13952) );
  OAI22_X1 U15905 ( .A1(n13953), .A2(n14088), .B1(n14562), .B2(n13952), .ZN(
        n13954) );
  AOI21_X1 U15906 ( .B1(n14140), .B2(n14595), .A(n13954), .ZN(n13955) );
  OAI211_X1 U15907 ( .C1(n14145), .C2(n14092), .A(n13956), .B(n13955), .ZN(
        P1_U3267) );
  AOI21_X1 U15908 ( .B1(n13961), .B2(n13958), .A(n13957), .ZN(n13959) );
  INV_X1 U15909 ( .A(n13959), .ZN(n14151) );
  OAI21_X1 U15910 ( .B1(n13962), .B2(n13961), .A(n13960), .ZN(n14149) );
  AOI21_X1 U15911 ( .B1(n13981), .B2(n13969), .A(n14575), .ZN(n13964) );
  NAND2_X1 U15912 ( .A1(n13964), .A2(n13963), .ZN(n14147) );
  NAND2_X1 U15913 ( .A1(n13965), .A2(n14586), .ZN(n13966) );
  NAND2_X1 U15914 ( .A1(n14146), .A2(n13966), .ZN(n13967) );
  MUX2_X1 U15915 ( .A(P1_REG2_REG_25__SCAN_IN), .B(n13967), .S(n14562), .Z(
        n13968) );
  AOI21_X1 U15916 ( .B1(n13969), .B2(n14585), .A(n13968), .ZN(n13970) );
  OAI21_X1 U15917 ( .B1(n14147), .B2(n14109), .A(n13970), .ZN(n13971) );
  AOI21_X1 U15918 ( .B1(n14149), .B2(n14063), .A(n13971), .ZN(n13972) );
  OAI21_X1 U15919 ( .B1(n14092), .B2(n14151), .A(n13972), .ZN(P1_U3268) );
  OAI21_X1 U15920 ( .B1(n13974), .B2(n13973), .A(n14625), .ZN(n13977) );
  OAI21_X1 U15921 ( .B1(n13977), .B2(n13976), .A(n13975), .ZN(n14154) );
  INV_X1 U15922 ( .A(n14154), .ZN(n13988) );
  OAI21_X1 U15923 ( .B1(n13980), .B2(n13979), .A(n13978), .ZN(n14156) );
  OAI211_X1 U15924 ( .C1(n14153), .C2(n6423), .A(n14591), .B(n13981), .ZN(
        n14152) );
  AOI22_X1 U15925 ( .A1(n13982), .A2(n14586), .B1(n14599), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n13985) );
  NAND2_X1 U15926 ( .A1(n13983), .A2(n14585), .ZN(n13984) );
  OAI211_X1 U15927 ( .C1(n14152), .C2(n14109), .A(n13985), .B(n13984), .ZN(
        n13986) );
  AOI21_X1 U15928 ( .B1(n14156), .B2(n14596), .A(n13986), .ZN(n13987) );
  OAI21_X1 U15929 ( .B1(n13988), .B2(n14599), .A(n13987), .ZN(P1_U3269) );
  XNOR2_X1 U15930 ( .A(n13989), .B(n13997), .ZN(n13991) );
  AOI21_X1 U15931 ( .B1(n13991), .B2(n14625), .A(n13990), .ZN(n14161) );
  AOI211_X1 U15932 ( .C1(n14159), .C2(n14002), .A(n14575), .B(n6423), .ZN(
        n14158) );
  INV_X1 U15933 ( .A(n13992), .ZN(n13993) );
  AOI22_X1 U15934 ( .A1(n14599), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n13993), 
        .B2(n14586), .ZN(n13994) );
  OAI21_X1 U15935 ( .B1(n13995), .B2(n14088), .A(n13994), .ZN(n13999) );
  XOR2_X1 U15936 ( .A(n13996), .B(n13997), .Z(n14162) );
  NOR2_X1 U15937 ( .A1(n14162), .A2(n14092), .ZN(n13998) );
  AOI211_X1 U15938 ( .C1(n14158), .C2(n14595), .A(n13999), .B(n13998), .ZN(
        n14000) );
  OAI21_X1 U15939 ( .B1(n14161), .B2(n14599), .A(n14000), .ZN(P1_U3270) );
  XNOR2_X1 U15940 ( .A(n14001), .B(n14010), .ZN(n14166) );
  INV_X1 U15941 ( .A(n14022), .ZN(n14004) );
  INV_X1 U15942 ( .A(n14002), .ZN(n14003) );
  AOI211_X1 U15943 ( .C1(n6934), .C2(n14004), .A(n14575), .B(n14003), .ZN(
        n14163) );
  AOI22_X1 U15944 ( .A1(n14599), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14005), 
        .B2(n14586), .ZN(n14006) );
  OAI21_X1 U15945 ( .B1(n14007), .B2(n14088), .A(n14006), .ZN(n14015) );
  OAI21_X1 U15946 ( .B1(n14010), .B2(n14009), .A(n14008), .ZN(n14013) );
  INV_X1 U15947 ( .A(n14011), .ZN(n14012) );
  AOI21_X1 U15948 ( .B1(n14013), .B2(n14625), .A(n14012), .ZN(n14165) );
  NOR2_X1 U15949 ( .A1(n14165), .A2(n14599), .ZN(n14014) );
  AOI211_X1 U15950 ( .C1(n14163), .C2(n14595), .A(n14015), .B(n14014), .ZN(
        n14016) );
  OAI21_X1 U15951 ( .B1(n14166), .B2(n14092), .A(n14016), .ZN(P1_U3271) );
  OAI21_X1 U15952 ( .B1(n14018), .B2(n14021), .A(n14017), .ZN(n14019) );
  INV_X1 U15953 ( .A(n14019), .ZN(n14173) );
  AOI21_X1 U15954 ( .B1(n6535), .B2(n14021), .A(n14020), .ZN(n14167) );
  NAND2_X1 U15955 ( .A1(n14167), .A2(n14063), .ZN(n14031) );
  AOI211_X1 U15956 ( .C1(n14170), .C2(n14023), .A(n14575), .B(n14022), .ZN(
        n14168) );
  INV_X1 U15957 ( .A(n14169), .ZN(n14025) );
  OAI22_X1 U15958 ( .A1(n14025), .A2(n14599), .B1(n14024), .B2(n14555), .ZN(
        n14026) );
  AOI21_X1 U15959 ( .B1(P1_REG2_REG_21__SCAN_IN), .B2(n14599), .A(n14026), 
        .ZN(n14027) );
  OAI21_X1 U15960 ( .B1(n14028), .B2(n14088), .A(n14027), .ZN(n14029) );
  AOI21_X1 U15961 ( .B1(n14168), .B2(n14595), .A(n14029), .ZN(n14030) );
  OAI211_X1 U15962 ( .C1(n14173), .C2(n14092), .A(n14031), .B(n14030), .ZN(
        P1_U3272) );
  AOI211_X1 U15963 ( .C1(n14041), .C2(n14033), .A(n14635), .B(n14032), .ZN(
        n14036) );
  INV_X1 U15964 ( .A(n14034), .ZN(n14035) );
  NOR2_X1 U15965 ( .A1(n14036), .A2(n14035), .ZN(n14177) );
  XNOR2_X1 U15966 ( .A(n14175), .B(n14052), .ZN(n14037) );
  NOR2_X1 U15967 ( .A1(n14037), .A2(n14575), .ZN(n14174) );
  AOI22_X1 U15968 ( .A1(n14599), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14038), 
        .B2(n14586), .ZN(n14039) );
  OAI21_X1 U15969 ( .B1(n14040), .B2(n14088), .A(n14039), .ZN(n14046) );
  NOR2_X1 U15970 ( .A1(n14042), .A2(n14041), .ZN(n14043) );
  OR2_X1 U15971 ( .A1(n14044), .A2(n14043), .ZN(n14178) );
  NOR2_X1 U15972 ( .A1(n14178), .A2(n14092), .ZN(n14045) );
  AOI211_X1 U15973 ( .C1(n14174), .C2(n14595), .A(n14046), .B(n14045), .ZN(
        n14047) );
  OAI21_X1 U15974 ( .B1(n14177), .B2(n14599), .A(n14047), .ZN(P1_U3273) );
  XNOR2_X1 U15975 ( .A(n14048), .B(n14050), .ZN(n14185) );
  OAI21_X1 U15976 ( .B1(n14051), .B2(n14050), .A(n14049), .ZN(n14183) );
  AOI21_X1 U15977 ( .B1(n14060), .B2(n14069), .A(n14575), .ZN(n14053) );
  NAND2_X1 U15978 ( .A1(n14053), .A2(n14052), .ZN(n14180) );
  INV_X1 U15979 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14058) );
  INV_X1 U15980 ( .A(n14179), .ZN(n14054) );
  NAND2_X1 U15981 ( .A1(n14054), .A2(n14562), .ZN(n14057) );
  NAND2_X1 U15982 ( .A1(n14055), .A2(n14586), .ZN(n14056) );
  OAI211_X1 U15983 ( .C1(n14562), .C2(n14058), .A(n14057), .B(n14056), .ZN(
        n14059) );
  AOI21_X1 U15984 ( .B1(n14060), .B2(n14585), .A(n14059), .ZN(n14061) );
  OAI21_X1 U15985 ( .B1(n14180), .B2(n14109), .A(n14061), .ZN(n14062) );
  AOI21_X1 U15986 ( .B1(n14183), .B2(n14063), .A(n14062), .ZN(n14064) );
  OAI21_X1 U15987 ( .B1(n14092), .B2(n14185), .A(n14064), .ZN(P1_U3274) );
  AOI211_X1 U15988 ( .C1(n14075), .C2(n14066), .A(n14635), .B(n14065), .ZN(
        n14068) );
  NOR2_X1 U15989 ( .A1(n14068), .A2(n14067), .ZN(n14189) );
  INV_X1 U15990 ( .A(n14069), .ZN(n14070) );
  AOI211_X1 U15991 ( .C1(n14187), .C2(n14071), .A(n14575), .B(n14070), .ZN(
        n14186) );
  INV_X1 U15992 ( .A(n14072), .ZN(n14073) );
  AOI22_X1 U15993 ( .A1(n14599), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14073), 
        .B2(n14586), .ZN(n14074) );
  OAI21_X1 U15994 ( .B1(n6936), .B2(n14088), .A(n14074), .ZN(n14078) );
  XNOR2_X1 U15995 ( .A(n14076), .B(n14075), .ZN(n14190) );
  NOR2_X1 U15996 ( .A1(n14190), .A2(n14092), .ZN(n14077) );
  AOI211_X1 U15997 ( .C1(n14186), .C2(n14595), .A(n14078), .B(n14077), .ZN(
        n14079) );
  OAI21_X1 U15998 ( .B1(n14189), .B2(n14599), .A(n14079), .ZN(P1_U3275) );
  AOI211_X1 U15999 ( .C1(n14090), .C2(n14080), .A(n14635), .B(n6562), .ZN(
        n14083) );
  INV_X1 U16000 ( .A(n14081), .ZN(n14082) );
  NOR2_X1 U16001 ( .A1(n14083), .A2(n14082), .ZN(n14194) );
  XNOR2_X1 U16002 ( .A(n14084), .B(n14192), .ZN(n14085) );
  NOR2_X1 U16003 ( .A1(n14085), .A2(n14575), .ZN(n14191) );
  AOI22_X1 U16004 ( .A1(n14599), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14086), 
        .B2(n14586), .ZN(n14087) );
  OAI21_X1 U16005 ( .B1(n14089), .B2(n14088), .A(n14087), .ZN(n14094) );
  XOR2_X1 U16006 ( .A(n14091), .B(n14090), .Z(n14195) );
  NOR2_X1 U16007 ( .A1(n14195), .A2(n14092), .ZN(n14093) );
  AOI211_X1 U16008 ( .C1(n14191), .C2(n14595), .A(n14094), .B(n14093), .ZN(
        n14095) );
  OAI21_X1 U16009 ( .B1(n14194), .B2(n14599), .A(n14095), .ZN(P1_U3276) );
  OAI211_X1 U16010 ( .C1(n14097), .C2(n14112), .A(n14096), .B(n14625), .ZN(
        n14487) );
  INV_X1 U16011 ( .A(n14487), .ZN(n14104) );
  OR2_X1 U16012 ( .A1(n14099), .A2(n14098), .ZN(n14103) );
  NAND2_X1 U16013 ( .A1(n14101), .A2(n14100), .ZN(n14102) );
  NAND2_X1 U16014 ( .A1(n14103), .A2(n14102), .ZN(n14480) );
  OAI21_X1 U16015 ( .B1(n14104), .B2(n14480), .A(n14562), .ZN(n14116) );
  OAI22_X1 U16016 ( .A1(n14562), .A2(n14105), .B1(n14466), .B2(n14555), .ZN(
        n14111) );
  AOI21_X1 U16017 ( .B1(n14481), .B2(n14106), .A(n14575), .ZN(n14108) );
  NAND2_X1 U16018 ( .A1(n14108), .A2(n14107), .ZN(n14485) );
  NOR2_X1 U16019 ( .A1(n14485), .A2(n14109), .ZN(n14110) );
  AOI211_X1 U16020 ( .C1(n14585), .C2(n14481), .A(n14111), .B(n14110), .ZN(
        n14115) );
  NAND2_X1 U16021 ( .A1(n14113), .A2(n14112), .ZN(n14482) );
  NAND3_X1 U16022 ( .A1(n14483), .A2(n14482), .A3(n14596), .ZN(n14114) );
  NAND3_X1 U16023 ( .A1(n14116), .A2(n14115), .A3(n14114), .ZN(P1_U3279) );
  OAI211_X1 U16024 ( .C1(n14118), .C2(n14686), .A(n14117), .B(n14119), .ZN(
        n14208) );
  MUX2_X1 U16025 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14208), .S(n14709), .Z(
        P1_U3559) );
  MUX2_X1 U16026 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14209), .S(n14709), .Z(
        P1_U3558) );
  MUX2_X1 U16027 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14210), .S(n14709), .Z(
        P1_U3557) );
  OAI211_X1 U16028 ( .C1(n14130), .C2(n14686), .A(n14129), .B(n14128), .ZN(
        n14131) );
  MUX2_X1 U16029 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14211), .S(n14709), .Z(
        P1_U3556) );
  AOI21_X1 U16030 ( .B1(n14652), .B2(n6701), .A(n14134), .ZN(n14136) );
  OAI211_X1 U16031 ( .C1(n14644), .C2(n14138), .A(n14137), .B(n14136), .ZN(
        n14212) );
  MUX2_X1 U16032 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14212), .S(n14709), .Z(
        P1_U3555) );
  INV_X1 U16033 ( .A(n14139), .ZN(n14141) );
  AOI211_X1 U16034 ( .C1(n14652), .C2(n14142), .A(n14141), .B(n14140), .ZN(
        n14143) );
  OAI211_X1 U16035 ( .C1(n14644), .C2(n14145), .A(n14144), .B(n14143), .ZN(
        n14213) );
  MUX2_X1 U16036 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14213), .S(n14709), .Z(
        P1_U3554) );
  OAI211_X1 U16037 ( .C1(n6930), .C2(n14686), .A(n14147), .B(n14146), .ZN(
        n14148) );
  AOI21_X1 U16038 ( .B1(n14149), .B2(n14625), .A(n14148), .ZN(n14150) );
  OAI21_X1 U16039 ( .B1(n14644), .B2(n14151), .A(n14150), .ZN(n14214) );
  MUX2_X1 U16040 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14214), .S(n14709), .Z(
        P1_U3553) );
  OAI21_X1 U16041 ( .B1(n14153), .B2(n14686), .A(n14152), .ZN(n14155) );
  AOI211_X1 U16042 ( .C1(n14683), .C2(n14156), .A(n14155), .B(n14154), .ZN(
        n14157) );
  INV_X1 U16043 ( .A(n14157), .ZN(n14215) );
  MUX2_X1 U16044 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14215), .S(n14709), .Z(
        P1_U3552) );
  AOI21_X1 U16045 ( .B1(n14652), .B2(n14159), .A(n14158), .ZN(n14160) );
  OAI211_X1 U16046 ( .C1(n14644), .C2(n14162), .A(n14161), .B(n14160), .ZN(
        n14216) );
  MUX2_X1 U16047 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14216), .S(n14709), .Z(
        P1_U3551) );
  AOI21_X1 U16048 ( .B1(n14652), .B2(n6934), .A(n14163), .ZN(n14164) );
  OAI211_X1 U16049 ( .C1(n14644), .C2(n14166), .A(n14165), .B(n14164), .ZN(
        n14217) );
  MUX2_X1 U16050 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14217), .S(n14709), .Z(
        P1_U3550) );
  NAND2_X1 U16051 ( .A1(n14167), .A2(n14625), .ZN(n14172) );
  AOI211_X1 U16052 ( .C1(n14652), .C2(n14170), .A(n14169), .B(n14168), .ZN(
        n14171) );
  OAI211_X1 U16053 ( .C1(n14644), .C2(n14173), .A(n14172), .B(n14171), .ZN(
        n14218) );
  MUX2_X1 U16054 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14218), .S(n14709), .Z(
        P1_U3549) );
  AOI21_X1 U16055 ( .B1(n14652), .B2(n14175), .A(n14174), .ZN(n14176) );
  OAI211_X1 U16056 ( .C1(n14644), .C2(n14178), .A(n14177), .B(n14176), .ZN(
        n14219) );
  MUX2_X1 U16057 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14219), .S(n14709), .Z(
        P1_U3548) );
  OAI211_X1 U16058 ( .C1(n14181), .C2(n14686), .A(n14180), .B(n14179), .ZN(
        n14182) );
  AOI21_X1 U16059 ( .B1(n14183), .B2(n14625), .A(n14182), .ZN(n14184) );
  OAI21_X1 U16060 ( .B1(n14644), .B2(n14185), .A(n14184), .ZN(n14220) );
  MUX2_X1 U16061 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14220), .S(n14709), .Z(
        P1_U3547) );
  AOI21_X1 U16062 ( .B1(n14652), .B2(n14187), .A(n14186), .ZN(n14188) );
  OAI211_X1 U16063 ( .C1(n14644), .C2(n14190), .A(n14189), .B(n14188), .ZN(
        n14221) );
  MUX2_X1 U16064 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14221), .S(n14709), .Z(
        P1_U3546) );
  AOI21_X1 U16065 ( .B1(n14652), .B2(n14192), .A(n14191), .ZN(n14193) );
  OAI211_X1 U16066 ( .C1(n14644), .C2(n14195), .A(n14194), .B(n14193), .ZN(
        n14222) );
  MUX2_X1 U16067 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14222), .S(n14709), .Z(
        P1_U3545) );
  AOI21_X1 U16068 ( .B1(n14652), .B2(n14197), .A(n14196), .ZN(n14198) );
  OAI211_X1 U16069 ( .C1(n14644), .C2(n14200), .A(n14199), .B(n14198), .ZN(
        n14223) );
  MUX2_X1 U16070 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14223), .S(n14709), .Z(
        P1_U3544) );
  OAI21_X1 U16071 ( .B1(n14202), .B2(n14686), .A(n14201), .ZN(n14203) );
  AOI211_X1 U16072 ( .C1(n14205), .C2(n14683), .A(n14204), .B(n14203), .ZN(
        n14206) );
  OAI21_X1 U16073 ( .B1(n14635), .B2(n14207), .A(n14206), .ZN(n14224) );
  MUX2_X1 U16074 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14224), .S(n14709), .Z(
        P1_U3543) );
  MUX2_X1 U16075 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14208), .S(n14693), .Z(
        P1_U3527) );
  MUX2_X1 U16076 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14209), .S(n14693), .Z(
        P1_U3526) );
  MUX2_X1 U16077 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14210), .S(n14693), .Z(
        P1_U3525) );
  MUX2_X1 U16078 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14211), .S(n14693), .Z(
        P1_U3524) );
  MUX2_X1 U16079 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14212), .S(n14693), .Z(
        P1_U3523) );
  MUX2_X1 U16080 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14213), .S(n14693), .Z(
        P1_U3522) );
  MUX2_X1 U16081 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14214), .S(n14693), .Z(
        P1_U3521) );
  MUX2_X1 U16082 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14215), .S(n14693), .Z(
        P1_U3520) );
  MUX2_X1 U16083 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14216), .S(n14693), .Z(
        P1_U3519) );
  MUX2_X1 U16084 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14217), .S(n14693), .Z(
        P1_U3518) );
  MUX2_X1 U16085 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14218), .S(n14693), .Z(
        P1_U3517) );
  MUX2_X1 U16086 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14219), .S(n14693), .Z(
        P1_U3516) );
  MUX2_X1 U16087 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14220), .S(n14693), .Z(
        P1_U3515) );
  MUX2_X1 U16088 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14221), .S(n14693), .Z(
        P1_U3513) );
  MUX2_X1 U16089 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14222), .S(n14693), .Z(
        P1_U3510) );
  MUX2_X1 U16090 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14223), .S(n14693), .Z(
        P1_U3507) );
  MUX2_X1 U16091 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14224), .S(n14693), .Z(
        P1_U3504) );
  NAND2_X1 U16092 ( .A1(n14226), .A2(n14225), .ZN(n14230) );
  NAND2_X1 U16093 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n14227) );
  OR3_X1 U16094 ( .A1(n14228), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14227), .ZN(
        n14229) );
  OAI211_X1 U16095 ( .C1(n14231), .C2(n14245), .A(n14230), .B(n14229), .ZN(
        P1_U3324) );
  OAI222_X1 U16096 ( .A1(n14244), .A2(n14234), .B1(n14233), .B2(P1_U3086), 
        .C1(n14232), .C2(n14245), .ZN(P1_U3325) );
  INV_X1 U16097 ( .A(n14235), .ZN(n14237) );
  OAI222_X1 U16098 ( .A1(n14244), .A2(n14237), .B1(n6415), .B2(P1_U3086), .C1(
        n14236), .C2(n14245), .ZN(P1_U3327) );
  OAI222_X1 U16099 ( .A1(n14245), .A2(n7103), .B1(n14244), .B2(n14239), .C1(
        P1_U3086), .C2(n6394), .ZN(P1_U3328) );
  OAI222_X1 U16100 ( .A1(n14244), .A2(n14241), .B1(n14240), .B2(P1_U3086), 
        .C1(n6709), .C2(n14245), .ZN(P1_U3329) );
  OAI222_X1 U16101 ( .A1(n14245), .A2(n6685), .B1(n14244), .B2(n14243), .C1(
        P1_U3086), .C2(n14242), .ZN(P1_U3330) );
  INV_X1 U16102 ( .A(n9760), .ZN(n14248) );
  OAI222_X1 U16103 ( .A1(n14244), .A2(n14249), .B1(n14248), .B2(P1_U3086), 
        .C1(n14246), .C2(n14245), .ZN(P1_U3331) );
  MUX2_X1 U16104 ( .A(n14251), .B(n14250), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16105 ( .A(n14252), .ZN(n14253) );
  MUX2_X1 U16106 ( .A(n14253), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16107 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14828) );
  XOR2_X1 U16108 ( .A(n14828), .B(n14254), .Z(SUB_1596_U62) );
  AOI21_X1 U16109 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14255) );
  OAI21_X1 U16110 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14255), 
        .ZN(U28) );
  INV_X1 U16111 ( .A(P1_RD_REG_SCAN_IN), .ZN(n14257) );
  OAI221_X1 U16112 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7423), .C2(n14257), .A(n14256), .ZN(U29) );
  AOI21_X1 U16113 ( .B1(n14260), .B2(n14259), .A(n14258), .ZN(n14261) );
  XOR2_X1 U16114 ( .A(n14261), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  INV_X1 U16115 ( .A(n14262), .ZN(n14263) );
  AOI22_X1 U16116 ( .A1(n14263), .A2(n14288), .B1(SI_9_), .B2(n14287), .ZN(
        n14264) );
  OAI21_X1 U16117 ( .B1(P3_U3151), .B2(n14896), .A(n14264), .ZN(P3_U3286) );
  INV_X1 U16118 ( .A(SI_10_), .ZN(n14265) );
  OAI22_X1 U16119 ( .A1(n14266), .A2(n14277), .B1(n14265), .B2(n14275), .ZN(
        n14267) );
  INV_X1 U16120 ( .A(n14267), .ZN(n14268) );
  OAI21_X1 U16121 ( .B1(P3_U3151), .B2(n14914), .A(n14268), .ZN(P3_U3285) );
  AOI22_X1 U16122 ( .A1(n14269), .A2(n14288), .B1(SI_11_), .B2(n14287), .ZN(
        n14270) );
  OAI21_X1 U16123 ( .B1(P3_U3151), .B2(n14931), .A(n14270), .ZN(P3_U3284) );
  OAI22_X1 U16124 ( .A1(n14272), .A2(n14277), .B1(n14271), .B2(n14275), .ZN(
        n14273) );
  INV_X1 U16125 ( .A(n14273), .ZN(n14274) );
  OAI21_X1 U16126 ( .B1(P3_U3151), .B2(n14949), .A(n14274), .ZN(P3_U3283) );
  OAI22_X1 U16127 ( .A1(n14278), .A2(n14277), .B1(n14276), .B2(n14275), .ZN(
        n14279) );
  INV_X1 U16128 ( .A(n14279), .ZN(n14280) );
  OAI21_X1 U16129 ( .B1(P3_U3151), .B2(n14967), .A(n14280), .ZN(P3_U3282) );
  XOR2_X1 U16130 ( .A(n14282), .B(n14281), .Z(SUB_1596_U57) );
  AOI22_X1 U16131 ( .A1(n14283), .A2(n14288), .B1(SI_14_), .B2(n14287), .ZN(
        n14284) );
  OAI21_X1 U16132 ( .B1(P3_U3151), .B2(n14986), .A(n14284), .ZN(P3_U3281) );
  AOI22_X1 U16133 ( .A1(n14285), .A2(n14288), .B1(SI_15_), .B2(n14287), .ZN(
        n14286) );
  OAI21_X1 U16134 ( .B1(P3_U3151), .B2(n14331), .A(n14286), .ZN(P3_U3280) );
  AOI22_X1 U16135 ( .A1(n14289), .A2(n14288), .B1(SI_16_), .B2(n14287), .ZN(
        n14290) );
  OAI21_X1 U16136 ( .B1(P3_U3151), .B2(n14349), .A(n14290), .ZN(P3_U3279) );
  XOR2_X1 U16137 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14291), .Z(SUB_1596_U55) );
  INV_X1 U16138 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14731) );
  XOR2_X1 U16139 ( .A(n14731), .B(n14292), .Z(SUB_1596_U54) );
  AOI21_X1 U16140 ( .B1(n14295), .B2(n14294), .A(n14293), .ZN(n14296) );
  XOR2_X1 U16141 ( .A(n14296), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  XNOR2_X1 U16142 ( .A(n14297), .B(n14299), .ZN(n14305) );
  OAI211_X1 U16143 ( .C1(n14300), .C2(n14299), .A(n14298), .B(n14625), .ZN(
        n14301) );
  OAI211_X1 U16144 ( .C1(n14305), .C2(n14568), .A(n14302), .B(n14301), .ZN(
        n14315) );
  INV_X1 U16145 ( .A(n14315), .ZN(n14312) );
  AOI222_X1 U16146 ( .A1(n14304), .A2(n14585), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14599), .C1(n14303), .C2(n14586), .ZN(n14311) );
  INV_X1 U16147 ( .A(n14305), .ZN(n14317) );
  INV_X1 U16148 ( .A(n14306), .ZN(n14308) );
  OAI211_X1 U16149 ( .C1(n14308), .C2(n14314), .A(n14591), .B(n14307), .ZN(
        n14313) );
  INV_X1 U16150 ( .A(n14313), .ZN(n14309) );
  AOI22_X1 U16151 ( .A1(n14317), .A2(n14577), .B1(n14595), .B2(n14309), .ZN(
        n14310) );
  OAI211_X1 U16152 ( .C1(n14599), .C2(n14312), .A(n14311), .B(n14310), .ZN(
        P1_U3281) );
  INV_X1 U16153 ( .A(n14656), .ZN(n14674) );
  OAI21_X1 U16154 ( .B1(n14314), .B2(n14686), .A(n14313), .ZN(n14316) );
  AOI211_X1 U16155 ( .C1(n14674), .C2(n14317), .A(n14316), .B(n14315), .ZN(
        n14319) );
  INV_X1 U16156 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U16157 ( .A1(n14693), .A2(n14319), .B1(n14318), .B2(n14691), .ZN(
        P1_U3495) );
  AOI22_X1 U16158 ( .A1(n14709), .A2(n14319), .B1(n11186), .B2(n14706), .ZN(
        P1_U3540) );
  AOI21_X1 U16159 ( .B1(n14322), .B2(n14321), .A(n14320), .ZN(n14323) );
  XOR2_X1 U16160 ( .A(n14323), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  AOI21_X1 U16161 ( .B1(n14326), .B2(n14325), .A(n14324), .ZN(n14340) );
  OAI21_X1 U16162 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14328), .A(n14327), 
        .ZN(n14333) );
  AOI21_X1 U16163 ( .B1(n14984), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n14329), 
        .ZN(n14330) );
  OAI21_X1 U16164 ( .B1(n14987), .B2(n14331), .A(n14330), .ZN(n14332) );
  AOI21_X1 U16165 ( .B1(n14333), .B2(n14989), .A(n14332), .ZN(n14339) );
  AOI21_X1 U16166 ( .B1(n14336), .B2(n14335), .A(n14334), .ZN(n14337) );
  OR2_X1 U16167 ( .A1(n14337), .A2(n14952), .ZN(n14338) );
  OAI211_X1 U16168 ( .C1(n14340), .C2(n14997), .A(n14339), .B(n14338), .ZN(
        P3_U3197) );
  AOI21_X1 U16169 ( .B1(n14343), .B2(n14342), .A(n14341), .ZN(n14360) );
  OAI21_X1 U16170 ( .B1(n14346), .B2(n14345), .A(n14344), .ZN(n14351) );
  AOI21_X1 U16171 ( .B1(n14984), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n14347), 
        .ZN(n14348) );
  OAI21_X1 U16172 ( .B1(n14987), .B2(n14349), .A(n14348), .ZN(n14350) );
  AOI21_X1 U16173 ( .B1(n14351), .B2(n14989), .A(n14350), .ZN(n14359) );
  INV_X1 U16174 ( .A(n14352), .ZN(n14353) );
  NOR2_X1 U16175 ( .A1(n14354), .A2(n14353), .ZN(n14356) );
  NAND2_X1 U16176 ( .A1(n14357), .A2(n14356), .ZN(n14355) );
  OAI211_X1 U16177 ( .C1(n14357), .C2(n14356), .A(n14991), .B(n14355), .ZN(
        n14358) );
  OAI211_X1 U16178 ( .C1(n14360), .C2(n14997), .A(n14359), .B(n14358), .ZN(
        P3_U3198) );
  AOI22_X1 U16179 ( .A1(n14865), .A2(n14361), .B1(n14984), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14375) );
  OAI21_X1 U16180 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14363), .A(n14362), 
        .ZN(n14368) );
  AOI211_X1 U16181 ( .C1(n14366), .C2(n14365), .A(n14364), .B(n14952), .ZN(
        n14367) );
  AOI21_X1 U16182 ( .B1(n14368), .B2(n14989), .A(n14367), .ZN(n14374) );
  NAND2_X1 U16183 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14373)
         );
  OAI221_X1 U16184 ( .B1(n14371), .B2(n14370), .C1(n14371), .C2(n14369), .A(
        n14385), .ZN(n14372) );
  NAND4_X1 U16185 ( .A1(n14375), .A2(n14374), .A3(n14373), .A4(n14372), .ZN(
        P3_U3199) );
  AOI22_X1 U16186 ( .A1(n14865), .A2(n14376), .B1(n14984), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14392) );
  OAI21_X1 U16187 ( .B1(n14379), .B2(n14378), .A(n14377), .ZN(n14384) );
  OAI21_X1 U16188 ( .B1(n14382), .B2(n14381), .A(n14380), .ZN(n14383) );
  AOI22_X1 U16189 ( .A1(n14384), .A2(n14989), .B1(n14991), .B2(n14383), .ZN(
        n14391) );
  OAI221_X1 U16190 ( .B1(n14388), .B2(n14387), .C1(n14388), .C2(n14386), .A(
        n14385), .ZN(n14389) );
  NAND4_X1 U16191 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        P3_U3200) );
  NOR2_X1 U16192 ( .A1(n14394), .A2(n14393), .ZN(n14409) );
  AOI21_X1 U16193 ( .B1(n14409), .B2(n15109), .A(n14395), .ZN(n14398) );
  AOI22_X1 U16194 ( .A1(n14407), .A2(n15003), .B1(P3_REG2_REG_31__SCAN_IN), 
        .B2(n15005), .ZN(n14396) );
  NAND2_X1 U16195 ( .A1(n14398), .A2(n14396), .ZN(P3_U3202) );
  AOI22_X1 U16196 ( .A1(n14411), .A2(n15003), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15005), .ZN(n14397) );
  NAND2_X1 U16197 ( .A1(n14398), .A2(n14397), .ZN(P3_U3203) );
  AOI21_X1 U16198 ( .B1(n15001), .B2(n14400), .A(n14399), .ZN(n14403) );
  AOI22_X1 U16199 ( .A1(n15003), .A2(n14401), .B1(P3_REG2_REG_12__SCAN_IN), 
        .B2(n15005), .ZN(n14402) );
  OAI21_X1 U16200 ( .B1(n14403), .B2(n15005), .A(n14402), .ZN(n14404) );
  INV_X1 U16201 ( .A(n14404), .ZN(n14405) );
  OAI21_X1 U16202 ( .B1(n14406), .B2(n15078), .A(n14405), .ZN(P3_U3221) );
  AOI21_X1 U16203 ( .B1(n14407), .B2(n14410), .A(n14409), .ZN(n14419) );
  INV_X1 U16204 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U16205 ( .A1(n15159), .A2(n14419), .B1(n14408), .B2(n9457), .ZN(
        P3_U3490) );
  AOI21_X1 U16206 ( .B1(n14411), .B2(n14410), .A(n14409), .ZN(n14421) );
  AOI22_X1 U16207 ( .A1(n15159), .A2(n14421), .B1(n14412), .B2(n9457), .ZN(
        P3_U3489) );
  NOR2_X1 U16208 ( .A1(n14413), .A2(n15076), .ZN(n14415) );
  AOI211_X1 U16209 ( .C1(n15136), .C2(n14416), .A(n14415), .B(n14414), .ZN(
        n14422) );
  INV_X1 U16210 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U16211 ( .A1(n15159), .A2(n14422), .B1(n14417), .B2(n9457), .ZN(
        P3_U3470) );
  AOI22_X1 U16212 ( .A1(n15143), .A2(n14419), .B1(n14418), .B2(n15142), .ZN(
        P3_U3458) );
  INV_X1 U16213 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14420) );
  AOI22_X1 U16214 ( .A1(n15143), .A2(n14421), .B1(n14420), .B2(n15142), .ZN(
        P3_U3457) );
  AOI22_X1 U16215 ( .A1(n15143), .A2(n14422), .B1(n8334), .B2(n15142), .ZN(
        P3_U3423) );
  OAI211_X1 U16216 ( .C1(n14425), .C2(n14849), .A(n14424), .B(n14423), .ZN(
        n14426) );
  AOI21_X1 U16217 ( .B1(n14427), .B2(n14440), .A(n14426), .ZN(n14449) );
  AOI22_X1 U16218 ( .A1(n14857), .A2(n14449), .B1(n7792), .B2(n8929), .ZN(
        P2_U3514) );
  NOR2_X1 U16219 ( .A1(n14429), .A2(n14428), .ZN(n14435) );
  OAI211_X1 U16220 ( .C1(n14432), .C2(n14849), .A(n14431), .B(n14430), .ZN(
        n14433) );
  AOI21_X1 U16221 ( .B1(n14435), .B2(n14434), .A(n14433), .ZN(n14452) );
  AOI22_X1 U16222 ( .A1(n14857), .A2(n14452), .B1(n7773), .B2(n8929), .ZN(
        P2_U3513) );
  OAI211_X1 U16223 ( .C1(n14438), .C2(n14849), .A(n14437), .B(n14436), .ZN(
        n14439) );
  AOI21_X1 U16224 ( .B1(n14441), .B2(n14440), .A(n14439), .ZN(n14454) );
  AOI22_X1 U16225 ( .A1(n14857), .A2(n14454), .B1(n11390), .B2(n8929), .ZN(
        P2_U3512) );
  INV_X1 U16226 ( .A(n14442), .ZN(n14447) );
  OAI21_X1 U16227 ( .B1(n14444), .B2(n14849), .A(n14443), .ZN(n14446) );
  AOI211_X1 U16228 ( .C1(n9151), .C2(n14447), .A(n14446), .B(n14445), .ZN(
        n14456) );
  AOI22_X1 U16229 ( .A1(n14857), .A2(n14456), .B1(n11387), .B2(n8929), .ZN(
        P2_U3511) );
  INV_X1 U16230 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U16231 ( .A1(n14854), .A2(n14449), .B1(n14448), .B2(n14450), .ZN(
        P2_U3475) );
  INV_X1 U16232 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U16233 ( .A1(n14457), .A2(n14452), .B1(n14451), .B2(n14450), .ZN(
        P2_U3472) );
  INV_X1 U16234 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14453) );
  AOI22_X1 U16235 ( .A1(n14457), .A2(n14454), .B1(n14453), .B2(n14450), .ZN(
        P2_U3469) );
  INV_X1 U16236 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14455) );
  AOI22_X1 U16237 ( .A1(n14457), .A2(n14456), .B1(n14455), .B2(n14450), .ZN(
        P2_U3466) );
  AND2_X1 U16238 ( .A1(n14459), .A2(n14458), .ZN(n14462) );
  OAI21_X1 U16239 ( .B1(n14462), .B2(n14461), .A(n14460), .ZN(n14463) );
  AOI222_X1 U16240 ( .A1(n14475), .A2(n14481), .B1(n14480), .B2(n14472), .C1(
        n14463), .C2(n14470), .ZN(n14465) );
  OAI211_X1 U16241 ( .C1(n14479), .C2(n14466), .A(n14465), .B(n14464), .ZN(
        P1_U3215) );
  OAI21_X1 U16242 ( .B1(n13587), .B2(n14468), .A(n14467), .ZN(n14469) );
  NAND2_X1 U16243 ( .A1(n7379), .A2(n14469), .ZN(n14471) );
  AOI222_X1 U16244 ( .A1(n14475), .A2(n14474), .B1(n14473), .B2(n14472), .C1(
        n14471), .C2(n14470), .ZN(n14477) );
  OAI211_X1 U16245 ( .C1(n14479), .C2(n14478), .A(n14477), .B(n14476), .ZN(
        P1_U3236) );
  AOI21_X1 U16246 ( .B1(n14481), .B2(n14652), .A(n14480), .ZN(n14486) );
  NAND3_X1 U16247 ( .A1(n14483), .A2(n14482), .A3(n14683), .ZN(n14484) );
  AOI22_X1 U16248 ( .A1(n14709), .A2(n14505), .B1(n14488), .B2(n14706), .ZN(
        P1_U3542) );
  INV_X1 U16249 ( .A(n14489), .ZN(n14496) );
  INV_X1 U16250 ( .A(n14490), .ZN(n14491) );
  OAI211_X1 U16251 ( .C1(n14493), .C2(n14686), .A(n14492), .B(n14491), .ZN(
        n14495) );
  AOI211_X1 U16252 ( .C1(n14496), .C2(n14683), .A(n14495), .B(n14494), .ZN(
        n14507) );
  AOI22_X1 U16253 ( .A1(n14709), .A2(n14507), .B1(n11290), .B2(n14706), .ZN(
        P1_U3541) );
  AND2_X1 U16254 ( .A1(n14497), .A2(n14683), .ZN(n14502) );
  OAI21_X1 U16255 ( .B1(n14499), .B2(n14686), .A(n14498), .ZN(n14500) );
  NOR3_X1 U16256 ( .A1(n14502), .A2(n14501), .A3(n14500), .ZN(n14508) );
  AOI22_X1 U16257 ( .A1(n14709), .A2(n14508), .B1(n14503), .B2(n14706), .ZN(
        P1_U3539) );
  INV_X1 U16258 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14504) );
  AOI22_X1 U16259 ( .A1(n14693), .A2(n14505), .B1(n14504), .B2(n14691), .ZN(
        P1_U3501) );
  INV_X1 U16260 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U16261 ( .A1(n14693), .A2(n14507), .B1(n14506), .B2(n14691), .ZN(
        P1_U3498) );
  AOI22_X1 U16262 ( .A1(n14693), .A2(n14508), .B1(n11177), .B2(n14691), .ZN(
        P1_U3492) );
  AOI21_X1 U16263 ( .B1(n14511), .B2(n14510), .A(n14509), .ZN(n14512) );
  XOR2_X1 U16264 ( .A(n14512), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  XOR2_X1 U16265 ( .A(n6961), .B(n14513), .Z(SUB_1596_U68) );
  AOI21_X1 U16266 ( .B1(n14516), .B2(n14515), .A(n14514), .ZN(n14517) );
  XOR2_X1 U16267 ( .A(n14517), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16268 ( .B1(n14520), .B2(n14519), .A(n14518), .ZN(n14521) );
  XOR2_X1 U16269 ( .A(n14521), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16270 ( .A1(n14523), .A2(n14522), .ZN(n14524) );
  XOR2_X1 U16271 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14524), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16272 ( .B1(n14527), .B2(n14526), .A(n14525), .ZN(n14528) );
  XOR2_X1 U16273 ( .A(n14528), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16274 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14530), .A(n14529), 
        .ZN(n14540) );
  AOI21_X1 U16275 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14532), .A(n14531), 
        .ZN(n14534) );
  OR2_X1 U16276 ( .A1(n14534), .A2(n14533), .ZN(n14538) );
  NAND2_X1 U16277 ( .A1(n14536), .A2(n14535), .ZN(n14537) );
  OAI211_X1 U16278 ( .C1(n14540), .C2(n14539), .A(n14538), .B(n14537), .ZN(
        n14541) );
  INV_X1 U16279 ( .A(n14541), .ZN(n14543) );
  OAI211_X1 U16280 ( .C1(n14545), .C2(n14544), .A(n14543), .B(n14542), .ZN(
        P1_U3258) );
  XNOR2_X1 U16281 ( .A(n14546), .B(n14549), .ZN(n14671) );
  AOI21_X1 U16282 ( .B1(n14547), .B2(n14666), .A(n14575), .ZN(n14548) );
  NAND2_X1 U16283 ( .A1(n14548), .A2(n6438), .ZN(n14667) );
  AOI21_X1 U16284 ( .B1(n14550), .B2(n14549), .A(n14635), .ZN(n14553) );
  AOI21_X1 U16285 ( .B1(n14553), .B2(n14552), .A(n14551), .ZN(n14668) );
  NOR2_X1 U16286 ( .A1(n14555), .A2(n14554), .ZN(n14556) );
  AOI21_X1 U16287 ( .B1(n14666), .B2(n14557), .A(n14556), .ZN(n14558) );
  OAI211_X1 U16288 ( .C1(n14559), .C2(n14667), .A(n14668), .B(n14558), .ZN(
        n14560) );
  AOI21_X1 U16289 ( .B1(n14561), .B2(n14671), .A(n14560), .ZN(n14563) );
  AOI22_X1 U16290 ( .A1(n14599), .A2(n10983), .B1(n14563), .B2(n14562), .ZN(
        P1_U3285) );
  OAI21_X1 U16291 ( .B1(n14565), .B2(n14566), .A(n14564), .ZN(n14571) );
  XNOR2_X1 U16292 ( .A(n14567), .B(n14566), .ZN(n14655) );
  NOR2_X1 U16293 ( .A1(n14655), .A2(n14568), .ZN(n14569) );
  AOI211_X1 U16294 ( .C1(n14625), .C2(n14571), .A(n14570), .B(n14569), .ZN(
        n14654) );
  INV_X1 U16295 ( .A(n14572), .ZN(n14573) );
  AOI222_X1 U16296 ( .A1(n14651), .A2(n14585), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n14599), .C1(n14573), .C2(n14586), .ZN(n14580) );
  INV_X1 U16297 ( .A(n14655), .ZN(n14578) );
  AOI211_X1 U16298 ( .C1(n14651), .C2(n14576), .A(n14575), .B(n14574), .ZN(
        n14650) );
  AOI22_X1 U16299 ( .A1(n14578), .A2(n14577), .B1(n14595), .B2(n14650), .ZN(
        n14579) );
  OAI211_X1 U16300 ( .C1(n14599), .C2(n14654), .A(n14580), .B(n14579), .ZN(
        P1_U3287) );
  XNOR2_X1 U16301 ( .A(n14582), .B(n14581), .ZN(n14584) );
  AOI21_X1 U16302 ( .B1(n14584), .B2(n14625), .A(n14583), .ZN(n14617) );
  AOI222_X1 U16303 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n14599), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14586), .C1(n14589), .C2(n14585), .ZN(
        n14598) );
  XNOR2_X1 U16304 ( .A(n14588), .B(n14587), .ZN(n14620) );
  NAND2_X1 U16305 ( .A1(n14590), .A2(n14589), .ZN(n14592) );
  NAND2_X1 U16306 ( .A1(n14592), .A2(n14591), .ZN(n14593) );
  NOR2_X1 U16307 ( .A1(n14594), .A2(n14593), .ZN(n14614) );
  AOI22_X1 U16308 ( .A1(n14596), .A2(n14620), .B1(n14595), .B2(n14614), .ZN(
        n14597) );
  OAI211_X1 U16309 ( .C1(n14599), .C2(n14617), .A(n14598), .B(n14597), .ZN(
        P1_U3291) );
  AND2_X1 U16310 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14603), .ZN(P1_U3294) );
  AND2_X1 U16311 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14603), .ZN(P1_U3295) );
  AND2_X1 U16312 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14603), .ZN(P1_U3296) );
  AND2_X1 U16313 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14603), .ZN(P1_U3297) );
  AND2_X1 U16314 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14603), .ZN(P1_U3298) );
  AND2_X1 U16315 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14603), .ZN(P1_U3299) );
  AND2_X1 U16316 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14603), .ZN(P1_U3300) );
  AND2_X1 U16317 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14603), .ZN(P1_U3301) );
  AND2_X1 U16318 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14603), .ZN(P1_U3302) );
  AND2_X1 U16319 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14603), .ZN(P1_U3303) );
  AND2_X1 U16320 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14603), .ZN(P1_U3304) );
  AND2_X1 U16321 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14603), .ZN(P1_U3305) );
  AND2_X1 U16322 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14603), .ZN(P1_U3306) );
  NOR2_X1 U16323 ( .A1(n14602), .A2(n14600), .ZN(P1_U3307) );
  AND2_X1 U16324 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14603), .ZN(P1_U3308) );
  AND2_X1 U16325 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14603), .ZN(P1_U3309) );
  NOR2_X1 U16326 ( .A1(n14602), .A2(n14601), .ZN(P1_U3310) );
  AND2_X1 U16327 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14603), .ZN(P1_U3311) );
  AND2_X1 U16328 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14603), .ZN(P1_U3312) );
  AND2_X1 U16329 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14603), .ZN(P1_U3313) );
  AND2_X1 U16330 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14603), .ZN(P1_U3314) );
  AND2_X1 U16331 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14603), .ZN(P1_U3315) );
  AND2_X1 U16332 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14603), .ZN(P1_U3316) );
  AND2_X1 U16333 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14603), .ZN(P1_U3317) );
  AND2_X1 U16334 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14603), .ZN(P1_U3318) );
  AND2_X1 U16335 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14603), .ZN(P1_U3319) );
  AND2_X1 U16336 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14603), .ZN(P1_U3320) );
  AND2_X1 U16337 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14603), .ZN(P1_U3321) );
  AND2_X1 U16338 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14603), .ZN(P1_U3322) );
  AND2_X1 U16339 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14603), .ZN(P1_U3323) );
  INV_X1 U16340 ( .A(n14613), .ZN(n14607) );
  NAND3_X1 U16341 ( .A1(n14605), .A2(n14625), .A3(n14604), .ZN(n14606) );
  OAI21_X1 U16342 ( .B1(n14607), .B2(n14656), .A(n14606), .ZN(n14612) );
  INV_X1 U16343 ( .A(n14608), .ZN(n14610) );
  OAI211_X1 U16344 ( .C1(n6591), .C2(n14686), .A(n14610), .B(n14609), .ZN(
        n14611) );
  AOI211_X1 U16345 ( .C1(n14675), .C2(n14613), .A(n14612), .B(n14611), .ZN(
        n14694) );
  AOI22_X1 U16346 ( .A1(n14693), .A2(n14694), .B1(n9707), .B2(n14691), .ZN(
        P1_U3462) );
  INV_X1 U16347 ( .A(n14614), .ZN(n14615) );
  OAI21_X1 U16348 ( .B1(n14616), .B2(n14686), .A(n14615), .ZN(n14619) );
  INV_X1 U16349 ( .A(n14617), .ZN(n14618) );
  AOI211_X1 U16350 ( .C1(n14620), .C2(n14683), .A(n14619), .B(n14618), .ZN(
        n14695) );
  AOI22_X1 U16351 ( .A1(n14693), .A2(n14695), .B1(n9746), .B2(n14691), .ZN(
        P1_U3465) );
  INV_X1 U16352 ( .A(n14628), .ZN(n14630) );
  OAI211_X1 U16353 ( .C1(n14623), .C2(n14686), .A(n14622), .B(n14621), .ZN(
        n14624) );
  AOI21_X1 U16354 ( .B1(n14626), .B2(n14625), .A(n14624), .ZN(n14627) );
  OAI21_X1 U16355 ( .B1(n14628), .B2(n14656), .A(n14627), .ZN(n14629) );
  AOI21_X1 U16356 ( .B1(n14675), .B2(n14630), .A(n14629), .ZN(n14696) );
  INV_X1 U16357 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14631) );
  AOI22_X1 U16358 ( .A1(n14693), .A2(n14696), .B1(n14631), .B2(n14691), .ZN(
        P1_U3468) );
  OAI211_X1 U16359 ( .C1(n14634), .C2(n14686), .A(n14633), .B(n14632), .ZN(
        n14638) );
  NOR2_X1 U16360 ( .A1(n14636), .A2(n14635), .ZN(n14637) );
  AOI211_X1 U16361 ( .C1(n14639), .C2(n14683), .A(n14638), .B(n14637), .ZN(
        n14697) );
  INV_X1 U16362 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U16363 ( .A1(n14693), .A2(n14697), .B1(n14640), .B2(n14691), .ZN(
        P1_U3471) );
  AND2_X1 U16364 ( .A1(n14641), .A2(n14652), .ZN(n14642) );
  NOR2_X1 U16365 ( .A1(n14643), .A2(n14642), .ZN(n14647) );
  OR2_X1 U16366 ( .A1(n14645), .A2(n14644), .ZN(n14646) );
  AND3_X1 U16367 ( .A1(n14648), .A2(n14647), .A3(n14646), .ZN(n14699) );
  INV_X1 U16368 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14649) );
  AOI22_X1 U16369 ( .A1(n14693), .A2(n14699), .B1(n14649), .B2(n14691), .ZN(
        P1_U3474) );
  AOI21_X1 U16370 ( .B1(n14652), .B2(n14651), .A(n14650), .ZN(n14653) );
  OAI211_X1 U16371 ( .C1(n14656), .C2(n14655), .A(n14654), .B(n14653), .ZN(
        n14657) );
  INV_X1 U16372 ( .A(n14657), .ZN(n14701) );
  INV_X1 U16373 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14658) );
  AOI22_X1 U16374 ( .A1(n14693), .A2(n14701), .B1(n14658), .B2(n14691), .ZN(
        P1_U3477) );
  NAND2_X1 U16375 ( .A1(n14659), .A2(n14674), .ZN(n14661) );
  OAI211_X1 U16376 ( .C1(n14662), .C2(n14686), .A(n14661), .B(n14660), .ZN(
        n14663) );
  NOR2_X1 U16377 ( .A1(n14664), .A2(n14663), .ZN(n14702) );
  INV_X1 U16378 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14665) );
  AOI22_X1 U16379 ( .A1(n14693), .A2(n14702), .B1(n14665), .B2(n14691), .ZN(
        P1_U3480) );
  INV_X1 U16380 ( .A(n14666), .ZN(n14669) );
  OAI211_X1 U16381 ( .C1(n14669), .C2(n14686), .A(n14668), .B(n14667), .ZN(
        n14670) );
  AOI21_X1 U16382 ( .B1(n14671), .B2(n14683), .A(n14670), .ZN(n14703) );
  INV_X1 U16383 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14672) );
  AOI22_X1 U16384 ( .A1(n14693), .A2(n14703), .B1(n14672), .B2(n14691), .ZN(
        P1_U3483) );
  OAI21_X1 U16385 ( .B1(n14675), .B2(n14674), .A(n14673), .ZN(n14676) );
  INV_X1 U16386 ( .A(n14676), .ZN(n14681) );
  OAI21_X1 U16387 ( .B1(n14678), .B2(n14686), .A(n14677), .ZN(n14679) );
  NOR3_X1 U16388 ( .A1(n14681), .A2(n14680), .A3(n14679), .ZN(n14705) );
  INV_X1 U16389 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14682) );
  AOI22_X1 U16390 ( .A1(n14693), .A2(n14705), .B1(n14682), .B2(n14691), .ZN(
        P1_U3486) );
  AND2_X1 U16391 ( .A1(n14684), .A2(n14683), .ZN(n14690) );
  OAI21_X1 U16392 ( .B1(n14687), .B2(n14686), .A(n14685), .ZN(n14688) );
  NOR3_X1 U16393 ( .A1(n14690), .A2(n14689), .A3(n14688), .ZN(n14708) );
  INV_X1 U16394 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14692) );
  AOI22_X1 U16395 ( .A1(n14693), .A2(n14708), .B1(n14692), .B2(n14691), .ZN(
        P1_U3489) );
  AOI22_X1 U16396 ( .A1(n14709), .A2(n14694), .B1(n10016), .B2(n14706), .ZN(
        P1_U3529) );
  AOI22_X1 U16397 ( .A1(n14709), .A2(n14695), .B1(n10015), .B2(n14706), .ZN(
        P1_U3530) );
  AOI22_X1 U16398 ( .A1(n14709), .A2(n14696), .B1(n10021), .B2(n14706), .ZN(
        P1_U3531) );
  AOI22_X1 U16399 ( .A1(n14709), .A2(n14697), .B1(n10024), .B2(n14706), .ZN(
        P1_U3532) );
  AOI22_X1 U16400 ( .A1(n14709), .A2(n14699), .B1(n14698), .B2(n14706), .ZN(
        P1_U3533) );
  AOI22_X1 U16401 ( .A1(n14709), .A2(n14701), .B1(n14700), .B2(n14706), .ZN(
        P1_U3534) );
  AOI22_X1 U16402 ( .A1(n14709), .A2(n14702), .B1(n10966), .B2(n14706), .ZN(
        P1_U3535) );
  AOI22_X1 U16403 ( .A1(n14709), .A2(n14703), .B1(n10979), .B2(n14706), .ZN(
        P1_U3536) );
  AOI22_X1 U16404 ( .A1(n14709), .A2(n14705), .B1(n14704), .B2(n14706), .ZN(
        P1_U3537) );
  AOI22_X1 U16405 ( .A1(n14709), .A2(n14708), .B1(n14707), .B2(n14706), .ZN(
        P1_U3538) );
  NOR2_X1 U16406 ( .A1(n14773), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI21_X1 U16407 ( .B1(n14776), .B2(P2_REG2_REG_0__SCAN_IN), .A(n14710), .ZN(
        n14714) );
  AOI22_X1 U16408 ( .A1(n14773), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14713) );
  OAI22_X1 U16409 ( .A1(n14816), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14822), .ZN(n14711) );
  OAI21_X1 U16410 ( .B1(n14819), .B2(n14711), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14712) );
  OAI211_X1 U16411 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14714), .A(n14713), .B(
        n14712), .ZN(P2_U3214) );
  NAND2_X1 U16412 ( .A1(n14716), .A2(n14715), .ZN(n14717) );
  NAND2_X1 U16413 ( .A1(n14718), .A2(n14717), .ZN(n14719) );
  NAND2_X1 U16414 ( .A1(n14719), .A2(n14779), .ZN(n14726) );
  NAND2_X1 U16415 ( .A1(n14721), .A2(n14720), .ZN(n14722) );
  NAND2_X1 U16416 ( .A1(n14723), .A2(n14722), .ZN(n14724) );
  NAND2_X1 U16417 ( .A1(n14724), .A2(n14776), .ZN(n14725) );
  OAI211_X1 U16418 ( .C1(n14807), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        n14728) );
  INV_X1 U16419 ( .A(n14728), .ZN(n14730) );
  OAI211_X1 U16420 ( .C1(n14731), .C2(n14827), .A(n14730), .B(n14729), .ZN(
        P2_U3223) );
  AND2_X1 U16421 ( .A1(n14733), .A2(n14732), .ZN(n14734) );
  OAI21_X1 U16422 ( .B1(n14735), .B2(n14734), .A(n14779), .ZN(n14745) );
  INV_X1 U16423 ( .A(n14736), .ZN(n14738) );
  NAND3_X1 U16424 ( .A1(n14739), .A2(n14738), .A3(n14737), .ZN(n14740) );
  NAND2_X1 U16425 ( .A1(n14741), .A2(n14740), .ZN(n14743) );
  AOI22_X1 U16426 ( .A1(n14743), .A2(n14776), .B1(n14742), .B2(n14819), .ZN(
        n14744) );
  AND2_X1 U16427 ( .A1(n14745), .A2(n14744), .ZN(n14747) );
  OAI211_X1 U16428 ( .C1(n6961), .C2(n14827), .A(n14747), .B(n14746), .ZN(
        P2_U3226) );
  OAI21_X1 U16429 ( .B1(n14807), .B2(n14749), .A(n14748), .ZN(n14750) );
  AOI21_X1 U16430 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n14773), .A(n14750), 
        .ZN(n14759) );
  OAI211_X1 U16431 ( .C1(n14753), .C2(n14752), .A(n14751), .B(n14779), .ZN(
        n14758) );
  OAI211_X1 U16432 ( .C1(n14756), .C2(n14755), .A(n14754), .B(n14776), .ZN(
        n14757) );
  NAND3_X1 U16433 ( .A1(n14759), .A2(n14758), .A3(n14757), .ZN(P2_U3227) );
  NOR2_X1 U16434 ( .A1(n14761), .A2(n14760), .ZN(n14762) );
  XOR2_X1 U16435 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n14762), .Z(n14770) );
  XNOR2_X1 U16436 ( .A(n14764), .B(n14763), .ZN(n14765) );
  NAND2_X1 U16437 ( .A1(n14765), .A2(n14779), .ZN(n14767) );
  OAI211_X1 U16438 ( .C1(n14768), .C2(n14827), .A(n14767), .B(n14766), .ZN(
        n14769) );
  AOI21_X1 U16439 ( .B1(n14770), .B2(n14776), .A(n14769), .ZN(n14771) );
  OAI21_X1 U16440 ( .B1(n14772), .B2(n14807), .A(n14771), .ZN(P2_U3228) );
  AOI22_X1 U16441 ( .A1(n14773), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14784) );
  NAND2_X1 U16442 ( .A1(n14819), .A2(n14774), .ZN(n14783) );
  OAI211_X1 U16443 ( .C1(n14777), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14776), 
        .B(n14775), .ZN(n14782) );
  OAI211_X1 U16444 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n14780), .A(n14779), 
        .B(n14778), .ZN(n14781) );
  NAND4_X1 U16445 ( .A1(n14784), .A2(n14783), .A3(n14782), .A4(n14781), .ZN(
        P2_U3229) );
  OAI21_X1 U16446 ( .B1(n14787), .B2(n14786), .A(n14785), .ZN(n14792) );
  OAI21_X1 U16447 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n14791) );
  OAI222_X1 U16448 ( .A1(n14807), .A2(n14793), .B1(n14816), .B2(n14792), .C1(
        n14822), .C2(n14791), .ZN(n14794) );
  INV_X1 U16449 ( .A(n14794), .ZN(n14796) );
  OAI211_X1 U16450 ( .C1(n14797), .C2(n14827), .A(n14796), .B(n14795), .ZN(
        P2_U3230) );
  OAI21_X1 U16451 ( .B1(n14800), .B2(n14799), .A(n14798), .ZN(n14805) );
  OAI21_X1 U16452 ( .B1(n14803), .B2(n14802), .A(n14801), .ZN(n14804) );
  OAI222_X1 U16453 ( .A1(n14807), .A2(n14806), .B1(n14816), .B2(n14805), .C1(
        n14822), .C2(n14804), .ZN(n14808) );
  INV_X1 U16454 ( .A(n14808), .ZN(n14810) );
  OAI211_X1 U16455 ( .C1(n14811), .C2(n14827), .A(n14810), .B(n14809), .ZN(
        P2_U3231) );
  OAI21_X1 U16456 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n14813), .A(n14812), 
        .ZN(n14823) );
  AOI21_X1 U16457 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14815), .A(n14814), 
        .ZN(n14817) );
  OR2_X1 U16458 ( .A1(n14817), .A2(n14816), .ZN(n14821) );
  NAND2_X1 U16459 ( .A1(n14819), .A2(n14818), .ZN(n14820) );
  OAI211_X1 U16460 ( .C1(n14823), .C2(n14822), .A(n14821), .B(n14820), .ZN(
        n14824) );
  INV_X1 U16461 ( .A(n14824), .ZN(n14826) );
  OAI211_X1 U16462 ( .C1(n14828), .C2(n14827), .A(n14826), .B(n14825), .ZN(
        P2_U3232) );
  NOR2_X1 U16463 ( .A1(n14837), .A2(n14829), .ZN(n14831) );
  AND2_X1 U16464 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14832), .ZN(P2_U3266) );
  AND2_X1 U16465 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14832), .ZN(P2_U3267) );
  AND2_X1 U16466 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14832), .ZN(P2_U3268) );
  AND2_X1 U16467 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14832), .ZN(P2_U3269) );
  AND2_X1 U16468 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14832), .ZN(P2_U3270) );
  NOR2_X1 U16469 ( .A1(n14831), .A2(n14830), .ZN(P2_U3271) );
  AND2_X1 U16470 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14832), .ZN(P2_U3272) );
  AND2_X1 U16471 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14832), .ZN(P2_U3273) );
  AND2_X1 U16472 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14832), .ZN(P2_U3274) );
  AND2_X1 U16473 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14832), .ZN(P2_U3275) );
  AND2_X1 U16474 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14832), .ZN(P2_U3276) );
  AND2_X1 U16475 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14832), .ZN(P2_U3277) );
  AND2_X1 U16476 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14832), .ZN(P2_U3278) );
  AND2_X1 U16477 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14832), .ZN(P2_U3279) );
  AND2_X1 U16478 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14832), .ZN(P2_U3280) );
  AND2_X1 U16479 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14832), .ZN(P2_U3281) );
  AND2_X1 U16480 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14832), .ZN(P2_U3282) );
  AND2_X1 U16481 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14832), .ZN(P2_U3283) );
  AND2_X1 U16482 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14832), .ZN(P2_U3284) );
  AND2_X1 U16483 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14832), .ZN(P2_U3285) );
  AND2_X1 U16484 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14832), .ZN(P2_U3286) );
  AND2_X1 U16485 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14832), .ZN(P2_U3287) );
  AND2_X1 U16486 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14832), .ZN(P2_U3288) );
  AND2_X1 U16487 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14832), .ZN(P2_U3289) );
  AND2_X1 U16488 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14832), .ZN(P2_U3290) );
  AND2_X1 U16489 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14832), .ZN(P2_U3291) );
  AND2_X1 U16490 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14832), .ZN(P2_U3292) );
  AND2_X1 U16491 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14832), .ZN(P2_U3293) );
  AND2_X1 U16492 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14832), .ZN(P2_U3294) );
  AND2_X1 U16493 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14832), .ZN(P2_U3295) );
  AOI22_X1 U16494 ( .A1(n14835), .A2(n14834), .B1(n14833), .B2(n14837), .ZN(
        P2_U3416) );
  AOI21_X1 U16495 ( .B1(n14838), .B2(n14837), .A(n14836), .ZN(P2_U3417) );
  INV_X1 U16496 ( .A(n14839), .ZN(n14845) );
  INV_X1 U16497 ( .A(n14840), .ZN(n14841) );
  OAI21_X1 U16498 ( .B1(n14842), .B2(n14849), .A(n14841), .ZN(n14844) );
  AOI211_X1 U16499 ( .C1(n9151), .C2(n14845), .A(n14844), .B(n14843), .ZN(
        n14855) );
  INV_X1 U16500 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14846) );
  AOI22_X1 U16501 ( .A1(n14854), .A2(n14855), .B1(n14846), .B2(n14450), .ZN(
        P2_U3454) );
  INV_X1 U16502 ( .A(n14847), .ZN(n14852) );
  OAI21_X1 U16503 ( .B1(n6944), .B2(n14849), .A(n14848), .ZN(n14851) );
  AOI211_X1 U16504 ( .C1(n9151), .C2(n14852), .A(n14851), .B(n14850), .ZN(
        n14856) );
  INV_X1 U16505 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14853) );
  AOI22_X1 U16506 ( .A1(n14854), .A2(n14856), .B1(n14853), .B2(n14450), .ZN(
        P2_U3460) );
  AOI22_X1 U16507 ( .A1(n14857), .A2(n14855), .B1(n9965), .B2(n8929), .ZN(
        P2_U3507) );
  AOI22_X1 U16508 ( .A1(n14857), .A2(n14856), .B1(n9978), .B2(n8929), .ZN(
        P2_U3509) );
  NOR2_X1 U16509 ( .A1(P3_U3897), .A2(n14984), .ZN(P3_U3150) );
  INV_X1 U16510 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n14872) );
  INV_X1 U16511 ( .A(n14858), .ZN(n14862) );
  AOI222_X1 U16512 ( .A1(n14862), .A2(n14861), .B1(n15083), .B2(n14860), .C1(
        n6906), .C2(n14859), .ZN(n14863) );
  OAI21_X1 U16513 ( .B1(n14864), .B2(n14872), .A(n14863), .ZN(P3_U3172) );
  NAND3_X1 U16514 ( .A1(n14997), .A2(n14877), .A3(n14952), .ZN(n14869) );
  NAND2_X1 U16515 ( .A1(n14869), .A2(n14868), .ZN(n14870) );
  OAI211_X1 U16516 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n14872), .A(n14871), .B(
        n14870), .ZN(P3_U3182) );
  XNOR2_X1 U16517 ( .A(n14874), .B(n14873), .ZN(n14883) );
  XOR2_X1 U16518 ( .A(P3_REG1_REG_5__SCAN_IN), .B(n14875), .Z(n14876) );
  NOR2_X1 U16519 ( .A1(n14877), .A2(n14876), .ZN(n14882) );
  AOI21_X1 U16520 ( .B1(n14879), .B2(n15037), .A(n14878), .ZN(n14880) );
  OAI22_X1 U16521 ( .A1(n14880), .A2(n14997), .B1(n6844), .B2(n14987), .ZN(
        n14881) );
  AOI211_X1 U16522 ( .C1(n14991), .C2(n14883), .A(n14882), .B(n14881), .ZN(
        n14885) );
  OAI211_X1 U16523 ( .C1(n14887), .C2(n14886), .A(n14885), .B(n14884), .ZN(
        P3_U3187) );
  AOI21_X1 U16524 ( .B1(n14890), .B2(n14889), .A(n14888), .ZN(n14905) );
  NOR2_X1 U16525 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14891), .ZN(n14899) );
  NAND2_X1 U16526 ( .A1(n14893), .A2(n14892), .ZN(n14894) );
  XNOR2_X1 U16527 ( .A(n14895), .B(n14894), .ZN(n14897) );
  OAI22_X1 U16528 ( .A1(n14897), .A2(n14952), .B1(n14896), .B2(n14987), .ZN(
        n14898) );
  AOI211_X1 U16529 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14984), .A(n14899), .B(
        n14898), .ZN(n14904) );
  OAI21_X1 U16530 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14901), .A(n14900), .ZN(
        n14902) );
  NAND2_X1 U16531 ( .A1(n14902), .A2(n14989), .ZN(n14903) );
  OAI211_X1 U16532 ( .C1(n14905), .C2(n14997), .A(n14904), .B(n14903), .ZN(
        P3_U3191) );
  AOI21_X1 U16533 ( .B1(n14908), .B2(n14907), .A(n14906), .ZN(n14923) );
  OAI21_X1 U16534 ( .B1(n14911), .B2(n14910), .A(n14909), .ZN(n14916) );
  AOI21_X1 U16535 ( .B1(n14984), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n14912), 
        .ZN(n14913) );
  OAI21_X1 U16536 ( .B1(n14987), .B2(n14914), .A(n14913), .ZN(n14915) );
  AOI21_X1 U16537 ( .B1(n14916), .B2(n14989), .A(n14915), .ZN(n14922) );
  OAI21_X1 U16538 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(n14920) );
  NAND2_X1 U16539 ( .A1(n14991), .A2(n14920), .ZN(n14921) );
  OAI211_X1 U16540 ( .C1(n14923), .C2(n14997), .A(n14922), .B(n14921), .ZN(
        P3_U3192) );
  AOI21_X1 U16541 ( .B1(n14926), .B2(n14925), .A(n14924), .ZN(n14940) );
  OAI21_X1 U16542 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n14928), .A(n14927), 
        .ZN(n14933) );
  AOI21_X1 U16543 ( .B1(n14984), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n14929), 
        .ZN(n14930) );
  OAI21_X1 U16544 ( .B1(n14987), .B2(n14931), .A(n14930), .ZN(n14932) );
  AOI21_X1 U16545 ( .B1(n14933), .B2(n14989), .A(n14932), .ZN(n14939) );
  OAI21_X1 U16546 ( .B1(n14936), .B2(n14935), .A(n14934), .ZN(n14937) );
  NAND2_X1 U16547 ( .A1(n14937), .A2(n14991), .ZN(n14938) );
  OAI211_X1 U16548 ( .C1(n14940), .C2(n14997), .A(n14939), .B(n14938), .ZN(
        P3_U3193) );
  AOI21_X1 U16549 ( .B1(n14943), .B2(n14942), .A(n14941), .ZN(n14959) );
  OAI21_X1 U16550 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n14951) );
  AOI21_X1 U16551 ( .B1(n14984), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n14947), 
        .ZN(n14948) );
  OAI21_X1 U16552 ( .B1(n14987), .B2(n14949), .A(n14948), .ZN(n14950) );
  AOI21_X1 U16553 ( .B1(n14951), .B2(n14989), .A(n14950), .ZN(n14958) );
  AOI21_X1 U16554 ( .B1(n14954), .B2(n14953), .A(n14952), .ZN(n14956) );
  NAND2_X1 U16555 ( .A1(n14956), .A2(n14955), .ZN(n14957) );
  OAI211_X1 U16556 ( .C1(n14959), .C2(n14997), .A(n14958), .B(n14957), .ZN(
        P3_U3194) );
  AOI21_X1 U16557 ( .B1(n14962), .B2(n14961), .A(n14960), .ZN(n14976) );
  OAI21_X1 U16558 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n14964), .A(n14963), 
        .ZN(n14969) );
  AOI21_X1 U16559 ( .B1(n14984), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n14965), 
        .ZN(n14966) );
  OAI21_X1 U16560 ( .B1(n14987), .B2(n14967), .A(n14966), .ZN(n14968) );
  AOI21_X1 U16561 ( .B1(n14969), .B2(n14989), .A(n14968), .ZN(n14975) );
  OAI21_X1 U16562 ( .B1(n14972), .B2(n14971), .A(n14970), .ZN(n14973) );
  NAND2_X1 U16563 ( .A1(n14973), .A2(n14991), .ZN(n14974) );
  OAI211_X1 U16564 ( .C1(n14976), .C2(n14997), .A(n14975), .B(n14974), .ZN(
        P3_U3195) );
  AOI21_X1 U16565 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n14998) );
  OAI21_X1 U16566 ( .B1(n14982), .B2(n14981), .A(n14980), .ZN(n14990) );
  AOI21_X1 U16567 ( .B1(n14984), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n14983), 
        .ZN(n14985) );
  OAI21_X1 U16568 ( .B1(n14987), .B2(n14986), .A(n14985), .ZN(n14988) );
  AOI21_X1 U16569 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14996) );
  OAI211_X1 U16570 ( .C1(n14994), .C2(n14993), .A(n14992), .B(n14991), .ZN(
        n14995) );
  OAI211_X1 U16571 ( .C1(n14998), .C2(n14997), .A(n14996), .B(n14995), .ZN(
        P3_U3196) );
  AOI21_X1 U16572 ( .B1(n15001), .B2(n15000), .A(n14999), .ZN(n15006) );
  AOI22_X1 U16573 ( .A1(n15003), .A2(n15002), .B1(P3_REG2_REG_10__SCAN_IN), 
        .B2(n15005), .ZN(n15004) );
  OAI21_X1 U16574 ( .B1(n15006), .B2(n15005), .A(n15004), .ZN(n15007) );
  INV_X1 U16575 ( .A(n15007), .ZN(n15008) );
  OAI21_X1 U16576 ( .B1(n15009), .B2(n15078), .A(n15008), .ZN(P3_U3223) );
  INV_X1 U16577 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n15023) );
  NOR2_X1 U16578 ( .A1(n15010), .A2(n15076), .ZN(n15135) );
  AOI22_X1 U16579 ( .A1(n15070), .A2(n15135), .B1(n15103), .B2(n15011), .ZN(
        n15022) );
  INV_X1 U16580 ( .A(n15012), .ZN(n15013) );
  AOI21_X1 U16581 ( .B1(n15018), .B2(n15014), .A(n15013), .ZN(n15015) );
  OAI222_X1 U16582 ( .A1(n15046), .A2(n15017), .B1(n15044), .B2(n15016), .C1(
        n15052), .C2(n15015), .ZN(n15134) );
  XNOR2_X1 U16583 ( .A(n15019), .B(n15018), .ZN(n15137) );
  AOI22_X1 U16584 ( .A1(n15134), .A2(n15109), .B1(n15137), .B2(n15020), .ZN(
        n15021) );
  OAI211_X1 U16585 ( .C1(n15023), .C2(n15109), .A(n15022), .B(n15021), .ZN(
        P3_U3225) );
  XNOR2_X1 U16586 ( .A(n15024), .B(n15026), .ZN(n15033) );
  INV_X1 U16587 ( .A(n15033), .ZN(n15124) );
  OAI21_X1 U16588 ( .B1(n15027), .B2(n15026), .A(n15025), .ZN(n15031) );
  OAI22_X1 U16589 ( .A1(n15029), .A2(n15044), .B1(n15028), .B2(n15046), .ZN(
        n15030) );
  AOI21_X1 U16590 ( .B1(n15031), .B2(n15089), .A(n15030), .ZN(n15032) );
  OAI21_X1 U16591 ( .B1(n15094), .B2(n15033), .A(n15032), .ZN(n15122) );
  AOI21_X1 U16592 ( .B1(n15097), .B2(n15124), .A(n15122), .ZN(n15038) );
  NOR2_X1 U16593 ( .A1(n15034), .A2(n15076), .ZN(n15123) );
  AOI22_X1 U16594 ( .A1(n15070), .A2(n15123), .B1(n15103), .B2(n15035), .ZN(
        n15036) );
  OAI221_X1 U16595 ( .B1(n15005), .B2(n15038), .C1(n15109), .C2(n15037), .A(
        n15036), .ZN(P3_U3228) );
  NOR2_X1 U16596 ( .A1(n15039), .A2(n15076), .ZN(n15120) );
  AOI22_X1 U16597 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n15005), .B1(n15070), 
        .B2(n15120), .ZN(n15056) );
  XNOR2_X1 U16598 ( .A(n15040), .B(n15041), .ZN(n15051) );
  XNOR2_X1 U16599 ( .A(n15043), .B(n15042), .ZN(n15121) );
  OAI22_X1 U16600 ( .A1(n15047), .A2(n15046), .B1(n15045), .B2(n15044), .ZN(
        n15048) );
  AOI21_X1 U16601 ( .B1(n15121), .B2(n15049), .A(n15048), .ZN(n15050) );
  OAI21_X1 U16602 ( .B1(n15052), .B2(n15051), .A(n15050), .ZN(n15119) );
  INV_X1 U16603 ( .A(n15121), .ZN(n15053) );
  NOR2_X1 U16604 ( .A1(n15053), .A2(n15106), .ZN(n15054) );
  OAI21_X1 U16605 ( .B1(n15119), .B2(n15054), .A(n15109), .ZN(n15055) );
  OAI211_X1 U16606 ( .C1(n15057), .C2(n15078), .A(n15056), .B(n15055), .ZN(
        P3_U3229) );
  INV_X1 U16607 ( .A(n15059), .ZN(n15064) );
  XNOR2_X1 U16608 ( .A(n15058), .B(n15064), .ZN(n15068) );
  INV_X1 U16609 ( .A(n15068), .ZN(n15118) );
  AOI22_X1 U16610 ( .A1(n15084), .A2(n15061), .B1(n15060), .B2(n15081), .ZN(
        n15067) );
  INV_X1 U16611 ( .A(n15062), .ZN(n15065) );
  OAI211_X1 U16612 ( .C1(n15065), .C2(n15064), .A(n15089), .B(n15063), .ZN(
        n15066) );
  OAI211_X1 U16613 ( .C1(n15068), .C2(n15094), .A(n15067), .B(n15066), .ZN(
        n15116) );
  AOI21_X1 U16614 ( .B1(n15097), .B2(n15118), .A(n15116), .ZN(n15073) );
  INV_X1 U16615 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n15072) );
  NOR2_X1 U16616 ( .A1(n15069), .A2(n15076), .ZN(n15117) );
  AOI22_X1 U16617 ( .A1(n15070), .A2(n15117), .B1(n15103), .B2(n8203), .ZN(
        n15071) );
  OAI221_X1 U16618 ( .B1(n15005), .B2(n15073), .C1(n15109), .C2(n15072), .A(
        n15071), .ZN(P3_U3230) );
  INV_X1 U16619 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15099) );
  XNOR2_X1 U16620 ( .A(n15075), .B(n15074), .ZN(n15095) );
  INV_X1 U16621 ( .A(n15095), .ZN(n15115) );
  NOR2_X1 U16622 ( .A1(n15077), .A2(n15076), .ZN(n15114) );
  INV_X1 U16623 ( .A(n15114), .ZN(n15080) );
  OAI22_X1 U16624 ( .A1(n15080), .A2(n15079), .B1(n15078), .B2(n9662), .ZN(
        n15096) );
  AOI22_X1 U16625 ( .A1(n15084), .A2(n15083), .B1(n15082), .B2(n15081), .ZN(
        n15093) );
  INV_X1 U16626 ( .A(n15085), .ZN(n15091) );
  AND3_X1 U16627 ( .A1(n15087), .A2(n15088), .A3(n15086), .ZN(n15090) );
  OAI21_X1 U16628 ( .B1(n15091), .B2(n15090), .A(n15089), .ZN(n15092) );
  OAI211_X1 U16629 ( .C1(n15095), .C2(n15094), .A(n15093), .B(n15092), .ZN(
        n15113) );
  AOI211_X1 U16630 ( .C1(n15097), .C2(n15115), .A(n15096), .B(n15113), .ZN(
        n15098) );
  AOI22_X1 U16631 ( .A1(n15005), .A2(n15099), .B1(n15098), .B2(n15109), .ZN(
        P3_U3231) );
  INV_X1 U16632 ( .A(n15100), .ZN(n15107) );
  AOI22_X1 U16633 ( .A1(n15103), .A2(P3_REG3_REG_1__SCAN_IN), .B1(n15102), 
        .B2(n15101), .ZN(n15104) );
  OAI211_X1 U16634 ( .C1(n15107), .C2(n15106), .A(n15105), .B(n15104), .ZN(
        n15108) );
  INV_X1 U16635 ( .A(n15108), .ZN(n15110) );
  AOI22_X1 U16636 ( .A1(n15005), .A2(n15111), .B1(n15110), .B2(n15109), .ZN(
        P3_U3232) );
  AOI22_X1 U16637 ( .A1(n15143), .A2(n15112), .B1(n8170), .B2(n15142), .ZN(
        P3_U3393) );
  AOI211_X1 U16638 ( .C1(n15115), .C2(n15140), .A(n15114), .B(n15113), .ZN(
        n15145) );
  AOI22_X1 U16639 ( .A1(n15143), .A2(n15145), .B1(n8191), .B2(n15142), .ZN(
        P3_U3396) );
  AOI211_X1 U16640 ( .C1(n15118), .C2(n15140), .A(n15117), .B(n15116), .ZN(
        n15146) );
  AOI22_X1 U16641 ( .A1(n15143), .A2(n15146), .B1(n8204), .B2(n15142), .ZN(
        P3_U3399) );
  AOI211_X1 U16642 ( .C1(n15121), .C2(n15140), .A(n15120), .B(n15119), .ZN(
        n15148) );
  AOI22_X1 U16643 ( .A1(n15143), .A2(n15148), .B1(n8218), .B2(n15142), .ZN(
        P3_U3402) );
  AOI211_X1 U16644 ( .C1(n15124), .C2(n15140), .A(n15123), .B(n15122), .ZN(
        n15150) );
  AOI22_X1 U16645 ( .A1(n15143), .A2(n15150), .B1(n8235), .B2(n15142), .ZN(
        P3_U3405) );
  INV_X1 U16646 ( .A(n15125), .ZN(n15127) );
  AOI211_X1 U16647 ( .C1(n15128), .C2(n15140), .A(n15127), .B(n15126), .ZN(
        n15152) );
  AOI22_X1 U16648 ( .A1(n15143), .A2(n15152), .B1(n8251), .B2(n15142), .ZN(
        P3_U3408) );
  INV_X1 U16649 ( .A(n15129), .ZN(n15133) );
  INV_X1 U16650 ( .A(n15130), .ZN(n15131) );
  AOI211_X1 U16651 ( .C1(n15133), .C2(n15140), .A(n15132), .B(n15131), .ZN(
        n15154) );
  AOI22_X1 U16652 ( .A1(n15143), .A2(n15154), .B1(n8267), .B2(n15142), .ZN(
        P3_U3411) );
  AOI211_X1 U16653 ( .C1(n15137), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        n15156) );
  AOI22_X1 U16654 ( .A1(n15143), .A2(n15156), .B1(n8283), .B2(n15142), .ZN(
        P3_U3414) );
  AOI211_X1 U16655 ( .C1(n15141), .C2(n15140), .A(n15139), .B(n15138), .ZN(
        n15158) );
  AOI22_X1 U16656 ( .A1(n15143), .A2(n15158), .B1(n8302), .B2(n15142), .ZN(
        P3_U3417) );
  INV_X1 U16657 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15144) );
  AOI22_X1 U16658 ( .A1(n15159), .A2(n15145), .B1(n15144), .B2(n9457), .ZN(
        P3_U3461) );
  AOI22_X1 U16659 ( .A1(n15159), .A2(n15146), .B1(n10321), .B2(n9457), .ZN(
        P3_U3462) );
  AOI22_X1 U16660 ( .A1(n15159), .A2(n15148), .B1(n15147), .B2(n9457), .ZN(
        P3_U3463) );
  INV_X1 U16661 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15149) );
  AOI22_X1 U16662 ( .A1(n15159), .A2(n15150), .B1(n15149), .B2(n9457), .ZN(
        P3_U3464) );
  AOI22_X1 U16663 ( .A1(n15159), .A2(n15152), .B1(n15151), .B2(n9457), .ZN(
        P3_U3465) );
  INV_X1 U16664 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U16665 ( .A1(n15159), .A2(n15154), .B1(n15153), .B2(n9457), .ZN(
        P3_U3466) );
  AOI22_X1 U16666 ( .A1(n15159), .A2(n15156), .B1(n15155), .B2(n9457), .ZN(
        P3_U3467) );
  AOI22_X1 U16667 ( .A1(n15159), .A2(n15158), .B1(n15157), .B2(n9457), .ZN(
        P3_U3468) );
  XNOR2_X1 U16668 ( .A(n15160), .B(n15161), .ZN(SUB_1596_U59) );
  XNOR2_X1 U16669 ( .A(n15162), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16670 ( .B1(n15164), .B2(n15163), .A(n15173), .ZN(SUB_1596_U53) );
  XNOR2_X1 U16671 ( .A(n15166), .B(n15165), .ZN(SUB_1596_U56) );
  OAI21_X1 U16672 ( .B1(n15169), .B2(n15168), .A(n15167), .ZN(n15171) );
  XOR2_X1 U16673 ( .A(n15171), .B(n15170), .Z(SUB_1596_U60) );
  XOR2_X1 U16674 ( .A(n15173), .B(n15172), .Z(SUB_1596_U5) );
  AND2_X1 U7241 ( .A1(n8154), .A2(n8155), .ZN(n6419) );
  BUF_X2 U7148 ( .A(n6419), .Z(n8606) );
  INV_X2 U7245 ( .A(n11178), .ZN(n12154) );
  AND2_X1 U7210 ( .A1(n14042), .A2(n14041), .ZN(n14044) );
  AND2_X1 U7139 ( .A1(n11211), .A2(n14687), .ZN(n11212) );
  CLKBUF_X1 U7153 ( .A(n12572), .Z(n6392) );
  CLKBUF_X1 U7178 ( .A(n13064), .Z(n6644) );
  OR2_X1 U7274 ( .A1(n14125), .A2(n6938), .ZN(n6453) );
  INV_X2 U7275 ( .A(n11992), .ZN(n6591) );
  XNOR2_X1 U7465 ( .A(n12249), .B(n8787), .ZN(n12358) );
  CLKBUF_X1 U7548 ( .A(n13008), .Z(n6399) );
  CLKBUF_X1 U7858 ( .A(n9791), .Z(n6415) );
endmodule

