

module b17_C_gen_AntiSAT_k_256_9 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332;

  NAND2_X1 U11242 ( .A1(n15480), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15479) );
  INV_X1 U11243 ( .A(n17393), .ZN(n18350) );
  NAND2_X1 U11244 ( .A1(n9947), .A2(n11966), .ZN(n12051) );
  OR2_X2 U11245 ( .A1(n11985), .A2(n11979), .ZN(n12064) );
  BUF_X1 U11246 ( .A(n12968), .Z(n15764) );
  INV_X2 U11247 ( .A(n17296), .ZN(n17276) );
  AND2_X1 U11248 ( .A1(n13278), .A2(n11619), .ZN(n11772) );
  AND2_X1 U11249 ( .A1(n13280), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11790) );
  AND2_X1 U11250 ( .A1(n11759), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11782) );
  INV_X1 U11251 ( .A(n13764), .ZN(n17304) );
  INV_X2 U11252 ( .A(n11300), .ZN(n17145) );
  INV_X2 U11253 ( .A(n17172), .ZN(n17243) );
  INV_X2 U11254 ( .A(n10327), .ZN(n17297) );
  CLKBUF_X2 U11256 ( .A(n9839), .Z(n10495) );
  NAND2_X1 U11257 ( .A1(n11718), .A2(n11717), .ZN(n11851) );
  NAND2_X1 U11258 ( .A1(n10118), .A2(n10116), .ZN(n11820) );
  AND2_X2 U11260 ( .A1(n15768), .A2(n15769), .ZN(n13275) );
  BUF_X2 U11261 ( .A(n10431), .Z(n11063) );
  AND2_X1 U11262 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15766) );
  AND2_X1 U11263 ( .A1(n13942), .A2(n13612), .ZN(n11109) );
  CLKBUF_X1 U11264 ( .A(n18505), .Z(n9798) );
  NOR2_X1 U11265 ( .A1(n18822), .A2(n18467), .ZN(n18505) );
  NOR2_X1 U11266 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11601) );
  CLKBUF_X2 U11267 ( .A(n11109), .Z(n11049) );
  AND2_X1 U11268 ( .A1(n10142), .A2(n9897), .ZN(n9949) );
  AND2_X1 U11269 ( .A1(n11853), .A2(n11837), .ZN(n11847) );
  NAND2_X2 U11271 ( .A1(n11886), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12360) );
  CLKBUF_X1 U11272 ( .A(n11758), .Z(n15772) );
  AND2_X1 U11273 ( .A1(n13278), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12080) );
  NAND2_X1 U11274 ( .A1(n14132), .A2(n12188), .ZN(n12810) );
  OR2_X2 U11275 ( .A1(n11985), .A2(n11975), .ZN(n12061) );
  OR2_X1 U11276 ( .A1(n11972), .A2(n11979), .ZN(n19588) );
  AND2_X1 U11277 ( .A1(n12956), .A2(n15764), .ZN(n11981) );
  NOR2_X1 U11278 ( .A1(n14762), .A2(n14759), .ZN(n15982) );
  INV_X1 U11279 ( .A(n12793), .ZN(n12795) );
  NAND2_X1 U11280 ( .A1(n11930), .A2(n11929), .ZN(n11947) );
  OR2_X1 U11281 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15818), .ZN(
        n13764) );
  INV_X2 U11282 ( .A(n11450), .ZN(n17293) );
  INV_X1 U11283 ( .A(n13764), .ZN(n9804) );
  AOI211_X1 U11284 ( .C1(n9808), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n11487), .B(n11486), .ZN(n18342) );
  NOR2_X1 U11285 ( .A1(n10155), .A2(n20274), .ZN(n10470) );
  AND2_X1 U11286 ( .A1(n14352), .A2(n10318), .ZN(n12672) );
  AND2_X1 U11287 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n12631), .ZN(
        n12947) );
  OAI211_X1 U11288 ( .C1(n12326), .C2(n12195), .A(n12194), .B(n12208), .ZN(
        n13515) );
  OR2_X1 U11289 ( .A1(n13554), .A2(n10209), .ZN(n15056) );
  NAND2_X1 U11290 ( .A1(n10050), .A2(n10049), .ZN(n16323) );
  OR2_X1 U11291 ( .A1(n13642), .A2(n13641), .ZN(n13644) );
  NOR2_X1 U11292 ( .A1(n18796), .A2(n18814), .ZN(n18271) );
  INV_X1 U11293 ( .A(n13566), .ZN(n12771) );
  XNOR2_X1 U11294 ( .A(n14959), .B(n12897), .ZN(n16210) );
  INV_X1 U11295 ( .A(n15680), .ZN(n14008) );
  NAND2_X1 U11296 ( .A1(n13515), .A2(n13516), .ZN(n13518) );
  AOI22_X1 U11297 ( .A1(n16089), .A2(n20260), .B1(n16173), .B2(n16088), .ZN(
        n16091) );
  XNOR2_X1 U11298 ( .A(n14975), .B(n14976), .ZN(n15514) );
  BUF_X1 U11299 ( .A(n15019), .Z(n9807) );
  AND2_X2 U11300 ( .A1(n10363), .A2(n10370), .ZN(n9799) );
  AND4_X1 U11301 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n9800) );
  AND4_X1 U11302 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n9801) );
  NAND2_X2 U11303 ( .A1(n10293), .A2(n10292), .ZN(n10643) );
  NOR3_X4 U11304 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n11308), .ZN(n11518) );
  INV_X2 U11305 ( .A(n11309), .ZN(n15798) );
  OR2_X2 U11306 ( .A1(n14750), .A2(n14749), .ZN(n14762) );
  AND2_X2 U11307 ( .A1(n11759), .A2(n11619), .ZN(n11788) );
  INV_X1 U11308 ( .A(n12584), .ZN(n9802) );
  AND2_X4 U11309 ( .A1(n11653), .A2(n11652), .ZN(n12584) );
  AND2_X4 U11310 ( .A1(n11873), .A2(n11887), .ZN(n11925) );
  AND4_X2 U11311 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10375) );
  AOI21_X2 U11312 ( .B1(n14329), .B2(n14327), .A(n14328), .ZN(n14638) );
  NAND2_X2 U11315 ( .A1(n11742), .A2(n11741), .ZN(n11839) );
  NAND2_X2 U11317 ( .A1(n10460), .A2(n10459), .ZN(n12643) );
  AND2_X2 U11318 ( .A1(n15768), .A2(n15769), .ZN(n9805) );
  AOI221_X2 U11320 ( .B1(n18047), .B2(n10076), .C1(n18063), .C2(n10076), .A(
        n18046), .ZN(n18071) );
  AOI22_X1 U11321 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14912), .B1(n14911), 
        .B2(n20054), .ZN(n15019) );
  XOR2_X2 U11322 ( .A(n11280), .B(n14754), .Z(n16086) );
  NAND2_X2 U11323 ( .A1(n12334), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11938) );
  OR2_X2 U11324 ( .A1(n12936), .A2(n19314), .ZN(n10325) );
  XNOR2_X2 U11325 ( .A(n11226), .B(n11216), .ZN(n13749) );
  NAND2_X2 U11326 ( .A1(n11215), .A2(n11214), .ZN(n11226) );
  NOR2_X2 U11327 ( .A1(n15187), .A2(n15186), .ZN(n15185) );
  NAND2_X2 U11328 ( .A1(n10221), .A2(n10220), .ZN(n12039) );
  NAND2_X2 U11329 ( .A1(n10011), .A2(n10468), .ZN(n10537) );
  OAI21_X2 U11330 ( .B1(n20338), .B2(n11239), .A(n11204), .ZN(n13723) );
  NAND2_X1 U11331 ( .A1(n14515), .A2(n14516), .ZN(n14488) );
  INV_X1 U11332 ( .A(n10012), .ZN(n14515) );
  NOR2_X1 U11333 ( .A1(n17393), .A2(n17387), .ZN(n17383) );
  AND2_X1 U11334 ( .A1(n10619), .A2(n10618), .ZN(n20410) );
  NAND2_X1 U11335 ( .A1(n10303), .A2(n10302), .ZN(n10584) );
  OR2_X1 U11336 ( .A1(n9981), .A2(n9980), .ZN(n17433) );
  NAND2_X1 U11337 ( .A1(n13651), .A2(n13447), .ZN(n20938) );
  AOI221_X1 U11338 ( .B1(n19008), .B2(n15817), .C1(n17541), .C2(n15817), .A(
        n15815), .ZN(n15909) );
  NAND2_X1 U11339 ( .A1(n11950), .A2(n11951), .ZN(n11954) );
  NAND2_X1 U11340 ( .A1(n9956), .A2(n11920), .ZN(n11950) );
  INV_X2 U11342 ( .A(n12501), .ZN(n11863) );
  AOI211_X1 U11343 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n11415), .B(n11414), .ZN(n17471) );
  NOR2_X2 U11344 ( .A1(n20287), .A2(n20281), .ZN(n13939) );
  INV_X1 U11345 ( .A(n10574), .ZN(n10469) );
  NOR2_X1 U11346 ( .A1(n10574), .A2(n10577), .ZN(n10816) );
  INV_X1 U11347 ( .A(n11839), .ZN(n11812) );
  INV_X1 U11348 ( .A(n11837), .ZN(n12174) );
  NAND2_X2 U11349 ( .A1(n9863), .A2(n9838), .ZN(n20274) );
  AND4_X1 U11350 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n9863) );
  AND4_X1 U11351 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10331) );
  AOI22_X1 U11352 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10434) );
  BUF_X2 U11353 ( .A(n9799), .Z(n10945) );
  CLKBUF_X1 U11354 ( .A(n10446), .Z(n11092) );
  INV_X4 U11355 ( .A(n11378), .ZN(n17307) );
  INV_X4 U11356 ( .A(n9858), .ZN(n17117) );
  BUF_X2 U11357 ( .A(n10407), .Z(n11110) );
  BUF_X2 U11358 ( .A(n10488), .Z(n10925) );
  CLKBUF_X2 U11359 ( .A(n11086), .Z(n11116) );
  CLKBUF_X2 U11360 ( .A(n10441), .Z(n11111) );
  BUF_X2 U11361 ( .A(n11117), .Z(n11027) );
  CLKBUF_X2 U11362 ( .A(n10412), .Z(n11087) );
  CLKBUF_X2 U11363 ( .A(n13269), .Z(n13279) );
  CLKBUF_X2 U11364 ( .A(n13869), .Z(n20941) );
  AND2_X2 U11365 ( .A1(n10369), .A2(n10368), .ZN(n10349) );
  INV_X4 U11366 ( .A(n11340), .ZN(n9808) );
  CLKBUF_X2 U11368 ( .A(n10421), .Z(n11028) );
  AND2_X1 U11369 ( .A1(n10322), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10370) );
  AND2_X2 U11370 ( .A1(n10324), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10368) );
  INV_X4 U11371 ( .A(n10328), .ZN(n9810) );
  INV_X1 U11372 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18962) );
  NAND2_X1 U11373 ( .A1(n10286), .A2(n9900), .ZN(n14636) );
  XNOR2_X1 U11374 ( .A(n14690), .B(n14871), .ZN(n14864) );
  NAND2_X1 U11375 ( .A1(n12671), .A2(n12674), .ZN(n14634) );
  AND2_X1 U11376 ( .A1(n14343), .A2(n14327), .ZN(n14655) );
  OAI21_X1 U11377 ( .B1(n15355), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15344), .ZN(n15534) );
  OR2_X1 U11378 ( .A1(n14328), .A2(n12673), .ZN(n12674) );
  AND3_X1 U11379 ( .A1(n10233), .A2(n12577), .A3(n10234), .ZN(n12779) );
  AND2_X1 U11380 ( .A1(n9961), .A2(n9960), .ZN(n15257) );
  AOI21_X1 U11381 ( .B1(n10151), .B2(n10150), .A(n9872), .ZN(n15651) );
  NOR2_X1 U11382 ( .A1(n12893), .A2(n12899), .ZN(n12790) );
  AOI21_X1 U11383 ( .B1(n14408), .B2(n14407), .A(n14406), .ZN(n14702) );
  OR2_X1 U11384 ( .A1(n15404), .A2(n9931), .ZN(n12893) );
  AOI21_X1 U11385 ( .B1(n14645), .B2(n14805), .A(n16036), .ZN(n14661) );
  AND2_X1 U11386 ( .A1(n10273), .A2(n10272), .ZN(n9843) );
  CLKBUF_X1 U11387 ( .A(n14364), .Z(n14365) );
  OR2_X1 U11388 ( .A1(n13216), .A2(n13215), .ZN(n10273) );
  NAND3_X1 U11389 ( .A1(n14704), .A2(n10097), .A3(n10287), .ZN(n14645) );
  NAND2_X1 U11390 ( .A1(n15672), .A2(n15668), .ZN(n15654) );
  NAND2_X1 U11391 ( .A1(n15162), .A2(n9862), .ZN(n13216) );
  NOR2_X2 U11392 ( .A1(n14488), .A2(n10022), .ZN(n9875) );
  INV_X1 U11393 ( .A(n14747), .ZN(n16006) );
  NAND2_X1 U11394 ( .A1(n9951), .A2(n12523), .ZN(n16292) );
  NAND2_X1 U11395 ( .A1(n14780), .A2(n11275), .ZN(n14747) );
  NAND2_X1 U11396 ( .A1(n15169), .A2(n13166), .ZN(n13190) );
  OR2_X1 U11397 ( .A1(n13165), .A2(n13164), .ZN(n13166) );
  OR2_X2 U11398 ( .A1(n14190), .A2(n11274), .ZN(n14780) );
  AND2_X1 U11399 ( .A1(n15179), .A2(n14993), .ZN(n15165) );
  NOR2_X1 U11400 ( .A1(n15183), .A2(n15178), .ZN(n15179) );
  NAND2_X1 U11401 ( .A1(n12443), .A2(n12442), .ZN(n15481) );
  NOR2_X1 U11402 ( .A1(n11285), .A2(n10102), .ZN(n10101) );
  NOR2_X1 U11403 ( .A1(n10774), .A2(n10015), .ZN(n10013) );
  AOI21_X1 U11404 ( .B1(n10300), .B2(n11274), .A(n9930), .ZN(n10299) );
  INV_X1 U11405 ( .A(n10300), .ZN(n10102) );
  AND2_X1 U11406 ( .A1(n10301), .A2(n11275), .ZN(n10300) );
  AND2_X1 U11407 ( .A1(n11435), .A2(n17994), .ZN(n17628) );
  AND2_X1 U11408 ( .A1(n12450), .A2(n9892), .ZN(n9841) );
  AOI211_X1 U11409 ( .C1(n20913), .C2(n20144), .A(n14069), .B(n14068), .ZN(
        n14070) );
  NOR2_X1 U11410 ( .A1(n15207), .A2(n15005), .ZN(n15195) );
  NAND2_X1 U11411 ( .A1(n15218), .A2(n9890), .ZN(n15207) );
  OAI21_X1 U11412 ( .B1(n12447), .B2(n12788), .A(n19152), .ZN(n12449) );
  NAND2_X1 U11413 ( .A1(n12089), .A2(n15741), .ZN(n15747) );
  NOR2_X2 U11414 ( .A1(n15226), .A2(n12389), .ZN(n15218) );
  AND3_X1 U11415 ( .A1(n11430), .A2(n11429), .A3(n11428), .ZN(n17639) );
  NAND2_X1 U11416 ( .A1(n10710), .A2(n10709), .ZN(n14102) );
  NAND2_X1 U11417 ( .A1(n15233), .A2(n15227), .ZN(n15226) );
  NOR2_X1 U11418 ( .A1(n14120), .A2(n14123), .ZN(n14121) );
  AOI21_X1 U11419 ( .B1(n10677), .B2(n10816), .A(n10676), .ZN(n13969) );
  XNOR2_X1 U11420 ( .A(n12092), .B(n12090), .ZN(n12437) );
  AND2_X1 U11421 ( .A1(n12129), .A2(n12090), .ZN(n10057) );
  AOI21_X1 U11422 ( .B1(n11231), .B2(n10816), .A(n10653), .ZN(n13882) );
  AND2_X1 U11423 ( .A1(n12127), .A2(n12126), .ZN(n12129) );
  NAND2_X1 U11424 ( .A1(n10668), .A2(n10095), .ZN(n11266) );
  NAND2_X1 U11425 ( .A1(n13781), .A2(n12995), .ZN(n13834) );
  AND2_X1 U11426 ( .A1(n10645), .A2(n10670), .ZN(n11231) );
  AND2_X1 U11427 ( .A1(n12088), .A2(n12087), .ZN(n12090) );
  NAND2_X1 U11428 ( .A1(n9967), .A2(n9965), .ZN(n13781) );
  NAND2_X1 U11429 ( .A1(n13839), .A2(n13836), .ZN(n13910) );
  NAND2_X1 U11430 ( .A1(n16506), .A2(n18175), .ZN(n18131) );
  AND2_X1 U11431 ( .A1(n12967), .A2(n13780), .ZN(n13789) );
  OR2_X1 U11432 ( .A1(n12992), .A2(n9968), .ZN(n9966) );
  NOR2_X2 U11433 ( .A1(n13840), .A2(n13841), .ZN(n13839) );
  INV_X1 U11434 ( .A(n10089), .ZN(n10293) );
  NAND2_X1 U11435 ( .A1(n12551), .A2(n12566), .ZN(n12519) );
  NAND2_X1 U11436 ( .A1(n13830), .A2(n13831), .ZN(n13840) );
  OAI21_X1 U11437 ( .B1(n11217), .B2(n10580), .A(n10306), .ZN(n13813) );
  NAND2_X1 U11438 ( .A1(n10027), .A2(n10601), .ZN(n10089) );
  OR2_X1 U11439 ( .A1(n12991), .A2(n12966), .ZN(n12967) );
  NAND2_X1 U11440 ( .A1(n11981), .A2(n11973), .ZN(n12055) );
  NOR2_X1 U11441 ( .A1(n13805), .A2(n13806), .ZN(n13830) );
  AND2_X1 U11442 ( .A1(n13506), .A2(n12985), .ZN(n13664) );
  OR2_X1 U11443 ( .A1(n12525), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U11444 ( .A1(n12965), .A2(n12964), .ZN(n12991) );
  AND2_X1 U11445 ( .A1(n12517), .A2(n12516), .ZN(n12529) );
  INV_X1 U11446 ( .A(n20410), .ZN(n10292) );
  NAND2_X1 U11447 ( .A1(n10584), .A2(n10541), .ZN(n10600) );
  NAND2_X1 U11448 ( .A1(n10584), .A2(n10583), .ZN(n20339) );
  NOR2_X1 U11449 ( .A1(n20417), .A2(n20288), .ZN(n20797) );
  NOR2_X1 U11450 ( .A1(n20417), .A2(n20303), .ZN(n20817) );
  NOR2_X1 U11451 ( .A1(n20417), .A2(n20231), .ZN(n20826) );
  NOR2_X1 U11452 ( .A1(n20417), .A2(n20295), .ZN(n20811) );
  NOR2_X1 U11453 ( .A1(n20417), .A2(n20227), .ZN(n20806) );
  NOR2_X1 U11454 ( .A1(n20417), .A2(n20283), .ZN(n20791) );
  NOR2_X1 U11455 ( .A1(n20417), .A2(n20276), .ZN(n20785) );
  NOR2_X1 U11456 ( .A1(n20417), .A2(n20267), .ZN(n20773) );
  NAND2_X1 U11457 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17427), .ZN(n17426) );
  AND2_X1 U11458 ( .A1(n12469), .A2(n10111), .ZN(n12517) );
  NAND2_X1 U11459 ( .A1(n12976), .A2(n12975), .ZN(n12982) );
  NOR2_X2 U11460 ( .A1(n17433), .A2(n17609), .ZN(n17427) );
  OR2_X1 U11461 ( .A1(n16452), .A2(n12974), .ZN(n11979) );
  NOR2_X1 U11462 ( .A1(n17192), .A2(n17176), .ZN(n17156) );
  NAND2_X1 U11463 ( .A1(n9955), .A2(n11924), .ZN(n10257) );
  OR2_X2 U11464 ( .A1(n13650), .A2(n12641), .ZN(n13651) );
  NAND2_X1 U11465 ( .A1(n10294), .A2(n10507), .ZN(n9976) );
  OR2_X1 U11466 ( .A1(n15909), .A2(n15908), .ZN(n9979) );
  AND2_X1 U11467 ( .A1(n11193), .A2(n11192), .ZN(n13686) );
  NOR2_X2 U11468 ( .A1(n19336), .A2(n19786), .ZN(n19337) );
  NOR2_X2 U11469 ( .A1(n19332), .A2(n19786), .ZN(n19333) );
  NOR2_X2 U11470 ( .A1(n19323), .A2(n19786), .ZN(n19324) );
  NOR2_X1 U11471 ( .A1(n17226), .A2(n17225), .ZN(n17222) );
  AND2_X1 U11472 ( .A1(n10537), .A2(n10536), .ZN(n10539) );
  OR2_X1 U11473 ( .A1(n12453), .A2(n12785), .ZN(n12566) );
  NAND2_X1 U11474 ( .A1(n11908), .A2(n11909), .ZN(n11951) );
  AND2_X1 U11475 ( .A1(n11899), .A2(n11898), .ZN(n11922) );
  INV_X2 U11476 ( .A(n13360), .ZN(n19263) );
  AOI21_X1 U11477 ( .B1(n11931), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11945), .ZN(n12343) );
  NOR2_X1 U11478 ( .A1(n11919), .A2(n11918), .ZN(n11920) );
  AOI21_X1 U11479 ( .B1(n11931), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11932), .ZN(n11946) );
  NAND2_X1 U11480 ( .A1(n10139), .A2(n11913), .ZN(n11931) );
  NAND2_X1 U11481 ( .A1(n11885), .A2(n15773), .ZN(n12334) );
  NAND2_X2 U11482 ( .A1(n19008), .A2(n17542), .ZN(n17608) );
  NAND2_X1 U11483 ( .A1(n10005), .A2(n10004), .ZN(n17934) );
  CLKBUF_X1 U11484 ( .A(n11901), .Z(n15755) );
  OR2_X1 U11485 ( .A1(n17954), .A2(n17955), .ZN(n10006) );
  NOR2_X1 U11486 ( .A1(n11883), .A2(n11882), .ZN(n11901) );
  INV_X1 U11487 ( .A(n11865), .ZN(n11886) );
  CLKBUF_X1 U11488 ( .A(n11877), .Z(n13351) );
  NAND2_X1 U11489 ( .A1(n12170), .A2(n11896), .ZN(n11913) );
  NOR2_X1 U11490 ( .A1(n14922), .A2(n15011), .ZN(n14943) );
  AND2_X1 U11491 ( .A1(n11891), .A2(n11892), .ZN(n11916) );
  AND2_X1 U11492 ( .A1(n11895), .A2(n11894), .ZN(n12170) );
  NAND2_X1 U11493 ( .A1(n11557), .A2(n17351), .ZN(n11533) );
  AND2_X1 U11494 ( .A1(n11359), .A2(n11358), .ZN(n17483) );
  OR2_X1 U11495 ( .A1(n13573), .A2(n13792), .ZN(n13705) );
  AOI211_X1 U11496 ( .C1(n11448), .C2(n11447), .A(n11553), .B(n11551), .ZN(
        n18772) );
  INV_X1 U11497 ( .A(n11848), .ZN(n11864) );
  NAND2_X1 U11498 ( .A1(n11329), .A2(n10332), .ZN(n17496) );
  NAND2_X1 U11499 ( .A1(n11765), .A2(n11808), .ZN(n16465) );
  INV_X1 U11500 ( .A(n18337), .ZN(n17351) );
  INV_X1 U11501 ( .A(n10470), .ZN(n14035) );
  NAND2_X1 U11502 ( .A1(n11847), .A2(n11838), .ZN(n11848) );
  AND3_X2 U11503 ( .A1(n11878), .A2(n11743), .A3(n10326), .ZN(n11873) );
  NOR2_X1 U11504 ( .A1(n9948), .A2(n11851), .ZN(n11814) );
  NAND2_X1 U11505 ( .A1(n20055), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20061) );
  AOI211_X2 U11506 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n11498), .B(n11497), .ZN(n18337) );
  NAND3_X1 U11507 ( .A1(n11345), .A2(n11344), .A3(n11343), .ZN(n17978) );
  AND2_X1 U11508 ( .A1(n10458), .A2(n13566), .ZN(n13698) );
  NAND2_X1 U11509 ( .A1(n9801), .A2(n9842), .ZN(n10017) );
  NAND2_X2 U11510 ( .A1(n10216), .A2(n10214), .ZN(n20055) );
  AND3_X1 U11511 ( .A1(n11328), .A2(n11327), .A3(n11326), .ZN(n10332) );
  INV_X2 U11512 ( .A(n12174), .ZN(n12785) );
  AOI211_X1 U11513 ( .C1(n9804), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n11335), .B(n11334), .ZN(n11345) );
  NOR2_X1 U11514 ( .A1(n11338), .A2(n11337), .ZN(n11344) );
  NAND2_X2 U11515 ( .A1(n10352), .A2(n10354), .ZN(n10574) );
  OR2_X2 U11516 ( .A1(n16581), .A2(n16533), .ZN(n16583) );
  AND2_X2 U11517 ( .A1(n10404), .A2(n10353), .ZN(n14162) );
  NAND2_X2 U11518 ( .A1(n10331), .A2(n10351), .ZN(n20281) );
  AND4_X1 U11519 ( .A1(n10382), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        n10352) );
  NAND2_X1 U11520 ( .A1(n10146), .A2(n10145), .ZN(n11837) );
  AND4_X1 U11521 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10404) );
  INV_X1 U11522 ( .A(n17219), .ZN(n17292) );
  AND4_X1 U11523 ( .A1(n10367), .A2(n10366), .A3(n10365), .A4(n10364), .ZN(
        n10376) );
  AND4_X1 U11524 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10378) );
  INV_X1 U11525 ( .A(n15772), .ZN(n9811) );
  AND2_X2 U11526 ( .A1(n13258), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11781) );
  AND2_X2 U11527 ( .A1(n13225), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11783) );
  NAND2_X1 U11528 ( .A1(n10008), .A2(n11302), .ZN(n17219) );
  NAND2_X2 U11529 ( .A1(n19020), .A2(n11561), .ZN(n16515) );
  OR2_X1 U11530 ( .A1(n11311), .A2(n11307), .ZN(n9858) );
  INV_X2 U11531 ( .A(n16619), .ZN(n16621) );
  OR2_X2 U11532 ( .A1(n11307), .A2(n11310), .ZN(n10327) );
  INV_X2 U11533 ( .A(n20068), .ZN(n20071) );
  BUF_X4 U11534 ( .A(n10431), .Z(n9812) );
  AND2_X2 U11535 ( .A1(n13578), .A2(n13942), .ZN(n10488) );
  AND2_X1 U11536 ( .A1(n10576), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10369) );
  AND2_X2 U11537 ( .A1(n10010), .A2(n10009), .ZN(n13942) );
  NAND2_X1 U11538 ( .A1(n18962), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U11539 ( .A1(n18972), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11310) );
  NAND2_X1 U11540 ( .A1(n18987), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11308) );
  NAND3_X1 U11541 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18980), .ZN(n11312) );
  NOR2_X1 U11542 ( .A1(n19286), .A2(n10185), .ZN(n10184) );
  NAND2_X1 U11543 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18802) );
  NAND2_X1 U11544 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11307) );
  NOR2_X4 U11545 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13578) );
  INV_X2 U11546 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15769) );
  CLKBUF_X1 U11548 ( .A(n19273), .Z(n9813) );
  NAND2_X1 U11549 ( .A1(n12429), .A2(n14012), .ZN(n19273) );
  AND2_X1 U11550 ( .A1(n14959), .A2(n14958), .ZN(n15496) );
  AND2_X2 U11551 ( .A1(n11955), .A2(n11954), .ZN(n12974) );
  NAND2_X1 U11552 ( .A1(n10263), .A2(n9975), .ZN(n10265) );
  NAND3_X2 U11553 ( .A1(n9800), .A2(n10437), .A3(n9831), .ZN(n10155) );
  NAND2_X1 U11554 ( .A1(n9949), .A2(n9950), .ZN(n12092) );
  NAND2_X1 U11555 ( .A1(n11815), .A2(n9802), .ZN(n11846) );
  XNOR2_X1 U11556 ( .A(n11954), .B(n11959), .ZN(n16452) );
  OR2_X2 U11557 ( .A1(n11965), .A2(n11984), .ZN(n12058) );
  AOI21_X1 U11558 ( .B1(n10235), .B2(n10238), .A(n15329), .ZN(n15331) );
  AND2_X4 U11559 ( .A1(n10368), .A2(n13941), .ZN(n10446) );
  AOI211_X2 U11560 ( .C1(n19282), .C2(n19098), .A(n16278), .B(n16277), .ZN(
        n16279) );
  NAND2_X2 U11561 ( .A1(n12835), .A2(n13504), .ZN(n12208) );
  NAND2_X4 U11562 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18794), .ZN(
        n11489) );
  AND2_X2 U11564 ( .A1(n14364), .A2(n14367), .ZN(n14352) );
  AND2_X1 U11565 ( .A1(n14404), .A2(n10309), .ZN(n14364) );
  NAND2_X1 U11566 ( .A1(n15481), .A2(n15482), .ZN(n9814) );
  CLKBUF_X1 U11567 ( .A(n14011), .Z(n9815) );
  INV_X1 U11568 ( .A(n16439), .ZN(n9816) );
  OAI21_X1 U11569 ( .B1(n15455), .B2(n15456), .A(n12541), .ZN(n9817) );
  NAND2_X1 U11570 ( .A1(n15481), .A2(n15482), .ZN(n12451) );
  NAND2_X1 U11571 ( .A1(n10643), .A2(n10620), .ZN(n9818) );
  CLKBUF_X1 U11572 ( .A(n14138), .Z(n9819) );
  NOR2_X1 U11573 ( .A1(n14762), .A2(n14759), .ZN(n9820) );
  OAI21_X1 U11574 ( .B1(n16006), .B2(n14770), .A(n14748), .ZN(n9821) );
  AND2_X1 U11575 ( .A1(n13942), .A2(n13612), .ZN(n9822) );
  INV_X1 U11576 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9823) );
  NAND2_X1 U11577 ( .A1(n10643), .A2(n10620), .ZN(n20520) );
  OAI21_X1 U11578 ( .B1(n16006), .B2(n14770), .A(n14748), .ZN(n15993) );
  OR2_X2 U11579 ( .A1(n11965), .A2(n11979), .ZN(n19471) );
  NOR2_X2 U11580 ( .A1(n14630), .A2(n14629), .ZN(n14631) );
  NOR2_X2 U11581 ( .A1(n15982), .A2(n14752), .ZN(n15986) );
  INV_X1 U11582 ( .A(n11938), .ZN(n11939) );
  OR2_X1 U11583 ( .A1(n11938), .A2(n13531), .ZN(n11929) );
  MUX2_X2 U11584 ( .A(n9820), .B(n15986), .S(n14753), .Z(n14754) );
  OAI21_X1 U11585 ( .B1(n15373), .B2(n15369), .A(n15370), .ZN(n15359) );
  NAND2_X1 U11586 ( .A1(n15373), .A2(n15370), .ZN(n10235) );
  NAND2_X2 U11587 ( .A1(n11273), .A2(n11272), .ZN(n14190) );
  NAND2_X1 U11588 ( .A1(n11238), .A2(n11237), .ZN(n14075) );
  AND4_X1 U11589 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n10377) );
  OAI21_X1 U11590 ( .B1(n12640), .B2(n12861), .A(n13705), .ZN(n10462) );
  NAND2_X4 U11591 ( .A1(n9944), .A2(n12169), .ZN(n11897) );
  XNOR2_X2 U11592 ( .A(n12039), .B(n10219), .ZN(n19274) );
  OAI21_X2 U11593 ( .B1(n15397), .B2(n15396), .A(n15395), .ZN(n15439) );
  NAND2_X2 U11594 ( .A1(n10534), .A2(n10467), .ZN(n10544) );
  BUF_X4 U11595 ( .A(n11643), .Z(n13258) );
  AND2_X2 U11596 ( .A1(n11852), .A2(n11839), .ZN(n10326) );
  NAND2_X4 U11597 ( .A1(n11730), .A2(n11729), .ZN(n11852) );
  OAI21_X2 U11598 ( .B1(n12451), .B2(n9864), .A(n10067), .ZN(n15696) );
  OAI21_X1 U11599 ( .B1(n12414), .B2(n14015), .A(n12036), .ZN(n19276) );
  NAND2_X2 U11600 ( .A1(n10062), .A2(n10064), .ZN(n15382) );
  OAI21_X2 U11601 ( .B1(n11250), .B2(n10285), .A(n10283), .ZN(n16016) );
  XNOR2_X2 U11602 ( .A(n13725), .B(n11212), .ZN(n13672) );
  OAI21_X2 U11603 ( .B1(n13692), .B2(n10462), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10534) );
  OAI21_X2 U11604 ( .B1(n12640), .B2(n12878), .A(n12643), .ZN(n13692) );
  OAI21_X1 U11605 ( .B1(n10591), .B2(n10297), .A(n10295), .ZN(n10530) );
  OAI21_X2 U11606 ( .B1(n15455), .B2(n15456), .A(n12541), .ZN(n15397) );
  OAI21_X2 U11607 ( .B1(n15654), .B2(n12496), .A(n15653), .ZN(n15455) );
  AND2_X4 U11608 ( .A1(n10370), .A2(n10368), .ZN(n10431) );
  NAND2_X1 U11609 ( .A1(n15669), .A2(n15667), .ZN(n15672) );
  OAI21_X2 U11610 ( .B1(n16292), .B2(n12483), .A(n16290), .ZN(n15669) );
  INV_X1 U11611 ( .A(n10432), .ZN(n9826) );
  INV_X1 U11612 ( .A(n10432), .ZN(n9827) );
  NAND2_X2 U11613 ( .A1(n13942), .A2(n10363), .ZN(n10432) );
  AND3_X4 U11614 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n11600), .ZN(n11748) );
  NAND2_X1 U11615 ( .A1(n10293), .A2(n10644), .ZN(n10670) );
  NOR2_X1 U11616 ( .A1(n20410), .A2(n10339), .ZN(n10644) );
  AND2_X1 U11617 ( .A1(n10528), .A2(n10527), .ZN(n10529) );
  NOR2_X1 U11618 ( .A1(n10274), .A2(n9896), .ZN(n9964) );
  AOI21_X1 U11619 ( .B1(n15813), .B2(n18772), .A(n13763), .ZN(n15907) );
  AOI21_X1 U11621 ( .B1(n13568), .B2(n13624), .A(n13698), .ZN(n10475) );
  NOR2_X1 U11622 ( .A1(n9806), .A2(n17351), .ZN(n11548) );
  NAND2_X1 U11623 ( .A1(n18314), .A2(n17393), .ZN(n11532) );
  NAND2_X1 U11624 ( .A1(n16629), .A2(n11543), .ZN(n15809) );
  NOR2_X1 U11625 ( .A1(n14342), .A2(n10321), .ZN(n10320) );
  INV_X1 U11626 ( .A(n14353), .ZN(n10321) );
  OR2_X1 U11627 ( .A1(n10024), .A2(n14460), .ZN(n10022) );
  INV_X1 U11628 ( .A(n11128), .ZN(n11102) );
  INV_X1 U11629 ( .A(n10600), .ZN(n10027) );
  AND3_X1 U11630 ( .A1(n12957), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20060), 
        .ZN(n13160) );
  INV_X1 U11631 ( .A(n13160), .ZN(n13213) );
  INV_X1 U11632 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10229) );
  OR2_X1 U11633 ( .A1(n12544), .A2(n15412), .ZN(n12545) );
  INV_X1 U11634 ( .A(n15464), .ZN(n10148) );
  INV_X1 U11635 ( .A(n12326), .ZN(n12298) );
  NAND2_X1 U11636 ( .A1(n12188), .A2(n12174), .ZN(n12326) );
  NOR2_X1 U11637 ( .A1(n11800), .A2(n11698), .ZN(n13347) );
  AND2_X1 U11638 ( .A1(n11697), .A2(n11696), .ZN(n11698) );
  INV_X1 U11639 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14248) );
  NOR2_X1 U11640 ( .A1(n11556), .A2(n18790), .ZN(n11541) );
  INV_X1 U11641 ( .A(n9803), .ZN(n11556) );
  INV_X1 U11642 ( .A(n15810), .ZN(n17502) );
  AOI21_X1 U11643 ( .B1(n15809), .B2(n18839), .A(n19006), .ZN(n15810) );
  NAND4_X1 U11644 ( .A1(n11544), .A2(n18337), .A3(n11531), .A4(n17503), .ZN(
        n17541) );
  AND2_X1 U11645 ( .A1(n10577), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11132) );
  NAND2_X1 U11646 ( .A1(n10530), .A2(n10527), .ZN(n10305) );
  NAND2_X1 U11647 ( .A1(n10018), .A2(n10540), .ZN(n11205) );
  AND2_X1 U11648 ( .A1(n12566), .A2(n14979), .ZN(n12787) );
  INV_X1 U11649 ( .A(n13886), .ZN(n10191) );
  NAND2_X1 U11650 ( .A1(n15165), .A2(n10123), .ZN(n12895) );
  NOR2_X1 U11651 ( .A1(n10126), .A2(n10124), .ZN(n10123) );
  OR2_X1 U11652 ( .A1(n10127), .A2(n15154), .ZN(n10126) );
  NAND2_X1 U11653 ( .A1(n10125), .A2(n15164), .ZN(n10124) );
  NAND2_X1 U11654 ( .A1(n12997), .A2(n10275), .ZN(n10274) );
  INV_X1 U11655 ( .A(n10276), .ZN(n10275) );
  AND2_X1 U11656 ( .A1(n19217), .A2(n14130), .ZN(n14131) );
  AND2_X1 U11657 ( .A1(n10277), .A2(n14176), .ZN(n9971) );
  AND2_X1 U11658 ( .A1(n10279), .A2(n10278), .ZN(n10277) );
  INV_X1 U11659 ( .A(n15203), .ZN(n10278) );
  NAND2_X1 U11660 ( .A1(n12344), .A2(n12343), .ZN(n12345) );
  NOR2_X1 U11661 ( .A1(n12889), .A2(n10226), .ZN(n10107) );
  INV_X1 U11662 ( .A(n10226), .ZN(n10109) );
  NAND2_X1 U11663 ( .A1(n15355), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15344) );
  INV_X1 U11664 ( .A(n15404), .ZN(n10259) );
  AND2_X1 U11665 ( .A1(n11832), .A2(n13493), .ZN(n12502) );
  NOR2_X1 U11666 ( .A1(n11693), .A2(n20061), .ZN(n11694) );
  INV_X1 U11667 ( .A(n11800), .ZN(n11693) );
  INV_X1 U11668 ( .A(n17432), .ZN(n9980) );
  OAI211_X1 U11669 ( .C1(n17172), .C2(n17241), .A(n11528), .B(n11527), .ZN(
        n13762) );
  XNOR2_X1 U11670 ( .A(n12895), .B(n12894), .ZN(n16211) );
  NAND2_X1 U11671 ( .A1(n11145), .A2(n11144), .ZN(n11150) );
  NOR2_X1 U11672 ( .A1(n14752), .A2(n11277), .ZN(n10301) );
  OR2_X1 U11673 ( .A1(n10640), .A2(n10639), .ZN(n11241) );
  NOR2_X1 U11674 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n11147), .ZN(
        n11180) );
  OR2_X1 U11675 ( .A1(n10617), .A2(n10616), .ZN(n11201) );
  AND2_X1 U11676 ( .A1(n10112), .A2(n12411), .ZN(n10111) );
  NAND2_X1 U11677 ( .A1(n10106), .A2(n10105), .ZN(n12400) );
  NAND2_X1 U11678 ( .A1(n12501), .A2(n11683), .ZN(n10105) );
  NAND2_X1 U11679 ( .A1(n12025), .A2(n11863), .ZN(n10106) );
  AND4_X1 U11680 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12149) );
  AND2_X1 U11681 ( .A1(n11630), .A2(n11629), .ZN(n11687) );
  NAND2_X1 U11682 ( .A1(n12956), .A2(n13549), .ZN(n11972) );
  NOR2_X1 U11683 ( .A1(n11851), .A2(n11820), .ZN(n11743) );
  OR2_X1 U11684 ( .A1(n11362), .A2(n17483), .ZN(n11375) );
  NOR4_X1 U11685 ( .A1(n18790), .A2(n13762), .A3(n11532), .A4(n11533), .ZN(
        n11539) );
  AOI21_X1 U11686 ( .B1(n18821), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11437), .ZN(n11443) );
  OAI22_X1 U11687 ( .A1(n18972), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18826), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11442) );
  NOR2_X1 U11688 ( .A1(n11557), .A2(n11556), .ZN(n11545) );
  OAI211_X1 U11689 ( .C1(n17296), .C2(n14243), .A(n10087), .B(n10086), .ZN(
        n10085) );
  NAND2_X1 U11690 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10087) );
  NAND2_X1 U11691 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10086) );
  NOR2_X1 U11692 ( .A1(n18350), .A2(n18327), .ZN(n11544) );
  AND2_X1 U11693 ( .A1(n10311), .A2(n10310), .ZN(n10309) );
  INV_X1 U11694 ( .A(n14379), .ZN(n10310) );
  INV_X1 U11695 ( .A(n10314), .ZN(n10313) );
  INV_X1 U11696 ( .A(n14525), .ZN(n10016) );
  NAND2_X1 U11697 ( .A1(n10698), .A2(n10671), .ZN(n11240) );
  AND2_X1 U11698 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10649), .ZN(
        n10673) );
  CLKBUF_X1 U11699 ( .A(n10621), .Z(n11104) );
  AOI21_X1 U11700 ( .B1(n14729), .B2(n10291), .A(n16053), .ZN(n10290) );
  INV_X1 U11701 ( .A(n11290), .ZN(n10291) );
  NAND2_X1 U11702 ( .A1(n14739), .A2(n10099), .ZN(n10097) );
  AND2_X1 U11703 ( .A1(n14740), .A2(n10290), .ZN(n10099) );
  NAND2_X1 U11704 ( .A1(n10290), .A2(n14751), .ZN(n10287) );
  NOR2_X1 U11705 ( .A1(n10170), .A2(n14518), .ZN(n10169) );
  INV_X1 U11706 ( .A(n14495), .ZN(n10170) );
  AND2_X1 U11707 ( .A1(n13566), .A2(n13709), .ZN(n12758) );
  NOR2_X1 U11708 ( .A1(n10699), .A2(n10096), .ZN(n10095) );
  AND2_X1 U11709 ( .A1(n16169), .A2(n14110), .ZN(n10172) );
  INV_X1 U11710 ( .A(n11249), .ZN(n10284) );
  NAND2_X1 U11711 ( .A1(n12771), .A2(n13709), .ZN(n12745) );
  INV_X1 U11712 ( .A(n13753), .ZN(n10162) );
  OR2_X1 U11713 ( .A1(n10505), .A2(n10504), .ZN(n11207) );
  INV_X1 U11714 ( .A(n11267), .ZN(n10522) );
  AND2_X1 U11715 ( .A1(n10589), .A2(n10296), .ZN(n10295) );
  INV_X1 U11716 ( .A(n10570), .ZN(n11264) );
  NAND2_X1 U11717 ( .A1(n14162), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10570) );
  NAND2_X1 U11718 ( .A1(n10607), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11176) );
  OR2_X1 U11719 ( .A1(n10534), .A2(n10543), .ZN(n10556) );
  XNOR2_X1 U11720 ( .A(n10535), .B(n10534), .ZN(n20378) );
  AND2_X1 U11721 ( .A1(n11633), .A2(n11632), .ZN(n11636) );
  NAND2_X1 U11722 ( .A1(n12572), .A2(n12571), .ZN(n14981) );
  NOR2_X1 U11723 ( .A1(n13215), .A2(n10272), .ZN(n10268) );
  AOI21_X1 U11724 ( .B1(n13110), .B2(n10264), .A(n9916), .ZN(n10263) );
  NAND2_X1 U11725 ( .A1(n15185), .A2(n10264), .ZN(n9975) );
  INV_X1 U11726 ( .A(n14995), .ZN(n10200) );
  NAND2_X1 U11727 ( .A1(n10196), .A2(n10195), .ZN(n10194) );
  INV_X1 U11728 ( .A(n15297), .ZN(n10195) );
  INV_X1 U11729 ( .A(n15026), .ZN(n10196) );
  AND2_X1 U11730 ( .A1(n13043), .A2(n15216), .ZN(n10279) );
  INV_X1 U11731 ( .A(n12798), .ZN(n12621) );
  NOR2_X1 U11732 ( .A1(n15024), .A2(n10130), .ZN(n10129) );
  INV_X1 U11733 ( .A(n15217), .ZN(n10130) );
  INV_X1 U11734 ( .A(n10242), .ZN(n10069) );
  INV_X1 U11735 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10185) );
  NAND2_X1 U11736 ( .A1(n15373), .A2(n10236), .ZN(n10231) );
  AND2_X1 U11737 ( .A1(n15370), .A2(n10240), .ZN(n10236) );
  OR2_X1 U11738 ( .A1(n10238), .A2(n10237), .ZN(n10232) );
  OR2_X1 U11739 ( .A1(n10136), .A2(n10135), .ZN(n10134) );
  INV_X1 U11740 ( .A(n13999), .ZN(n10135) );
  NAND2_X1 U11741 ( .A1(n12369), .A2(n13896), .ZN(n10136) );
  OR2_X1 U11742 ( .A1(n10212), .A2(n15080), .ZN(n10211) );
  NAND2_X1 U11743 ( .A1(n10213), .A2(n13557), .ZN(n10212) );
  INV_X1 U11744 ( .A(n13553), .ZN(n10213) );
  NOR2_X1 U11745 ( .A1(n15702), .A2(n10244), .ZN(n10243) );
  INV_X1 U11746 ( .A(n12461), .ZN(n10244) );
  BUF_X1 U11747 ( .A(n12360), .Z(n12793) );
  OR2_X1 U11748 ( .A1(n12154), .A2(n12153), .ZN(n12160) );
  NOR2_X1 U11749 ( .A1(n12125), .A2(n12124), .ZN(n12404) );
  INV_X1 U11750 ( .A(n12038), .ZN(n10221) );
  NAND2_X1 U11751 ( .A1(n10142), .A2(n12026), .ZN(n12037) );
  OR2_X1 U11752 ( .A1(n11834), .A2(n11833), .ZN(n15770) );
  NAND2_X1 U11753 ( .A1(n12973), .A2(n12972), .ZN(n12988) );
  NAND2_X1 U11754 ( .A1(n11723), .A2(n11619), .ZN(n11730) );
  NOR2_X1 U11755 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11301) );
  INV_X1 U11756 ( .A(n9806), .ZN(n11557) );
  NOR2_X1 U11757 ( .A1(n17779), .A2(n17988), .ZN(n11432) );
  AND2_X1 U11758 ( .A1(n11434), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10254) );
  NOR2_X1 U11759 ( .A1(n11433), .A2(n11432), .ZN(n10255) );
  NOR2_X1 U11760 ( .A1(n9992), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9991) );
  INV_X1 U11761 ( .A(n10346), .ZN(n9992) );
  XNOR2_X1 U11762 ( .A(n11362), .B(n11360), .ZN(n11361) );
  INV_X1 U11763 ( .A(n17483), .ZN(n11360) );
  INV_X1 U11764 ( .A(n17496), .ZN(n11572) );
  XNOR2_X1 U11765 ( .A(n17496), .B(n11317), .ZN(n11347) );
  AND2_X1 U11766 ( .A1(n11530), .A2(n11529), .ZN(n9988) );
  INV_X1 U11767 ( .A(n18327), .ZN(n18790) );
  NAND2_X1 U11768 ( .A1(n15809), .A2(n17541), .ZN(n18788) );
  NOR2_X1 U11769 ( .A1(n10463), .A2(n12849), .ZN(n13597) );
  NOR2_X1 U11770 ( .A1(n20938), .A2(n12854), .ZN(n20117) );
  INV_X1 U11771 ( .A(n10474), .ZN(n10482) );
  INV_X1 U11772 ( .A(n13686), .ZN(n13678) );
  AND2_X1 U11773 ( .A1(n14659), .A2(n10621), .ZN(n11058) );
  NAND2_X1 U11774 ( .A1(n14352), .A2(n14353), .ZN(n14341) );
  NAND2_X1 U11775 ( .A1(n10288), .A2(n14751), .ZN(n14704) );
  NAND2_X1 U11776 ( .A1(n10673), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10693) );
  AOI21_X1 U11777 ( .B1(n10581), .B2(n10308), .A(n10307), .ZN(n10306) );
  INV_X1 U11778 ( .A(n10599), .ZN(n10307) );
  INV_X1 U11779 ( .A(n13862), .ZN(n13563) );
  INV_X1 U11780 ( .A(n13709), .ZN(n12857) );
  NOR3_X1 U11781 ( .A1(n9857), .A2(n10163), .A3(n14330), .ZN(n14332) );
  OR2_X1 U11782 ( .A1(n13714), .A2(n13703), .ZN(n16070) );
  OR3_X1 U11783 ( .A1(n15958), .A2(n14903), .A3(n14527), .ZN(n14528) );
  NOR2_X1 U11784 ( .A1(n16147), .A2(n14185), .ZN(n15960) );
  NOR2_X1 U11785 ( .A1(n14097), .A2(n14096), .ZN(n16170) );
  AND2_X2 U11786 ( .A1(n20274), .A2(n10155), .ZN(n13709) );
  AND2_X1 U11787 ( .A1(n12771), .A2(n12704), .ZN(n13862) );
  INV_X1 U11788 ( .A(n11205), .ZN(n10302) );
  NAND2_X1 U11789 ( .A1(n13602), .A2(n13601), .ZN(n15846) );
  INV_X1 U11790 ( .A(n20074), .ZN(n13690) );
  NOR2_X1 U11791 ( .A1(n20417), .A2(n20654), .ZN(n20584) );
  OR2_X1 U11792 ( .A1(n20339), .A2(n20338), .ZN(n20703) );
  NAND2_X1 U11793 ( .A1(n20339), .A2(n14150), .ZN(n20626) );
  NAND2_X1 U11794 ( .A1(n11217), .A2(n10292), .ZN(n20777) );
  NOR2_X1 U11795 ( .A1(n12169), .A2(n16438), .ZN(n13397) );
  AND2_X1 U11796 ( .A1(n12519), .A2(n9852), .ZN(n12565) );
  NAND2_X1 U11797 ( .A1(n12519), .A2(n9906), .ZN(n12559) );
  AND2_X1 U11798 ( .A1(n12471), .A2(n12470), .ZN(n15052) );
  INV_X1 U11799 ( .A(n19183), .ZN(n19134) );
  NAND2_X1 U11800 ( .A1(n9966), .A2(n12993), .ZN(n9965) );
  NAND2_X1 U11801 ( .A1(n10273), .A2(n10271), .ZN(n15159) );
  AND2_X1 U11802 ( .A1(n13109), .A2(n13137), .ZN(n13110) );
  INV_X1 U11803 ( .A(n15230), .ZN(n9962) );
  NAND2_X1 U11804 ( .A1(n15218), .A2(n10129), .ZN(n15205) );
  NAND2_X1 U11805 ( .A1(n10042), .A2(n10258), .ZN(n10041) );
  AND2_X1 U11806 ( .A1(n9914), .A2(n10121), .ZN(n13797) );
  NAND2_X1 U11807 ( .A1(n12783), .A2(n10109), .ZN(n10108) );
  NOR2_X1 U11808 ( .A1(n12890), .A2(n12888), .ZN(n10224) );
  XNOR2_X1 U11809 ( .A(n12789), .B(n14912), .ZN(n10226) );
  INV_X1 U11810 ( .A(n9951), .ZN(n12548) );
  INV_X1 U11811 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9941) );
  OAI21_X1 U11812 ( .B1(n10147), .B2(n10051), .A(n9928), .ZN(n9943) );
  AND2_X1 U11813 ( .A1(n15231), .A2(n14090), .ZN(n15233) );
  AND2_X1 U11814 ( .A1(n12300), .A2(n12299), .ZN(n15037) );
  AND2_X1 U11815 ( .A1(n10245), .A2(n10243), .ZN(n16325) );
  OR2_X1 U11816 ( .A1(n12473), .A2(n15707), .ZN(n16309) );
  NAND2_X1 U11817 ( .A1(n15463), .A2(n12162), .ZN(n12508) );
  NAND2_X1 U11818 ( .A1(n10052), .A2(n10147), .ZN(n15463) );
  NAND2_X1 U11819 ( .A1(n12159), .A2(n10045), .ZN(n10052) );
  INV_X1 U11820 ( .A(n15712), .ZN(n10045) );
  NAND2_X1 U11821 ( .A1(n15712), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15713) );
  AND2_X1 U11822 ( .A1(n12788), .A2(n12298), .ZN(n12233) );
  XNOR2_X1 U11823 ( .A(n12988), .B(n12986), .ZN(n13663) );
  AND2_X1 U11824 ( .A1(n12221), .A2(n12220), .ZN(n13886) );
  NOR2_X2 U11825 ( .A1(n11846), .A2(n9945), .ZN(n11876) );
  NAND2_X1 U11826 ( .A1(n11847), .A2(n9948), .ZN(n9945) );
  NAND2_X1 U11827 ( .A1(n12974), .A2(n12978), .ZN(n12976) );
  INV_X1 U11828 ( .A(n16495), .ZN(n13493) );
  NAND2_X1 U11829 ( .A1(n19987), .A2(n19586), .ZN(n19559) );
  NAND2_X1 U11830 ( .A1(n20015), .A2(n19994), .ZN(n19624) );
  NAND2_X1 U11831 ( .A1(n9865), .A2(n10344), .ZN(n10144) );
  OR2_X1 U11832 ( .A1(n19987), .A2(n20031), .ZN(n19755) );
  OAI21_X2 U11833 ( .B1(n19995), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12628), 
        .ZN(n19836) );
  INV_X1 U11834 ( .A(n20007), .ZN(n20002) );
  INV_X1 U11835 ( .A(n19836), .ZN(n19786) );
  NOR2_X1 U11836 ( .A1(n19008), .A2(n17503), .ZN(n11543) );
  NOR2_X1 U11837 ( .A1(n10074), .A2(n10077), .ZN(n10073) );
  INV_X1 U11838 ( .A(n18772), .ZN(n10077) );
  INV_X1 U11839 ( .A(n10075), .ZN(n10074) );
  OR2_X1 U11840 ( .A1(n16715), .A2(n16894), .ZN(n10038) );
  XOR2_X1 U11841 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n12924), .Z(
        n16985) );
  INV_X1 U11842 ( .A(n11516), .ZN(n9984) );
  OR2_X1 U11843 ( .A1(n11517), .A2(n9986), .ZN(n9985) );
  NAND2_X1 U11844 ( .A1(n9987), .A2(n9870), .ZN(n9986) );
  INV_X1 U11845 ( .A(n11311), .ZN(n10008) );
  INV_X1 U11846 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17120) );
  INV_X1 U11847 ( .A(n11314), .ZN(n10001) );
  NAND2_X1 U11848 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10003) );
  OR2_X1 U11849 ( .A1(n17307), .A2(n17162), .ZN(n10338) );
  AND2_X1 U11850 ( .A1(n17276), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11305) );
  NOR3_X1 U11851 ( .A1(n15907), .A2(n17503), .A3(n16646), .ZN(n15908) );
  AOI21_X1 U11852 ( .B1(n17191), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n11323), .ZN(n11327) );
  NOR2_X1 U11853 ( .A1(n17242), .A2(n17184), .ZN(n11323) );
  AND2_X1 U11854 ( .A1(n10251), .A2(n10250), .ZN(n11320) );
  NAND2_X1 U11855 ( .A1(n11392), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10251) );
  NOR2_X1 U11856 ( .A1(n12925), .A2(n17975), .ZN(n16498) );
  NOR2_X1 U11857 ( .A1(n17768), .A2(n17772), .ZN(n17758) );
  NOR2_X1 U11858 ( .A1(n17872), .A2(n16850), .ZN(n17809) );
  NAND2_X1 U11859 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16966) );
  INV_X1 U11860 ( .A(n19008), .ZN(n16646) );
  NOR2_X1 U11861 ( .A1(n12912), .A2(n15827), .ZN(n12919) );
  NAND2_X1 U11862 ( .A1(n9867), .A2(n11421), .ZN(n9993) );
  OR2_X1 U11863 ( .A1(n11422), .A2(n18116), .ZN(n11421) );
  INV_X1 U11864 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17842) );
  INV_X1 U11865 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10246) );
  NOR2_X1 U11866 ( .A1(n17918), .A2(n18246), .ZN(n17917) );
  XNOR2_X1 U11867 ( .A(n17496), .B(n18968), .ZN(n17970) );
  NOR2_X1 U11868 ( .A1(n18987), .A2(n18802), .ZN(n18794) );
  OAI21_X1 U11869 ( .B1(n15815), .B2(n17502), .A(n15814), .ZN(n18813) );
  NAND2_X1 U11870 ( .A1(n15871), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20074) );
  INV_X1 U11871 ( .A(n20107), .ZN(n20152) );
  INV_X1 U11872 ( .A(n20155), .ZN(n20130) );
  INV_X1 U11873 ( .A(n13559), .ZN(n20731) );
  AND2_X1 U11874 ( .A1(n11130), .A2(n11082), .ZN(n14651) );
  XNOR2_X1 U11875 ( .A(n10092), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14816) );
  NAND2_X1 U11876 ( .A1(n10094), .A2(n10093), .ZN(n10092) );
  CLKBUF_X1 U11877 ( .A(n13608), .Z(n13609) );
  INV_X1 U11878 ( .A(n20526), .ZN(n20547) );
  AND2_X1 U11879 ( .A1(n13345), .A2(n14963), .ZN(n14955) );
  AND2_X1 U11880 ( .A1(n13397), .A2(n13493), .ZN(n20052) );
  INV_X1 U11881 ( .A(n20031), .ZN(n19586) );
  NAND2_X1 U11882 ( .A1(n15246), .A2(n15247), .ZN(n16221) );
  NAND2_X1 U11883 ( .A1(n19256), .A2(n13418), .ZN(n19225) );
  AOI21_X1 U11884 ( .B1(n16211), .B2(n19282), .A(n12940), .ZN(n12941) );
  AOI21_X1 U11885 ( .B1(n14971), .B2(n19282), .A(n12636), .ZN(n12637) );
  AOI21_X1 U11886 ( .B1(n15531), .B2(n19282), .A(n15356), .ZN(n9939) );
  OAI21_X1 U11887 ( .B1(n16221), .B2(n19301), .A(n10204), .ZN(n10203) );
  AND2_X1 U11888 ( .A1(n10207), .A2(n10205), .ZN(n10204) );
  NOR2_X1 U11889 ( .A1(n15505), .A2(n10206), .ZN(n10205) );
  OR2_X1 U11890 ( .A1(n15509), .A2(n15508), .ZN(n10207) );
  NAND2_X1 U11891 ( .A1(n15506), .A2(n16412), .ZN(n10208) );
  INV_X1 U11892 ( .A(n16383), .ZN(n15688) );
  INV_X1 U11893 ( .A(n19303), .ZN(n16413) );
  NAND2_X1 U11894 ( .A1(n12502), .A2(n12172), .ZN(n19301) );
  NAND2_X1 U11895 ( .A1(n12502), .A2(n20040), .ZN(n19303) );
  OR2_X1 U11896 ( .A1(n16444), .A2(n12958), .ZN(n19995) );
  INV_X1 U11897 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16473) );
  NAND2_X1 U11898 ( .A1(n19023), .A2(n17503), .ZN(n19021) );
  INV_X1 U11899 ( .A(n16672), .ZN(n10037) );
  OR2_X1 U11900 ( .A1(n16675), .A2(n16674), .ZN(n10035) );
  NOR2_X1 U11901 ( .A1(n16680), .A2(n16681), .ZN(n16679) );
  INV_X1 U11902 ( .A(n17023), .ZN(n17016) );
  NOR2_X2 U11903 ( .A1(n17471), .A2(n17983), .ZN(n17852) );
  INV_X1 U11904 ( .A(n17972), .ZN(n17983) );
  INV_X1 U11905 ( .A(n17962), .ZN(n17984) );
  NOR2_X2 U11906 ( .A1(n18287), .A2(n16518), .ZN(n18194) );
  AOI21_X2 U11907 ( .B1(n13307), .B2(n13306), .A(n18846), .ZN(n18293) );
  AOI211_X1 U11908 ( .C1(n18779), .C2(n13304), .A(n13303), .B(n15812), .ZN(
        n13307) );
  AND2_X1 U11909 ( .A1(n11956), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10230) );
  INV_X1 U11910 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10322) );
  INV_X1 U11911 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10177) );
  OAI22_X1 U11912 ( .A1(n12007), .A2(n19588), .B1(n12045), .B2(n13177), .ZN(
        n12010) );
  OAI22_X1 U11913 ( .A1(n12067), .A2(n12008), .B1(n12044), .B2(n13169), .ZN(
        n12009) );
  AND2_X1 U11914 ( .A1(n13269), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11706) );
  AND2_X1 U11915 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11705) );
  AND2_X1 U11916 ( .A1(n11760), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11763) );
  OR2_X1 U11917 ( .A1(n10689), .A2(n10688), .ZN(n11258) );
  NAND2_X1 U11918 ( .A1(n13677), .A2(n10154), .ZN(n13679) );
  NAND2_X1 U11919 ( .A1(n11109), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10372) );
  NOR2_X1 U11920 ( .A1(n12422), .A2(n12416), .ZN(n12415) );
  INV_X1 U11921 ( .A(n15174), .ZN(n10264) );
  NOR2_X1 U11922 ( .A1(n11852), .A2(n11851), .ZN(n11838) );
  OR2_X1 U11923 ( .A1(n12086), .A2(n12085), .ZN(n12403) );
  OR2_X1 U11924 ( .A1(n11796), .A2(n11795), .ZN(n12003) );
  NAND2_X1 U11925 ( .A1(n10058), .A2(n10057), .ZN(n12154) );
  INV_X1 U11926 ( .A(n12092), .ZN(n10058) );
  INV_X1 U11927 ( .A(n10138), .ZN(n10137) );
  OAI211_X1 U11928 ( .C1(n12360), .C2(n15139), .A(n11888), .B(n11889), .ZN(
        n10138) );
  INV_X1 U11929 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12977) );
  OR2_X1 U11930 ( .A1(n11664), .A2(n11663), .ZN(n12025) );
  AND2_X1 U11931 ( .A1(n12173), .A2(n12958), .ZN(n12188) );
  NAND2_X1 U11932 ( .A1(n11881), .A2(n11880), .ZN(n11882) );
  NAND2_X1 U11933 ( .A1(n11879), .A2(n19341), .ZN(n11881) );
  AND2_X1 U11934 ( .A1(n11684), .A2(n11683), .ZN(n11695) );
  AOI22_X1 U11935 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11758), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U11936 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13225), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11712) );
  NOR2_X1 U11937 ( .A1(n17480), .A2(n11375), .ZN(n11391) );
  OAI21_X1 U11938 ( .B1(n18332), .B2(n9824), .A(n11544), .ZN(n11546) );
  AND2_X1 U11939 ( .A1(n18332), .A2(n11545), .ZN(n11531) );
  AND2_X1 U11940 ( .A1(n10320), .A2(n10319), .ZN(n10318) );
  INV_X1 U11941 ( .A(n14329), .ZN(n10319) );
  AND2_X1 U11942 ( .A1(n11004), .A2(n10980), .ZN(n10311) );
  INV_X1 U11943 ( .A(n14408), .ZN(n10980) );
  NAND2_X1 U11944 ( .A1(n10312), .A2(n14474), .ZN(n10024) );
  AND2_X1 U11945 ( .A1(n10853), .A2(n10834), .ZN(n10314) );
  NOR2_X1 U11946 ( .A1(n14108), .A2(n14146), .ZN(n10315) );
  OR2_X1 U11947 ( .A1(n10164), .A2(n10166), .ZN(n10163) );
  NAND2_X1 U11948 ( .A1(n10165), .A2(n14344), .ZN(n10164) );
  INV_X1 U11949 ( .A(n14368), .ZN(n10165) );
  INV_X1 U11950 ( .A(n14354), .ZN(n10166) );
  AND2_X1 U11951 ( .A1(n14451), .A2(n10176), .ZN(n10175) );
  INV_X1 U11952 ( .A(n14439), .ZN(n10176) );
  NAND2_X1 U11953 ( .A1(n11281), .A2(n14751), .ZN(n11289) );
  NAND2_X1 U11954 ( .A1(n12736), .A2(n10169), .ZN(n10168) );
  NAND2_X1 U11955 ( .A1(n11231), .A2(n11230), .ZN(n11234) );
  INV_X1 U11956 ( .A(n12758), .ZN(n12768) );
  OR2_X1 U11957 ( .A1(n10520), .A2(n10519), .ZN(n11206) );
  AOI21_X1 U11958 ( .B1(n13565), .B2(n20274), .A(n10282), .ZN(n13569) );
  NOR2_X1 U11959 ( .A1(n11176), .A2(n11239), .ZN(n11179) );
  NOR2_X1 U11960 ( .A1(n10607), .A2(n20936), .ZN(n11163) );
  AOI21_X1 U11961 ( .B1(n11181), .B2(n11148), .A(n11180), .ZN(n12649) );
  INV_X1 U11962 ( .A(n20281), .ZN(n10452) );
  INV_X1 U11963 ( .A(n13963), .ZN(n14161) );
  AOI21_X1 U11964 ( .B1(n20935), .B2(n16190), .A(n20905), .ZN(n13963) );
  AND2_X1 U11965 ( .A1(n10421), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10021) );
  OR2_X1 U11966 ( .A1(n12520), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12551) );
  AND2_X1 U11967 ( .A1(n9844), .A2(n9902), .ZN(n10112) );
  NAND2_X1 U11968 ( .A1(n12469), .A2(n9844), .ZN(n12485) );
  OR2_X1 U11969 ( .A1(n12453), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12406) );
  NOR2_X1 U11970 ( .A1(n12445), .A2(n12444), .ZN(n12456) );
  NAND2_X1 U11971 ( .A1(n12439), .A2(n12438), .ZN(n12445) );
  AND2_X1 U11972 ( .A1(n12415), .A2(n12430), .ZN(n12439) );
  NAND2_X1 U11973 ( .A1(n10104), .A2(n10103), .ZN(n12416) );
  NAND2_X1 U11974 ( .A1(n12785), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10103) );
  OR2_X1 U11975 ( .A1(n12400), .A2(n12785), .ZN(n10104) );
  INV_X1 U11976 ( .A(n14976), .ZN(n10125) );
  INV_X1 U11977 ( .A(n12625), .ZN(n10127) );
  INV_X1 U11978 ( .A(n15153), .ZN(n10267) );
  INV_X1 U11979 ( .A(n12990), .ZN(n9968) );
  INV_X1 U11980 ( .A(n11938), .ZN(n9954) );
  CLKBUF_X1 U11981 ( .A(n13084), .Z(n13246) );
  INV_X1 U11982 ( .A(n10265), .ZN(n13165) );
  AND2_X1 U11983 ( .A1(n14919), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14916) );
  NOR2_X1 U11984 ( .A1(n15447), .A2(n10181), .ZN(n10180) );
  NOR2_X1 U11985 ( .A1(n16344), .A2(n10188), .ZN(n10187) );
  INV_X1 U11986 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10188) );
  INV_X1 U11987 ( .A(n14927), .ZN(n14923) );
  AND3_X1 U11988 ( .A1(n11645), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11644), .ZN(n11646) );
  AND2_X1 U11989 ( .A1(n11647), .A2(n11619), .ZN(n11648) );
  AOI22_X1 U11990 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9805), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11649) );
  AND2_X1 U11991 ( .A1(n10241), .A2(n10239), .ZN(n10238) );
  NAND2_X1 U11992 ( .A1(n15369), .A2(n15370), .ZN(n10239) );
  NOR2_X1 U11993 ( .A1(n15520), .A2(n10281), .ZN(n10280) );
  AND4_X1 U11994 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(
        n12151) );
  AND4_X1 U11995 ( .A1(n12136), .A2(n12135), .A3(n12134), .A4(n12133), .ZN(
        n12152) );
  AND4_X1 U11996 ( .A1(n12144), .A2(n12143), .A3(n12142), .A4(n12141), .ZN(
        n12150) );
  NAND2_X1 U11997 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n10261), .ZN(
        n10260) );
  NOR2_X1 U11998 ( .A1(n10262), .A2(n12509), .ZN(n10261) );
  NAND2_X1 U11999 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10262) );
  AND2_X1 U12000 ( .A1(n16327), .A2(n10243), .ZN(n10242) );
  NOR2_X1 U12001 ( .A1(n15712), .A2(n10051), .ZN(n10047) );
  OR2_X1 U12002 ( .A1(n11778), .A2(n11777), .ZN(n12027) );
  OR2_X1 U12003 ( .A1(n12002), .A2(n12001), .ZN(n12399) );
  NOR2_X1 U12004 ( .A1(n13213), .A2(n12977), .ZN(n12983) );
  NAND2_X1 U12005 ( .A1(n12959), .A2(n12958), .ZN(n12979) );
  AND2_X1 U12006 ( .A1(n11689), .A2(n11688), .ZN(n11800) );
  NAND2_X1 U12007 ( .A1(n9947), .A2(n11956), .ZN(n12045) );
  INV_X1 U12008 ( .A(n11979), .ZN(n11980) );
  AND2_X1 U12009 ( .A1(n11743), .A2(n10326), .ZN(n11765) );
  NOR3_X1 U12010 ( .A1(n11548), .A2(n11547), .A3(n11546), .ZN(n13298) );
  NAND2_X1 U12011 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n9987) );
  NAND2_X1 U12012 ( .A1(n11548), .A2(n11541), .ZN(n13761) );
  NAND2_X1 U12013 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10250) );
  OR2_X1 U12014 ( .A1(n17877), .A2(n15827), .ZN(n9995) );
  NAND2_X1 U12015 ( .A1(n11391), .A2(n11566), .ZN(n11405) );
  OAI21_X1 U12016 ( .B1(n17917), .B2(n10248), .A(n10247), .ZN(n17780) );
  NAND2_X1 U12017 ( .A1(n17908), .A2(n10249), .ZN(n10247) );
  OR2_X1 U12018 ( .A1(n11390), .A2(n11404), .ZN(n10248) );
  INV_X1 U12019 ( .A(n17978), .ZN(n11573) );
  NOR2_X1 U12020 ( .A1(n10076), .A2(n16646), .ZN(n10075) );
  NOR2_X1 U12021 ( .A1(n15811), .A2(n18805), .ZN(n18803) );
  NAND2_X1 U12022 ( .A1(n14282), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10083) );
  AOI21_X1 U12023 ( .B1(n17297), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n10085), .ZN(n10084) );
  INV_X1 U12024 ( .A(n11453), .ZN(n10088) );
  NOR2_X1 U12025 ( .A1(n11546), .A2(n18789), .ZN(n15813) );
  INV_X1 U12026 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15951) );
  NAND2_X1 U12027 ( .A1(n15941), .A2(n20146), .ZN(n20131) );
  OR2_X1 U12028 ( .A1(n20117), .A2(n20834), .ZN(n14032) );
  NAND2_X1 U12029 ( .A1(n20148), .A2(n12875), .ZN(n20115) );
  AND2_X1 U12030 ( .A1(n12714), .A2(n12713), .ZN(n14185) );
  NOR2_X1 U12031 ( .A1(n15974), .A2(n13792), .ZN(n13796) );
  AND2_X1 U12032 ( .A1(n13653), .A2(n13652), .ZN(n20180) );
  INV_X1 U12033 ( .A(n13453), .ZN(n13629) );
  NOR2_X1 U12034 ( .A1(n11079), .A2(n14657), .ZN(n11080) );
  OR2_X1 U12035 ( .A1(n11021), .A2(n14683), .ZN(n11023) );
  OR2_X1 U12036 ( .A1(n11023), .A2(n11022), .ZN(n11079) );
  AND2_X1 U12037 ( .A1(n10999), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11000) );
  NAND2_X1 U12038 ( .A1(n11000), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11021) );
  NAND2_X1 U12039 ( .A1(n10937), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10998) );
  CLKBUF_X1 U12040 ( .A(n14404), .Z(n14405) );
  NOR2_X1 U12041 ( .A1(n10902), .A2(n14732), .ZN(n10903) );
  NAND2_X1 U12042 ( .A1(n10903), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10935) );
  NAND2_X1 U12043 ( .A1(n10870), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10902) );
  AND2_X1 U12044 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n10869), .ZN(
        n10870) );
  INV_X1 U12045 ( .A(n10868), .ZN(n10869) );
  AND2_X1 U12046 ( .A1(n10867), .A2(n10866), .ZN(n14507) );
  NOR2_X1 U12047 ( .A1(n10836), .A2(n14493), .ZN(n10837) );
  OR2_X1 U12048 ( .A1(n10799), .A2(n15951), .ZN(n10804) );
  AND3_X1 U12049 ( .A1(n10803), .A2(n10802), .A3(n10801), .ZN(n14525) );
  AND2_X1 U12050 ( .A1(n10755), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10756) );
  NAND2_X1 U12051 ( .A1(n10773), .A2(n10772), .ZN(n14619) );
  NOR2_X1 U12052 ( .A1(n10751), .A2(n20097), .ZN(n10755) );
  NAND2_X1 U12053 ( .A1(n10725), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10751) );
  AND2_X1 U12054 ( .A1(n10703), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10725) );
  INV_X1 U12055 ( .A(n10708), .ZN(n10709) );
  INV_X1 U12056 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10692) );
  NOR2_X1 U12057 ( .A1(n10693), .A2(n10692), .ZN(n10703) );
  CLKBUF_X1 U12058 ( .A(n14057), .Z(n14058) );
  INV_X1 U12059 ( .A(n11240), .ZN(n10677) );
  NOR2_X1 U12060 ( .A1(n10623), .A2(n10622), .ZN(n10649) );
  INV_X1 U12061 ( .A(n13812), .ZN(n10597) );
  OR2_X2 U12062 ( .A1(n13686), .A2(n20074), .ZN(n13650) );
  AND2_X1 U12063 ( .A1(n14821), .A2(n14828), .ZN(n10091) );
  NOR3_X1 U12064 ( .A1(n9857), .A2(n10166), .A3(n14368), .ZN(n14356) );
  INV_X1 U12065 ( .A(n10290), .ZN(n9973) );
  NOR2_X1 U12066 ( .A1(n9857), .A2(n14368), .ZN(n14369) );
  AND2_X1 U12067 ( .A1(n10287), .A2(n16042), .ZN(n10098) );
  NOR2_X1 U12068 ( .A1(n14425), .A2(n14410), .ZN(n14411) );
  NAND2_X1 U12069 ( .A1(n14465), .A2(n10173), .ZN(n14425) );
  AND2_X1 U12070 ( .A1(n10175), .A2(n10174), .ZN(n10173) );
  INV_X1 U12071 ( .A(n14423), .ZN(n10174) );
  NAND2_X1 U12072 ( .A1(n14465), .A2(n10175), .ZN(n14441) );
  NAND2_X1 U12073 ( .A1(n14465), .A2(n14451), .ZN(n14453) );
  NOR2_X1 U12074 ( .A1(n9832), .A2(n14463), .ZN(n14465) );
  AND2_X1 U12075 ( .A1(n12729), .A2(n12728), .ZN(n14495) );
  NOR2_X1 U12076 ( .A1(n14528), .A2(n10167), .ZN(n15923) );
  INV_X1 U12077 ( .A(n10169), .ZN(n10167) );
  NOR2_X1 U12078 ( .A1(n14528), .A2(n14518), .ZN(n14519) );
  AND2_X1 U12079 ( .A1(n12720), .A2(n12719), .ZN(n14903) );
  AND3_X1 U12080 ( .A1(n11264), .A2(n11230), .A3(n11267), .ZN(n11265) );
  INV_X1 U12081 ( .A(n16144), .ZN(n10171) );
  NAND2_X1 U12082 ( .A1(n20906), .A2(n20936), .ZN(n11198) );
  NAND2_X1 U12083 ( .A1(n16170), .A2(n10172), .ZN(n16145) );
  AOI21_X1 U12084 ( .B1(n14056), .B2(n10284), .A(n9874), .ZN(n10283) );
  INV_X1 U12085 ( .A(n14056), .ZN(n10285) );
  AND2_X1 U12086 ( .A1(n16170), .A2(n16169), .ZN(n16172) );
  NAND2_X1 U12087 ( .A1(n10158), .A2(n10162), .ZN(n14097) );
  NOR2_X1 U12088 ( .A1(n10159), .A2(n13752), .ZN(n10158) );
  INV_X1 U12089 ( .A(n14077), .ZN(n10160) );
  NAND2_X1 U12090 ( .A1(n10162), .A2(n9920), .ZN(n14078) );
  INV_X1 U12091 ( .A(n13752), .ZN(n10157) );
  NOR2_X1 U12092 ( .A1(n13918), .A2(n13752), .ZN(n10161) );
  OR2_X1 U12093 ( .A1(n13752), .A2(n13753), .ZN(n13919) );
  INV_X1 U12094 ( .A(n15888), .ZN(n14803) );
  NAND2_X1 U12095 ( .A1(n13715), .A2(n20264), .ZN(n16160) );
  NAND2_X1 U12096 ( .A1(n13691), .A2(n13690), .ZN(n13714) );
  OAI21_X1 U12097 ( .B1(n11176), .B2(n20271), .A(n10510), .ZN(n10589) );
  NAND2_X1 U12098 ( .A1(n10089), .A2(n20410), .ZN(n10620) );
  INV_X1 U12099 ( .A(n13624), .ZN(n13580) );
  NAND2_X1 U12100 ( .A1(n10552), .A2(n10551), .ZN(n13635) );
  AND2_X1 U12101 ( .A1(n20521), .A2(n9818), .ZN(n20382) );
  INV_X1 U12102 ( .A(n20382), .ZN(n20383) );
  INV_X1 U12103 ( .A(n20273), .ZN(n20300) );
  AOI22_X1 U12104 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10400) );
  NAND2_X1 U12105 ( .A1(n16001), .A2(n14153), .ZN(n20304) );
  AOI21_X1 U12106 ( .B1(n20696), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20417), 
        .ZN(n20779) );
  CLKBUF_X1 U12107 ( .A(n12640), .Z(n12641) );
  NAND2_X1 U12108 ( .A1(n10215), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10214) );
  NAND2_X1 U12109 ( .A1(n10217), .A2(n11619), .ZN(n10216) );
  AND2_X1 U12110 ( .A1(n14916), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14948) );
  NAND2_X1 U12111 ( .A1(n12519), .A2(n12549), .ZN(n12556) );
  NAND2_X1 U12112 ( .A1(n12529), .A2(n12593), .ZN(n12520) );
  INV_X1 U12113 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15011) );
  NAND2_X1 U12114 ( .A1(n14934), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14937) );
  NAND2_X1 U12115 ( .A1(n12469), .A2(n12407), .ZN(n12481) );
  AND2_X1 U12116 ( .A1(n12463), .A2(n12366), .ZN(n12465) );
  AND2_X1 U12117 ( .A1(n12465), .A2(n13914), .ZN(n12468) );
  AND2_X1 U12118 ( .A1(n13347), .A2(n13493), .ZN(n14963) );
  INV_X1 U12119 ( .A(n10270), .ZN(n10269) );
  AOI21_X1 U12120 ( .B1(n10270), .B2(n10268), .A(n10267), .ZN(n10266) );
  NAND2_X1 U12121 ( .A1(n13215), .A2(n10272), .ZN(n10270) );
  XNOR2_X1 U12122 ( .A(n10265), .B(n13164), .ZN(n15171) );
  NAND2_X1 U12123 ( .A1(n13908), .A2(n12186), .ZN(n10276) );
  NAND2_X1 U12124 ( .A1(n10198), .A2(n15261), .ZN(n10197) );
  NAND2_X1 U12125 ( .A1(n15161), .A2(n15163), .ZN(n15162) );
  AND2_X1 U12126 ( .A1(n12824), .A2(n12823), .ZN(n14995) );
  NAND2_X1 U12127 ( .A1(n10201), .A2(n12820), .ZN(n15276) );
  INV_X1 U12128 ( .A(n15569), .ZN(n10201) );
  NAND2_X1 U12129 ( .A1(n10193), .A2(n15009), .ZN(n10192) );
  INV_X1 U12130 ( .A(n10194), .ZN(n10193) );
  NOR2_X1 U12131 ( .A1(n15316), .A2(n10194), .ZN(n15299) );
  OR2_X1 U12132 ( .A1(n13027), .A2(n13026), .ZN(n15216) );
  AND2_X1 U12133 ( .A1(n12331), .A2(n12330), .ZN(n12332) );
  NAND2_X1 U12134 ( .A1(n14008), .A2(n12329), .ZN(n14129) );
  AND2_X1 U12135 ( .A1(n14124), .A2(n14125), .ZN(n12329) );
  AND2_X1 U12136 ( .A1(n11837), .A2(n11852), .ZN(n14132) );
  CLKBUF_X1 U12137 ( .A(n14121), .Z(n14122) );
  NAND2_X1 U12138 ( .A1(n13537), .A2(n10189), .ZN(n13976) );
  AND2_X1 U12139 ( .A1(n12215), .A2(n10190), .ZN(n10189) );
  AND2_X1 U12140 ( .A1(n10191), .A2(n13979), .ZN(n10190) );
  INV_X1 U12141 ( .A(n13342), .ZN(n19318) );
  NAND2_X1 U12142 ( .A1(n14916), .A2(n9849), .ZN(n14947) );
  NOR2_X1 U12143 ( .A1(n14942), .A2(n10178), .ZN(n14919) );
  NAND2_X1 U12144 ( .A1(n14943), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14942) );
  NAND2_X1 U12145 ( .A1(n14939), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14922) );
  INV_X1 U12146 ( .A(n15204), .ZN(n10128) );
  AND2_X1 U12147 ( .A1(n14934), .A2(n10179), .ZN(n14939) );
  AND2_X1 U12148 ( .A1(n9845), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10179) );
  NAND2_X1 U12149 ( .A1(n14934), .A2(n9845), .ZN(n14938) );
  INV_X1 U12150 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15447) );
  NOR2_X1 U12151 ( .A1(n15650), .A2(n15641), .ZN(n10055) );
  NOR2_X1 U12152 ( .A1(n14935), .A2(n16281), .ZN(n14934) );
  NAND2_X1 U12153 ( .A1(n14932), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14935) );
  NOR2_X1 U12154 ( .A1(n16300), .A2(n14933), .ZN(n14932) );
  NOR2_X1 U12155 ( .A1(n13910), .A2(n10134), .ZN(n14043) );
  INV_X1 U12156 ( .A(n10068), .ZN(n10067) );
  OAI21_X1 U12157 ( .B1(n9841), .B2(n9864), .A(n12476), .ZN(n10068) );
  AND2_X1 U12158 ( .A1(n14923), .A2(n10186), .ZN(n14930) );
  AND2_X1 U12159 ( .A1(n9840), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10186) );
  NAND2_X1 U12160 ( .A1(n14923), .A2(n9840), .ZN(n14931) );
  NAND2_X1 U12161 ( .A1(n14923), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14929) );
  AND2_X1 U12162 ( .A1(n10183), .A2(n9898), .ZN(n14928) );
  AND2_X1 U12163 ( .A1(n12355), .A2(n12354), .ZN(n13806) );
  NAND2_X1 U12164 ( .A1(n10183), .A2(n10184), .ZN(n14925) );
  NAND2_X1 U12165 ( .A1(n10121), .A2(n10120), .ZN(n13805) );
  AND3_X1 U12166 ( .A1(n12345), .A2(n12348), .A3(n13798), .ZN(n10120) );
  NOR2_X1 U12167 ( .A1(n14924), .A2(n19286), .ZN(n14926) );
  AND2_X1 U12168 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14021) );
  INV_X1 U12169 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15136) );
  INV_X1 U12170 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15126) );
  AOI21_X1 U12171 ( .B1(n16210), .B2(n16387), .A(n12898), .ZN(n12902) );
  INV_X1 U12172 ( .A(n15507), .ZN(n10206) );
  AND2_X1 U12173 ( .A1(n15547), .A2(n12843), .ZN(n15493) );
  AND2_X1 U12174 ( .A1(n19051), .A2(n12543), .ZN(n15412) );
  NAND2_X1 U12175 ( .A1(n12803), .A2(n15314), .ZN(n15316) );
  OR2_X1 U12176 ( .A1(n15316), .A2(n15026), .ZN(n15298) );
  OR2_X1 U12177 ( .A1(n12538), .A2(n15604), .ZN(n15423) );
  NOR2_X1 U12178 ( .A1(n10054), .A2(n15450), .ZN(n10053) );
  INV_X1 U12179 ( .A(n10055), .ZN(n10054) );
  OR2_X1 U12180 ( .A1(n19062), .A2(n12539), .ZN(n15436) );
  NAND2_X1 U12181 ( .A1(n15664), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15642) );
  NOR2_X1 U12182 ( .A1(n10134), .A2(n10133), .ZN(n10132) );
  INV_X1 U12183 ( .A(n14042), .ZN(n10133) );
  NAND2_X1 U12184 ( .A1(n10245), .A2(n10242), .ZN(n16310) );
  NOR2_X1 U12185 ( .A1(n13910), .A2(n10136), .ZN(n14000) );
  NOR2_X1 U12186 ( .A1(n13910), .A2(n13911), .ZN(n13909) );
  NAND2_X1 U12187 ( .A1(n10210), .A2(n13660), .ZN(n10209) );
  INV_X1 U12188 ( .A(n10211), .ZN(n10210) );
  OR2_X1 U12189 ( .A1(n13554), .A2(n10212), .ZN(n15079) );
  NOR2_X1 U12190 ( .A1(n16406), .A2(n16408), .ZN(n16393) );
  AND2_X1 U12191 ( .A1(n12363), .A2(n12362), .ZN(n13841) );
  NAND2_X1 U12192 ( .A1(n13978), .A2(n12230), .ZN(n13501) );
  XNOR2_X1 U12193 ( .A(n12449), .B(n12448), .ZN(n15482) );
  OAI21_X1 U12194 ( .B1(n19273), .B2(n19272), .A(n12436), .ZN(n15735) );
  INV_X1 U12195 ( .A(n12037), .ZN(n10220) );
  XNOR2_X1 U12196 ( .A(n11947), .B(n11946), .ZN(n11948) );
  INV_X1 U12197 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13531) );
  XNOR2_X1 U12198 ( .A(n12982), .B(n12983), .ZN(n13508) );
  AND2_X1 U12199 ( .A1(n13538), .A2(n13537), .ZN(n15127) );
  NOR2_X1 U12200 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15765) );
  INV_X1 U12201 ( .A(n20003), .ZN(n19698) );
  NOR2_X1 U12202 ( .A1(n19316), .A2(n19317), .ZN(n19357) );
  NOR2_X1 U12203 ( .A1(n19318), .A2(n19317), .ZN(n19356) );
  INV_X1 U12204 ( .A(n11851), .ZN(n19347) );
  OR2_X1 U12205 ( .A1(n19987), .A2(n19586), .ZN(n19783) );
  NAND2_X1 U12206 ( .A1(n19466), .A2(n20022), .ZN(n19832) );
  INV_X1 U12207 ( .A(n19356), .ZN(n19364) );
  INV_X1 U12208 ( .A(n19357), .ZN(n19366) );
  NOR2_X1 U12209 ( .A1(n19533), .A2(n16478), .ZN(n16485) );
  AOI21_X1 U12210 ( .B1(n16715), .B2(n17630), .A(n16894), .ZN(n16693) );
  NOR2_X1 U12211 ( .A1(n16693), .A2(n17613), .ZN(n16692) );
  AND2_X1 U12212 ( .A1(n10033), .A2(n16931), .ZN(n16739) );
  NOR2_X1 U12213 ( .A1(n16739), .A2(n17664), .ZN(n16738) );
  NOR2_X1 U12214 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16910), .ZN(n16897) );
  NAND2_X1 U12215 ( .A1(n17097), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n17083) );
  NAND2_X1 U12216 ( .A1(n17156), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n17032) );
  NAND2_X1 U12217 ( .A1(n18799), .A2(n11301), .ZN(n17242) );
  OAI211_X1 U12218 ( .C1(n11489), .C2(n18335), .A(n11372), .B(n11371), .ZN(
        n11568) );
  AND2_X1 U12219 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11337) );
  NOR2_X1 U12220 ( .A1(n11340), .A2(n14248), .ZN(n11341) );
  NOR2_X1 U12221 ( .A1(n18337), .A2(n11557), .ZN(n18815) );
  OAI211_X1 U12222 ( .C1(n17307), .C2(n14248), .A(n11508), .B(n11507), .ZN(
        n17503) );
  AOI22_X1 U12223 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11508) );
  AOI211_X1 U12224 ( .C1(n9810), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n11506), .B(n11505), .ZN(n11507) );
  NOR2_X1 U12225 ( .A1(n17540), .A2(n17502), .ZN(n17521) );
  NOR2_X1 U12226 ( .A1(n17541), .A2(n17540), .ZN(n17542) );
  NAND2_X1 U12227 ( .A1(n17640), .A2(n9847), .ZN(n12925) );
  NAND2_X1 U12228 ( .A1(n17640), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17622) );
  AND2_X1 U12229 ( .A1(n17758), .A2(n10028), .ZN(n17680) );
  AND2_X1 U12230 ( .A1(n9846), .A2(n9918), .ZN(n10028) );
  NAND2_X1 U12231 ( .A1(n17758), .A2(n9846), .ZN(n17698) );
  NOR2_X1 U12232 ( .A1(n17737), .A2(n10030), .ZN(n10029) );
  NAND2_X1 U12233 ( .A1(n17758), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17735) );
  NAND2_X1 U12234 ( .A1(n17809), .A2(n9887), .ZN(n17768) );
  NAND2_X1 U12235 ( .A1(n17916), .A2(n9894), .ZN(n17872) );
  AND2_X1 U12236 ( .A1(n17916), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17906) );
  INV_X1 U12237 ( .A(n16966), .ZN(n17945) );
  NAND2_X1 U12238 ( .A1(n9996), .A2(n9994), .ZN(n12918) );
  AND2_X1 U12239 ( .A1(n9995), .A2(n9999), .ZN(n9994) );
  NAND2_X1 U12240 ( .A1(n12911), .A2(n17779), .ZN(n9996) );
  NAND2_X1 U12241 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18967), .ZN(
        n9999) );
  AOI21_X1 U12242 ( .B1(n12914), .B2(n17877), .A(n12920), .ZN(n12915) );
  NOR2_X1 U12243 ( .A1(n12911), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12917) );
  NOR2_X1 U12244 ( .A1(n15879), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15878) );
  NAND2_X1 U12245 ( .A1(n11435), .A2(n9997), .ZN(n12911) );
  NOR2_X1 U12246 ( .A1(n9998), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9997) );
  INV_X1 U12247 ( .A(n16512), .ZN(n9998) );
  NAND2_X1 U12248 ( .A1(n10252), .A2(n17638), .ZN(n12912) );
  NOR2_X1 U12249 ( .A1(n11433), .A2(n9912), .ZN(n10252) );
  INV_X1 U12250 ( .A(n11432), .ZN(n10253) );
  INV_X1 U12251 ( .A(n17628), .ZN(n16514) );
  NOR2_X1 U12252 ( .A1(n13313), .A2(n18131), .ZN(n17985) );
  OR2_X1 U12253 ( .A1(n17660), .A2(n17877), .ZN(n11429) );
  NAND2_X1 U12254 ( .A1(n9990), .A2(n9989), .ZN(n17671) );
  NAND2_X1 U12255 ( .A1(n11426), .A2(n17877), .ZN(n9989) );
  NOR2_X1 U12256 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17711), .ZN(
        n17704) );
  INV_X1 U12257 ( .A(n17710), .ZN(n10256) );
  INV_X1 U12258 ( .A(n11422), .ZN(n18124) );
  AND2_X1 U12259 ( .A1(n17857), .A2(n9924), .ZN(n17803) );
  NAND2_X1 U12260 ( .A1(n18177), .A2(n18114), .ZN(n17792) );
  NAND2_X1 U12261 ( .A1(n17857), .A2(n9854), .ZN(n17829) );
  NOR2_X1 U12262 ( .A1(n18786), .A2(n11541), .ZN(n10082) );
  NAND2_X1 U12263 ( .A1(n18801), .A2(n15811), .ZN(n18796) );
  INV_X1 U12264 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18212) );
  XNOR2_X1 U12265 ( .A(n17780), .B(n11416), .ZN(n17891) );
  NOR2_X1 U12266 ( .A1(n11582), .A2(n17919), .ZN(n17899) );
  NAND2_X1 U12267 ( .A1(n17942), .A2(n9866), .ZN(n10004) );
  NOR2_X1 U12268 ( .A1(n18775), .A2(n13308), .ZN(n13303) );
  AOI21_X1 U12269 ( .B1(n11553), .B2(n11552), .A(n11551), .ZN(n18779) );
  NOR2_X1 U12270 ( .A1(n13309), .A2(n13308), .ZN(n18776) );
  INV_X1 U12271 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18821) );
  INV_X1 U12272 ( .A(n11540), .ZN(n18792) );
  INV_X1 U12273 ( .A(n11307), .ZN(n18799) );
  INV_X1 U12274 ( .A(n18803), .ZN(n15817) );
  NAND3_X1 U12275 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15818) );
  INV_X1 U12276 ( .A(n17503), .ZN(n18314) );
  AOI211_X1 U12277 ( .C1(n17228), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n11476), .B(n11475), .ZN(n18322) );
  AND2_X1 U12278 ( .A1(n9935), .A2(n9933), .ZN(n18327) );
  NOR2_X1 U12279 ( .A1(n11466), .A2(n9934), .ZN(n9933) );
  INV_X1 U12280 ( .A(n11465), .ZN(n9935) );
  AND2_X1 U12281 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n9934) );
  INV_X1 U12282 ( .A(n13762), .ZN(n18332) );
  NAND2_X1 U12283 ( .A1(n11561), .A2(n18312), .ZN(n18356) );
  AOI21_X1 U12284 ( .B1(n18271), .B2(n10073), .A(n9833), .ZN(n18782) );
  INV_X1 U12285 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U12286 ( .A1(n14035), .A2(n12771), .ZN(n14315) );
  NAND2_X1 U12287 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20940) );
  OR2_X1 U12288 ( .A1(n20117), .A2(n20661), .ZN(n20098) );
  NOR2_X2 U12289 ( .A1(n14032), .A2(n14031), .ZN(n20127) );
  INV_X1 U12290 ( .A(n14030), .ZN(n14031) );
  INV_X1 U12291 ( .A(n20098), .ZN(n20139) );
  OR2_X1 U12292 ( .A1(n14036), .A2(n12860), .ZN(n20155) );
  INV_X1 U12293 ( .A(n20127), .ZN(n20142) );
  OR2_X1 U12294 ( .A1(n14036), .A2(n12879), .ZN(n20107) );
  NAND2_X1 U12295 ( .A1(n12877), .A2(n10152), .ZN(n12879) );
  INV_X1 U12296 ( .A(n10153), .ZN(n10152) );
  INV_X1 U12297 ( .A(n20115), .ZN(n20106) );
  INV_X1 U12298 ( .A(n14532), .ZN(n20176) );
  OR2_X1 U12299 ( .A1(n12675), .A2(n12857), .ZN(n12676) );
  OR2_X1 U12300 ( .A1(n15974), .A2(n13795), .ZN(n14597) );
  AND2_X1 U12301 ( .A1(n13796), .A2(n14153), .ZN(n15977) );
  INV_X1 U12302 ( .A(n14624), .ZN(n15978) );
  INV_X1 U12303 ( .A(n14597), .ZN(n15976) );
  NAND2_X2 U12304 ( .A1(n12654), .A2(n13690), .ZN(n15974) );
  NAND2_X1 U12305 ( .A1(n12653), .A2(n12652), .ZN(n12654) );
  OR2_X1 U12306 ( .A1(n15976), .A2(n13796), .ZN(n14622) );
  INV_X1 U12307 ( .A(n15974), .ZN(n14611) );
  OR2_X1 U12308 ( .A1(n20223), .A2(n20274), .ZN(n20212) );
  NOR2_X2 U12309 ( .A1(n13651), .A2(n13630), .ZN(n20248) );
  INV_X1 U12310 ( .A(n20212), .ZN(n20251) );
  NAND2_X1 U12311 ( .A1(n14341), .A2(n14342), .ZN(n14343) );
  INV_X1 U12312 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14657) );
  OAI21_X1 U12313 ( .B1(n14365), .B2(n14367), .A(n14366), .ZN(n14675) );
  NAND2_X1 U12314 ( .A1(n10289), .A2(n14729), .ZN(n14705) );
  NAND2_X1 U12315 ( .A1(n14738), .A2(n11290), .ZN(n10289) );
  INV_X1 U12316 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14732) );
  INV_X1 U12317 ( .A(n16022), .ZN(n16024) );
  INV_X1 U12318 ( .A(n16029), .ZN(n16015) );
  XNOR2_X1 U12319 ( .A(n12859), .B(n12858), .ZN(n14790) );
  NOR2_X1 U12320 ( .A1(n14636), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14630) );
  OR2_X1 U12321 ( .A1(n14332), .A2(n14331), .ZN(n14832) );
  NOR2_X1 U12322 ( .A1(n14794), .A2(n15901), .ZN(n16055) );
  OR2_X1 U12323 ( .A1(n11198), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16162) );
  NAND2_X1 U12324 ( .A1(n11250), .A2(n11249), .ZN(n14055) );
  OR2_X1 U12325 ( .A1(n13714), .A2(n13948), .ZN(n20264) );
  INV_X1 U12326 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20696) );
  NOR2_X2 U12327 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20698) );
  INV_X1 U12328 ( .A(n20698), .ZN(n20920) );
  NOR2_X1 U12329 ( .A1(n13686), .A2(n20661), .ZN(n20905) );
  AND2_X1 U12330 ( .A1(n13605), .A2(n13604), .ZN(n20909) );
  OAI21_X1 U12331 ( .B1(n20433), .B2(n20418), .A(n20736), .ZN(n20436) );
  OAI211_X1 U12332 ( .C1(n20545), .C2(n20661), .A(n20584), .B(n20530), .ZN(
        n20548) );
  INV_X1 U12333 ( .A(n20588), .ZN(n20613) );
  INV_X1 U12334 ( .A(n20649), .ZN(n20690) );
  OAI211_X1 U12335 ( .C1(n20762), .C2(n20737), .A(n20736), .B(n20735), .ZN(
        n20766) );
  INV_X1 U12336 ( .A(n20665), .ZN(n20786) );
  INV_X1 U12337 ( .A(n20353), .ZN(n20792) );
  OR2_X1 U12338 ( .A1(n20777), .A2(n20626), .ZN(n20803) );
  INV_X1 U12339 ( .A(n20596), .ZN(n20798) );
  INV_X1 U12340 ( .A(n20683), .ZN(n20818) );
  INV_X1 U12341 ( .A(n20803), .ZN(n20828) );
  AND2_X1 U12342 ( .A1(n20834), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15871) );
  INV_X1 U12343 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20661) );
  NAND2_X1 U12344 ( .A1(n12579), .A2(n9853), .ZN(n12784) );
  NAND2_X1 U12345 ( .A1(n14950), .A2(n14949), .ZN(n16198) );
  NAND2_X1 U12346 ( .A1(n12579), .A2(n12578), .ZN(n12780) );
  NAND2_X1 U12347 ( .A1(n16238), .A2(n16239), .ZN(n16237) );
  AND2_X1 U12348 ( .A1(n12567), .A2(n12787), .ZN(n16236) );
  OR2_X1 U12349 ( .A1(n12565), .A2(n12563), .ZN(n15003) );
  NAND2_X1 U12350 ( .A1(n14992), .A2(n15362), .ZN(n14991) );
  INV_X1 U12351 ( .A(n19193), .ZN(n19163) );
  AND2_X1 U12352 ( .A1(n10115), .A2(n12560), .ZN(n16248) );
  NAND2_X1 U12353 ( .A1(n15838), .A2(n15839), .ZN(n15837) );
  AND2_X1 U12354 ( .A1(n12530), .A2(n12532), .ZN(n15018) );
  INV_X1 U12355 ( .A(n19186), .ZN(n19102) );
  INV_X1 U12356 ( .A(n19181), .ZN(n19166) );
  AND2_X1 U12357 ( .A1(n9913), .A2(n13537), .ZN(n13980) );
  NAND2_X1 U12358 ( .A1(n16200), .A2(n14956), .ZN(n19183) );
  INV_X1 U12359 ( .A(n19891), .ZN(n19190) );
  OR2_X1 U12360 ( .A1(n12310), .A2(n12309), .ZN(n14088) );
  OR2_X1 U12361 ( .A1(n12297), .A2(n12296), .ZN(n14086) );
  OR2_X1 U12362 ( .A1(n12269), .A2(n12268), .ZN(n14004) );
  AND2_X1 U12363 ( .A1(n13843), .A2(n13842), .ZN(n12995) );
  INV_X2 U12364 ( .A(n15235), .ZN(n15221) );
  INV_X1 U12365 ( .A(n15237), .ZN(n15224) );
  AND2_X2 U12366 ( .A1(n13292), .A2(n13493), .ZN(n15235) );
  NAND2_X1 U12367 ( .A1(n10271), .A2(n9843), .ZN(n9961) );
  NAND2_X1 U12368 ( .A1(n15159), .A2(n15158), .ZN(n9960) );
  NOR2_X1 U12369 ( .A1(n15185), .A2(n13110), .ZN(n15175) );
  AND2_X1 U12370 ( .A1(n14131), .A2(n19318), .ZN(n19200) );
  AND2_X1 U12371 ( .A1(n14131), .A2(n19316), .ZN(n19197) );
  NAND2_X1 U12372 ( .A1(n13497), .A2(n13496), .ZN(n19217) );
  NAND2_X1 U12373 ( .A1(n9969), .A2(n12990), .ZN(n13783) );
  NAND2_X1 U12374 ( .A1(n13789), .A2(n13788), .ZN(n9969) );
  INV_X1 U12375 ( .A(n19198), .ZN(n15310) );
  AND2_X1 U12376 ( .A1(n19217), .A2(n19369), .ZN(n19198) );
  INV_X1 U12377 ( .A(n19217), .ZN(n19203) );
  INV_X1 U12378 ( .A(n15327), .ZN(n16268) );
  OAI21_X1 U12379 ( .B1(n13416), .B2(n13415), .A(n13490), .ZN(n13417) );
  INV_X2 U12380 ( .A(n19225), .ZN(n19254) );
  AND2_X2 U12381 ( .A1(n14955), .A2(n12173), .ZN(n19266) );
  XNOR2_X1 U12382 ( .A(n12949), .B(n12948), .ZN(n14911) );
  NAND2_X1 U12383 ( .A1(n12947), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12949) );
  XNOR2_X1 U12384 ( .A(n12800), .B(n12799), .ZN(n16205) );
  AND2_X1 U12385 ( .A1(n15205), .A2(n15025), .ZN(n15617) );
  INV_X1 U12386 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19286) );
  NAND2_X1 U12387 ( .A1(n10121), .A2(n12345), .ZN(n13785) );
  NAND2_X1 U12388 ( .A1(n13349), .A2(n12629), .ZN(n19285) );
  INV_X1 U12389 ( .A(n19317), .ZN(n19282) );
  AND2_X1 U12391 ( .A1(n19285), .A2(n13386), .ZN(n19270) );
  INV_X1 U12392 ( .A(n19270), .ZN(n16366) );
  INV_X1 U12393 ( .A(n19285), .ZN(n16355) );
  NAND3_X1 U12394 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20007), .A3(n19836), 
        .ZN(n19317) );
  NAND2_X1 U12395 ( .A1(n16205), .A2(n16412), .ZN(n10122) );
  NAND2_X1 U12396 ( .A1(n10226), .A2(n12783), .ZN(n10225) );
  OAI21_X1 U12397 ( .B1(n10224), .B2(n10109), .A(n10108), .ZN(n10223) );
  NAND2_X1 U12398 ( .A1(n12892), .A2(n10107), .ZN(n10222) );
  OAI21_X1 U12399 ( .B1(n12510), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12893), .ZN(n15488) );
  NAND2_X1 U12400 ( .A1(n9860), .A2(n10065), .ZN(n10064) );
  INV_X1 U12401 ( .A(n9893), .ZN(n10065) );
  NAND2_X1 U12402 ( .A1(n10063), .A2(n9893), .ZN(n10066) );
  NAND2_X1 U12403 ( .A1(n15389), .A2(n15387), .ZN(n10063) );
  NAND2_X1 U12404 ( .A1(n10060), .A2(n12159), .ZN(n10059) );
  INV_X1 U12405 ( .A(n9943), .ZN(n9942) );
  NOR2_X1 U12406 ( .A1(n15712), .A2(n10051), .ZN(n10060) );
  NAND2_X1 U12407 ( .A1(n15664), .A2(n10053), .ZN(n10056) );
  NAND2_X1 U12408 ( .A1(n19303), .A2(n13524), .ZN(n10150) );
  AND2_X1 U12409 ( .A1(n13529), .A2(n15641), .ZN(n10149) );
  NAND2_X1 U12410 ( .A1(n10245), .A2(n12461), .ZN(n15701) );
  NAND2_X1 U12411 ( .A1(n15713), .A2(n12159), .ZN(n15465) );
  INV_X1 U12412 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15738) );
  INV_X1 U12413 ( .A(n19314), .ZN(n19296) );
  OR2_X1 U12414 ( .A1(n12982), .A2(n13514), .ZN(n20031) );
  INV_X1 U12415 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20019) );
  NAND2_X1 U12416 ( .A1(n13662), .A2(n13665), .ZN(n20015) );
  INV_X1 U12417 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15906) );
  INV_X1 U12418 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15761) );
  CLKBUF_X1 U12419 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n19998) );
  INV_X1 U12420 ( .A(n20022), .ZN(n19994) );
  INV_X1 U12421 ( .A(n20015), .ZN(n19466) );
  XNOR2_X1 U12422 ( .A(n13788), .B(n13789), .ZN(n19987) );
  INV_X1 U12423 ( .A(n11846), .ZN(n13410) );
  NOR2_X1 U12424 ( .A1(n19624), .A2(n19526), .ZN(n19401) );
  INV_X1 U12425 ( .A(n19478), .ZN(n19495) );
  INV_X1 U12426 ( .A(n19518), .ZN(n19521) );
  OAI21_X1 U12427 ( .B1(n19505), .B2(n19504), .A(n19503), .ZN(n19522) );
  OAI21_X1 U12428 ( .B1(n19505), .B2(n19501), .A(n19500), .ZN(n19523) );
  OR2_X1 U12429 ( .A1(n19531), .A2(n19530), .ZN(n19556) );
  NOR2_X1 U12430 ( .A1(n19832), .A2(n19526), .ZN(n19582) );
  NAND2_X1 U12431 ( .A1(n19596), .A2(n19595), .ZN(n19613) );
  OR2_X1 U12432 ( .A1(n19783), .A2(n19624), .ZN(n19645) );
  INV_X1 U12433 ( .A(n19632), .ZN(n19649) );
  NOR2_X1 U12434 ( .A1(n19755), .A2(n19698), .ZN(n19722) );
  OAI22_X1 U12435 ( .A1(n15260), .A2(n19366), .B1(n15259), .B2(n19364), .ZN(
        n19760) );
  OAI22_X1 U12436 ( .A1(n14551), .A2(n19366), .B1(n19340), .B2(n19364), .ZN(
        n19764) );
  OAI22_X1 U12437 ( .A1(n14535), .A2(n19366), .B1(n19358), .B2(n19364), .ZN(
        n19774) );
  AND2_X1 U12438 ( .A1(n19790), .A2(n19789), .ZN(n19801) );
  OAI22_X1 U12439 ( .A1(n14560), .A2(n19366), .B1(n19331), .B2(n19364), .ZN(
        n19800) );
  OAI22_X1 U12440 ( .A1(n14540), .A2(n19366), .B1(n19352), .B2(n19364), .ZN(
        n19811) );
  OR2_X1 U12441 ( .A1(n19755), .A2(n19754), .ZN(n19818) );
  OAI21_X1 U12442 ( .B1(n19795), .B2(n19794), .A(n19793), .ZN(n19822) );
  INV_X1 U12443 ( .A(n19801), .ZN(n19823) );
  INV_X1 U12444 ( .A(n19818), .ZN(n19820) );
  INV_X1 U12445 ( .A(n19880), .ZN(n19826) );
  INV_X1 U12446 ( .A(n19665), .ZN(n19838) );
  INV_X1 U12447 ( .A(n19763), .ZN(n19848) );
  OAI22_X1 U12448 ( .A1(n20296), .A2(n19366), .B1(n19351), .B2(n19364), .ZN(
        n19866) );
  INV_X1 U12449 ( .A(n19679), .ZN(n19872) );
  OR2_X1 U12450 ( .A1(n19783), .A2(n19832), .ZN(n19885) );
  OAI22_X1 U12451 ( .A1(n19363), .A2(n19366), .B1(n19362), .B2(n19364), .ZN(
        n19880) );
  NAND2_X1 U12452 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11831), .ZN(n16495) );
  OAI21_X1 U12453 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n20054), .ZN(n16490) );
  INV_X1 U12454 ( .A(n15122), .ZN(n19891) );
  INV_X1 U12455 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20054) );
  AND2_X1 U12456 ( .A1(n16484), .A2(n16483), .ZN(n19890) );
  INV_X1 U12457 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n12958) );
  NOR2_X1 U12458 ( .A1(n18778), .A2(n17540), .ZN(n19023) );
  INV_X1 U12459 ( .A(n19023), .ZN(n19019) );
  NAND2_X1 U12460 ( .A1(n19004), .A2(n18779), .ZN(n17540) );
  NAND2_X1 U12461 ( .A1(n10072), .A2(n10070), .ZN(n16630) );
  INV_X1 U12462 ( .A(n10071), .ZN(n10070) );
  OR2_X1 U12463 ( .A1(n18271), .A2(n9833), .ZN(n10072) );
  OAI21_X1 U12464 ( .B1(n10073), .B2(n9833), .A(n19004), .ZN(n10071) );
  INV_X1 U12465 ( .A(n10038), .ZN(n16702) );
  AND2_X1 U12466 ( .A1(n10038), .A2(n17630), .ZN(n16701) );
  INV_X1 U12467 ( .A(n16999), .ZN(n17025) );
  CLKBUF_X1 U12468 ( .A(n16985), .Z(n16894) );
  NOR2_X1 U12469 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16861), .ZN(n16846) );
  NOR2_X1 U12470 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16960), .ZN(n16943) );
  NAND2_X1 U12471 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17028), .ZN(n16965) );
  INV_X1 U12472 ( .A(n16965), .ZN(n17011) );
  NAND3_X1 U12473 ( .A1(n16976), .A2(n19019), .A3(n18844), .ZN(n17028) );
  NAND2_X1 U12474 ( .A1(n17088), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17079) );
  NOR2_X1 U12475 ( .A1(n17083), .A2(n17035), .ZN(n17088) );
  NOR2_X1 U12476 ( .A1(n17092), .A2(n16753), .ZN(n17097) );
  NOR2_X1 U12477 ( .A1(n17221), .A2(n17206), .ZN(n17193) );
  NAND2_X1 U12478 ( .A1(n17193), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n17192) );
  NAND2_X1 U12479 ( .A1(n17322), .A2(n14212), .ZN(n17226) );
  AND2_X1 U12480 ( .A1(n17344), .A2(n9936), .ZN(n17322) );
  INV_X1 U12481 ( .A(n13775), .ZN(n9936) );
  INV_X1 U12482 ( .A(n17341), .ZN(n17324) );
  NAND2_X1 U12483 ( .A1(n11515), .A2(n9983), .ZN(n17393) );
  NOR2_X1 U12484 ( .A1(n9985), .A2(n9984), .ZN(n9983) );
  NAND2_X1 U12485 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(P3_EAX_REG_29__SCAN_IN), 
        .ZN(n9982) );
  NOR2_X1 U12486 ( .A1(n17373), .A2(n17566), .ZN(n17368) );
  NOR3_X1 U12487 ( .A1(n17373), .A2(n17566), .A3(n17568), .ZN(n17356) );
  NOR3_X1 U12488 ( .A1(n17393), .A2(n17426), .A3(n17546), .ZN(n17418) );
  NOR2_X2 U12489 ( .A1(n9806), .A2(n17488), .ZN(n17424) );
  NOR2_X2 U12490 ( .A1(n17351), .A2(n17488), .ZN(n17425) );
  AND2_X1 U12491 ( .A1(n19004), .A2(n9978), .ZN(n9977) );
  INV_X1 U12492 ( .A(n17431), .ZN(n9978) );
  NOR2_X1 U12493 ( .A1(n17431), .A2(n17486), .ZN(n17473) );
  AOI211_X1 U12494 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n11387), .B(n11386), .ZN(n17476) );
  NOR2_X1 U12495 ( .A1(n11357), .A2(n10333), .ZN(n11358) );
  NOR2_X1 U12496 ( .A1(n11306), .A2(n11305), .ZN(n11316) );
  AOI211_X1 U12497 ( .C1(n14282), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n10002), .B(n10001), .ZN(n10000) );
  NAND2_X1 U12498 ( .A1(n9824), .A2(n15911), .ZN(n17490) );
  NAND2_X1 U12499 ( .A1(n9979), .A2(n19004), .ZN(n17494) );
  AOI211_X1 U12500 ( .C1(n9810), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n11322), .B(n11321), .ZN(n11329) );
  INV_X1 U12501 ( .A(n17494), .ZN(n15911) );
  NOR2_X1 U12502 ( .A1(n9824), .A2(n17488), .ZN(n17498) );
  INV_X1 U12503 ( .A(n17490), .ZN(n17497) );
  CLKBUF_X1 U12504 ( .A(n17605), .Z(n17597) );
  NOR2_X1 U12505 ( .A1(n19008), .A2(n17597), .ZN(n17598) );
  OAI21_X1 U12506 ( .B1(n19008), .B2(n19009), .A(n17542), .ZN(n17605) );
  NOR2_X1 U12508 ( .A1(n17653), .A2(n17654), .ZN(n17640) );
  OAI21_X1 U12509 ( .B1(n17703), .B2(n10081), .A(n10078), .ZN(n17650) );
  AOI21_X1 U12510 ( .B1(n9830), .B2(n17871), .A(n9923), .ZN(n10078) );
  INV_X1 U12511 ( .A(n18348), .ZN(n18708) );
  OAI21_X1 U12512 ( .B1(n10081), .B2(n18177), .A(n16506), .ZN(n10080) );
  OAI21_X1 U12513 ( .B1(n17885), .B2(n17871), .A(n9830), .ZN(n17867) );
  NOR2_X1 U12514 ( .A1(n16966), .A2(n16971), .ZN(n17916) );
  INV_X1 U12515 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16984) );
  INV_X1 U12516 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17960) );
  NOR2_X2 U12517 ( .A1(n16646), .A2(n16630), .ZN(n17962) );
  NOR2_X1 U12518 ( .A1(n17946), .A2(n18855), .ZN(n17976) );
  NOR2_X2 U12519 ( .A1(n16630), .A2(n19008), .ZN(n17972) );
  INV_X1 U12520 ( .A(n17966), .ZN(n17971) );
  INV_X1 U12521 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17975) );
  INV_X1 U12522 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18966) );
  OAI21_X1 U12523 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19003), .A(n16630), 
        .ZN(n17979) );
  NAND2_X1 U12524 ( .A1(n11421), .A2(n9891), .ZN(n17757) );
  NAND2_X1 U12525 ( .A1(n18271), .A2(n18809), .ZN(n18235) );
  NOR2_X1 U12526 ( .A1(n18137), .A2(n17819), .ZN(n18144) );
  AND2_X1 U12527 ( .A1(n17857), .A2(n9919), .ZN(n17840) );
  INV_X1 U12528 ( .A(n18814), .ZN(n18804) );
  NOR2_X1 U12529 ( .A1(n17917), .A2(n11390), .ZN(n17909) );
  AND2_X1 U12530 ( .A1(n10006), .A2(n9836), .ZN(n17943) );
  INV_X1 U12531 ( .A(n18236), .ZN(n18289) );
  INV_X1 U12532 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18819) );
  INV_X1 U12533 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18826) );
  AOI211_X1 U12534 ( .C1(n19004), .C2(n18813), .A(n18313), .B(n15816), .ZN(
        n18988) );
  INV_X1 U12535 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18783) );
  INV_X1 U12536 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18330) );
  INV_X1 U12537 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18340) );
  INV_X1 U12538 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18345) );
  NOR2_X1 U12539 ( .A1(n18337), .A2(n18349), .ZN(n18691) );
  NOR2_X1 U12540 ( .A1(n18350), .A2(n18349), .ZN(n18765) );
  INV_X1 U12541 ( .A(n17006), .ZN(n18852) );
  NOR2_X1 U12542 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n11561), .ZN(n18851) );
  INV_X1 U12543 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18954) );
  OAI211_X1 U12544 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18873), .B(n18939), .ZN(n19006) );
  INV_X1 U12545 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18873) );
  NAND2_X1 U12546 ( .A1(n18873), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18997) );
  INV_X1 U12547 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21289) );
  INV_X1 U12548 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21130) );
  CLKBUF_X1 U12549 ( .A(n16612), .Z(n16616) );
  OAI21_X1 U12550 ( .B1(n14816), .B2(n9970), .A(n9873), .ZN(P1_U2968) );
  INV_X1 U12551 ( .A(n11296), .ZN(n9970) );
  NAND2_X1 U12552 ( .A1(n9959), .A2(n9957), .ZN(P2_U2860) );
  INV_X1 U12553 ( .A(n9958), .ZN(n9957) );
  NAND2_X1 U12554 ( .A1(n15257), .A2(n15224), .ZN(n9959) );
  OAI21_X1 U12555 ( .B1(n15514), .B2(n15221), .A(n15160), .ZN(n9958) );
  NAND2_X1 U12556 ( .A1(n12937), .A2(n16361), .ZN(n12945) );
  NAND2_X1 U12557 ( .A1(n9940), .A2(n9937), .ZN(P2_U2988) );
  INV_X1 U12558 ( .A(n9938), .ZN(n9937) );
  OAI21_X1 U12559 ( .B1(n15534), .B2(n19277), .A(n9939), .ZN(n9938) );
  OAI21_X1 U12560 ( .B1(n12955), .B2(n19314), .A(n10227), .ZN(P2_U3015) );
  INV_X1 U12561 ( .A(n10228), .ZN(n10227) );
  OAI21_X1 U12562 ( .B1(n12946), .B2(n19303), .A(n10061), .ZN(n10228) );
  AND2_X1 U12563 ( .A1(n12848), .A2(n10122), .ZN(n10061) );
  NAND2_X1 U12564 ( .A1(n10208), .A2(n10202), .ZN(n15510) );
  INV_X1 U12565 ( .A(n10203), .ZN(n10202) );
  AOI21_X1 U12566 ( .B1(n10036), .B2(n17006), .A(n10035), .ZN(n16678) );
  XNOR2_X1 U12567 ( .A(n16671), .B(n10037), .ZN(n10036) );
  AOI21_X1 U12568 ( .B1(n13327), .B2(n17852), .A(n12934), .ZN(n12935) );
  OAI211_X1 U12569 ( .C1(n13325), .C2(n18302), .A(n13324), .B(n13323), .ZN(
        n13326) );
  NOR2_X2 U12570 ( .A1(n17014), .A2(n11310), .ZN(n11392) );
  NAND2_X1 U12572 ( .A1(n10835), .A2(n10834), .ZN(n14490) );
  INV_X1 U12573 ( .A(n9830), .ZN(n10081) );
  INV_X1 U12574 ( .A(n10017), .ZN(n14169) );
  AND4_X2 U12575 ( .A1(n10322), .A2(n10324), .A3(n10323), .A4(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9839) );
  INV_X1 U12576 ( .A(n12222), .ZN(n10219) );
  AND3_X1 U12577 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9828) );
  AND2_X1 U12578 ( .A1(n18271), .A2(n10075), .ZN(n9829) );
  INV_X1 U12579 ( .A(n11610), .ZN(n11992) );
  OR2_X1 U12580 ( .A1(n17984), .A2(n17816), .ZN(n9830) );
  AND3_X1 U12581 ( .A1(n10440), .A2(n10438), .A3(n10439), .ZN(n9831) );
  OR3_X1 U12582 ( .A1(n14528), .A2(n10168), .A3(n14477), .ZN(n9832) );
  AND2_X1 U12583 ( .A1(n13298), .A2(n13303), .ZN(n9833) );
  OR2_X1 U12584 ( .A1(n15404), .A2(n10262), .ZN(n15378) );
  NAND2_X1 U12585 ( .A1(n14615), .A2(n14616), .ZN(n14524) );
  NOR2_X1 U12586 ( .A1(n15569), .A2(n10199), .ZN(n9834) );
  NAND2_X1 U12587 ( .A1(n10259), .A2(n10261), .ZN(n9835) );
  OR2_X1 U12588 ( .A1(n18270), .A2(n11347), .ZN(n9836) );
  NOR2_X1 U12589 ( .A1(n14488), .A2(n10024), .ZN(n9837) );
  AND4_X1 U12590 ( .A1(n10449), .A2(n10020), .A3(n10447), .A4(n10448), .ZN(
        n9838) );
  INV_X1 U12591 ( .A(n12162), .ZN(n10051) );
  AND2_X1 U12592 ( .A1(n10187), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9840) );
  AND4_X1 U12593 ( .A1(n10394), .A2(n10393), .A3(n10392), .A4(n10391), .ZN(
        n9842) );
  NAND2_X1 U12594 ( .A1(n18980), .A2(n18987), .ZN(n17014) );
  NAND2_X1 U12595 ( .A1(n20055), .A2(n12584), .ZN(n12501) );
  INV_X1 U12596 ( .A(n10450), .ZN(n10461) );
  INV_X1 U12597 ( .A(n10023), .ZN(n14475) );
  NAND2_X1 U12598 ( .A1(n9963), .A2(n9964), .ZN(n14087) );
  NAND2_X1 U12599 ( .A1(n14174), .A2(n10279), .ZN(n15202) );
  NAND2_X1 U12600 ( .A1(n15199), .A2(n15200), .ZN(n15191) );
  NAND2_X1 U12601 ( .A1(n14174), .A2(n15216), .ZN(n15210) );
  AND2_X1 U12602 ( .A1(n12407), .A2(n9907), .ZN(n9844) );
  AND2_X1 U12603 ( .A1(n10180), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9845) );
  AND2_X1 U12604 ( .A1(n10029), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9846) );
  INV_X1 U12605 ( .A(n10669), .ZN(n10096) );
  AND2_X1 U12606 ( .A1(n9828), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9847) );
  AND2_X1 U12607 ( .A1(n9964), .A2(n9962), .ZN(n9848) );
  AND2_X1 U12608 ( .A1(n13280), .A2(n11619), .ZN(n13033) );
  AND2_X1 U12609 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9849) );
  AND2_X1 U12610 ( .A1(n9906), .A2(n10113), .ZN(n9850) );
  AND2_X1 U12611 ( .A1(n9849), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9851) );
  AND2_X1 U12612 ( .A1(n9850), .A2(n15172), .ZN(n9852) );
  AND2_X1 U12613 ( .A1(n12578), .A2(n9921), .ZN(n9853) );
  AND2_X1 U12614 ( .A1(n9919), .A2(n17842), .ZN(n9854) );
  OR2_X1 U12615 ( .A1(n10260), .A2(n15546), .ZN(n9855) );
  OR2_X1 U12616 ( .A1(n9855), .A2(n9929), .ZN(n9856) );
  OR2_X1 U12617 ( .A1(n14396), .A2(n14381), .ZN(n9857) );
  INV_X1 U12618 ( .A(n12835), .ZN(n12813) );
  NAND2_X1 U12619 ( .A1(n12469), .A2(n10112), .ZN(n9859) );
  NAND2_X1 U12620 ( .A1(n10059), .A2(n9942), .ZN(n15417) );
  NAND2_X1 U12621 ( .A1(n9814), .A2(n9841), .ZN(n10245) );
  INV_X1 U12622 ( .A(n10079), .ZN(n17778) );
  AOI21_X1 U12623 ( .B1(n17885), .B2(n9830), .A(n10080), .ZN(n10079) );
  NAND2_X1 U12624 ( .A1(n9814), .A2(n12450), .ZN(n15467) );
  XNOR2_X1 U12625 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n12554), .ZN(
        n9860) );
  NAND2_X1 U12626 ( .A1(n11981), .A2(n11966), .ZN(n12067) );
  NAND2_X1 U12627 ( .A1(n14404), .A2(n10311), .ZN(n14378) );
  NAND2_X1 U12628 ( .A1(n14404), .A2(n10980), .ZN(n14390) );
  NOR2_X1 U12629 ( .A1(n15191), .A2(n15192), .ZN(n13109) );
  NAND2_X1 U12630 ( .A1(n12174), .A2(n12957), .ZN(n12193) );
  NAND2_X1 U12631 ( .A1(n12508), .A2(n15609), .ZN(n15428) );
  OR3_X1 U12632 ( .A1(n17373), .A2(n17566), .A3(n9982), .ZN(n9861) );
  OR2_X1 U12633 ( .A1(n13192), .A2(n13191), .ZN(n9862) );
  OR2_X1 U12634 ( .A1(n16313), .A2(n10069), .ZN(n9864) );
  INV_X1 U12635 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19151) );
  NAND2_X1 U12636 ( .A1(n10835), .A2(n10314), .ZN(n14506) );
  NAND2_X1 U12637 ( .A1(n15355), .A2(n10280), .ZN(n15337) );
  AND3_X1 U12638 ( .A1(n11747), .A2(n11619), .A3(n11746), .ZN(n9865) );
  INV_X1 U12639 ( .A(n10432), .ZN(n10406) );
  NAND2_X1 U12640 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11361), .ZN(
        n9866) );
  AND2_X1 U12641 ( .A1(n17766), .A2(n9991), .ZN(n9867) );
  INV_X2 U12642 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11619) );
  OR2_X1 U12643 ( .A1(n9857), .A2(n10163), .ZN(n9868) );
  NOR2_X1 U12644 ( .A1(n15404), .A2(n9856), .ZN(n12510) );
  XNOR2_X1 U12645 ( .A(n13190), .B(n13191), .ZN(n15161) );
  NAND2_X1 U12646 ( .A1(n14619), .A2(n10774), .ZN(n14615) );
  AND2_X1 U12647 ( .A1(n10056), .A2(n15629), .ZN(n9869) );
  OR2_X1 U12648 ( .A1(n14488), .A2(n10025), .ZN(n10023) );
  INV_X1 U12649 ( .A(n9974), .ZN(n14738) );
  NAND2_X1 U12650 ( .A1(n14739), .A2(n14740), .ZN(n9974) );
  OR2_X1 U12651 ( .A1(n17307), .A2(n17057), .ZN(n9870) );
  INV_X1 U12652 ( .A(n9972), .ZN(n14660) );
  AOI21_X1 U12653 ( .B1(n9974), .B2(n14729), .A(n9973), .ZN(n9972) );
  INV_X1 U12654 ( .A(n14162), .ZN(n13706) );
  AND2_X1 U12655 ( .A1(n11642), .A2(n11641), .ZN(n9871) );
  NAND2_X1 U12656 ( .A1(n12519), .A2(n9850), .ZN(n10115) );
  NAND2_X1 U12657 ( .A1(n15664), .A2(n10055), .ZN(n10151) );
  OR2_X1 U12658 ( .A1(n15662), .A2(n10149), .ZN(n9872) );
  INV_X1 U12659 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11600) );
  AND2_X1 U12660 ( .A1(n11298), .A2(n11297), .ZN(n9873) );
  AND2_X1 U12661 ( .A1(n11255), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9874) );
  INV_X1 U12662 ( .A(n18805), .ZN(n18801) );
  OR2_X1 U12663 ( .A1(n18788), .A2(n9988), .ZN(n18805) );
  OR2_X1 U12664 ( .A1(n14975), .A2(n14976), .ZN(n9876) );
  NOR2_X1 U12665 ( .A1(n15404), .A2(n10260), .ZN(n9877) );
  AND2_X1 U12666 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9878) );
  INV_X1 U12667 ( .A(n10271), .ZN(n15151) );
  NAND2_X1 U12668 ( .A1(n13216), .A2(n13215), .ZN(n10271) );
  AND3_X1 U12669 ( .A1(n11452), .A2(n10084), .A3(n10083), .ZN(n9879) );
  NOR3_X1 U12670 ( .A1(n14975), .A2(n14976), .A3(n15154), .ZN(n9880) );
  AND2_X1 U12671 ( .A1(n9878), .A2(n10184), .ZN(n9881) );
  AND2_X1 U12672 ( .A1(n9860), .A2(n15387), .ZN(n9882) );
  INV_X1 U12673 ( .A(n11404), .ZN(n10249) );
  INV_X1 U12674 ( .A(n12447), .ZN(n12130) );
  NAND2_X1 U12675 ( .A1(n12128), .A2(n12154), .ZN(n12447) );
  AND2_X1 U12676 ( .A1(n11812), .A2(n9948), .ZN(n11884) );
  INV_X1 U12677 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10324) );
  INV_X1 U12678 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18980) );
  OR2_X1 U12679 ( .A1(n11599), .A2(n11598), .ZN(P3_U2801) );
  INV_X1 U12680 ( .A(n10816), .ZN(n10308) );
  NAND2_X1 U12681 ( .A1(n10452), .A2(n20287), .ZN(n13562) );
  AND3_X1 U12682 ( .A1(n14057), .A2(n14102), .A3(n10315), .ZN(n14147) );
  AND2_X1 U12683 ( .A1(n14121), .A2(n14176), .ZN(n14174) );
  AND2_X1 U12684 ( .A1(n14121), .A2(n9971), .ZN(n15199) );
  NAND2_X1 U12685 ( .A1(n15218), .A2(n15217), .ZN(n15023) );
  AND2_X1 U12686 ( .A1(n17857), .A2(n18198), .ZN(n9884) );
  INV_X1 U12687 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20012) );
  AND2_X1 U12688 ( .A1(n14934), .A2(n10180), .ZN(n9885) );
  AND2_X1 U12689 ( .A1(n14923), .A2(n10187), .ZN(n9886) );
  INV_X1 U12690 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10010) );
  NOR2_X1 U12691 ( .A1(n14129), .A2(n12332), .ZN(n12803) );
  NAND2_X1 U12692 ( .A1(n14057), .A2(n14102), .ZN(n14101) );
  INV_X1 U12693 ( .A(n10336), .ZN(n12993) );
  NAND2_X1 U12694 ( .A1(n9952), .A2(n11229), .ZN(n13901) );
  AND2_X1 U12695 ( .A1(n17807), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9887) );
  INV_X1 U12696 ( .A(n17703), .ZN(n17885) );
  NOR2_X1 U12697 ( .A1(n13310), .A2(n17983), .ZN(n17703) );
  NOR2_X1 U12698 ( .A1(n13554), .A2(n10211), .ZN(n9888) );
  NAND2_X1 U12699 ( .A1(n12437), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15748) );
  INV_X1 U12700 ( .A(n15748), .ZN(n10042) );
  NOR2_X1 U12701 ( .A1(n14091), .A2(n14092), .ZN(n14090) );
  INV_X2 U12702 ( .A(n10432), .ZN(n10983) );
  NOR2_X1 U12703 ( .A1(n13554), .A2(n13553), .ZN(n9889) );
  AND2_X1 U12704 ( .A1(n10129), .A2(n10128), .ZN(n9890) );
  AND2_X1 U12705 ( .A1(n17766), .A2(n10346), .ZN(n9891) );
  AND2_X1 U12706 ( .A1(n15469), .A2(n15715), .ZN(n9892) );
  OR2_X1 U12707 ( .A1(n12553), .A2(n12812), .ZN(n9893) );
  NOR2_X1 U12708 ( .A1(n15197), .A2(n15184), .ZN(n12604) );
  INV_X1 U12709 ( .A(n11427), .ZN(n17727) );
  NAND2_X1 U12710 ( .A1(n9993), .A2(n17779), .ZN(n11427) );
  AND2_X1 U12711 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9894) );
  INV_X1 U12712 ( .A(n14108), .ZN(n10316) );
  AND4_X1 U12713 ( .A1(n10724), .A2(n10723), .A3(n10722), .A4(n10721), .ZN(
        n14108) );
  NAND2_X1 U12714 ( .A1(n14438), .A2(n14421), .ZN(n9895) );
  NAND2_X1 U12715 ( .A1(n14086), .A2(n14088), .ZN(n9896) );
  INV_X1 U12716 ( .A(n10015), .ZN(n10014) );
  NAND2_X1 U12717 ( .A1(n10016), .A2(n14616), .ZN(n10015) );
  NOR2_X1 U12718 ( .A1(n14507), .A2(n10313), .ZN(n10312) );
  INV_X1 U12719 ( .A(n13908), .ZN(n12996) );
  OR2_X1 U12720 ( .A1(n12255), .A2(n12254), .ZN(n13908) );
  AND3_X1 U12721 ( .A1(n12004), .A2(n12026), .A3(n12222), .ZN(n9897) );
  AND2_X1 U12722 ( .A1(n10184), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9898) );
  AND2_X1 U12723 ( .A1(n12805), .A2(n12804), .ZN(n15026) );
  AND2_X1 U12724 ( .A1(n10315), .A2(n14184), .ZN(n9899) );
  AND2_X1 U12725 ( .A1(n11294), .A2(n14839), .ZN(n9900) );
  NOR2_X1 U12726 ( .A1(n15175), .A2(n15174), .ZN(n9901) );
  OR2_X1 U12727 ( .A1(n13508), .A2(n13507), .ZN(n13506) );
  NAND2_X1 U12728 ( .A1(n12785), .A2(n12408), .ZN(n9902) );
  AND2_X1 U12729 ( .A1(n10014), .A2(n10772), .ZN(n9903) );
  AND2_X1 U12730 ( .A1(n10172), .A2(n10171), .ZN(n9904) );
  NAND2_X1 U12731 ( .A1(n19016), .A2(n15813), .ZN(n18809) );
  INV_X1 U12732 ( .A(n18809), .ZN(n10076) );
  NOR2_X1 U12733 ( .A1(n13834), .A2(n10276), .ZN(n13895) );
  NOR2_X1 U12734 ( .A1(n13834), .A2(n10274), .ZN(n14002) );
  OR2_X1 U12735 ( .A1(n11625), .A2(n11624), .ZN(n12222) );
  INV_X1 U12736 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10576) );
  INV_X1 U12737 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10009) );
  NAND2_X1 U12738 ( .A1(n17640), .A2(n9828), .ZN(n9905) );
  AND2_X1 U12739 ( .A1(n12549), .A2(n10114), .ZN(n9906) );
  INV_X1 U12740 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20028) );
  NAND2_X1 U12741 ( .A1(n12785), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n9907) );
  AND2_X1 U12742 ( .A1(n13537), .A2(n12215), .ZN(n9908) );
  NAND2_X1 U12743 ( .A1(n10019), .A2(n10538), .ZN(n20312) );
  NAND2_X1 U12744 ( .A1(n9963), .A2(n9848), .ZN(n14120) );
  INV_X1 U12745 ( .A(n17779), .ZN(n17877) );
  NAND2_X1 U12746 ( .A1(n16519), .A2(n13310), .ZN(n17779) );
  OR2_X1 U12747 ( .A1(n14528), .A2(n10168), .ZN(n9909) );
  NOR2_X1 U12748 ( .A1(n17909), .A2(n17908), .ZN(n9910) );
  INV_X1 U12749 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U12750 ( .A1(n14916), .A2(n9851), .ZN(n10182) );
  NAND2_X1 U12751 ( .A1(n9979), .A2(n9977), .ZN(n9981) );
  AND2_X1 U12752 ( .A1(n9963), .A2(n12186), .ZN(n9911) );
  NAND2_X1 U12753 ( .A1(n10254), .A2(n10253), .ZN(n9912) );
  AND2_X1 U12754 ( .A1(n12215), .A2(n10191), .ZN(n9913) );
  AND2_X2 U12755 ( .A1(n20274), .A2(n20287), .ZN(n13566) );
  AND2_X1 U12756 ( .A1(n12345), .A2(n12348), .ZN(n9914) );
  AND2_X1 U12757 ( .A1(n9851), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9915) );
  INV_X1 U12758 ( .A(n10199), .ZN(n10198) );
  NAND2_X1 U12759 ( .A1(n12820), .A2(n10200), .ZN(n10199) );
  INV_X1 U12760 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20936) );
  AND2_X1 U12761 ( .A1(n13137), .A2(n13136), .ZN(n9916) );
  NOR2_X1 U12762 ( .A1(n16172), .A2(n16171), .ZN(n9917) );
  INV_X1 U12763 ( .A(n18846), .ZN(n19004) );
  NAND2_X2 U12764 ( .A1(n15768), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15774) );
  AND2_X1 U12765 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9918) );
  AND2_X1 U12766 ( .A1(n18198), .A2(n10246), .ZN(n9919) );
  AND3_X1 U12767 ( .A1(n10157), .A2(n13925), .A3(n10156), .ZN(n9920) );
  OR2_X1 U12768 ( .A1(n12174), .A2(n12624), .ZN(n9921) );
  INV_X1 U12769 ( .A(n13918), .ZN(n10156) );
  INV_X1 U12770 ( .A(n15158), .ZN(n10272) );
  AND2_X1 U12771 ( .A1(n10162), .A2(n10161), .ZN(n9922) );
  NAND2_X1 U12772 ( .A1(n18000), .A2(n16506), .ZN(n9923) );
  AND2_X1 U12773 ( .A1(n9854), .A2(n17819), .ZN(n9924) );
  AND2_X1 U12774 ( .A1(n9853), .A2(n10110), .ZN(n9925) );
  INV_X1 U12775 ( .A(n17701), .ZN(n10007) );
  INV_X1 U12776 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10178) );
  AND2_X1 U12777 ( .A1(n12665), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14609)
         );
  AND2_X1 U12778 ( .A1(n17758), .A2(n10029), .ZN(n9926) );
  AND4_X1 U12779 ( .A1(n16085), .A2(n14794), .A3(n11291), .A4(n14884), .ZN(
        n9927) );
  AND2_X1 U12780 ( .A1(n15609), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9928) );
  NAND2_X1 U12781 ( .A1(n10280), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9929) );
  INV_X1 U12782 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10114) );
  INV_X1 U12783 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10113) );
  INV_X1 U12784 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10110) );
  NAND3_X1 U12785 ( .A1(n11279), .A2(n11278), .A3(n11280), .ZN(n9930) );
  INV_X1 U12786 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10281) );
  INV_X1 U12787 ( .A(n10240), .ZN(n10237) );
  AND2_X1 U12788 ( .A1(n15520), .A2(n15508), .ZN(n10240) );
  OR2_X1 U12789 ( .A1(n9856), .A2(n15492), .ZN(n9931) );
  INV_X1 U12790 ( .A(n16380), .ZN(n10048) );
  INV_X1 U12791 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10181) );
  INV_X1 U12792 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10030) );
  AND2_X1 U12793 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9932) );
  OAI22_X2 U12794 ( .A1(n14560), .A2(n20306), .B1(n20272), .B2(n20304), .ZN(
        n20787) );
  OAI22_X2 U12795 ( .A1(n19363), .A2(n20306), .B1(n21021), .B2(n20304), .ZN(
        n20827) );
  NOR3_X2 U12796 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18849), .A3(
        n18401), .ZN(n18371) );
  NOR3_X2 U12797 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18849), .A3(
        n18467), .ZN(n18462) );
  NOR4_X2 U12798 ( .A1(n16085), .A2(n16121), .A3(n16109), .A4(n16078), .ZN(
        n15889) );
  OAI22_X2 U12799 ( .A1(n14540), .A2(n20306), .B1(n20293), .B2(n20304), .ZN(
        n20754) );
  OAI22_X2 U12800 ( .A1(n20268), .A2(n20306), .B1(n21073), .B2(n20304), .ZN(
        n20781) );
  NAND2_X1 U12801 ( .A1(n16001), .A2(n14609), .ZN(n20306) );
  NOR3_X2 U12802 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18849), .A3(
        n18558), .ZN(n18553) );
  INV_X2 U12803 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18987) );
  NAND4_X2 U12804 ( .A1(n18980), .A2(n18972), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17296) );
  OR2_X1 U12805 ( .A1(n15539), .A2(n19278), .ZN(n9940) );
  NOR2_X2 U12806 ( .A1(n15404), .A2(n9855), .ZN(n15355) );
  OR2_X2 U12807 ( .A1(n15417), .A2(n9941), .ZN(n15404) );
  AND2_X2 U12808 ( .A1(n11874), .A2(n13344), .ZN(n12169) );
  NAND2_X1 U12809 ( .A1(n11873), .A2(n20055), .ZN(n13344) );
  NAND2_X1 U12810 ( .A1(n13412), .A2(n11815), .ZN(n11874) );
  AND3_X2 U12811 ( .A1(n11814), .A2(n11875), .A3(n11813), .ZN(n13412) );
  NAND2_X1 U12812 ( .A1(n11876), .A2(n11875), .ZN(n9944) );
  NAND2_X1 U12813 ( .A1(n12341), .A2(n9946), .ZN(n10121) );
  XNOR2_X2 U12814 ( .A(n12341), .B(n9946), .ZN(n12956) );
  XNOR2_X2 U12815 ( .A(n12342), .B(n12343), .ZN(n9946) );
  XNOR2_X2 U12816 ( .A(n12038), .B(n12037), .ZN(n12414) );
  NAND2_X2 U12817 ( .A1(n9950), .A2(n12004), .ZN(n12038) );
  OR2_X2 U12818 ( .A1(n12006), .A2(n12005), .ZN(n9950) );
  NAND2_X2 U12819 ( .A1(n9947), .A2(n11973), .ZN(n12046) );
  NAND2_X1 U12820 ( .A1(n10230), .A2(n9947), .ZN(n11957) );
  INV_X2 U12821 ( .A(n11972), .ZN(n9947) );
  XNOR2_X2 U12822 ( .A(n12158), .B(n12156), .ZN(n15712) );
  NAND2_X2 U12823 ( .A1(n15479), .A2(n12132), .ZN(n12158) );
  NAND2_X1 U12824 ( .A1(n11897), .A2(n12173), .ZN(n11885) );
  INV_X2 U12825 ( .A(n11820), .ZN(n9948) );
  AOI21_X2 U12826 ( .B1(n15425), .B2(n15423), .A(n15398), .ZN(n15415) );
  AND2_X2 U12827 ( .A1(n15439), .A2(n15436), .ZN(n15425) );
  OR2_X2 U12828 ( .A1(n15696), .A2(n15693), .ZN(n9951) );
  NAND2_X1 U12829 ( .A1(n13851), .A2(n13852), .ZN(n9952) );
  NAND2_X1 U12830 ( .A1(n9953), .A2(n11227), .ZN(n13851) );
  NAND2_X1 U12831 ( .A1(n13748), .A2(n13749), .ZN(n9953) );
  NAND2_X1 U12832 ( .A1(n9954), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n9956) );
  NAND2_X1 U12833 ( .A1(n11949), .A2(n11954), .ZN(n9955) );
  XNOR2_X1 U12834 ( .A(n11922), .B(n11921), .ZN(n11949) );
  OAI21_X2 U12835 ( .B1(n11938), .B2(n15783), .A(n10137), .ZN(n11921) );
  INV_X1 U12836 ( .A(n13834), .ZN(n9963) );
  NAND3_X1 U12837 ( .A1(n13789), .A2(n12993), .A3(n13788), .ZN(n9967) );
  NAND2_X2 U12838 ( .A1(n11288), .A2(n11289), .ZN(n14739) );
  XNOR2_X2 U12839 ( .A(n9976), .B(n10589), .ZN(n20338) );
  INV_X2 U12840 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18972) );
  INV_X1 U12841 ( .A(n9981), .ZN(n17466) );
  INV_X1 U12842 ( .A(n17356), .ZN(n17361) );
  NAND3_X1 U12843 ( .A1(n9867), .A2(n11421), .A3(n11426), .ZN(n9990) );
  INV_X1 U12844 ( .A(n9993), .ZN(n17756) );
  NAND3_X1 U12845 ( .A1(n10329), .A2(n10000), .A3(n11316), .ZN(n11317) );
  NAND3_X1 U12846 ( .A1(n11315), .A2(n11313), .A3(n10003), .ZN(n10002) );
  NAND3_X1 U12847 ( .A1(n10006), .A2(n9836), .A3(n9866), .ZN(n10005) );
  NOR2_X1 U12848 ( .A1(n17943), .A2(n17942), .ZN(n17941) );
  INV_X1 U12849 ( .A(n10006), .ZN(n17953) );
  AND2_X1 U12850 ( .A1(n11422), .A2(n10007), .ZN(n17710) );
  NOR2_X2 U12851 ( .A1(n17792), .A2(n18112), .ZN(n11422) );
  AND2_X2 U12852 ( .A1(n13942), .A2(n10368), .ZN(n10412) );
  XNOR2_X2 U12853 ( .A(n10537), .B(n10483), .ZN(n10591) );
  NAND2_X1 U12854 ( .A1(n10544), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10011) );
  AOI21_X1 U12855 ( .B1(n10773), .B2(n9903), .A(n10013), .ZN(n10012) );
  AND2_X2 U12856 ( .A1(n10395), .A2(n10017), .ZN(n10477) );
  NAND4_X1 U12857 ( .A1(n10469), .A2(n13706), .A3(n10450), .A4(n10017), .ZN(
        n13624) );
  NAND2_X1 U12858 ( .A1(n10017), .A2(n10574), .ZN(n13792) );
  AND2_X1 U12859 ( .A1(n14169), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10672) );
  NAND2_X1 U12860 ( .A1(n10017), .A2(n13706), .ZN(n10430) );
  NAND2_X1 U12861 ( .A1(n10461), .A2(n10017), .ZN(n13795) );
  OAI21_X1 U12862 ( .B1(n13680), .B2(n10574), .A(n10017), .ZN(n13564) );
  NAND2_X1 U12863 ( .A1(n20179), .A2(n10017), .ZN(n14532) );
  NAND2_X1 U12864 ( .A1(n20312), .A2(n10558), .ZN(n13559) );
  NAND3_X1 U12865 ( .A1(n20312), .A2(n10558), .A3(n20936), .ZN(n10018) );
  INV_X1 U12866 ( .A(n20378), .ZN(n10019) );
  AOI21_X1 U12867 ( .B1(n10983), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n10021), .ZN(n10020) );
  INV_X1 U12868 ( .A(n14488), .ZN(n10835) );
  INV_X1 U12869 ( .A(n10312), .ZN(n10025) );
  XNOR2_X2 U12870 ( .A(n10026), .B(n10573), .ZN(n10601) );
  OAI22_X2 U12871 ( .A1(n13608), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11220), 
        .B2(n10570), .ZN(n10026) );
  INV_X1 U12872 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10032) );
  INV_X1 U12873 ( .A(n10034), .ZN(n16746) );
  INV_X1 U12874 ( .A(n10033), .ZN(n16745) );
  NAND2_X1 U12875 ( .A1(n10034), .A2(n17681), .ZN(n10033) );
  OR2_X1 U12876 ( .A1(n16760), .A2(n16985), .ZN(n10034) );
  NOR2_X1 U12877 ( .A1(n16679), .A2(n16985), .ZN(n16671) );
  OR2_X2 U12878 ( .A1(n15764), .A2(n12956), .ZN(n11985) );
  NAND3_X1 U12879 ( .A1(n13549), .A2(n10039), .A3(n11973), .ZN(n12044) );
  INV_X1 U12880 ( .A(n12956), .ZN(n10039) );
  NAND2_X2 U12881 ( .A1(n15746), .A2(n15747), .ZN(n15745) );
  NAND2_X1 U12882 ( .A1(n12043), .A2(n12042), .ZN(n15746) );
  NAND2_X1 U12883 ( .A1(n10044), .A2(n15745), .ZN(n10040) );
  NAND3_X1 U12884 ( .A1(n15746), .A2(n12447), .A3(n15747), .ZN(n10043) );
  AND2_X1 U12885 ( .A1(n12130), .A2(n15748), .ZN(n10044) );
  AND2_X1 U12886 ( .A1(n10046), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10050) );
  NAND4_X2 U12887 ( .A1(n10049), .A2(n10046), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A4(n10048), .ZN(n16316) );
  OR2_X2 U12888 ( .A1(n10147), .A2(n10051), .ZN(n10046) );
  INV_X1 U12890 ( .A(n10151), .ZN(n15459) );
  NAND2_X2 U12891 ( .A1(n12158), .A2(n12157), .ZN(n12159) );
  INV_X1 U12892 ( .A(n12090), .ZN(n12091) );
  NAND2_X1 U12893 ( .A1(n15389), .A2(n9882), .ZN(n10062) );
  NOR2_X1 U12894 ( .A1(n10066), .A2(n9860), .ZN(n15575) );
  OAI21_X2 U12895 ( .B1(n12414), .B2(n12788), .A(n15114), .ZN(n12427) );
  OAI21_X2 U12896 ( .B1(n18805), .B2(n10082), .A(n11540), .ZN(n18814) );
  AOI21_X2 U12897 ( .B1(n11538), .B2(n18790), .A(n13300), .ZN(n11540) );
  NAND3_X1 U12898 ( .A1(n10088), .A2(n11454), .A3(n9879), .ZN(n11455) );
  INV_X1 U12899 ( .A(n14636), .ZN(n10090) );
  NOR2_X2 U12900 ( .A1(n14635), .A2(n11295), .ZN(n14629) );
  NAND2_X1 U12901 ( .A1(n10090), .A2(n10091), .ZN(n10093) );
  NAND2_X1 U12902 ( .A1(n14629), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10094) );
  NAND2_X1 U12903 ( .A1(n10668), .A2(n10669), .ZN(n10698) );
  NAND3_X1 U12904 ( .A1(n11266), .A2(n11251), .A3(n11230), .ZN(n11254) );
  NAND2_X1 U12906 ( .A1(n20274), .A2(n20266), .ZN(n14028) );
  NAND3_X1 U12907 ( .A1(n14704), .A2(n10097), .A3(n10098), .ZN(n14676) );
  NAND2_X1 U12908 ( .A1(n14138), .A2(n11271), .ZN(n11273) );
  NAND2_X1 U12909 ( .A1(n10100), .A2(n16017), .ZN(n14138) );
  NAND2_X1 U12910 ( .A1(n16016), .A2(n16018), .ZN(n10100) );
  AOI21_X2 U12911 ( .B1(n14780), .B2(n10101), .A(n10343), .ZN(n11288) );
  AND2_X1 U12912 ( .A1(n12579), .A2(n9925), .ZN(n12786) );
  INV_X1 U12913 ( .A(n10115), .ZN(n12562) );
  NOR2_X4 U12914 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16446) );
  NAND2_X1 U12915 ( .A1(n10117), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10116) );
  NAND4_X1 U12916 ( .A1(n11605), .A2(n11602), .A3(n11603), .A4(n11604), .ZN(
        n10117) );
  NAND2_X1 U12917 ( .A1(n10119), .A2(n11619), .ZN(n10118) );
  NAND4_X1 U12918 ( .A1(n11609), .A2(n11607), .A3(n11608), .A4(n11606), .ZN(
        n10119) );
  NAND2_X1 U12919 ( .A1(n15165), .A2(n15164), .ZN(n14975) );
  INV_X1 U12920 ( .A(n13910), .ZN(n10131) );
  NAND2_X1 U12921 ( .A1(n10131), .A2(n10132), .ZN(n14091) );
  NAND2_X1 U12922 ( .A1(n10140), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U12923 ( .A1(n11916), .A2(n10141), .ZN(n10140) );
  NAND2_X1 U12924 ( .A1(n11893), .A2(n11863), .ZN(n10141) );
  NAND4_X1 U12925 ( .A1(n12023), .A2(n12021), .A3(n12022), .A4(n12024), .ZN(
        n10142) );
  NAND2_X2 U12926 ( .A1(n10144), .A2(n10143), .ZN(n12957) );
  NAND3_X1 U12927 ( .A1(n10341), .A2(n11752), .A3(n11751), .ZN(n10143) );
  NAND4_X1 U12928 ( .A1(n11763), .A2(n11761), .A3(n11762), .A4(n11764), .ZN(
        n10145) );
  NAND4_X1 U12929 ( .A1(n11757), .A2(n11756), .A3(n11755), .A4(n11754), .ZN(
        n10146) );
  AOI21_X2 U12930 ( .B1(n12159), .B2(n15719), .A(n10148), .ZN(n10147) );
  NAND2_X1 U12931 ( .A1(n10155), .A2(n20281), .ZN(n13560) );
  AND2_X1 U12932 ( .A1(n13706), .A2(n10155), .ZN(n10607) );
  NAND2_X1 U12933 ( .A1(n12678), .A2(n10155), .ZN(n12704) );
  NAND2_X1 U12934 ( .A1(n12878), .A2(n10155), .ZN(n13453) );
  OAI21_X1 U12935 ( .B1(n12878), .B2(n21166), .A(n10155), .ZN(n10153) );
  NAND2_X1 U12936 ( .A1(n13572), .A2(n10155), .ZN(n12640) );
  AND2_X1 U12937 ( .A1(n13684), .A2(n10155), .ZN(n13567) );
  AND2_X1 U12938 ( .A1(n13792), .A2(n10155), .ZN(n10154) );
  NAND2_X1 U12939 ( .A1(n20180), .A2(n10155), .ZN(n13880) );
  NAND3_X1 U12940 ( .A1(n10160), .A2(n10156), .A3(n13925), .ZN(n10159) );
  NAND2_X1 U12941 ( .A1(n16170), .A2(n9904), .ZN(n16147) );
  AND2_X2 U12942 ( .A1(n10177), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10363) );
  NAND2_X1 U12943 ( .A1(n14916), .A2(n9915), .ZN(n14913) );
  INV_X1 U12944 ( .A(n10182), .ZN(n14914) );
  INV_X1 U12945 ( .A(n14924), .ZN(n10183) );
  NAND2_X1 U12946 ( .A1(n10183), .A2(n9881), .ZN(n14927) );
  NAND2_X1 U12947 ( .A1(n13533), .A2(n13534), .ZN(n13537) );
  NOR2_X1 U12948 ( .A1(n15316), .A2(n10192), .ZN(n15008) );
  NOR2_X2 U12949 ( .A1(n15569), .A2(n10197), .ZN(n14983) );
  NAND3_X1 U12950 ( .A1(n11636), .A2(n11635), .A3(n11634), .ZN(n10215) );
  NAND3_X1 U12951 ( .A1(n10218), .A2(n11640), .A3(n11639), .ZN(n10217) );
  AND2_X1 U12952 ( .A1(n11637), .A2(n11638), .ZN(n10218) );
  OAI211_X1 U12953 ( .C1(n12892), .C2(n10225), .A(n10223), .B(n10222), .ZN(
        n12955) );
  AND3_X4 U12954 ( .A1(n10229), .A2(n11600), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13280) );
  NAND3_X1 U12955 ( .A1(n10232), .A2(n15334), .A3(n10231), .ZN(n10233) );
  NAND3_X1 U12956 ( .A1(n10235), .A2(n10238), .A3(n9932), .ZN(n10234) );
  AND2_X1 U12957 ( .A1(n15353), .A2(n15358), .ZN(n10241) );
  NAND2_X2 U12958 ( .A1(n17639), .A2(n17649), .ZN(n17638) );
  NAND2_X1 U12959 ( .A1(n10255), .A2(n17638), .ZN(n11435) );
  AND3_X1 U12960 ( .A1(n10255), .A2(n17638), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17627) );
  AND2_X2 U12961 ( .A1(n11427), .A2(n10256), .ZN(n17752) );
  NAND2_X1 U12962 ( .A1(n10257), .A2(n11934), .ZN(n11937) );
  XNOR2_X1 U12963 ( .A(n11948), .B(n10257), .ZN(n12968) );
  OAI21_X1 U12964 ( .B1(n12092), .B2(n12091), .A(n10258), .ZN(n12128) );
  INV_X1 U12965 ( .A(n12129), .ZN(n10258) );
  NOR2_X1 U12966 ( .A1(n15404), .A2(n15405), .ZN(n15386) );
  OAI21_X1 U12967 ( .B1(n13216), .B2(n10269), .A(n10266), .ZN(n15146) );
  AND2_X4 U12968 ( .A1(n10363), .A2(n13941), .ZN(n11068) );
  AND2_X2 U12969 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13941) );
  NAND2_X1 U12970 ( .A1(n10429), .A2(n14162), .ZN(n13568) );
  NOR2_X1 U12971 ( .A1(n12771), .A2(n10429), .ZN(n10282) );
  AND2_X2 U12972 ( .A1(n10477), .A2(n10405), .ZN(n10429) );
  NAND2_X1 U12973 ( .A1(n14662), .A2(n14838), .ZN(n14635) );
  INV_X1 U12974 ( .A(n14662), .ZN(n10286) );
  NAND2_X1 U12975 ( .A1(n14671), .A2(n11293), .ZN(n14662) );
  NAND3_X1 U12976 ( .A1(n11288), .A2(n9927), .A3(n11289), .ZN(n10288) );
  NAND2_X1 U12977 ( .A1(n10591), .A2(n20936), .ZN(n10294) );
  NAND2_X1 U12978 ( .A1(n10507), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10296) );
  INV_X1 U12979 ( .A(n10507), .ZN(n10297) );
  NAND2_X1 U12980 ( .A1(n14190), .A2(n10300), .ZN(n10298) );
  NAND2_X1 U12981 ( .A1(n10298), .A2(n10299), .ZN(n11281) );
  INV_X1 U12982 ( .A(n10582), .ZN(n10303) );
  NAND2_X1 U12983 ( .A1(n10304), .A2(n10541), .ZN(n10582) );
  NAND2_X1 U12984 ( .A1(n10530), .A2(n10529), .ZN(n10541) );
  NAND2_X1 U12985 ( .A1(n10305), .A2(n10526), .ZN(n10304) );
  XNOR2_X2 U12987 ( .A(n10600), .B(n10601), .ZN(n11217) );
  AND3_X2 U12988 ( .A1(n14057), .A2(n14102), .A3(n9899), .ZN(n10760) );
  NAND3_X1 U12989 ( .A1(n14057), .A2(n14102), .A3(n10316), .ZN(n10317) );
  INV_X1 U12990 ( .A(n10317), .ZN(n14107) );
  NAND2_X1 U12991 ( .A1(n14352), .A2(n10320), .ZN(n14327) );
  INV_X1 U12992 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10323) );
  INV_X1 U12993 ( .A(n9807), .ZN(n15758) );
  INV_X1 U12994 ( .A(n12909), .ZN(n12910) );
  INV_X1 U12995 ( .A(n12943), .ZN(n12944) );
  OAI21_X1 U12996 ( .B1(n12942), .B2(n19277), .A(n12941), .ZN(n12943) );
  NAND2_X1 U12997 ( .A1(n11981), .A2(n11980), .ZN(n12050) );
  AOI211_X2 U12998 ( .C1(n15502), .C2(n16413), .A(n15501), .B(n15500), .ZN(
        n15503) );
  OAI22_X1 U12999 ( .A1(n12977), .A2(n12064), .B1(n12050), .B2(n11982), .ZN(
        n11983) );
  NAND2_X1 U13000 ( .A1(n13810), .A2(n10599), .ZN(n13855) );
  INV_X1 U13001 ( .A(n13562), .ZN(n10428) );
  NOR2_X1 U13002 ( .A1(n12055), .A2(n13123), .ZN(n11987) );
  NAND2_X1 U13003 ( .A1(n11981), .A2(n11956), .ZN(n12047) );
  AOI21_X2 U13004 ( .B1(n12555), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15382), .ZN(n15373) );
  AND2_X2 U13005 ( .A1(n10370), .A2(n13612), .ZN(n10350) );
  OR2_X1 U13006 ( .A1(n12946), .A2(n19277), .ZN(n12954) );
  OR4_X2 U13007 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(n18987), .ZN(n10328) );
  OR2_X2 U13008 ( .A1(n15974), .A2(n13793), .ZN(n14624) );
  AND2_X1 U13009 ( .A1(n11299), .A2(n10338), .ZN(n10329) );
  OR2_X1 U13010 ( .A1(n20179), .A2(n14319), .ZN(n10330) );
  AND2_X1 U13011 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10333) );
  AND2_X1 U13012 ( .A1(n11851), .A2(n11852), .ZN(n10334) );
  INV_X2 U13013 ( .A(n18997), .ZN(n18936) );
  OR2_X1 U13014 ( .A1(n13325), .A2(n17984), .ZN(n10335) );
  INV_X1 U13015 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20097) );
  OR2_X1 U13016 ( .A1(n13213), .A2(n11613), .ZN(n10336) );
  AND3_X1 U13017 ( .A1(n18139), .A2(n11418), .A3(n18112), .ZN(n10337) );
  INV_X1 U13018 ( .A(n14489), .ZN(n10834) );
  AND2_X1 U13019 ( .A1(n10642), .A2(n10641), .ZN(n10339) );
  INV_X1 U13020 ( .A(n17488), .ZN(n17408) );
  NAND2_X2 U13021 ( .A1(n15911), .A2(n17393), .ZN(n17488) );
  NAND2_X2 U13022 ( .A1(n20179), .A2(n14169), .ZN(n14521) );
  OR2_X1 U13023 ( .A1(n15488), .A2(n19277), .ZN(n10340) );
  NAND2_X1 U13024 ( .A1(n17693), .A2(n17979), .ZN(n17721) );
  AND3_X1 U13025 ( .A1(n11750), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11749), .ZN(n10341) );
  NAND2_X1 U13026 ( .A1(n20274), .A2(n10450), .ZN(n11239) );
  INV_X1 U13027 ( .A(n11317), .ZN(n17489) );
  OR2_X1 U13028 ( .A1(n12535), .A2(n15456), .ZN(n10342) );
  INV_X1 U13029 ( .A(n11984), .ZN(n11966) );
  OR2_X1 U13030 ( .A1(n14749), .A2(n14770), .ZN(n10343) );
  AND2_X1 U13031 ( .A1(n11745), .A2(n11744), .ZN(n10344) );
  NAND2_X1 U13032 ( .A1(n12817), .A2(n12816), .ZN(n10345) );
  INV_X1 U13033 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20617) );
  OR2_X1 U13034 ( .A1(n17779), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10346) );
  NAND2_X1 U13035 ( .A1(n12585), .A2(n20060), .ZN(n19278) );
  BUF_X1 U13036 ( .A(n11812), .Z(n19341) );
  AND2_X1 U13037 ( .A1(n11135), .A2(n20698), .ZN(n16025) );
  INV_X1 U13038 ( .A(n20179), .ZN(n14530) );
  AND2_X2 U13039 ( .A1(n12677), .A2(n13690), .ZN(n20179) );
  OR2_X1 U13040 ( .A1(n13650), .A2(n15859), .ZN(n20080) );
  INV_X1 U13041 ( .A(n16515), .ZN(n18199) );
  NAND2_X1 U13042 ( .A1(n17344), .A2(n17393), .ZN(n17336) );
  NOR2_X1 U13043 ( .A1(n20578), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10347) );
  INV_X1 U13044 ( .A(n12187), .ZN(n12811) );
  AND2_X1 U13045 ( .A1(n13294), .A2(n13293), .ZN(n10348) );
  INV_X1 U13046 ( .A(n11975), .ZN(n11956) );
  INV_X1 U13047 ( .A(n10350), .ZN(n13938) );
  AND4_X1 U13048 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10351) );
  INV_X1 U13049 ( .A(n10672), .ZN(n10707) );
  AND4_X1 U13050 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n10353) );
  AND4_X1 U13051 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10354) );
  AND2_X2 U13052 ( .A1(n10369), .A2(n13612), .ZN(n10407) );
  OR2_X1 U13053 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11143), .ZN(
        n11142) );
  NAND2_X1 U13054 ( .A1(n11848), .A2(n11812), .ZN(n11840) );
  OR2_X1 U13055 ( .A1(n11160), .A2(n11161), .ZN(n11141) );
  NAND2_X1 U13056 ( .A1(n10450), .A2(n10574), .ZN(n10451) );
  INV_X1 U13057 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13940) );
  OAI21_X1 U13058 ( .B1(n11671), .B2(n11628), .A(n11669), .ZN(n11667) );
  OAI22_X1 U13059 ( .A1(n13170), .A2(n12054), .B1(n12055), .B2(n13179), .ZN(
        n12011) );
  OAI22_X1 U13060 ( .A1(n11960), .A2(n12058), .B1(n12061), .B2(n13112), .ZN(
        n11961) );
  AOI22_X1 U13061 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13275), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11739) );
  OR2_X1 U13062 ( .A1(n10993), .A2(n10992), .ZN(n11005) );
  NAND2_X1 U13063 ( .A1(n10452), .A2(n10451), .ZN(n10453) );
  INV_X1 U13064 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U13065 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U13066 ( .A1(n11675), .A2(n11627), .ZN(n11671) );
  OR2_X1 U13067 ( .A1(n11667), .A2(n11665), .ZN(n11630) );
  AND2_X1 U13068 ( .A1(n11753), .A2(n11619), .ZN(n11756) );
  AND2_X1 U13069 ( .A1(n11181), .A2(n11180), .ZN(n12647) );
  INV_X1 U13070 ( .A(n15925), .ZN(n10853) );
  INV_X1 U13071 ( .A(n14392), .ZN(n11004) );
  OAI21_X1 U13072 ( .B1(n10707), .B2(n10706), .A(n10705), .ZN(n10708) );
  INV_X1 U13073 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10622) );
  OR2_X1 U13074 ( .A1(n10494), .A2(n10493), .ZN(n11267) );
  OR2_X1 U13075 ( .A1(n10665), .A2(n10664), .ZN(n11244) );
  NAND2_X1 U13076 ( .A1(n13792), .A2(n10430), .ZN(n10455) );
  AOI21_X1 U13077 ( .B1(n11150), .B2(n11149), .A(n11146), .ZN(n11181) );
  INV_X1 U13078 ( .A(n15212), .ZN(n13043) );
  NAND2_X1 U13079 ( .A1(n12360), .A2(n15761), .ZN(n11900) );
  NAND2_X1 U13080 ( .A1(n11735), .A2(n11619), .ZN(n11742) );
  OR2_X1 U13081 ( .A1(n11442), .A2(n11443), .ZN(n11438) );
  INV_X1 U13082 ( .A(n10935), .ZN(n10936) );
  NAND2_X1 U13083 ( .A1(n10760), .A2(n10759), .ZN(n10774) );
  INV_X1 U13084 ( .A(n10998), .ZN(n10999) );
  INV_X1 U13085 ( .A(n14450), .ZN(n10920) );
  INV_X1 U13086 ( .A(n14621), .ZN(n10772) );
  AND2_X1 U13087 ( .A1(n10691), .A2(n10690), .ZN(n10699) );
  INV_X1 U13088 ( .A(n12745), .ZN(n12762) );
  INV_X1 U13089 ( .A(n11239), .ZN(n11230) );
  NOR2_X1 U13090 ( .A1(n10569), .A2(n10568), .ZN(n11220) );
  INV_X1 U13091 ( .A(n11176), .ZN(n11185) );
  AND2_X1 U13092 ( .A1(n14004), .A2(n14003), .ZN(n12997) );
  INV_X1 U13093 ( .A(n12904), .ZN(n12905) );
  INV_X1 U13094 ( .A(n12003), .ZN(n12209) );
  INV_X1 U13095 ( .A(n11518), .ZN(n11450) );
  INV_X1 U13096 ( .A(n16522), .ZN(n11592) );
  AND2_X1 U13097 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11403), .ZN(
        n11404) );
  INV_X1 U13098 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17146) );
  INV_X1 U13099 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17045) );
  AND2_X1 U13100 ( .A1(n10936), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10937) );
  OR2_X1 U13101 ( .A1(n10553), .A2(n10554), .ZN(n10551) );
  AND3_X1 U13102 ( .A1(n13580), .A2(n10428), .A3(n13709), .ZN(n13696) );
  OR2_X1 U13103 ( .A1(n11130), .A2(n14639), .ZN(n11136) );
  NAND2_X1 U13104 ( .A1(n13580), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11128) );
  NAND2_X1 U13105 ( .A1(n10819), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10836) );
  INV_X1 U13106 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11143) );
  OR2_X1 U13107 ( .A1(n13958), .A2(n13957), .ZN(n15856) );
  INV_X1 U13108 ( .A(n14913), .ZN(n12631) );
  NAND2_X1 U13109 ( .A1(n12456), .A2(n12454), .ZN(n12453) );
  AND2_X1 U13110 ( .A1(n13159), .A2(n13158), .ZN(n13162) );
  AND2_X1 U13111 ( .A1(n20054), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12978) );
  INV_X1 U13112 ( .A(n15329), .ZN(n12577) );
  NOR2_X1 U13113 ( .A1(n12546), .A2(n12545), .ZN(n12547) );
  INV_X2 U13114 ( .A(n12153), .ZN(n12788) );
  INV_X1 U13116 ( .A(n15752), .ZN(n16451) );
  INV_X1 U13117 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14243) );
  INV_X1 U13118 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17258) );
  INV_X1 U13119 ( .A(n12913), .ZN(n12920) );
  AND2_X1 U13120 ( .A1(n17877), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11434) );
  NAND2_X1 U13121 ( .A1(n18026), .A2(n11425), .ZN(n11426) );
  INV_X1 U13122 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U13123 ( .A1(n10606), .A2(n10605), .ZN(n20411) );
  AND2_X1 U13124 ( .A1(n12703), .A2(n12702), .ZN(n16169) );
  INV_X1 U13125 ( .A(n13651), .ZN(n13628) );
  XNOR2_X1 U13126 ( .A(n11138), .B(n12880), .ZN(n14030) );
  NAND2_X1 U13127 ( .A1(n11080), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11130) );
  INV_X1 U13128 ( .A(n10621), .ZN(n11041) );
  NOR2_X1 U13129 ( .A1(n10804), .A2(n14774), .ZN(n10819) );
  AND2_X1 U13130 ( .A1(n14751), .A2(n11287), .ZN(n14770) );
  AOI21_X1 U13131 ( .B1(n11251), .B2(n10816), .A(n10697), .ZN(n14059) );
  INV_X1 U13132 ( .A(n16025), .ZN(n13814) );
  AND2_X1 U13133 ( .A1(n12761), .A2(n12760), .ZN(n14368) );
  AND2_X1 U13134 ( .A1(n12749), .A2(n12748), .ZN(n14423) );
  AND2_X1 U13135 ( .A1(n12727), .A2(n12726), .ZN(n14518) );
  OR2_X1 U13136 ( .A1(n13714), .A2(n13697), .ZN(n15888) );
  INV_X1 U13137 ( .A(n13935), .ZN(n13951) );
  INV_X1 U13138 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20655) );
  OR2_X1 U13139 ( .A1(n20919), .A2(n20703), .ZN(n20576) );
  OR2_X1 U13140 ( .A1(n20919), .A2(n20626), .ZN(n20649) );
  NOR2_X1 U13141 ( .A1(n20580), .A2(n20417), .ZN(n20736) );
  INV_X1 U13142 ( .A(n20338), .ZN(n14150) );
  NAND2_X1 U13143 ( .A1(n16194), .A2(n14161), .ZN(n20273) );
  NAND2_X1 U13144 ( .A1(n11846), .A2(n12501), .ZN(n11877) );
  NOR2_X1 U13145 ( .A1(n11825), .A2(n11694), .ZN(n16444) );
  AND2_X1 U13146 ( .A1(n12807), .A2(n12806), .ZN(n15297) );
  OR2_X1 U13147 ( .A1(n20052), .A2(n14965), .ZN(n19181) );
  OR2_X1 U13148 ( .A1(n12282), .A2(n12281), .ZN(n14003) );
  AND2_X1 U13149 ( .A1(n13351), .A2(n20057), .ZN(n13495) );
  OAI21_X1 U13150 ( .B1(n13341), .B2(n13340), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13342) );
  OR2_X1 U13151 ( .A1(n19095), .A2(n12494), .ZN(n15652) );
  AND3_X1 U13152 ( .A1(n12272), .A2(n12271), .A3(n12270), .ZN(n15057) );
  AND3_X1 U13153 ( .A1(n12191), .A2(n12190), .A3(n12189), .ZN(n15080) );
  NAND2_X1 U13154 ( .A1(n20056), .A2(n12627), .ZN(n12628) );
  AND2_X1 U13155 ( .A1(n20015), .A2(n20022), .ZN(n20003) );
  NAND2_X1 U13156 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19836), .ZN(n19368) );
  INV_X1 U13157 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16478) );
  AOI21_X1 U13158 ( .B1(n11443), .B2(n11442), .A(n11441), .ZN(n11553) );
  NOR2_X1 U13159 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16792), .ZN(n16781) );
  NOR2_X1 U13160 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16818), .ZN(n16803) );
  NOR2_X1 U13161 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16883), .ZN(n16876) );
  NOR2_X1 U13162 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16939), .ZN(n16920) );
  INV_X1 U13163 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17257) );
  INV_X1 U13164 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17241) );
  INV_X1 U13165 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17220) );
  INV_X1 U13166 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17116) );
  INV_X1 U13167 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17610) );
  NAND2_X1 U13168 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17680), .ZN(
        n17653) );
  INV_X1 U13169 ( .A(n17771), .ZN(n17736) );
  NOR2_X1 U13170 ( .A1(n17824), .A2(n17813), .ZN(n17807) );
  INV_X1 U13171 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17849) );
  NAND2_X1 U13172 ( .A1(n13311), .A2(n18150), .ZN(n13324) );
  NOR2_X1 U13173 ( .A1(n17902), .A2(n11405), .ZN(n16519) );
  NAND2_X1 U13174 ( .A1(n11590), .A2(n17878), .ZN(n18175) );
  INV_X1 U13175 ( .A(n17471), .ZN(n13310) );
  NOR2_X1 U13176 ( .A1(n11342), .A2(n11341), .ZN(n11343) );
  INV_X1 U13177 ( .A(n18356), .ZN(n18673) );
  OAI21_X1 U13178 ( .B1(n14790), .B2(n20155), .A(n12884), .ZN(n12885) );
  INV_X1 U13179 ( .A(n20134), .ZN(n20138) );
  NOR2_X2 U13180 ( .A1(n14032), .A2(n14030), .ZN(n20123) );
  OAI21_X1 U13181 ( .B1(n14818), .B2(n14521), .A(n10330), .ZN(n12775) );
  INV_X1 U13182 ( .A(n14521), .ZN(n20175) );
  AOI21_X1 U13183 ( .B1(n14476), .B2(n10023), .A(n9837), .ZN(n14745) );
  NAND2_X1 U13184 ( .A1(n10837), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10868) );
  NAND2_X1 U13185 ( .A1(n10756), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10799) );
  OR3_X1 U13186 ( .A1(n14835), .A2(n14812), .A3(n14821), .ZN(n14824) );
  AND2_X1 U13187 ( .A1(n16055), .A2(n14795), .ZN(n16037) );
  AND2_X1 U13188 ( .A1(n16043), .A2(n14804), .ZN(n14868) );
  INV_X1 U13189 ( .A(n20258), .ZN(n16173) );
  INV_X1 U13190 ( .A(n16182), .ZN(n20260) );
  NAND2_X1 U13191 ( .A1(n20936), .A2(n14161), .ZN(n20417) );
  NOR2_X1 U13192 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20906) );
  AND2_X1 U13193 ( .A1(n20382), .A2(n20647), .ZN(n20334) );
  OAI21_X1 U13194 ( .B1(n20346), .B2(n20345), .A(n20344), .ZN(n20374) );
  NOR2_X2 U13195 ( .A1(n20383), .A2(n20728), .ZN(n20405) );
  NOR2_X2 U13196 ( .A1(n20383), .A2(n20626), .ZN(n20435) );
  AND2_X1 U13197 ( .A1(n20498), .A2(n20444), .ZN(n20488) );
  AND2_X1 U13198 ( .A1(n20498), .A2(n20466), .ZN(n20516) );
  AND2_X1 U13199 ( .A1(n11217), .A2(n20410), .ZN(n20498) );
  NOR2_X1 U13200 ( .A1(n20339), .A2(n14150), .ZN(n20647) );
  INV_X1 U13201 ( .A(n20576), .ZN(n20612) );
  NAND2_X1 U13202 ( .A1(n20916), .A2(n20521), .ZN(n20919) );
  INV_X1 U13203 ( .A(n20727), .ZN(n20689) );
  NOR2_X2 U13204 ( .A1(n20777), .A2(n20703), .ZN(n20765) );
  INV_X1 U13205 ( .A(n20364), .ZN(n20812) );
  NAND2_X1 U13206 ( .A1(n20339), .A2(n20338), .ZN(n20728) );
  INV_X1 U13207 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20852) );
  INV_X1 U13208 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20837) );
  AND2_X1 U13209 ( .A1(n14963), .A2(n16482), .ZN(n19168) );
  OR2_X1 U13210 ( .A1(n13664), .A2(n13663), .ZN(n13665) );
  INV_X1 U13211 ( .A(n19157), .ZN(n19188) );
  OR2_X1 U13212 ( .A1(n12243), .A2(n12242), .ZN(n13843) );
  NAND2_X1 U13213 ( .A1(n13506), .A2(n13509), .ZN(n20022) );
  AND2_X1 U13214 ( .A1(n19217), .A2(n14132), .ZN(n16266) );
  AND2_X1 U13215 ( .A1(n19217), .A2(n13499), .ZN(n19213) );
  AND2_X1 U13216 ( .A1(n15207), .A2(n15206), .ZN(n19057) );
  INV_X1 U13217 ( .A(n19277), .ZN(n16350) );
  INV_X1 U13218 ( .A(n19278), .ZN(n16361) );
  AND2_X1 U13219 ( .A1(n11868), .A2(n15785), .ZN(n19271) );
  INV_X1 U13220 ( .A(n19301), .ZN(n16387) );
  INV_X1 U13221 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15783) );
  NOR2_X2 U13222 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20007) );
  NOR2_X1 U13223 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15785) );
  OAI21_X1 U13224 ( .B1(n19328), .B2(n19327), .A(n19326), .ZN(n19372) );
  OAI21_X1 U13225 ( .B1(n19441), .B2(n19440), .A(n19439), .ZN(n19458) );
  NOR2_X1 U13226 ( .A1(n19559), .A2(n19698), .ZN(n19494) );
  NAND2_X1 U13227 ( .A1(n19987), .A2(n20031), .ZN(n19526) );
  INV_X1 U13228 ( .A(n19552), .ZN(n19555) );
  INV_X1 U13229 ( .A(n19617), .ZN(n19609) );
  OAI21_X1 U13230 ( .B1(n19628), .B2(n19627), .A(n19626), .ZN(n19648) );
  INV_X1 U13231 ( .A(n19660), .ZN(n19682) );
  AND2_X1 U13232 ( .A1(n19692), .A2(n19691), .ZN(n19714) );
  OAI21_X1 U13233 ( .B1(n19741), .B2(n12958), .A(n19726), .ZN(n19743) );
  NAND2_X1 U13234 ( .A1(n19466), .A2(n19994), .ZN(n19754) );
  NOR2_X2 U13235 ( .A1(n19755), .A2(n19832), .ZN(n19881) );
  AND3_X1 U13236 ( .A1(n19029), .A2(n19971), .A3(n19028), .ZN(n20062) );
  INV_X1 U13237 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19913) );
  NOR2_X1 U13238 ( .A1(n18803), .A2(n18788), .ZN(n18778) );
  NOR2_X1 U13239 ( .A1(n17025), .A2(n16661), .ZN(n16696) );
  NOR2_X1 U13240 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16752), .ZN(n16723) );
  NOR2_X1 U13241 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16770), .ZN(n16759) );
  NOR2_X1 U13242 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16839), .ZN(n16825) );
  NOR2_X2 U13243 ( .A1(n19021), .A2(n18838), .ZN(n16999) );
  INV_X1 U13244 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16908) );
  INV_X1 U13245 ( .A(n17028), .ZN(n17019) );
  NOR2_X1 U13246 ( .A1(n16778), .A2(n17129), .ZN(n17098) );
  NAND2_X1 U13247 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17222), .ZN(n17221) );
  NAND2_X1 U13248 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17383), .ZN(n17382) );
  NOR2_X1 U13249 ( .A1(n17550), .A2(n17414), .ZN(n17409) );
  OAI211_X1 U13250 ( .C1(n17296), .C2(n18582), .A(n11402), .B(n11401), .ZN(
        n17903) );
  OR2_X1 U13251 ( .A1(n11597), .A2(n11596), .ZN(n11598) );
  NOR3_X2 U13252 ( .A1(n17946), .A2(P3_STATEBS16_REG_SCAN_IN), .A3(n18966), 
        .ZN(n17828) );
  INV_X1 U13253 ( .A(n17979), .ZN(n17946) );
  INV_X1 U13254 ( .A(n18176), .ZN(n18125) );
  AND2_X1 U13255 ( .A1(n16515), .A2(n18074), .ZN(n18082) );
  INV_X1 U13256 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18112) );
  INV_X1 U13257 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17819) );
  INV_X1 U13258 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18210) );
  INV_X1 U13259 ( .A(n18302), .ZN(n18277) );
  NOR3_X1 U13260 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19007), .ZN(n18613) );
  NOR2_X1 U13261 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18954), .ZN(
        n18981) );
  NAND2_X1 U13262 ( .A1(n18673), .A2(n18613), .ZN(n18348) );
  CLKBUF_X1 U13263 ( .A(n18699), .Z(n18675) );
  CLKBUF_X1 U13264 ( .A(n18419), .Z(n18415) );
  INV_X1 U13265 ( .A(n18444), .ZN(n18435) );
  INV_X1 U13266 ( .A(n18489), .ZN(n18482) );
  INV_X1 U13267 ( .A(n18646), .ZN(n18664) );
  AND2_X1 U13268 ( .A1(n18708), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18725) );
  INV_X1 U13269 ( .A(n18744), .ZN(n18763) );
  INV_X1 U13270 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18840) );
  INV_X1 U13271 ( .A(n19318), .ZN(n19316) );
  INV_X1 U13272 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21137) );
  INV_X1 U13273 ( .A(n12885), .ZN(n12886) );
  INV_X1 U13274 ( .A(n20123), .ZN(n20099) );
  INV_X1 U13275 ( .A(n20157), .ZN(n14071) );
  NAND2_X1 U13276 ( .A1(n13796), .A2(n14607), .ZN(n15981) );
  INV_X1 U13277 ( .A(n20158), .ZN(n13927) );
  INV_X1 U13278 ( .A(n14622), .ZN(n14610) );
  INV_X1 U13279 ( .A(n20180), .ZN(n20210) );
  AND2_X1 U13280 ( .A1(n13861), .A2(n13860), .ZN(n20288) );
  INV_X1 U13281 ( .A(n20248), .ZN(n20253) );
  NAND2_X1 U13282 ( .A1(n16029), .A2(n13726), .ZN(n16022) );
  NAND2_X1 U13283 ( .A1(n20080), .A2(n11196), .ZN(n16029) );
  OR2_X1 U13284 ( .A1(n13714), .A2(n13708), .ZN(n20258) );
  OR2_X1 U13285 ( .A1(n13714), .A2(n13695), .ZN(n16182) );
  OAI21_X1 U13286 ( .B1(n13964), .B2(n16195), .A(n20417), .ZN(n20923) );
  INV_X1 U13287 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20271) );
  NAND2_X1 U13288 ( .A1(n20382), .A2(n20444), .ZN(n20372) );
  AOI22_X1 U13289 ( .A1(n20342), .A2(n20345), .B1(n20580), .B2(n10347), .ZN(
        n20377) );
  AOI22_X1 U13290 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20385), .B1(n20388), 
        .B2(n20384), .ZN(n20409) );
  NAND2_X1 U13291 ( .A1(n20498), .A2(n20647), .ZN(n20464) );
  AOI22_X1 U13292 ( .A1(n20471), .A2(n20468), .B1(n20654), .B2(n10347), .ZN(
        n20492) );
  NAND2_X1 U13293 ( .A1(n20498), .A2(n20493), .ZN(n20526) );
  NAND2_X1 U13294 ( .A1(n20522), .A2(n20647), .ZN(n20575) );
  AOI22_X1 U13295 ( .A1(n20587), .A2(n20583), .B1(n20580), .B2(n20579), .ZN(
        n20616) );
  OR2_X1 U13296 ( .A1(n20919), .A2(n20728), .ZN(n20646) );
  INV_X1 U13297 ( .A(n20785), .ZN(n20669) );
  INV_X1 U13298 ( .A(n20817), .ZN(n20687) );
  OR2_X1 U13299 ( .A1(n20777), .A2(n20648), .ZN(n20727) );
  INV_X1 U13300 ( .A(n20706), .ZN(n20790) );
  OR2_X1 U13301 ( .A1(n20777), .A2(n20728), .ZN(n20832) );
  INV_X1 U13302 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20834) );
  INV_X1 U13303 ( .A(n20903), .ZN(n20899) );
  INV_X1 U13304 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21299) );
  INV_X1 U13305 ( .A(n20864), .ZN(n20881) );
  NAND2_X1 U13306 ( .A1(n20837), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20944) );
  INV_X1 U13307 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19029) );
  NAND2_X1 U13308 ( .A1(n12513), .A2(n13493), .ZN(n13349) );
  OR3_X1 U13309 ( .A1(n14951), .A2(n19897), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19157) );
  OR3_X1 U13310 ( .A1(n14951), .A2(n16201), .A3(n14910), .ZN(n19186) );
  INV_X1 U13311 ( .A(n19168), .ZN(n19179) );
  OR2_X1 U13312 ( .A1(n15221), .A2(n19369), .ZN(n15237) );
  INV_X1 U13313 ( .A(n19213), .ZN(n14010) );
  AND2_X1 U13314 ( .A1(n15310), .A2(n15327), .ZN(n19206) );
  NAND2_X1 U13315 ( .A1(n19217), .A2(n13504), .ZN(n15327) );
  OR2_X1 U13316 ( .A1(n19256), .A2(n20061), .ZN(n19219) );
  NAND2_X1 U13317 ( .A1(n13417), .A2(n20062), .ZN(n19256) );
  INV_X1 U13318 ( .A(n19266), .ZN(n13490) );
  AOI21_X1 U13319 ( .B1(n16205), .B2(n19282), .A(n12952), .ZN(n12953) );
  INV_X1 U13320 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16281) );
  INV_X1 U13321 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16300) );
  NAND2_X1 U13322 ( .A1(n12585), .A2(n12173), .ZN(n19277) );
  OR2_X1 U13323 ( .A1(n15454), .A2(n19314), .ZN(n12503) );
  INV_X1 U13324 ( .A(n16412), .ZN(n19308) );
  INV_X1 U13325 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20036) );
  INV_X1 U13326 ( .A(n19999), .ZN(n19996) );
  INV_X1 U13327 ( .A(n19401), .ZN(n19398) );
  OR2_X1 U13328 ( .A1(n19526), .A2(n19698), .ZN(n19462) );
  AND2_X1 U13329 ( .A1(n19470), .A2(n19469), .ZN(n19478) );
  INV_X1 U13330 ( .A(n19494), .ZN(n19491) );
  OR2_X1 U13331 ( .A1(n19526), .A2(n19754), .ZN(n19518) );
  OR2_X1 U13332 ( .A1(n19559), .A2(n19754), .ZN(n19552) );
  INV_X1 U13333 ( .A(n19582), .ZN(n19580) );
  OR2_X1 U13334 ( .A1(n19559), .A2(n19832), .ZN(n19617) );
  AND2_X1 U13335 ( .A1(n19623), .A2(n19622), .ZN(n19632) );
  OR2_X1 U13336 ( .A1(n19755), .A2(n19624), .ZN(n19660) );
  OR2_X1 U13337 ( .A1(n19783), .A2(n19698), .ZN(n19718) );
  INV_X1 U13338 ( .A(n19722), .ZN(n19746) );
  AND2_X1 U13339 ( .A1(n19750), .A2(n19749), .ZN(n19782) );
  INV_X1 U13340 ( .A(n19866), .ZN(n19814) );
  INV_X1 U13341 ( .A(n19800), .ZN(n19846) );
  INV_X1 U13342 ( .A(n19774), .ZN(n19875) );
  INV_X1 U13343 ( .A(n19890), .ZN(n19888) );
  INV_X1 U13344 ( .A(n19985), .ZN(n19896) );
  NAND2_X1 U13345 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19029), .ZN(n20068) );
  INV_X1 U13346 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19007) );
  INV_X1 U13347 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17813) );
  INV_X1 U13348 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17314) );
  INV_X1 U13349 ( .A(n17024), .ZN(n17013) );
  INV_X1 U13350 ( .A(n17336), .ZN(n17341) );
  NOR2_X1 U13351 ( .A1(n13775), .A2(n17338), .ZN(n17328) );
  INV_X1 U13352 ( .A(n17424), .ZN(n17407) );
  INV_X1 U13353 ( .A(n17498), .ZN(n17493) );
  NAND2_X1 U13354 ( .A1(n17521), .A2(n17503), .ZN(n17520) );
  INV_X1 U13355 ( .A(n17521), .ZN(n17539) );
  INV_X1 U13356 ( .A(n17852), .ZN(n17880) );
  NOR2_X1 U13357 ( .A1(n17642), .A2(n17828), .ZN(n17966) );
  NAND2_X1 U13358 ( .A1(n16515), .A2(n18287), .ZN(n18236) );
  INV_X1 U13359 ( .A(n18194), .ZN(n18223) );
  INV_X1 U13360 ( .A(n18293), .ZN(n18287) );
  INV_X1 U13361 ( .A(n14206), .ZN(n19003) );
  INV_X1 U13362 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18830) );
  INV_X1 U13363 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18325) );
  INV_X1 U13364 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18335) );
  INV_X1 U13365 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18397) );
  INV_X1 U13366 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18568) );
  INV_X1 U13367 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18582) );
  INV_X1 U13368 ( .A(n18740), .ZN(n18656) );
  INV_X1 U13369 ( .A(n18755), .ZN(n18662) );
  INV_X1 U13370 ( .A(n18690), .ZN(n18704) );
  INV_X1 U13371 ( .A(n18691), .ZN(n18752) );
  NAND2_X1 U13372 ( .A1(n18851), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18846) );
  INV_X1 U13373 ( .A(n18951), .ZN(n18948) );
  INV_X1 U13374 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18881) );
  CLKBUF_X1 U13375 ( .A(n18933), .Z(n18934) );
  NOR2_X1 U13376 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13343), .ZN(n16612)
         );
  INV_X1 U13377 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19218) );
  INV_X1 U13378 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19918) );
  OAI21_X1 U13379 ( .B1(n14634), .B2(n14532), .A(n12776), .ZN(P1_U2842) );
  NAND2_X1 U13380 ( .A1(n10340), .A2(n12639), .ZN(P2_U2985) );
  NAND2_X1 U13381 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10358) );
  NAND2_X1 U13382 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10357) );
  NAND2_X1 U13383 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10356) );
  NAND2_X1 U13384 ( .A1(n10446), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10355) );
  NAND2_X1 U13385 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10362) );
  AND2_X2 U13386 ( .A1(n10369), .A2(n13578), .ZN(n11086) );
  NAND2_X1 U13387 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10361) );
  NAND2_X1 U13388 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10360) );
  AND2_X2 U13389 ( .A1(n13612), .A2(n13941), .ZN(n10421) );
  NAND2_X1 U13390 ( .A1(n10421), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10359) );
  NAND2_X1 U13391 ( .A1(n10431), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10367) );
  AND2_X2 U13392 ( .A1(n10363), .A2(n10369), .ZN(n11117) );
  NAND2_X1 U13393 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10366) );
  NAND2_X1 U13394 ( .A1(n9839), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10365) );
  NAND2_X1 U13395 ( .A1(n10488), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10364) );
  NAND2_X1 U13396 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10374) );
  NAND2_X1 U13397 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10373) );
  AND2_X2 U13398 ( .A1(n13578), .A2(n13941), .ZN(n10441) );
  NAND2_X1 U13399 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10371) );
  NAND4_X4 U13400 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10450) );
  AOI22_X1 U13401 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n9839), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13402 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10349), .B1(
        n11109), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13403 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n9799), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13404 ( .A1(n9827), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10421), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13405 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10407), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13406 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13407 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10431), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13408 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10383) );
  NAND2_X1 U13409 ( .A1(n10461), .A2(n10574), .ZN(n10395) );
  AOI22_X1 U13410 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13411 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13412 ( .A1(n10431), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13413 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10421), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13414 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13415 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13416 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11109), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U13417 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13418 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13419 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13420 ( .A1(n10431), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13421 ( .A1(n10406), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10421), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13422 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13423 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13424 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10401) );
  AND2_X2 U13425 ( .A1(n10450), .A2(n14162), .ZN(n10458) );
  NAND2_X1 U13426 ( .A1(n10458), .A2(n10469), .ZN(n10405) );
  INV_X1 U13427 ( .A(n10432), .ZN(n10955) );
  AOI22_X1 U13428 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13429 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11109), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13430 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13431 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13432 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13433 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13434 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10421), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13435 ( .A1(n9827), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U13436 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10419) );
  AOI22_X1 U13437 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U13438 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10417) );
  NAND4_X1 U13439 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n10427) );
  AOI22_X1 U13440 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13441 ( .A1(n9839), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U13442 ( .A1(n10446), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10423) );
  AOI22_X1 U13443 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10421), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10422) );
  NAND4_X1 U13444 ( .A1(n10425), .A2(n10424), .A3(n10423), .A4(n10422), .ZN(
        n10426) );
  OR2_X2 U13445 ( .A1(n10427), .A2(n10426), .ZN(n20287) );
  NAND2_X1 U13446 ( .A1(n10429), .A2(n10428), .ZN(n11195) );
  NOR2_X2 U13447 ( .A1(n11195), .A2(n10455), .ZN(n13572) );
  AOI22_X1 U13448 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13449 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13450 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10421), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13451 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13452 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13453 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10438) );
  BUF_X4 U13454 ( .A(n10349), .Z(n11093) );
  AOI22_X1 U13455 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13456 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9839), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13457 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U13458 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11109), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13459 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13460 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U13461 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13462 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U13463 ( .A1(n13624), .A2(n20287), .ZN(n10457) );
  INV_X1 U13464 ( .A(n10458), .ZN(n10454) );
  OAI21_X1 U13465 ( .B1(n10454), .B2(n13680), .A(n10453), .ZN(n10456) );
  NAND3_X1 U13466 ( .A1(n10457), .A2(n10456), .A3(n10455), .ZN(n10463) );
  INV_X1 U13467 ( .A(n10463), .ZN(n10460) );
  AND2_X1 U13468 ( .A1(n10470), .A2(n10458), .ZN(n10459) );
  XNOR2_X1 U13469 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12861) );
  NAND3_X1 U13470 ( .A1(n13939), .A2(n10470), .A3(n10461), .ZN(n13573) );
  OAI211_X1 U13471 ( .C1(n13453), .C2(n14162), .A(n13560), .B(n14028), .ZN(
        n10479) );
  NOR2_X1 U13472 ( .A1(n10479), .A2(n13939), .ZN(n10465) );
  NAND2_X1 U13473 ( .A1(n10463), .A2(n20266), .ZN(n10464) );
  NAND3_X1 U13474 ( .A1(n10475), .A2(n10465), .A3(n10464), .ZN(n10466) );
  NAND2_X1 U13475 ( .A1(n10466), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10467) );
  MUX2_X1 U13476 ( .A(n11198), .B(n15871), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10468) );
  INV_X1 U13477 ( .A(n20287), .ZN(n12678) );
  AOI21_X1 U13478 ( .B1(n10469), .B2(n10450), .A(n12678), .ZN(n10473) );
  INV_X1 U13479 ( .A(n20906), .ZN(n10471) );
  NOR2_X1 U13480 ( .A1(n10471), .A2(n20936), .ZN(n10472) );
  NAND2_X1 U13481 ( .A1(n13939), .A2(n10469), .ZN(n13699) );
  OAI211_X1 U13482 ( .C1(n10473), .C2(n14315), .A(n10472), .B(n13699), .ZN(
        n10474) );
  INV_X1 U13483 ( .A(n10475), .ZN(n10476) );
  NAND2_X1 U13484 ( .A1(n10476), .A2(n20274), .ZN(n10481) );
  NAND2_X1 U13485 ( .A1(n10463), .A2(n10470), .ZN(n13571) );
  NOR2_X1 U13486 ( .A1(n10477), .A2(n13453), .ZN(n10478) );
  NOR2_X1 U13487 ( .A1(n10479), .A2(n10478), .ZN(n10480) );
  NAND4_X1 U13488 ( .A1(n10482), .A2(n10481), .A3(n13571), .A4(n10480), .ZN(
        n10536) );
  INV_X1 U13489 ( .A(n10536), .ZN(n10483) );
  AOI22_X1 U13490 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13491 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13492 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13493 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U13494 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10494) );
  AOI22_X1 U13495 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13496 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13497 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10421), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13498 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10489) );
  NAND4_X1 U13499 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10493) );
  AOI22_X1 U13500 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13501 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13502 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13503 ( .A1(n10495), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10421), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10496) );
  NAND4_X1 U13504 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10505) );
  AOI22_X1 U13505 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13506 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11110), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13507 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U13508 ( .A1(n11049), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10500) );
  NAND4_X1 U13509 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10504) );
  XNOR2_X1 U13510 ( .A(n10522), .B(n11207), .ZN(n10506) );
  NAND2_X1 U13511 ( .A1(n10506), .A2(n11264), .ZN(n10507) );
  NAND2_X1 U13512 ( .A1(n20266), .A2(n11207), .ZN(n10508) );
  OAI211_X1 U13513 ( .C1(n10522), .C2(n13706), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n10508), .ZN(n10509) );
  INV_X1 U13514 ( .A(n10509), .ZN(n10510) );
  NAND2_X1 U13515 ( .A1(n11264), .A2(n11267), .ZN(n10527) );
  INV_X1 U13516 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10525) );
  NAND2_X1 U13517 ( .A1(n20266), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10571) );
  INV_X1 U13518 ( .A(n10571), .ZN(n10521) );
  AOI22_X1 U13519 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13520 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13521 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13522 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10511) );
  NAND4_X1 U13523 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n10520) );
  AOI22_X1 U13524 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13525 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13526 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13527 ( .A1(n9827), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10515) );
  NAND4_X1 U13528 ( .A1(n10518), .A2(n10517), .A3(n10516), .A4(n10515), .ZN(
        n10519) );
  NAND2_X1 U13529 ( .A1(n10521), .A2(n11206), .ZN(n10524) );
  NAND2_X1 U13530 ( .A1(n11264), .A2(n10522), .ZN(n10523) );
  OAI211_X1 U13531 ( .C1(n11176), .C2(n10525), .A(n10524), .B(n10523), .ZN(
        n10526) );
  INV_X1 U13532 ( .A(n10526), .ZN(n10528) );
  NAND2_X1 U13533 ( .A1(n10544), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10533) );
  NAND2_X1 U13534 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10546) );
  OAI21_X1 U13535 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10546), .ZN(n20578) );
  OR2_X1 U13536 ( .A1(n15871), .A2(n20655), .ZN(n10542) );
  OAI21_X1 U13537 ( .B1(n11198), .B2(n20578), .A(n10542), .ZN(n10531) );
  INV_X1 U13538 ( .A(n10531), .ZN(n10532) );
  NAND2_X1 U13539 ( .A1(n10533), .A2(n10532), .ZN(n10535) );
  INV_X1 U13540 ( .A(n10539), .ZN(n10538) );
  NAND2_X2 U13541 ( .A1(n20378), .A2(n10539), .ZN(n10558) );
  NAND2_X1 U13542 ( .A1(n11264), .A2(n11206), .ZN(n10540) );
  AND2_X1 U13543 ( .A1(n10542), .A2(n13940), .ZN(n10543) );
  NAND2_X1 U13544 ( .A1(n10558), .A2(n10556), .ZN(n10552) );
  NAND2_X1 U13545 ( .A1(n10544), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10550) );
  INV_X1 U13546 ( .A(n11198), .ZN(n10548) );
  INV_X1 U13547 ( .A(n10546), .ZN(n10545) );
  NAND2_X1 U13548 ( .A1(n10545), .A2(n11143), .ZN(n20618) );
  NAND2_X1 U13549 ( .A1(n10546), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10547) );
  NAND2_X1 U13550 ( .A1(n20618), .A2(n10547), .ZN(n14155) );
  NAND2_X1 U13551 ( .A1(n10548), .A2(n14155), .ZN(n10549) );
  NAND2_X1 U13552 ( .A1(n10550), .A2(n10549), .ZN(n10553) );
  NOR2_X1 U13553 ( .A1(n15871), .A2(n11143), .ZN(n10554) );
  INV_X1 U13554 ( .A(n10553), .ZN(n10557) );
  INV_X1 U13555 ( .A(n10554), .ZN(n10555) );
  NAND4_X1 U13556 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        n10559) );
  NAND2_X1 U13557 ( .A1(n13635), .A2(n10559), .ZN(n13608) );
  AOI22_X1 U13558 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13559 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13560 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13561 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10560) );
  NAND4_X1 U13562 ( .A1(n10563), .A2(n10562), .A3(n10561), .A4(n10560), .ZN(
        n10569) );
  INV_X2 U13563 ( .A(n13938), .ZN(n11108) );
  AOI22_X1 U13564 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13565 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13566 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13567 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10564) );
  NAND4_X1 U13568 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10568) );
  INV_X1 U13569 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20286) );
  OAI22_X1 U13570 ( .A1(n11176), .A2(n20286), .B1(n10571), .B2(n11220), .ZN(
        n10572) );
  INV_X1 U13571 ( .A(n10572), .ZN(n10573) );
  INV_X2 U13572 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n10577) );
  INV_X1 U13573 ( .A(n13792), .ZN(n10575) );
  NAND2_X1 U13574 ( .A1(n10575), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10628) );
  NOR2_X2 U13575 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10621) );
  XNOR2_X1 U13576 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14297) );
  AOI21_X1 U13577 ( .B1(n11104), .B2(n14297), .A(n11132), .ZN(n10579) );
  NAND2_X1 U13578 ( .A1(n10672), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10578) );
  OAI211_X1 U13579 ( .C1(n10628), .C2(n10009), .A(n10579), .B(n10578), .ZN(
        n10580) );
  INV_X1 U13580 ( .A(n10580), .ZN(n10581) );
  NAND2_X1 U13581 ( .A1(n11132), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10599) );
  INV_X1 U13582 ( .A(n13813), .ZN(n10598) );
  NAND2_X1 U13583 ( .A1(n10582), .A2(n11205), .ZN(n10583) );
  NAND2_X1 U13584 ( .A1(n20339), .A2(n10816), .ZN(n10588) );
  AOI22_X1 U13585 ( .A1(n10672), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n10577), .ZN(n10586) );
  INV_X1 U13586 ( .A(n10628), .ZN(n10646) );
  NAND2_X1 U13587 ( .A1(n10646), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10585) );
  AND2_X1 U13588 ( .A1(n10586), .A2(n10585), .ZN(n10587) );
  NAND2_X1 U13589 ( .A1(n10588), .A2(n10587), .ZN(n13742) );
  NAND2_X1 U13590 ( .A1(n20338), .A2(n10469), .ZN(n10590) );
  NAND2_X1 U13591 ( .A1(n10590), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13719) );
  NAND2_X1 U13592 ( .A1(n10577), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10593) );
  NAND2_X1 U13593 ( .A1(n10672), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10592) );
  OAI211_X1 U13594 ( .C1(n10628), .C2(n10323), .A(n10593), .B(n10592), .ZN(
        n10594) );
  AOI21_X1 U13595 ( .B1(n10591), .B2(n10816), .A(n10594), .ZN(n10595) );
  OR2_X1 U13596 ( .A1(n13719), .A2(n10595), .ZN(n13720) );
  INV_X1 U13597 ( .A(n10595), .ZN(n13721) );
  OR2_X1 U13598 ( .A1(n13721), .A2(n11041), .ZN(n10596) );
  NAND2_X1 U13599 ( .A1(n13720), .A2(n10596), .ZN(n13741) );
  NAND2_X1 U13600 ( .A1(n13742), .A2(n13741), .ZN(n13812) );
  NAND2_X1 U13601 ( .A1(n10598), .A2(n10597), .ZN(n13810) );
  NAND2_X1 U13602 ( .A1(n10544), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10606) );
  NOR3_X1 U13603 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11143), .A3(
        n20655), .ZN(n20499) );
  NAND2_X1 U13604 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20499), .ZN(
        n20494) );
  NAND2_X1 U13605 ( .A1(n20617), .A2(n20494), .ZN(n10603) );
  NAND3_X1 U13606 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20776) );
  INV_X1 U13607 ( .A(n20776), .ZN(n10602) );
  NAND2_X1 U13608 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10602), .ZN(
        n20770) );
  NAND2_X1 U13609 ( .A1(n10603), .A2(n20770), .ZN(n20523) );
  OAI22_X1 U13610 ( .A1(n11198), .A2(n20523), .B1(n15871), .B2(n20617), .ZN(
        n10604) );
  INV_X1 U13611 ( .A(n10604), .ZN(n10605) );
  XNOR2_X2 U13612 ( .A(n13635), .B(n20411), .ZN(n20913) );
  NAND2_X1 U13613 ( .A1(n20913), .A2(n20936), .ZN(n10619) );
  AOI22_X1 U13614 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13615 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13616 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10609) );
  INV_X1 U13617 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20292) );
  AOI22_X1 U13618 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10608) );
  NAND4_X1 U13619 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10617) );
  AOI22_X1 U13620 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13621 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13622 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13623 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10612) );
  NAND4_X1 U13624 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10616) );
  AOI22_X1 U13625 ( .A1(n11163), .A2(n11201), .B1(n11185), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10618) );
  NAND2_X1 U13626 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10623) );
  INV_X1 U13627 ( .A(n10623), .ZN(n10625) );
  INV_X1 U13628 ( .A(n10649), .ZN(n10624) );
  OAI21_X1 U13629 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10625), .A(
        n10624), .ZN(n14067) );
  AOI22_X1 U13630 ( .A1(n11104), .A2(n14067), .B1(n11132), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10627) );
  NAND2_X1 U13631 ( .A1(n10672), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10626) );
  OAI211_X1 U13632 ( .C1(n10628), .C2(n10010), .A(n10627), .B(n10626), .ZN(
        n10629) );
  INV_X1 U13633 ( .A(n10629), .ZN(n10630) );
  OAI21_X1 U13634 ( .B1(n9818), .B2(n10308), .A(n10630), .ZN(n13854) );
  NAND2_X1 U13635 ( .A1(n13855), .A2(n13854), .ZN(n13853) );
  INV_X1 U13636 ( .A(n13853), .ZN(n10655) );
  AOI22_X1 U13637 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13638 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13639 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13640 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10631) );
  NAND4_X1 U13641 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10640) );
  AOI22_X1 U13642 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13643 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13644 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13645 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10635) );
  NAND4_X1 U13646 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n10639) );
  NAND2_X1 U13647 ( .A1(n11163), .A2(n11241), .ZN(n10642) );
  NAND2_X1 U13648 ( .A1(n11185), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10641) );
  NAND2_X1 U13649 ( .A1(n10643), .A2(n10339), .ZN(n10645) );
  NAND2_X1 U13650 ( .A1(n10646), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10652) );
  INV_X1 U13651 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10647) );
  AOI21_X1 U13652 ( .B1(n10647), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10648) );
  AOI21_X1 U13653 ( .B1(n10672), .B2(P1_EAX_REG_4__SCAN_IN), .A(n10648), .ZN(
        n10651) );
  NOR2_X1 U13654 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10649), .ZN(
        n10650) );
  NOR2_X1 U13655 ( .A1(n10673), .A2(n10650), .ZN(n13903) );
  AOI22_X1 U13656 ( .A1(n10652), .A2(n10651), .B1(n11104), .B2(n13903), .ZN(
        n10653) );
  INV_X1 U13657 ( .A(n13882), .ZN(n10654) );
  NAND2_X1 U13658 ( .A1(n10655), .A2(n10654), .ZN(n13881) );
  INV_X1 U13659 ( .A(n13881), .ZN(n10679) );
  INV_X1 U13660 ( .A(n10670), .ZN(n10668) );
  AOI22_X1 U13661 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13662 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13663 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10657) );
  INV_X1 U13664 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20299) );
  AOI22_X1 U13665 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10656) );
  NAND4_X1 U13666 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n10665) );
  AOI22_X1 U13667 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13668 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13669 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13670 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10660) );
  NAND4_X1 U13671 ( .A1(n10663), .A2(n10662), .A3(n10661), .A4(n10660), .ZN(
        n10664) );
  NAND2_X1 U13672 ( .A1(n11163), .A2(n11244), .ZN(n10667) );
  NAND2_X1 U13673 ( .A1(n11185), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10666) );
  NAND2_X1 U13674 ( .A1(n10667), .A2(n10666), .ZN(n10669) );
  NAND2_X1 U13675 ( .A1(n10670), .A2(n10096), .ZN(n10671) );
  INV_X1 U13676 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n10675) );
  OAI21_X1 U13677 ( .B1(n10673), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n10693), .ZN(n16023) );
  AOI22_X1 U13678 ( .A1(n16023), .A2(n11104), .B1(n11132), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10674) );
  OAI21_X1 U13679 ( .B1(n10707), .B2(n10675), .A(n10674), .ZN(n10676) );
  INV_X1 U13680 ( .A(n13969), .ZN(n10678) );
  NAND2_X1 U13681 ( .A1(n10679), .A2(n10678), .ZN(n13968) );
  AOI22_X1 U13682 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13683 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13684 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13685 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10680) );
  NAND4_X1 U13686 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(
        n10689) );
  AOI22_X1 U13687 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13688 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13689 ( .A1(n10495), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13690 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10684) );
  NAND4_X1 U13691 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10688) );
  NAND2_X1 U13692 ( .A1(n11163), .A2(n11258), .ZN(n10691) );
  NAND2_X1 U13693 ( .A1(n11185), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10690) );
  NAND2_X1 U13694 ( .A1(n10698), .A2(n10699), .ZN(n11251) );
  INV_X1 U13695 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10696) );
  AND2_X1 U13696 ( .A1(n10693), .A2(n10692), .ZN(n10694) );
  OR2_X1 U13697 ( .A1(n10694), .A2(n10703), .ZN(n20120) );
  AOI22_X1 U13698 ( .A1(n20120), .A2(n10621), .B1(n11132), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10695) );
  OAI21_X1 U13699 ( .B1(n10707), .B2(n10696), .A(n10695), .ZN(n10697) );
  NOR2_X2 U13700 ( .A1(n13968), .A2(n14059), .ZN(n14057) );
  INV_X1 U13701 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10701) );
  NAND2_X1 U13702 ( .A1(n11163), .A2(n11267), .ZN(n10700) );
  OAI21_X1 U13703 ( .B1(n10701), .B2(n11176), .A(n10700), .ZN(n10702) );
  XNOR2_X1 U13704 ( .A(n11266), .B(n10702), .ZN(n11256) );
  NAND2_X1 U13705 ( .A1(n11256), .A2(n10816), .ZN(n10710) );
  INV_X1 U13706 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10706) );
  NOR2_X1 U13707 ( .A1(n10703), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10704) );
  OR2_X1 U13708 ( .A1(n10725), .A2(n10704), .ZN(n20110) );
  AOI22_X1 U13709 ( .A1(n20110), .A2(n11104), .B1(n11132), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13710 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13711 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13712 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13713 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10711) );
  NAND4_X1 U13714 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n10720) );
  AOI22_X1 U13715 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13716 ( .A1(n10431), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13717 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13718 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10715) );
  NAND4_X1 U13719 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10719) );
  OAI21_X1 U13720 ( .B1(n10720), .B2(n10719), .A(n10816), .ZN(n10724) );
  NAND2_X1 U13721 ( .A1(n10672), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10723) );
  XNOR2_X1 U13722 ( .A(n10725), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14142) );
  NAND2_X1 U13723 ( .A1(n14142), .A2(n10621), .ZN(n10722) );
  NAND2_X1 U13724 ( .A1(n11132), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10721) );
  XNOR2_X1 U13725 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10751), .ZN(
        n20096) );
  INV_X1 U13726 ( .A(n20096), .ZN(n10740) );
  AOI22_X1 U13727 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9812), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13728 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13729 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13730 ( .A1(n11049), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10726) );
  NAND4_X1 U13731 ( .A1(n10729), .A2(n10728), .A3(n10727), .A4(n10726), .ZN(
        n10735) );
  AOI22_X1 U13732 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13733 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13734 ( .A1(n10495), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13735 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10730) );
  NAND4_X1 U13736 ( .A1(n10733), .A2(n10732), .A3(n10731), .A4(n10730), .ZN(
        n10734) );
  NOR2_X1 U13737 ( .A1(n10735), .A2(n10734), .ZN(n10738) );
  NAND2_X1 U13738 ( .A1(n10672), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10737) );
  NAND2_X1 U13739 ( .A1(n11132), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10736) );
  OAI211_X1 U13740 ( .C1(n10308), .C2(n10738), .A(n10737), .B(n10736), .ZN(
        n10739) );
  AOI21_X1 U13741 ( .B1(n10740), .B2(n11104), .A(n10739), .ZN(n14146) );
  AOI22_X1 U13742 ( .A1(n10431), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13743 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13744 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13745 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10741) );
  NAND4_X1 U13746 ( .A1(n10744), .A2(n10743), .A3(n10742), .A4(n10741), .ZN(
        n10750) );
  AOI22_X1 U13747 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13748 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13749 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13750 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10745) );
  NAND4_X1 U13751 ( .A1(n10748), .A2(n10747), .A3(n10746), .A4(n10745), .ZN(
        n10749) );
  NOR2_X1 U13752 ( .A1(n10750), .A2(n10749), .ZN(n10754) );
  XNOR2_X1 U13753 ( .A(n10755), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14785) );
  NAND2_X1 U13754 ( .A1(n14785), .A2(n10621), .ZN(n10753) );
  AOI22_X1 U13755 ( .A1(n10672), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n11132), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10752) );
  OAI211_X1 U13756 ( .C1(n10754), .C2(n10308), .A(n10753), .B(n10752), .ZN(
        n14184) );
  NAND2_X1 U13757 ( .A1(n10672), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n10758) );
  OAI21_X1 U13758 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10756), .A(
        n10799), .ZN(n16014) );
  AOI22_X1 U13759 ( .A1(n10621), .A2(n16014), .B1(n11132), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10757) );
  NAND2_X1 U13760 ( .A1(n10758), .A2(n10757), .ZN(n10759) );
  OAI21_X1 U13761 ( .B1(n10760), .B2(n10759), .A(n10774), .ZN(n14618) );
  INV_X1 U13762 ( .A(n14618), .ZN(n10773) );
  AOI22_X1 U13763 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9812), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13764 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13765 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13766 ( .A1(n11049), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10761) );
  NAND4_X1 U13767 ( .A1(n10764), .A2(n10763), .A3(n10762), .A4(n10761), .ZN(
        n10770) );
  AOI22_X1 U13768 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11110), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13769 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U13770 ( .A1(n10495), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13771 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10765) );
  NAND4_X1 U13772 ( .A1(n10768), .A2(n10767), .A3(n10766), .A4(n10765), .ZN(
        n10769) );
  OR2_X1 U13773 ( .A1(n10770), .A2(n10769), .ZN(n10771) );
  NAND2_X1 U13774 ( .A1(n10816), .A2(n10771), .ZN(n14621) );
  AOI22_X1 U13775 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9812), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13776 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13777 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13778 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10775) );
  NAND4_X1 U13779 ( .A1(n10778), .A2(n10777), .A3(n10776), .A4(n10775), .ZN(
        n10784) );
  AOI22_X1 U13780 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U13781 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10781) );
  AOI22_X1 U13782 ( .A1(n9839), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U13783 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10779) );
  NAND4_X1 U13784 ( .A1(n10782), .A2(n10781), .A3(n10780), .A4(n10779), .ZN(
        n10783) );
  NOR2_X1 U13785 ( .A1(n10784), .A2(n10783), .ZN(n10788) );
  XNOR2_X1 U13786 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10799), .ZN(
        n16000) );
  INV_X1 U13787 ( .A(n16000), .ZN(n10785) );
  AOI22_X1 U13788 ( .A1(n11132), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n10621), .B2(n10785), .ZN(n10787) );
  NAND2_X1 U13789 ( .A1(n10672), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10786) );
  OAI211_X1 U13790 ( .C1(n10308), .C2(n10788), .A(n10787), .B(n10786), .ZN(
        n14616) );
  AOI22_X1 U13791 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9812), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13792 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13793 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13794 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10789) );
  NAND4_X1 U13795 ( .A1(n10792), .A2(n10791), .A3(n10790), .A4(n10789), .ZN(
        n10798) );
  AOI22_X1 U13796 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13797 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13798 ( .A1(n10495), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13799 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10793) );
  NAND4_X1 U13800 ( .A1(n10796), .A2(n10795), .A3(n10794), .A4(n10793), .ZN(
        n10797) );
  OAI21_X1 U13801 ( .B1(n10798), .B2(n10797), .A(n10816), .ZN(n10803) );
  XNOR2_X1 U13802 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10804), .ZN(
        n15947) );
  INV_X1 U13803 ( .A(n11132), .ZN(n10864) );
  INV_X1 U13804 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14774) );
  OAI22_X1 U13805 ( .A1(n15947), .A2(n11041), .B1(n10864), .B2(n14774), .ZN(
        n10800) );
  INV_X1 U13806 ( .A(n10800), .ZN(n10802) );
  NAND2_X1 U13807 ( .A1(n10672), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10801) );
  XOR2_X1 U13808 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n10819), .Z(
        n15996) );
  AOI22_X1 U13809 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13810 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11093), .B1(
        n11110), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13811 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11108), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13812 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10805) );
  NAND4_X1 U13813 ( .A1(n10808), .A2(n10807), .A3(n10806), .A4(n10805), .ZN(
        n10814) );
  AOI22_X1 U13814 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13815 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11087), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U13816 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13817 ( .A1(n9839), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10809) );
  NAND4_X1 U13818 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(
        n10813) );
  OR2_X1 U13819 ( .A1(n10814), .A2(n10813), .ZN(n10815) );
  AOI22_X1 U13820 ( .A1(n10816), .A2(n10815), .B1(n11132), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10818) );
  NAND2_X1 U13821 ( .A1(n10672), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10817) );
  OAI211_X1 U13822 ( .C1(n15996), .C2(n11041), .A(n10818), .B(n10817), .ZN(
        n14516) );
  XNOR2_X1 U13823 ( .A(n10836), .B(n14493), .ZN(n14765) );
  AOI22_X1 U13824 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10431), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13825 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13826 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13827 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10820) );
  NAND4_X1 U13828 ( .A1(n10823), .A2(n10822), .A3(n10821), .A4(n10820), .ZN(
        n10829) );
  AOI22_X1 U13829 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13830 ( .A1(n10495), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13831 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13832 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10824) );
  NAND4_X1 U13833 ( .A1(n10827), .A2(n10826), .A3(n10825), .A4(n10824), .ZN(
        n10828) );
  NOR2_X1 U13834 ( .A1(n10829), .A2(n10828), .ZN(n10832) );
  NAND2_X1 U13835 ( .A1(n10672), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10831) );
  NAND2_X1 U13836 ( .A1(n11132), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10830) );
  OAI211_X1 U13837 ( .C1(n10308), .C2(n10832), .A(n10831), .B(n10830), .ZN(
        n10833) );
  AOI21_X1 U13838 ( .B1(n14765), .B2(n10621), .A(n10833), .ZN(n14489) );
  OR2_X1 U13839 ( .A1(n10837), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10838) );
  NAND2_X1 U13840 ( .A1(n10838), .A2(n10868), .ZN(n15991) );
  AOI22_X1 U13841 ( .A1(n10431), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13842 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11110), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13843 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13844 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10839) );
  NAND4_X1 U13845 ( .A1(n10842), .A2(n10841), .A3(n10840), .A4(n10839), .ZN(
        n10848) );
  AOI22_X1 U13846 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13847 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13848 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13849 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10843) );
  NAND4_X1 U13850 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10847) );
  NOR2_X1 U13851 ( .A1(n10848), .A2(n10847), .ZN(n10851) );
  OAI21_X1 U13852 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21137), .A(
        n10577), .ZN(n10850) );
  NAND2_X1 U13853 ( .A1(n10672), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n10849) );
  OAI211_X1 U13854 ( .C1(n11128), .C2(n10851), .A(n10850), .B(n10849), .ZN(
        n10852) );
  OAI21_X1 U13855 ( .B1(n15991), .B2(n11041), .A(n10852), .ZN(n15925) );
  AOI22_X1 U13856 ( .A1(n10495), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13857 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13858 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13859 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10854) );
  NAND4_X1 U13860 ( .A1(n10857), .A2(n10856), .A3(n10855), .A4(n10854), .ZN(
        n10863) );
  AOI22_X1 U13861 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U13862 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U13863 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13864 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10858) );
  NAND4_X1 U13865 ( .A1(n10861), .A2(n10860), .A3(n10859), .A4(n10858), .ZN(
        n10862) );
  OAI21_X1 U13866 ( .B1(n10863), .B2(n10862), .A(n11102), .ZN(n10867) );
  XNOR2_X1 U13867 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10868), .ZN(
        n15914) );
  INV_X1 U13868 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15912) );
  OAI22_X1 U13869 ( .A1(n15914), .A2(n11041), .B1(n10864), .B2(n15912), .ZN(
        n10865) );
  AOI21_X1 U13870 ( .B1(n10672), .B2(P1_EAX_REG_17__SCAN_IN), .A(n10865), .ZN(
        n10866) );
  INV_X1 U13871 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10872) );
  INV_X1 U13872 ( .A(n10870), .ZN(n10871) );
  NAND2_X1 U13873 ( .A1(n10872), .A2(n10871), .ZN(n10873) );
  NAND2_X1 U13874 ( .A1(n10902), .A2(n10873), .ZN(n14743) );
  AOI22_X1 U13875 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13876 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11110), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13877 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U13878 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10874) );
  NAND4_X1 U13879 ( .A1(n10877), .A2(n10876), .A3(n10875), .A4(n10874), .ZN(
        n10883) );
  AOI22_X1 U13880 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13881 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13882 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13883 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10878) );
  NAND4_X1 U13884 ( .A1(n10881), .A2(n10880), .A3(n10879), .A4(n10878), .ZN(
        n10882) );
  NOR2_X1 U13885 ( .A1(n10883), .A2(n10882), .ZN(n10885) );
  AOI22_X1 U13886 ( .A1(n10672), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n10577), .ZN(n10884) );
  OAI21_X1 U13887 ( .B1(n11128), .B2(n10885), .A(n10884), .ZN(n10886) );
  MUX2_X1 U13888 ( .A(n14743), .B(n10886), .S(n11041), .Z(n14474) );
  AOI22_X1 U13889 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13890 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U13891 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U13892 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10887) );
  NAND4_X1 U13893 ( .A1(n10890), .A2(n10889), .A3(n10888), .A4(n10887), .ZN(
        n10896) );
  AOI22_X1 U13894 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13895 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13896 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13897 ( .A1(n11049), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10891) );
  NAND4_X1 U13898 ( .A1(n10894), .A2(n10893), .A3(n10892), .A4(n10891), .ZN(
        n10895) );
  NOR2_X1 U13899 ( .A1(n10896), .A2(n10895), .ZN(n10899) );
  AOI21_X1 U13900 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14732), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10897) );
  AOI21_X1 U13901 ( .B1(n10672), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10897), .ZN(
        n10898) );
  OAI21_X1 U13902 ( .B1(n11128), .B2(n10899), .A(n10898), .ZN(n10901) );
  XNOR2_X1 U13903 ( .A(n10902), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14736) );
  NAND2_X1 U13904 ( .A1(n14736), .A2(n10621), .ZN(n10900) );
  NAND2_X1 U13905 ( .A1(n10901), .A2(n10900), .ZN(n14460) );
  INV_X1 U13906 ( .A(n10903), .ZN(n10904) );
  INV_X1 U13907 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14723) );
  NAND2_X1 U13908 ( .A1(n10904), .A2(n14723), .ZN(n10905) );
  AND2_X1 U13909 ( .A1(n10935), .A2(n10905), .ZN(n14727) );
  AOI22_X1 U13910 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13911 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U13912 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U13913 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10906) );
  NAND4_X1 U13914 ( .A1(n10909), .A2(n10908), .A3(n10907), .A4(n10906), .ZN(
        n10915) );
  AOI22_X1 U13915 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13916 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13917 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13918 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10910) );
  NAND4_X1 U13919 ( .A1(n10913), .A2(n10912), .A3(n10911), .A4(n10910), .ZN(
        n10914) );
  OR2_X1 U13920 ( .A1(n10915), .A2(n10914), .ZN(n10918) );
  INV_X1 U13921 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n10916) );
  OAI22_X1 U13922 ( .A1(n10707), .A2(n10916), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14723), .ZN(n10917) );
  AOI21_X1 U13923 ( .B1(n11102), .B2(n10918), .A(n10917), .ZN(n10919) );
  MUX2_X1 U13924 ( .A(n14727), .B(n10919), .S(n11041), .Z(n14450) );
  NAND2_X1 U13925 ( .A1(n9875), .A2(n10920), .ZN(n14419) );
  INV_X1 U13926 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14442) );
  XNOR2_X1 U13927 ( .A(n10935), .B(n14442), .ZN(n14716) );
  AOI22_X1 U13928 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U13929 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13930 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13931 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10921) );
  NAND4_X1 U13932 ( .A1(n10924), .A2(n10923), .A3(n10922), .A4(n10921), .ZN(
        n10931) );
  AOI22_X1 U13933 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13934 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13935 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13936 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10926) );
  NAND4_X1 U13937 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n10930) );
  NOR2_X1 U13938 ( .A1(n10931), .A2(n10930), .ZN(n10933) );
  AOI22_X1 U13939 ( .A1(n10672), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n10577), .ZN(n10932) );
  OAI21_X1 U13940 ( .B1(n11128), .B2(n10933), .A(n10932), .ZN(n10934) );
  MUX2_X1 U13941 ( .A(n14716), .B(n10934), .S(n11041), .Z(n14438) );
  INV_X1 U13942 ( .A(n10937), .ZN(n10939) );
  INV_X1 U13943 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10938) );
  NAND2_X1 U13944 ( .A1(n10939), .A2(n10938), .ZN(n10940) );
  NAND2_X1 U13945 ( .A1(n10998), .A2(n10940), .ZN(n14708) );
  AOI22_X1 U13946 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13947 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n11108), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13948 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13949 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10941) );
  NAND4_X1 U13950 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n10951) );
  AOI22_X1 U13951 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U13952 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n11110), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13953 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13954 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11068), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10946) );
  NAND4_X1 U13955 ( .A1(n10949), .A2(n10948), .A3(n10947), .A4(n10946), .ZN(
        n10950) );
  NOR2_X1 U13956 ( .A1(n10951), .A2(n10950), .ZN(n10953) );
  AOI22_X1 U13957 ( .A1(n10672), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10577), .ZN(n10952) );
  OAI21_X1 U13958 ( .B1(n11128), .B2(n10953), .A(n10952), .ZN(n10954) );
  MUX2_X1 U13959 ( .A(n14708), .B(n10954), .S(n11041), .Z(n14421) );
  NOR2_X2 U13960 ( .A1(n14419), .A2(n9895), .ZN(n14404) );
  AOI22_X1 U13961 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13962 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13963 ( .A1(n10431), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13964 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10956) );
  NAND4_X1 U13965 ( .A1(n10959), .A2(n10958), .A3(n10957), .A4(n10956), .ZN(
        n10965) );
  AOI22_X1 U13966 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U13967 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U13968 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13969 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10960) );
  NAND4_X1 U13970 ( .A1(n10963), .A2(n10962), .A3(n10961), .A4(n10960), .ZN(
        n10964) );
  NOR2_X1 U13971 ( .A1(n10965), .A2(n10964), .ZN(n10981) );
  AOI22_X1 U13972 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U13973 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U13974 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U13975 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10966) );
  NAND4_X1 U13976 ( .A1(n10969), .A2(n10968), .A3(n10967), .A4(n10966), .ZN(
        n10975) );
  AOI22_X1 U13977 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U13978 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U13979 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U13980 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10970) );
  NAND4_X1 U13981 ( .A1(n10973), .A2(n10972), .A3(n10971), .A4(n10970), .ZN(
        n10974) );
  NOR2_X1 U13982 ( .A1(n10975), .A2(n10974), .ZN(n10982) );
  XOR2_X1 U13983 ( .A(n10981), .B(n10982), .Z(n10978) );
  INV_X1 U13984 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n10976) );
  INV_X1 U13985 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14409) );
  OAI22_X1 U13986 ( .A1(n10707), .A2(n10976), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14409), .ZN(n10977) );
  AOI21_X1 U13987 ( .B1(n10978), .B2(n11102), .A(n10977), .ZN(n10979) );
  XNOR2_X1 U13988 ( .A(n10998), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14698) );
  MUX2_X1 U13989 ( .A(n10979), .B(n14698), .S(n10621), .Z(n14408) );
  NOR2_X1 U13990 ( .A1(n10982), .A2(n10981), .ZN(n11006) );
  AOI22_X1 U13991 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U13992 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U13993 ( .A1(n10431), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U13994 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10984) );
  NAND4_X1 U13995 ( .A1(n10987), .A2(n10986), .A3(n10985), .A4(n10984), .ZN(
        n10993) );
  AOI22_X1 U13996 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U13997 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U13998 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U13999 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10988) );
  NAND4_X1 U14000 ( .A1(n10991), .A2(n10990), .A3(n10989), .A4(n10988), .ZN(
        n10992) );
  INV_X1 U14001 ( .A(n11005), .ZN(n10994) );
  XNOR2_X1 U14002 ( .A(n11006), .B(n10994), .ZN(n10997) );
  INV_X1 U14003 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n10995) );
  INV_X1 U14004 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14692) );
  OAI22_X1 U14005 ( .A1(n10707), .A2(n10995), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14692), .ZN(n10996) );
  AOI21_X1 U14006 ( .B1(n10997), .B2(n11102), .A(n10996), .ZN(n11003) );
  INV_X1 U14007 ( .A(n11000), .ZN(n11001) );
  NAND2_X1 U14008 ( .A1(n11001), .A2(n14692), .ZN(n11002) );
  AND2_X1 U14009 ( .A1(n11021), .A2(n11002), .ZN(n14694) );
  MUX2_X1 U14010 ( .A(n11003), .B(n14694), .S(n10621), .Z(n14392) );
  NAND2_X1 U14011 ( .A1(n11006), .A2(n11005), .ZN(n11025) );
  AOI22_X1 U14012 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U14013 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U14014 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U14015 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11007) );
  NAND4_X1 U14016 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n11016) );
  AOI22_X1 U14017 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U14018 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14019 ( .A1(n10431), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U14020 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11011) );
  NAND4_X1 U14021 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(
        n11015) );
  NOR2_X1 U14022 ( .A1(n11016), .A2(n11015), .ZN(n11026) );
  XOR2_X1 U14023 ( .A(n11025), .B(n11026), .Z(n11019) );
  INV_X1 U14024 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n11017) );
  INV_X1 U14025 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14683) );
  OAI22_X1 U14026 ( .A1(n10707), .A2(n11017), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14683), .ZN(n11018) );
  AOI21_X1 U14027 ( .B1(n11019), .B2(n11102), .A(n11018), .ZN(n11020) );
  XNOR2_X1 U14028 ( .A(n11021), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14681) );
  MUX2_X1 U14029 ( .A(n11020), .B(n14681), .S(n11104), .Z(n14379) );
  INV_X1 U14030 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11022) );
  NAND2_X1 U14031 ( .A1(n11023), .A2(n11022), .ZN(n11024) );
  NAND2_X1 U14032 ( .A1(n11079), .A2(n11024), .ZN(n14668) );
  NOR2_X1 U14033 ( .A1(n11026), .A2(n11025), .ZN(n11044) );
  AOI22_X1 U14034 ( .A1(n11027), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U14035 ( .A1(n11116), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U14036 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U14037 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11029) );
  NAND4_X1 U14038 ( .A1(n11032), .A2(n11031), .A3(n11030), .A4(n11029), .ZN(
        n11038) );
  AOI22_X1 U14039 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U14040 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14041 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U14042 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11033) );
  NAND4_X1 U14043 ( .A1(n11036), .A2(n11035), .A3(n11034), .A4(n11033), .ZN(
        n11037) );
  OR2_X1 U14044 ( .A1(n11038), .A2(n11037), .ZN(n11043) );
  XNOR2_X1 U14045 ( .A(n11044), .B(n11043), .ZN(n11040) );
  AOI22_X1 U14046 ( .A1(n10672), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n10577), .ZN(n11039) );
  OAI21_X1 U14047 ( .B1(n11040), .B2(n11128), .A(n11039), .ZN(n11042) );
  MUX2_X1 U14048 ( .A(n14668), .B(n11042), .S(n11041), .Z(n14367) );
  NAND2_X1 U14049 ( .A1(n11044), .A2(n11043), .ZN(n11061) );
  AOI22_X1 U14050 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U14051 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U14052 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U14053 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11045) );
  NAND4_X1 U14054 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(
        n11055) );
  AOI22_X1 U14055 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14056 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11052) );
  AOI22_X1 U14057 ( .A1(n9839), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11051) );
  AOI22_X1 U14058 ( .A1(n11049), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11050) );
  NAND4_X1 U14059 ( .A1(n11053), .A2(n11052), .A3(n11051), .A4(n11050), .ZN(
        n11054) );
  NOR2_X1 U14060 ( .A1(n11055), .A2(n11054), .ZN(n11062) );
  XOR2_X1 U14061 ( .A(n11061), .B(n11062), .Z(n11056) );
  NAND2_X1 U14062 ( .A1(n11056), .A2(n11102), .ZN(n11060) );
  AOI21_X1 U14063 ( .B1(n14657), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11057) );
  AOI21_X1 U14064 ( .B1(n10672), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11057), .ZN(
        n11059) );
  XNOR2_X1 U14065 ( .A(n11079), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14659) );
  AOI21_X1 U14066 ( .B1(n11060), .B2(n11059), .A(n11058), .ZN(n14353) );
  NOR2_X1 U14067 ( .A1(n11062), .A2(n11061), .ZN(n11085) );
  AOI22_X1 U14068 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10945), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14069 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10495), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14070 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14071 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11064) );
  NAND4_X1 U14072 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n11074) );
  AOI22_X1 U14073 ( .A1(n11108), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14074 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14075 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14076 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11069) );
  NAND4_X1 U14077 ( .A1(n11072), .A2(n11071), .A3(n11070), .A4(n11069), .ZN(
        n11073) );
  OR2_X1 U14078 ( .A1(n11074), .A2(n11073), .ZN(n11084) );
  INV_X1 U14079 ( .A(n11084), .ZN(n11075) );
  XNOR2_X1 U14080 ( .A(n11085), .B(n11075), .ZN(n11078) );
  INV_X1 U14081 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n11076) );
  INV_X1 U14082 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14653) );
  OAI22_X1 U14083 ( .A1(n10707), .A2(n11076), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14653), .ZN(n11077) );
  AOI21_X1 U14084 ( .B1(n11078), .B2(n11102), .A(n11077), .ZN(n11083) );
  INV_X1 U14085 ( .A(n11080), .ZN(n11081) );
  NAND2_X1 U14086 ( .A1(n11081), .A2(n14653), .ZN(n11082) );
  MUX2_X1 U14087 ( .A(n11083), .B(n14651), .S(n11104), .Z(n14342) );
  NAND2_X1 U14088 ( .A1(n11085), .A2(n11084), .ZN(n11106) );
  AOI22_X1 U14089 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10431), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U14090 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11108), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14091 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14092 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11088) );
  NAND4_X1 U14093 ( .A1(n11091), .A2(n11090), .A3(n11089), .A4(n11088), .ZN(
        n11099) );
  AOI22_X1 U14094 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14095 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U14096 ( .A1(n10495), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11095) );
  AOI22_X1 U14097 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11094) );
  NAND4_X1 U14098 ( .A1(n11097), .A2(n11096), .A3(n11095), .A4(n11094), .ZN(
        n11098) );
  NOR2_X1 U14099 ( .A1(n11099), .A2(n11098), .ZN(n11107) );
  XOR2_X1 U14100 ( .A(n11106), .B(n11107), .Z(n11103) );
  INV_X1 U14101 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n11100) );
  INV_X1 U14102 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14639) );
  OAI22_X1 U14103 ( .A1(n10707), .A2(n11100), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14639), .ZN(n11101) );
  AOI21_X1 U14104 ( .B1(n11103), .B2(n11102), .A(n11101), .ZN(n11105) );
  XNOR2_X1 U14105 ( .A(n11130), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14641) );
  MUX2_X1 U14106 ( .A(n11105), .B(n14641), .S(n11104), .Z(n14329) );
  NOR2_X1 U14107 ( .A1(n11107), .A2(n11106), .ZN(n11126) );
  AOI22_X1 U14108 ( .A1(n10945), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11108), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11115) );
  AOI22_X1 U14109 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11049), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14110 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11111), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14111 ( .A1(n10495), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11112) );
  NAND4_X1 U14112 ( .A1(n11115), .A2(n11114), .A3(n11113), .A4(n11112), .ZN(
        n11124) );
  AOI22_X1 U14113 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11116), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11122) );
  AOI22_X1 U14114 ( .A1(n11117), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10446), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11121) );
  AOI22_X1 U14115 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11120) );
  AOI22_X1 U14116 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11119) );
  NAND4_X1 U14117 ( .A1(n11122), .A2(n11121), .A3(n11120), .A4(n11119), .ZN(
        n11123) );
  NOR2_X1 U14118 ( .A1(n11124), .A2(n11123), .ZN(n11125) );
  XOR2_X1 U14119 ( .A(n11126), .B(n11125), .Z(n11129) );
  AOI22_X1 U14120 ( .A1(n10672), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n10577), .ZN(n11127) );
  OAI21_X1 U14121 ( .B1(n11129), .B2(n11128), .A(n11127), .ZN(n11131) );
  INV_X1 U14122 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14318) );
  XNOR2_X1 U14123 ( .A(n11136), .B(n14318), .ZN(n14627) );
  MUX2_X1 U14124 ( .A(n11131), .B(n14627), .S(n10621), .Z(n12673) );
  NAND2_X1 U14125 ( .A1(n12672), .A2(n12673), .ZN(n12671) );
  AOI22_X1 U14126 ( .A1(n10672), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11132), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11133) );
  INV_X1 U14127 ( .A(n11133), .ZN(n11134) );
  XNOR2_X2 U14128 ( .A(n12671), .B(n11134), .ZN(n12855) );
  AND3_X1 U14129 ( .A1(n20936), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U14130 ( .A1(n12855), .A2(n16025), .ZN(n11298) );
  INV_X1 U14131 ( .A(n11136), .ZN(n11137) );
  NAND2_X1 U14132 ( .A1(n11137), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11138) );
  INV_X1 U14133 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12880) );
  NAND2_X1 U14134 ( .A1(n20655), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11140) );
  NAND2_X1 U14135 ( .A1(n13940), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11139) );
  NAND2_X1 U14136 ( .A1(n11140), .A2(n11139), .ZN(n11160) );
  NAND2_X1 U14137 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20696), .ZN(
        n11161) );
  NAND2_X1 U14138 ( .A1(n11141), .A2(n11140), .ZN(n11152) );
  NAND2_X1 U14139 ( .A1(n11152), .A2(n11142), .ZN(n11145) );
  NAND2_X1 U14140 ( .A1(n11143), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11144) );
  MUX2_X1 U14141 ( .A(n20617), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11149) );
  NOR2_X1 U14142 ( .A1(n9823), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11146) );
  NAND2_X1 U14143 ( .A1(n11147), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11148) );
  NAND2_X1 U14144 ( .A1(n11179), .A2(n12649), .ZN(n11193) );
  NAND2_X1 U14145 ( .A1(n12649), .A2(n11163), .ZN(n11191) );
  XNOR2_X1 U14146 ( .A(n11150), .B(n11149), .ZN(n12645) );
  NAND2_X1 U14147 ( .A1(n12878), .A2(n10450), .ZN(n11164) );
  NAND2_X1 U14148 ( .A1(n14035), .A2(n11164), .ZN(n11157) );
  INV_X1 U14149 ( .A(n11157), .ZN(n11175) );
  MUX2_X1 U14150 ( .A(n11143), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11151) );
  XNOR2_X1 U14151 ( .A(n11152), .B(n11151), .ZN(n12646) );
  INV_X1 U14152 ( .A(n12646), .ZN(n11153) );
  AND2_X1 U14153 ( .A1(n11163), .A2(n11153), .ZN(n11154) );
  INV_X1 U14154 ( .A(n11154), .ZN(n11174) );
  AOI211_X1 U14155 ( .C1(n12646), .C2(n11185), .A(n11154), .B(n11157), .ZN(
        n11173) );
  INV_X1 U14156 ( .A(n11161), .ZN(n11155) );
  AOI21_X1 U14157 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n10323), .A(
        n11155), .ZN(n11156) );
  AND2_X1 U14158 ( .A1(n11163), .A2(n11156), .ZN(n11159) );
  OAI21_X1 U14159 ( .B1(n20266), .B2(n10454), .A(n11156), .ZN(n11158) );
  OAI22_X1 U14160 ( .A1(n11179), .A2(n11159), .B1(n11158), .B2(n11157), .ZN(
        n11167) );
  INV_X1 U14161 ( .A(n11167), .ZN(n11171) );
  XNOR2_X1 U14162 ( .A(n11161), .B(n11160), .ZN(n12644) );
  NOR2_X1 U14163 ( .A1(n10450), .A2(n20936), .ZN(n11162) );
  AOI22_X1 U14164 ( .A1(n11185), .A2(n12644), .B1(n11164), .B2(n11165), .ZN(
        n11168) );
  INV_X1 U14165 ( .A(n11168), .ZN(n11170) );
  INV_X1 U14166 ( .A(n11165), .ZN(n11166) );
  NAND2_X1 U14167 ( .A1(n11166), .A2(n20274), .ZN(n11183) );
  AOI22_X1 U14168 ( .A1(n12644), .A2(n11183), .B1(n11168), .B2(n11167), .ZN(
        n11169) );
  AOI21_X1 U14169 ( .B1(n11171), .B2(n11170), .A(n11169), .ZN(n11172) );
  OAI22_X1 U14170 ( .A1(n11175), .A2(n11174), .B1(n11173), .B2(n11172), .ZN(
        n11178) );
  NAND2_X1 U14171 ( .A1(n11176), .A2(n12645), .ZN(n11177) );
  AOI22_X1 U14172 ( .A1(n11179), .A2(n12645), .B1(n11178), .B2(n11177), .ZN(
        n11188) );
  INV_X1 U14173 ( .A(n12647), .ZN(n11182) );
  NOR2_X1 U14174 ( .A1(n11185), .A2(n11182), .ZN(n11187) );
  INV_X1 U14175 ( .A(n11183), .ZN(n11184) );
  NAND3_X1 U14176 ( .A1(n11185), .A2(n11184), .A3(n12647), .ZN(n11186) );
  OAI21_X1 U14177 ( .B1(n11188), .B2(n11187), .A(n11186), .ZN(n11189) );
  AOI21_X1 U14178 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20936), .A(
        n11189), .ZN(n11190) );
  NAND2_X1 U14179 ( .A1(n11191), .A2(n11190), .ZN(n11192) );
  AND2_X1 U14180 ( .A1(n13624), .A2(n20266), .ZN(n11194) );
  NOR2_X1 U14181 ( .A1(n11195), .A2(n11194), .ZN(n13596) );
  NAND2_X1 U14182 ( .A1(n13596), .A2(n10458), .ZN(n15859) );
  NAND2_X1 U14183 ( .A1(n20920), .A2(n11198), .ZN(n20939) );
  NAND2_X1 U14184 ( .A1(n20939), .A2(n20936), .ZN(n11196) );
  NAND2_X1 U14185 ( .A1(n21137), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11197) );
  NAND2_X1 U14186 ( .A1(n20936), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15867) );
  NAND2_X1 U14187 ( .A1(n11197), .A2(n15867), .ZN(n13726) );
  INV_X1 U14188 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21028) );
  NOR2_X1 U14189 ( .A1(n16162), .A2(n21028), .ZN(n14798) );
  AOI21_X1 U14190 ( .B1(n16015), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14798), .ZN(n11199) );
  OAI21_X1 U14191 ( .B1(n14030), .B2(n16022), .A(n11199), .ZN(n11200) );
  INV_X1 U14192 ( .A(n11200), .ZN(n11297) );
  NAND2_X1 U14193 ( .A1(n11207), .A2(n11206), .ZN(n11219) );
  NAND2_X1 U14194 ( .A1(n11219), .A2(n11220), .ZN(n11218) );
  NAND2_X1 U14195 ( .A1(n11218), .A2(n11201), .ZN(n11243) );
  OAI211_X1 U14196 ( .C1(n11201), .C2(n11218), .A(n11243), .B(n13629), .ZN(
        n11202) );
  OAI21_X2 U14197 ( .B1(n20520), .B2(n11239), .A(n11202), .ZN(n11228) );
  INV_X1 U14198 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13917) );
  XNOR2_X1 U14199 ( .A(n11228), .B(n13917), .ZN(n13852) );
  NAND2_X1 U14200 ( .A1(n20266), .A2(n20287), .ZN(n11221) );
  OAI21_X1 U14201 ( .B1(n13453), .B2(n11207), .A(n11221), .ZN(n11203) );
  INV_X1 U14202 ( .A(n11203), .ZN(n11204) );
  NAND2_X2 U14203 ( .A1(n13723), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13725) );
  OR2_X1 U14204 ( .A1(n11205), .A2(n12878), .ZN(n11211) );
  XNOR2_X1 U14205 ( .A(n11207), .B(n11206), .ZN(n11208) );
  OAI211_X1 U14206 ( .C1(n11208), .C2(n13453), .A(n10428), .B(n10450), .ZN(
        n11209) );
  INV_X1 U14207 ( .A(n11209), .ZN(n11210) );
  NAND2_X1 U14208 ( .A1(n11211), .A2(n11210), .ZN(n11212) );
  NAND2_X1 U14209 ( .A1(n13672), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11215) );
  INV_X1 U14210 ( .A(n11212), .ZN(n11213) );
  OR2_X1 U14211 ( .A1(n13725), .A2(n11213), .ZN(n11214) );
  INV_X1 U14212 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11216) );
  NAND2_X1 U14213 ( .A1(n11217), .A2(n11230), .ZN(n11225) );
  OAI21_X1 U14214 ( .B1(n11220), .B2(n11219), .A(n11218), .ZN(n11223) );
  INV_X1 U14215 ( .A(n11221), .ZN(n11222) );
  AOI21_X1 U14216 ( .B1(n11223), .B2(n13629), .A(n11222), .ZN(n11224) );
  NAND2_X1 U14217 ( .A1(n11225), .A2(n11224), .ZN(n13748) );
  NAND2_X1 U14218 ( .A1(n11226), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11227) );
  NAND2_X1 U14219 ( .A1(n11228), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11229) );
  XNOR2_X1 U14220 ( .A(n11243), .B(n11241), .ZN(n11232) );
  NAND2_X1 U14221 ( .A1(n11232), .A2(n13629), .ZN(n11233) );
  NAND2_X1 U14222 ( .A1(n11234), .A2(n11233), .ZN(n11236) );
  INV_X1 U14223 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11235) );
  XNOR2_X1 U14224 ( .A(n11236), .B(n11235), .ZN(n13902) );
  NAND2_X1 U14225 ( .A1(n13901), .A2(n13902), .ZN(n11238) );
  NAND2_X1 U14226 ( .A1(n11236), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11237) );
  OR2_X1 U14227 ( .A1(n11240), .A2(n11239), .ZN(n11247) );
  INV_X1 U14228 ( .A(n11241), .ZN(n11242) );
  NOR2_X1 U14229 ( .A1(n11243), .A2(n11242), .ZN(n11245) );
  NAND2_X1 U14230 ( .A1(n11245), .A2(n11244), .ZN(n11257) );
  OAI211_X1 U14231 ( .C1(n11245), .C2(n11244), .A(n11257), .B(n13629), .ZN(
        n11246) );
  NAND2_X1 U14232 ( .A1(n11247), .A2(n11246), .ZN(n11248) );
  INV_X1 U14233 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16155) );
  XNOR2_X1 U14234 ( .A(n11248), .B(n16155), .ZN(n14076) );
  NAND2_X1 U14235 ( .A1(n14075), .A2(n14076), .ZN(n11250) );
  NAND2_X1 U14236 ( .A1(n11248), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11249) );
  XNOR2_X1 U14237 ( .A(n11257), .B(n11258), .ZN(n11252) );
  NAND2_X1 U14238 ( .A1(n11252), .A2(n13629), .ZN(n11253) );
  NAND2_X1 U14239 ( .A1(n11254), .A2(n11253), .ZN(n11255) );
  INV_X1 U14240 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16165) );
  XNOR2_X1 U14241 ( .A(n11255), .B(n16165), .ZN(n14056) );
  NAND2_X1 U14242 ( .A1(n11256), .A2(n11230), .ZN(n11262) );
  INV_X1 U14243 ( .A(n11257), .ZN(n11259) );
  NAND2_X1 U14244 ( .A1(n11259), .A2(n11258), .ZN(n11269) );
  XNOR2_X1 U14245 ( .A(n11269), .B(n11267), .ZN(n11260) );
  NAND2_X1 U14246 ( .A1(n11260), .A2(n13629), .ZN(n11261) );
  NAND2_X1 U14247 ( .A1(n11262), .A2(n11261), .ZN(n11263) );
  OR2_X1 U14248 ( .A1(n11263), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16018) );
  NAND2_X1 U14249 ( .A1(n11263), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16017) );
  NAND2_X4 U14250 ( .A1(n11266), .A2(n11265), .ZN(n14729) );
  NAND2_X1 U14251 ( .A1(n13629), .A2(n11267), .ZN(n11268) );
  OR2_X1 U14252 ( .A1(n11269), .A2(n11268), .ZN(n11270) );
  NAND2_X1 U14253 ( .A1(n14729), .A2(n11270), .ZN(n14139) );
  OR2_X1 U14254 ( .A1(n14139), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11271) );
  NAND2_X1 U14255 ( .A1(n14139), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11272) );
  INV_X1 U14256 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16152) );
  NOR2_X1 U14257 ( .A1(n14729), .A2(n16152), .ZN(n11274) );
  NAND2_X1 U14258 ( .A1(n14729), .A2(n16152), .ZN(n11275) );
  INV_X1 U14259 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11280) );
  AND2_X1 U14260 ( .A1(n14729), .A2(n11280), .ZN(n11277) );
  INV_X1 U14261 ( .A(n14729), .ZN(n11294) );
  INV_X1 U14262 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11279) );
  NAND2_X1 U14263 ( .A1(n11294), .A2(n11279), .ZN(n14753) );
  NAND2_X1 U14264 ( .A1(n14729), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14265 ( .A1(n14753), .A2(n11276), .ZN(n15983) );
  INV_X1 U14266 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11278) );
  NAND2_X1 U14267 ( .A1(n14729), .A2(n11278), .ZN(n15984) );
  NAND2_X1 U14268 ( .A1(n15983), .A2(n15984), .ZN(n14752) );
  INV_X2 U14269 ( .A(n14729), .ZN(n14751) );
  NAND2_X1 U14270 ( .A1(n14751), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15992) );
  INV_X1 U14271 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16121) );
  NAND2_X1 U14272 ( .A1(n14729), .A2(n16121), .ZN(n11282) );
  NAND2_X1 U14273 ( .A1(n15992), .A2(n11282), .ZN(n14771) );
  INV_X1 U14274 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14889) );
  NAND2_X1 U14275 ( .A1(n14729), .A2(n14889), .ZN(n14888) );
  NAND2_X1 U14276 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11283) );
  NAND2_X1 U14277 ( .A1(n14729), .A2(n11283), .ZN(n14769) );
  NAND2_X1 U14278 ( .A1(n14888), .A2(n14769), .ZN(n11284) );
  NOR2_X1 U14279 ( .A1(n14771), .A2(n11284), .ZN(n14748) );
  NAND2_X1 U14280 ( .A1(n14748), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11285) );
  NAND2_X1 U14281 ( .A1(n14751), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11286) );
  NAND2_X1 U14282 ( .A1(n15992), .A2(n11286), .ZN(n14749) );
  NOR2_X1 U14283 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14885) );
  NAND2_X1 U14284 ( .A1(n14885), .A2(n14889), .ZN(n11287) );
  XNOR2_X1 U14285 ( .A(n14729), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14740) );
  NAND2_X1 U14286 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14866) );
  INV_X1 U14287 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14884) );
  NOR2_X1 U14288 ( .A1(n14866), .A2(n14884), .ZN(n11290) );
  INV_X1 U14289 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16085) );
  INV_X1 U14290 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14794) );
  INV_X1 U14291 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11291) );
  INV_X1 U14292 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14857) );
  INV_X1 U14293 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14871) );
  NAND2_X1 U14294 ( .A1(n14857), .A2(n14871), .ZN(n11292) );
  OAI21_X1 U14295 ( .B1(n14676), .B2(n11292), .A(n14751), .ZN(n14671) );
  NAND3_X1 U14296 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14805) );
  INV_X1 U14297 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16036) );
  NAND2_X1 U14298 ( .A1(n14660), .A2(n14729), .ZN(n14677) );
  NAND2_X1 U14299 ( .A1(n14661), .A2(n14677), .ZN(n11293) );
  NOR2_X1 U14300 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14839) );
  AND2_X1 U14301 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14838) );
  NAND2_X1 U14302 ( .A1(n14729), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11295) );
  INV_X1 U14303 ( .A(n20080), .ZN(n11296) );
  INV_X1 U14304 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U14305 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11299) );
  NOR2_X4 U14306 ( .A1(n18962), .A2(n11312), .ZN(n11378) );
  INV_X1 U14307 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17162) );
  OR3_X2 U14308 ( .A1(n18962), .A2(n18972), .A3(n17014), .ZN(n11340) );
  INV_X2 U14309 ( .A(n17242), .ZN(n11331) );
  AOI22_X1 U14310 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11331), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11304) );
  NOR2_X2 U14311 ( .A1(n11308), .A2(n11310), .ZN(n11300) );
  INV_X1 U14312 ( .A(n17014), .ZN(n11302) );
  NAND2_X2 U14313 ( .A1(n11302), .A2(n11301), .ZN(n11376) );
  INV_X4 U14314 ( .A(n11376), .ZN(n17298) );
  AOI22_X1 U14315 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11303) );
  OAI211_X1 U14316 ( .C1(n11489), .C2(n18325), .A(n11304), .B(n11303), .ZN(
        n11306) );
  AOI22_X1 U14317 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11518), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11315) );
  NOR2_X2 U14318 ( .A1(n11311), .A2(n11308), .ZN(n11309) );
  AOI22_X1 U14319 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11392), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11314) );
  INV_X2 U14320 ( .A(n17219), .ZN(n14282) );
  OR2_X2 U14321 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11312), .ZN(
        n17172) );
  NAND2_X1 U14322 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11313) );
  AOI22_X1 U14323 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11378), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11318) );
  OAI21_X1 U14324 ( .B1(n17296), .B2(n18568), .A(n11318), .ZN(n11322) );
  INV_X1 U14325 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18320) );
  AOI22_X1 U14326 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11518), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11319) );
  OAI211_X1 U14327 ( .C1(n11489), .C2(n18320), .A(n11320), .B(n11319), .ZN(
        n11321) );
  AOI22_X1 U14328 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11328) );
  INV_X4 U14329 ( .A(n15798), .ZN(n17191) );
  INV_X1 U14330 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17184) );
  INV_X1 U14331 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U14332 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11324) );
  OAI21_X1 U14333 ( .B1(n10327), .B2(n17181), .A(n11324), .ZN(n11325) );
  INV_X1 U14334 ( .A(n11325), .ZN(n11326) );
  INV_X1 U14335 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18968) );
  NOR2_X1 U14336 ( .A1(n17496), .A2(n18968), .ZN(n11346) );
  INV_X1 U14337 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18317) );
  AOI22_X1 U14338 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11330) );
  OAI21_X1 U14339 ( .B1(n11489), .B2(n18317), .A(n11330), .ZN(n11335) );
  INV_X1 U14340 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18565) );
  AOI22_X1 U14341 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14342 ( .A1(n11309), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11518), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11332) );
  OAI211_X1 U14343 ( .C1(n17296), .C2(n18565), .A(n11333), .B(n11332), .ZN(
        n11334) );
  INV_X1 U14344 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U14345 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11392), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11336) );
  OAI21_X1 U14346 ( .B1(n9858), .B2(n17203), .A(n11336), .ZN(n11338) );
  INV_X4 U14347 ( .A(n17145), .ZN(n17228) );
  AOI22_X1 U14348 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11339) );
  INV_X1 U14349 ( .A(n11339), .ZN(n11342) );
  NAND2_X1 U14350 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17978), .ZN(
        n17977) );
  NOR2_X1 U14351 ( .A1(n17977), .A2(n17970), .ZN(n17969) );
  NOR2_X1 U14352 ( .A1(n11346), .A2(n17969), .ZN(n17955) );
  XNOR2_X1 U14353 ( .A(n18270), .B(n11347), .ZN(n17954) );
  NAND2_X1 U14354 ( .A1(n17496), .A2(n11317), .ZN(n11362) );
  AOI22_X1 U14355 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11392), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11354) );
  INV_X1 U14356 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18385) );
  AOI22_X1 U14357 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9804), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11348) );
  OAI21_X1 U14358 ( .B1(n10328), .B2(n18385), .A(n11348), .ZN(n11352) );
  AOI22_X1 U14359 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14360 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11349) );
  OAI211_X1 U14361 ( .C1(n11489), .C2(n18330), .A(n11350), .B(n11349), .ZN(
        n11351) );
  AOI211_X1 U14362 ( .C1(n17276), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n11352), .B(n11351), .ZN(n11353) );
  OAI211_X1 U14363 ( .C1(n17307), .C2(n17258), .A(n11354), .B(n11353), .ZN(
        n11355) );
  INV_X1 U14364 ( .A(n11355), .ZN(n11359) );
  AOI22_X1 U14365 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11356) );
  OAI21_X1 U14366 ( .B1(n11340), .B2(n17257), .A(n11356), .ZN(n11357) );
  XNOR2_X1 U14367 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11361), .ZN(
        n17942) );
  AOI22_X1 U14368 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11372) );
  INV_X1 U14369 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18575) );
  AOI22_X1 U14370 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14371 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11363) );
  OAI211_X1 U14372 ( .C1(n17296), .C2(n18575), .A(n11364), .B(n11363), .ZN(
        n11370) );
  AOI22_X1 U14373 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14374 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14375 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11366) );
  NAND2_X1 U14376 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11365) );
  NAND4_X1 U14377 ( .A1(n11368), .A2(n11367), .A3(n11366), .A4(n11365), .ZN(
        n11369) );
  AOI211_X1 U14378 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n11370), .B(n11369), .ZN(n11371) );
  XNOR2_X1 U14379 ( .A(n11375), .B(n11568), .ZN(n11373) );
  XNOR2_X1 U14380 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11373), .ZN(
        n17933) );
  NOR2_X1 U14381 ( .A1(n17934), .A2(n17933), .ZN(n17932) );
  AND2_X1 U14382 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11373), .ZN(
        n11374) );
  NOR2_X1 U14383 ( .A1(n17932), .A2(n11374), .ZN(n11389) );
  INV_X1 U14384 ( .A(n11568), .ZN(n17480) );
  AOI22_X1 U14385 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11377) );
  OAI21_X1 U14386 ( .B1(n11376), .B2(n17120), .A(n11377), .ZN(n11387) );
  AOI22_X1 U14387 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14388 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11379) );
  OAI21_X1 U14389 ( .B1(n11489), .B2(n18340), .A(n11379), .ZN(n11383) );
  INV_X1 U14390 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18578) );
  AOI22_X1 U14391 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14392 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11380) );
  OAI211_X1 U14393 ( .C1(n17296), .C2(n18578), .A(n11381), .B(n11380), .ZN(
        n11382) );
  AOI211_X1 U14394 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n11383), .B(n11382), .ZN(n11384) );
  OAI211_X1 U14395 ( .C1(n9858), .C2(n17116), .A(n11385), .B(n11384), .ZN(
        n11386) );
  XOR2_X1 U14396 ( .A(n11391), .B(n17476), .Z(n11388) );
  XNOR2_X1 U14397 ( .A(n11389), .B(n11388), .ZN(n17918) );
  INV_X1 U14398 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18246) );
  NOR2_X1 U14399 ( .A1(n11389), .A2(n11388), .ZN(n11390) );
  INV_X1 U14400 ( .A(n17476), .ZN(n11566) );
  AOI22_X1 U14401 ( .A1(n9804), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11378), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11402) );
  INV_X1 U14402 ( .A(n11392), .ZN(n17291) );
  INV_X2 U14403 ( .A(n17291), .ZN(n15791) );
  AOI22_X1 U14404 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14405 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11393) );
  OAI211_X1 U14406 ( .C1(n11489), .C2(n18345), .A(n11394), .B(n11393), .ZN(
        n11400) );
  AOI22_X1 U14407 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14408 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14409 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11396) );
  NAND2_X1 U14410 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11395) );
  NAND4_X1 U14411 ( .A1(n11398), .A2(n11397), .A3(n11396), .A4(n11395), .ZN(
        n11399) );
  AOI211_X1 U14412 ( .C1(n9810), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n11400), .B(n11399), .ZN(n11401) );
  XNOR2_X1 U14413 ( .A(n11405), .B(n17903), .ZN(n11403) );
  XNOR2_X1 U14414 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n11403), .ZN(
        n17908) );
  INV_X1 U14415 ( .A(n17903), .ZN(n17902) );
  INV_X1 U14416 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U14417 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11406) );
  OAI21_X1 U14418 ( .B1(n11340), .B2(n17057), .A(n11406), .ZN(n11415) );
  AOI22_X1 U14419 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11413) );
  INV_X1 U14420 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14258) );
  AOI22_X1 U14421 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11378), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11407) );
  OAI21_X1 U14422 ( .B1(n17296), .B2(n14258), .A(n11407), .ZN(n11411) );
  INV_X1 U14423 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18354) );
  AOI22_X1 U14424 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14425 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11408) );
  OAI211_X1 U14426 ( .C1(n11489), .C2(n18354), .A(n11409), .B(n11408), .ZN(
        n11410) );
  AOI211_X1 U14427 ( .C1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n9810), .A(
        n11411), .B(n11410), .ZN(n11412) );
  OAI211_X1 U14428 ( .C1(n17172), .C2(n17220), .A(n11413), .B(n11412), .ZN(
        n11414) );
  OAI21_X1 U14429 ( .B1(n16519), .B2(n13310), .A(n17779), .ZN(n11416) );
  NOR2_X1 U14430 ( .A1(n17891), .A2(n18210), .ZN(n17890) );
  NOR2_X1 U14431 ( .A1(n17780), .A2(n11416), .ZN(n11417) );
  NOR2_X2 U14432 ( .A1(n17890), .A2(n11417), .ZN(n11420) );
  NAND2_X1 U14433 ( .A1(n11420), .A2(n18212), .ZN(n17870) );
  NOR2_X2 U14434 ( .A1(n17870), .A2(n17877), .ZN(n17857) );
  INV_X1 U14435 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18198) );
  INV_X1 U14436 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18139) );
  INV_X1 U14437 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U14438 ( .A1(n17803), .A2(n10337), .ZN(n11419) );
  NAND2_X1 U14439 ( .A1(n11419), .A2(n17779), .ZN(n17766) );
  NOR2_X2 U14440 ( .A1(n11420), .A2(n18212), .ZN(n18177) );
  NAND2_X1 U14441 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18182) );
  NOR2_X1 U14442 ( .A1(n18182), .A2(n17842), .ZN(n18155) );
  NAND2_X1 U14443 ( .A1(n18155), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18137) );
  NAND2_X1 U14444 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18144), .ZN(
        n18086) );
  INV_X1 U14445 ( .A(n18086), .ZN(n18114) );
  INV_X1 U14446 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18116) );
  NAND2_X1 U14447 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17701) );
  INV_X1 U14448 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17751) );
  INV_X1 U14449 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18052) );
  NAND2_X1 U14450 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18062) );
  NOR3_X1 U14451 ( .A1(n17751), .A2(n18052), .A3(n18062), .ZN(n17702) );
  NAND2_X1 U14452 ( .A1(n17702), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11423) );
  NOR2_X1 U14453 ( .A1(n17752), .A2(n11423), .ZN(n17677) );
  NOR2_X1 U14454 ( .A1(n17701), .A2(n11423), .ZN(n18007) );
  INV_X1 U14455 ( .A(n18007), .ZN(n17986) );
  INV_X1 U14456 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17691) );
  NOR2_X1 U14457 ( .A1(n17986), .A2(n17691), .ZN(n17672) );
  NAND2_X1 U14458 ( .A1(n11422), .A2(n17672), .ZN(n18026) );
  NAND2_X1 U14459 ( .A1(n17779), .A2(n17751), .ZN(n17750) );
  NOR2_X1 U14460 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17750), .ZN(
        n11424) );
  INV_X1 U14461 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18050) );
  NAND2_X1 U14462 ( .A1(n11424), .A2(n18050), .ZN(n17711) );
  INV_X1 U14463 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18059) );
  NAND3_X1 U14464 ( .A1(n17704), .A2(n18059), .A3(n17691), .ZN(n11425) );
  INV_X1 U14465 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17676) );
  NAND2_X1 U14466 ( .A1(n17671), .A2(n17676), .ZN(n17670) );
  NAND3_X1 U14467 ( .A1(n17677), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17670), .ZN(n11431) );
  NAND2_X1 U14468 ( .A1(n11431), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11430) );
  INV_X1 U14469 ( .A(n17670), .ZN(n17660) );
  INV_X1 U14470 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18008) );
  NAND2_X1 U14471 ( .A1(n17877), .A2(n18008), .ZN(n11428) );
  INV_X1 U14472 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17649) );
  NAND2_X1 U14473 ( .A1(n17877), .A2(n11431), .ZN(n17659) );
  INV_X1 U14474 ( .A(n17659), .ZN(n11433) );
  NAND2_X1 U14475 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11558) );
  INV_X1 U14476 ( .A(n11558), .ZN(n17988) );
  INV_X1 U14477 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17994) );
  NOR2_X1 U14478 ( .A1(n17877), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16512) );
  NAND2_X1 U14479 ( .A1(n12912), .A2(n12911), .ZN(n11436) );
  XNOR2_X1 U14480 ( .A(n11436), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15831) );
  OAI22_X1 U14481 ( .A1(n18980), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18821), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U14482 ( .A1(n18819), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11549) );
  NOR2_X1 U14483 ( .A1(n11550), .A2(n11549), .ZN(n11437) );
  OAI21_X1 U14484 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18972), .A(
        n11438), .ZN(n11439) );
  OAI22_X1 U14485 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18830), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11439), .ZN(n11445) );
  NOR2_X1 U14486 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18830), .ZN(
        n11440) );
  NAND2_X1 U14487 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11439), .ZN(
        n11444) );
  AOI22_X1 U14488 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11445), .B1(
        n11440), .B2(n11444), .ZN(n11448) );
  OAI21_X1 U14489 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18819), .A(
        n11549), .ZN(n11554) );
  NOR2_X1 U14490 ( .A1(n11550), .A2(n11554), .ZN(n11447) );
  OAI21_X1 U14491 ( .B1(n11443), .B2(n11442), .A(n11448), .ZN(n11441) );
  AND2_X1 U14492 ( .A1(n11444), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11446) );
  OAI22_X1 U14493 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18783), .B1(
        n11446), .B2(n11445), .ZN(n11551) );
  AOI22_X1 U14494 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11449) );
  OAI21_X1 U14495 ( .B1(n17145), .B2(n18568), .A(n11449), .ZN(n11456) );
  INV_X1 U14496 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U14497 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11454) );
  INV_X1 U14498 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18723) );
  AOI22_X1 U14499 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11451) );
  OAI21_X1 U14500 ( .B1(n11489), .B2(n18723), .A(n11451), .ZN(n11453) );
  AOI22_X1 U14501 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11452) );
  AOI211_X4 U14502 ( .C1(n9808), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n11456), .B(n11455), .ZN(n19008) );
  AOI22_X1 U14503 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11457) );
  OAI21_X1 U14504 ( .B1(n11376), .B2(n18330), .A(n11457), .ZN(n11466) );
  AOI22_X1 U14505 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14506 ( .A1(n17276), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11458) );
  OAI21_X1 U14507 ( .B1(n17307), .B2(n17257), .A(n11458), .ZN(n11462) );
  INV_X1 U14508 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18737) );
  AOI22_X1 U14509 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14510 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11459) );
  OAI211_X1 U14511 ( .C1(n11489), .C2(n18737), .A(n11460), .B(n11459), .ZN(
        n11461) );
  AOI211_X1 U14512 ( .C1(n9804), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n11462), .B(n11461), .ZN(n11463) );
  OAI211_X1 U14513 ( .C1(n17242), .C2(n17146), .A(n11464), .B(n11463), .ZN(
        n11465) );
  AOI22_X1 U14514 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11467) );
  OAI21_X1 U14515 ( .B1(n11376), .B2(n18325), .A(n11467), .ZN(n11476) );
  INV_X1 U14516 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14279) );
  AOI22_X1 U14517 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11474) );
  INV_X1 U14518 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14274) );
  AOI22_X1 U14519 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11468) );
  OAI21_X1 U14520 ( .B1(n17296), .B2(n14274), .A(n11468), .ZN(n11472) );
  INV_X1 U14521 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18730) );
  AOI22_X1 U14522 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11518), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14523 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11469) );
  OAI211_X1 U14524 ( .C1(n11489), .C2(n18730), .A(n11470), .B(n11469), .ZN(
        n11471) );
  AOI211_X1 U14525 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n11472), .B(n11471), .ZN(n11473) );
  OAI211_X1 U14526 ( .C1(n15798), .C2(n14279), .A(n11474), .B(n11473), .ZN(
        n11475) );
  AOI22_X1 U14527 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11477) );
  OAI21_X1 U14528 ( .B1(n11376), .B2(n18345), .A(n11477), .ZN(n11487) );
  AOI22_X1 U14529 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11485) );
  INV_X1 U14530 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14531 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11478) );
  OAI21_X1 U14532 ( .B1(n13764), .B2(n11479), .A(n11478), .ZN(n11483) );
  INV_X1 U14533 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18759) );
  AOI22_X1 U14534 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14535 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11480) );
  OAI211_X1 U14536 ( .C1(n11489), .C2(n18759), .A(n11481), .B(n11480), .ZN(
        n11482) );
  AOI211_X1 U14537 ( .C1(n17276), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n11483), .B(n11482), .ZN(n11484) );
  OAI211_X1 U14538 ( .C1(n17307), .C2(n17045), .A(n11485), .B(n11484), .ZN(
        n11486) );
  AOI22_X1 U14539 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11488) );
  OAI21_X1 U14540 ( .B1(n11376), .B2(n18340), .A(n11488), .ZN(n11498) );
  INV_X1 U14541 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U14542 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11496) );
  INV_X1 U14543 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14221) );
  AOI22_X1 U14544 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9809), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11490) );
  OAI21_X1 U14545 ( .B1(n17296), .B2(n14221), .A(n11490), .ZN(n11494) );
  AOI22_X1 U14546 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U14547 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11518), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11491) );
  OAI211_X1 U14548 ( .C1(n10328), .C2(n17120), .A(n11492), .B(n11491), .ZN(
        n11493) );
  AOI211_X1 U14549 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n11494), .B(n11493), .ZN(n11495) );
  OAI211_X1 U14550 ( .C1(n17242), .C2(n17114), .A(n11496), .B(n11495), .ZN(
        n11497) );
  NOR2_X1 U14551 ( .A1(n13761), .A2(n16646), .ZN(n11530) );
  INV_X1 U14552 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18716) );
  AOI22_X1 U14553 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14554 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11499) );
  OAI211_X1 U14555 ( .C1(n11489), .C2(n18716), .A(n11500), .B(n11499), .ZN(
        n11506) );
  AOI22_X1 U14556 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14557 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14558 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11502) );
  NAND2_X1 U14559 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11501) );
  NAND4_X1 U14560 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11505) );
  AOI22_X1 U14561 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17117), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17292), .ZN(n11509) );
  OAI21_X1 U14562 ( .B1(n18397), .B2(n11450), .A(n11509), .ZN(n11517) );
  AOI22_X1 U14563 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n15791), .ZN(n11516) );
  INV_X1 U14564 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18771) );
  AOI22_X1 U14565 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n9810), .ZN(n11510) );
  OAI21_X1 U14566 ( .B1(n18771), .B2(n11489), .A(n11510), .ZN(n11514) );
  INV_X1 U14567 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U14568 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14569 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17297), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11511) );
  OAI211_X1 U14570 ( .C1(n17296), .C2(n17054), .A(n11512), .B(n11511), .ZN(
        n11513) );
  AOI211_X1 U14571 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n11514), .B(n11513), .ZN(n11515) );
  INV_X1 U14572 ( .A(n11532), .ZN(n11529) );
  AOI22_X1 U14573 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11528) );
  INV_X1 U14574 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14291) );
  AOI22_X1 U14575 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14576 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11519) );
  OAI211_X1 U14577 ( .C1(n17296), .C2(n14291), .A(n11520), .B(n11519), .ZN(
        n11526) );
  AOI22_X1 U14578 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14579 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14580 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9809), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11522) );
  NAND2_X1 U14581 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11521) );
  NAND4_X1 U14582 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11525) );
  AOI211_X1 U14583 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n11526), .B(n11525), .ZN(n11527) );
  NAND2_X1 U14584 ( .A1(n11539), .A2(n11556), .ZN(n13299) );
  NAND2_X1 U14585 ( .A1(n17541), .A2(n13299), .ZN(n16629) );
  NOR2_X1 U14586 ( .A1(n18337), .A2(n11556), .ZN(n13297) );
  NOR2_X1 U14587 ( .A1(n18314), .A2(n16646), .ZN(n11542) );
  OAI21_X1 U14588 ( .B1(n18350), .B2(n9824), .A(n11542), .ZN(n13301) );
  OAI21_X1 U14589 ( .B1(n11531), .B2(n13297), .A(n13301), .ZN(n11538) );
  NOR2_X1 U14590 ( .A1(n11556), .A2(n11533), .ZN(n13305) );
  NOR2_X1 U14591 ( .A1(n11531), .A2(n13305), .ZN(n11537) );
  AOI22_X1 U14592 ( .A1(n18327), .A2(n11532), .B1(n18332), .B2(n9824), .ZN(
        n11536) );
  NAND2_X1 U14593 ( .A1(n17393), .A2(n11533), .ZN(n11534) );
  OR2_X1 U14594 ( .A1(n11556), .A2(n11543), .ZN(n11547) );
  AOI22_X1 U14595 ( .A1(n11534), .A2(n13762), .B1(n11547), .B2(n11533), .ZN(
        n11535) );
  OAI211_X1 U14596 ( .C1(n11537), .C2(n17503), .A(n11536), .B(n11535), .ZN(
        n13300) );
  NAND2_X1 U14597 ( .A1(n11539), .A2(n11540), .ZN(n15811) );
  NOR2_X1 U14598 ( .A1(n19008), .A2(n11544), .ZN(n18786) );
  NOR2_X1 U14599 ( .A1(n11543), .A2(n11542), .ZN(n19016) );
  NAND2_X1 U14600 ( .A1(n11545), .A2(n13762), .ZN(n18789) );
  INV_X1 U14601 ( .A(n11553), .ZN(n11555) );
  XOR2_X1 U14602 ( .A(n11550), .B(n11549), .Z(n11552) );
  OAI21_X1 U14603 ( .B1(n11555), .B2(n11554), .A(n18779), .ZN(n18775) );
  NOR2_X1 U14604 ( .A1(n19008), .A2(n11556), .ZN(n13296) );
  NAND2_X1 U14605 ( .A1(n13296), .A2(n11557), .ZN(n13308) );
  NAND2_X1 U14606 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18009) );
  NOR2_X1 U14607 ( .A1(n18009), .A2(n11558), .ZN(n17992) );
  NAND2_X1 U14608 ( .A1(n18007), .A2(n17992), .ZN(n13313) );
  INV_X1 U14609 ( .A(n13313), .ZN(n13318) );
  NAND2_X1 U14610 ( .A1(n11422), .A2(n13318), .ZN(n17991) );
  NAND2_X1 U14611 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11591) );
  NOR2_X1 U14612 ( .A1(n17991), .A2(n11591), .ZN(n16524) );
  NOR2_X1 U14613 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16524), .ZN(
        n11559) );
  INV_X1 U14614 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15827) );
  NOR2_X1 U14615 ( .A1(n11591), .A2(n15827), .ZN(n16508) );
  INV_X1 U14616 ( .A(n16508), .ZN(n13312) );
  NOR2_X1 U14617 ( .A1(n17991), .A2(n13312), .ZN(n15821) );
  OR2_X1 U14618 ( .A1(n17885), .A2(n15821), .ZN(n16499) );
  OAI22_X1 U14619 ( .A1(n15831), .A2(n17880), .B1(n11559), .B2(n16499), .ZN(
        n11599) );
  INV_X1 U14620 ( .A(n18981), .ZN(n11560) );
  OAI221_X1 U14621 ( .B1(n18840), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n18966), .A(n11560), .ZN(n18312) );
  INV_X1 U14622 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16971) );
  NAND2_X1 U14623 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17873) );
  NOR3_X1 U14624 ( .A1(n17873), .A2(n16908), .A3(n17849), .ZN(n17794) );
  NAND2_X1 U14625 ( .A1(n17794), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16850) );
  INV_X1 U14626 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17824) );
  NAND2_X1 U14627 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17772) );
  NAND2_X1 U14628 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17737) );
  NAND2_X1 U14629 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17654) );
  INV_X1 U14630 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16650) );
  NAND2_X1 U14631 ( .A1(n18708), .A2(n12925), .ZN(n11593) );
  NAND2_X1 U14632 ( .A1(n18966), .A2(n18954), .ZN(n18956) );
  NOR2_X1 U14633 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18956), .ZN(n19020) );
  INV_X2 U14634 ( .A(n16515), .ZN(n18296) );
  NAND2_X1 U14635 ( .A1(n18296), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n15829) );
  NOR2_X1 U14636 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18840), .ZN(n17693) );
  AOI21_X1 U14637 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n14206)
         );
  NOR2_X1 U14638 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17721), .ZN(
        n12927) );
  NOR2_X1 U14639 ( .A1(n17975), .A2(n9905), .ZN(n16649) );
  INV_X1 U14640 ( .A(n16649), .ZN(n11562) );
  AOI21_X1 U14641 ( .B1(n10032), .B2(n11562), .A(n16498), .ZN(n16681) );
  OAI21_X1 U14642 ( .B1(n12927), .B2(n17828), .A(n16681), .ZN(n11563) );
  OAI211_X1 U14643 ( .C1(n11593), .C2(n9905), .A(n15829), .B(n11563), .ZN(
        n11597) );
  NOR2_X1 U14644 ( .A1(n18086), .A2(n18112), .ZN(n16506) );
  NOR2_X1 U14645 ( .A1(n11572), .A2(n11573), .ZN(n11570) );
  NOR2_X1 U14646 ( .A1(n11570), .A2(n11317), .ZN(n11569) );
  NOR2_X1 U14647 ( .A1(n17483), .A2(n11569), .ZN(n11567) );
  NAND2_X1 U14648 ( .A1(n11567), .A2(n11568), .ZN(n11565) );
  NOR2_X1 U14649 ( .A1(n17476), .A2(n11565), .ZN(n17900) );
  NAND2_X1 U14650 ( .A1(n17900), .A2(n17903), .ZN(n11564) );
  NOR2_X1 U14651 ( .A1(n17471), .A2(n11564), .ZN(n11589) );
  XNOR2_X1 U14652 ( .A(n13310), .B(n11564), .ZN(n11585) );
  XNOR2_X1 U14653 ( .A(n11566), .B(n11565), .ZN(n11581) );
  AND2_X1 U14654 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11581), .ZN(
        n11582) );
  XOR2_X1 U14655 ( .A(n11568), .B(n11567), .Z(n11579) );
  AND2_X1 U14656 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11579), .ZN(
        n11580) );
  INV_X1 U14657 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18251) );
  XNOR2_X1 U14658 ( .A(n17483), .B(n11569), .ZN(n11577) );
  NOR2_X1 U14659 ( .A1(n18251), .A2(n11577), .ZN(n11578) );
  XOR2_X1 U14660 ( .A(n11317), .B(n11570), .Z(n11575) );
  NOR2_X1 U14661 ( .A1(n11575), .A2(n18270), .ZN(n11576) );
  INV_X1 U14662 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18984) );
  NOR2_X1 U14663 ( .A1(n11572), .A2(n18984), .ZN(n11574) );
  NAND3_X1 U14664 ( .A1(n11573), .A2(n11572), .A3(n18984), .ZN(n11571) );
  OAI221_X1 U14665 ( .B1(n11574), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n11573), .C2(n11572), .A(n11571), .ZN(n17958) );
  XNOR2_X1 U14666 ( .A(n18270), .B(n11575), .ZN(n17957) );
  NOR2_X1 U14667 ( .A1(n17958), .A2(n17957), .ZN(n17956) );
  NOR2_X1 U14668 ( .A1(n11576), .A2(n17956), .ZN(n17940) );
  XNOR2_X1 U14669 ( .A(n18251), .B(n11577), .ZN(n17939) );
  NOR2_X1 U14670 ( .A1(n17940), .A2(n17939), .ZN(n17938) );
  NOR2_X1 U14671 ( .A1(n11578), .A2(n17938), .ZN(n17929) );
  XNOR2_X1 U14672 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11579), .ZN(
        n17928) );
  NOR2_X1 U14673 ( .A1(n17929), .A2(n17928), .ZN(n17927) );
  NOR2_X1 U14674 ( .A1(n11580), .A2(n17927), .ZN(n17921) );
  XNOR2_X1 U14675 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11581), .ZN(
        n17920) );
  NOR2_X1 U14676 ( .A1(n17921), .A2(n17920), .ZN(n17919) );
  INV_X1 U14677 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17901) );
  INV_X1 U14678 ( .A(n17900), .ZN(n17898) );
  XOR2_X1 U14679 ( .A(n17903), .B(n17898), .Z(n11583) );
  AOI222_X1 U14680 ( .A1(n17899), .A2(n17901), .B1(n17899), .B2(n11583), .C1(
        n17901), .C2(n11583), .ZN(n11586) );
  NOR2_X1 U14681 ( .A1(n11585), .A2(n11586), .ZN(n17892) );
  NOR2_X1 U14682 ( .A1(n17892), .A2(n18210), .ZN(n11584) );
  NAND2_X1 U14683 ( .A1(n11589), .A2(n11584), .ZN(n11590) );
  INV_X1 U14684 ( .A(n11584), .ZN(n11588) );
  AND2_X1 U14685 ( .A1(n11586), .A2(n11585), .ZN(n17893) );
  AOI21_X1 U14686 ( .B1(n11589), .B2(n11588), .A(n17893), .ZN(n11587) );
  OAI21_X1 U14687 ( .B1(n11589), .B2(n11588), .A(n11587), .ZN(n17879) );
  NAND2_X1 U14688 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17879), .ZN(
        n17878) );
  NAND2_X1 U14689 ( .A1(n16508), .A2(n17985), .ZN(n15823) );
  NAND2_X1 U14690 ( .A1(n17962), .A2(n15823), .ZN(n16500) );
  INV_X1 U14691 ( .A(n11591), .ZN(n13319) );
  NAND2_X1 U14692 ( .A1(n13319), .A2(n17985), .ZN(n16522) );
  NOR2_X1 U14693 ( .A1(n11592), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11595) );
  INV_X1 U14694 ( .A(n17693), .ZN(n17980) );
  OAI211_X1 U14695 ( .C1(n16649), .C2(n17980), .A(n17979), .B(n11593), .ZN(
        n12926) );
  NAND2_X1 U14696 ( .A1(n12926), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11594) );
  OAI21_X1 U14697 ( .B1(n16500), .B2(n11595), .A(n11594), .ZN(n11596) );
  AOI22_X1 U14698 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11604) );
  AND2_X4 U14699 ( .A1(n15766), .A2(n15761), .ZN(n11759) );
  AND2_X4 U14700 ( .A1(n11601), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13278) );
  AOI22_X1 U14701 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11603) );
  AND2_X4 U14702 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15768) );
  INV_X1 U14703 ( .A(n15774), .ZN(n13225) );
  AND2_X4 U14704 ( .A1(n16446), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11643) );
  AND2_X4 U14705 ( .A1(n16446), .A2(n15769), .ZN(n13269) );
  AOI22_X1 U14706 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14707 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14708 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14709 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14710 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11758), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11606) );
  NAND2_X2 U14711 ( .A1(n20071), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19971) );
  NOR2_X1 U14712 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19906) );
  INV_X1 U14713 ( .A(n19906), .ZN(n19028) );
  NAND2_X1 U14714 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20057) );
  NAND2_X1 U14715 ( .A1(n20062), .A2(n20057), .ZN(n13402) );
  INV_X1 U14716 ( .A(n13402), .ZN(n14952) );
  NAND2_X1 U14717 ( .A1(n11820), .A2(n14952), .ZN(n11830) );
  AND2_X2 U14718 ( .A1(n13258), .A2(n11619), .ZN(n13101) );
  AND2_X2 U14719 ( .A1(n13279), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12258) );
  AOI22_X1 U14720 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14721 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11617) );
  AND2_X2 U14722 ( .A1(n13275), .A2(n11619), .ZN(n11767) );
  AND2_X2 U14723 ( .A1(n13275), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12175) );
  AOI22_X1 U14724 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11616) );
  INV_X1 U14725 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11613) );
  INV_X2 U14726 ( .A(n15774), .ZN(n11758) );
  INV_X1 U14727 ( .A(n11783), .ZN(n11612) );
  AND2_X1 U14728 ( .A1(n11758), .A2(n11619), .ZN(n11610) );
  INV_X1 U14729 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11611) );
  OAI22_X1 U14730 ( .A1(n11613), .A2(n11612), .B1(n11992), .B2(n11611), .ZN(
        n11614) );
  INV_X1 U14731 ( .A(n11614), .ZN(n11615) );
  NAND4_X1 U14732 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11625) );
  AND2_X2 U14733 ( .A1(n11748), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13032) );
  AOI22_X1 U14734 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11623) );
  AND2_X2 U14735 ( .A1(n13279), .A2(n11619), .ZN(n11658) );
  AOI22_X1 U14736 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11622) );
  AND2_X2 U14737 ( .A1(n11748), .A2(n11619), .ZN(n11789) );
  AOI22_X1 U14738 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14739 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12080), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11620) );
  NAND4_X1 U14740 ( .A1(n11623), .A2(n11622), .A3(n11621), .A4(n11620), .ZN(
        n11624) );
  MUX2_X1 U14741 ( .A(n20028), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11676) );
  NAND2_X1 U14742 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20036), .ZN(
        n11673) );
  INV_X1 U14743 ( .A(n11673), .ZN(n11626) );
  NAND2_X1 U14744 ( .A1(n11676), .A2(n11626), .ZN(n11675) );
  NAND2_X1 U14745 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20028), .ZN(
        n11627) );
  NAND2_X1 U14746 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20019), .ZN(
        n11668) );
  INV_X1 U14747 ( .A(n11668), .ZN(n11628) );
  NAND2_X1 U14748 ( .A1(n15769), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11669) );
  MUX2_X1 U14749 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n20012), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11665) );
  NAND2_X1 U14750 ( .A1(n20012), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11629) );
  NOR2_X1 U14751 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15906), .ZN(
        n11631) );
  NAND2_X1 U14752 ( .A1(n11687), .A2(n11631), .ZN(n11684) );
  AOI22_X1 U14753 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14754 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14755 ( .A1(n13258), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14756 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11758), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14757 ( .A1(n13258), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14758 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14759 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14760 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13225), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14761 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11758), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14762 ( .A1(n13269), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11641) );
  BUF_X4 U14763 ( .A(n11643), .Z(n13084) );
  AOI22_X1 U14764 ( .A1(n13084), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11759), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14765 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11644) );
  NAND2_X1 U14766 ( .A1(n9871), .A2(n11646), .ZN(n11653) );
  AOI22_X1 U14767 ( .A1(n13084), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14768 ( .A1(n13280), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14769 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11748), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14770 ( .A1(n11651), .A2(n11650), .A3(n11649), .A4(n11648), .ZN(
        n11652) );
  MUX2_X1 U14771 ( .A(n12222), .B(n11684), .S(n12501), .Z(n12402) );
  AOI22_X1 U14772 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14773 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14774 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11655) );
  INV_X1 U14775 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U14776 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11610), .B1(
        n11783), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11654) );
  NAND4_X1 U14777 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11664) );
  AOI22_X1 U14778 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14779 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14780 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14781 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12080), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11659) );
  NAND4_X1 U14782 ( .A1(n11662), .A2(n11661), .A3(n11660), .A4(n11659), .ZN(
        n11663) );
  INV_X1 U14783 ( .A(n11665), .ZN(n11666) );
  XNOR2_X1 U14784 ( .A(n11667), .B(n11666), .ZN(n11683) );
  NAND2_X1 U14785 ( .A1(n12402), .A2(n12400), .ZN(n11766) );
  NAND2_X1 U14786 ( .A1(n11766), .A2(n12501), .ZN(n11691) );
  NAND2_X1 U14787 ( .A1(n20061), .A2(n20060), .ZN(n11672) );
  NAND2_X1 U14788 ( .A1(n11669), .A2(n11668), .ZN(n11670) );
  XNOR2_X1 U14789 ( .A(n11671), .B(n11670), .ZN(n11797) );
  MUX2_X1 U14790 ( .A(n11672), .B(n12501), .S(n11797), .Z(n11682) );
  INV_X4 U14791 ( .A(n12584), .ZN(n12173) );
  INV_X1 U14792 ( .A(n11797), .ZN(n11680) );
  OAI21_X1 U14793 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20036), .A(
        n11673), .ZN(n11700) );
  INV_X1 U14794 ( .A(n11700), .ZN(n11779) );
  INV_X1 U14795 ( .A(n11676), .ZN(n11674) );
  NAND2_X1 U14796 ( .A1(n11674), .A2(n11673), .ZN(n11780) );
  AND2_X1 U14797 ( .A1(n11780), .A2(n11675), .ZN(n11697) );
  OAI211_X1 U14798 ( .C1(n20060), .C2(n11779), .A(n11815), .B(n11697), .ZN(
        n11679) );
  NAND2_X1 U14799 ( .A1(n11676), .A2(n11779), .ZN(n11677) );
  NAND2_X1 U14800 ( .A1(n11863), .A2(n11677), .ZN(n11678) );
  OAI211_X1 U14801 ( .C1(n11846), .C2(n11680), .A(n11679), .B(n11678), .ZN(
        n11681) );
  NAND2_X1 U14802 ( .A1(n11682), .A2(n11681), .ZN(n11685) );
  NAND2_X1 U14803 ( .A1(n11685), .A2(n11695), .ZN(n11690) );
  NAND2_X1 U14804 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15906), .ZN(
        n11686) );
  NAND2_X1 U14805 ( .A1(n11687), .A2(n11686), .ZN(n11689) );
  NAND2_X1 U14806 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16473), .ZN(
        n11688) );
  AOI21_X1 U14807 ( .B1(n11691), .B2(n11690), .A(n11800), .ZN(n11692) );
  MUX2_X1 U14808 ( .A(n16473), .B(n11692), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n11825) );
  OR2_X1 U14809 ( .A1(n16444), .A2(n12173), .ZN(n13416) );
  NAND2_X1 U14810 ( .A1(n11695), .A2(n11797), .ZN(n11699) );
  INV_X1 U14811 ( .A(n11699), .ZN(n11696) );
  OAI21_X1 U14812 ( .B1(n11700), .B2(n11699), .A(n13347), .ZN(n11701) );
  INV_X1 U14813 ( .A(n11701), .ZN(n11704) );
  AND2_X1 U14814 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11702) );
  NAND2_X1 U14815 ( .A1(n19998), .A2(n11702), .ZN(n11703) );
  NAND2_X1 U14816 ( .A1(n11703), .A2(n16473), .ZN(n13409) );
  INV_X1 U14817 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13350) );
  OAI21_X1 U14818 ( .B1(n13032), .B2(n13409), .A(n13350), .ZN(n16486) );
  MUX2_X1 U14819 ( .A(n11704), .B(n16486), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20044) );
  NOR2_X1 U14820 ( .A1(n11706), .A2(n11705), .ZN(n11710) );
  AOI22_X1 U14821 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14822 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14823 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11758), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11707) );
  NAND4_X1 U14824 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(
        n11711) );
  NAND2_X1 U14825 ( .A1(n11711), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11718) );
  AOI22_X1 U14826 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14827 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14828 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11713) );
  NAND4_X1 U14829 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11716) );
  NAND2_X1 U14830 ( .A1(n11716), .A2(n11619), .ZN(n11717) );
  AOI22_X1 U14831 ( .A1(n13084), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U14832 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11748), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14833 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14834 ( .A1(n11758), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9805), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11719) );
  NAND4_X1 U14835 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n11723) );
  AOI22_X1 U14836 ( .A1(n11758), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13275), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14837 ( .A1(n13084), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14838 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14839 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11724) );
  NAND4_X1 U14840 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n11728) );
  NAND2_X1 U14841 ( .A1(n11728), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11729) );
  AOI22_X1 U14842 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14843 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14844 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14845 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11758), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11731) );
  NAND4_X1 U14846 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n11735) );
  AOI22_X1 U14847 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14848 ( .A1(n13258), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14849 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11736) );
  NAND4_X1 U14850 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n11740) );
  NAND2_X1 U14851 ( .A1(n11740), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11741) );
  AOI22_X1 U14852 ( .A1(n11758), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9805), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U14853 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14854 ( .A1(n13084), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U14855 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U14856 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14857 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14858 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13225), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14859 ( .A1(n13258), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14860 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11758), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14861 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14862 ( .A1(n13258), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14863 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14864 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13225), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14865 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14866 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14867 ( .A1(n13084), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11761) );
  NOR2_X2 U14868 ( .A1(n12957), .A2(n11837), .ZN(n11813) );
  NOR2_X1 U14869 ( .A1(n16465), .A2(n12173), .ZN(n11824) );
  INV_X1 U14870 ( .A(n11766), .ZN(n11802) );
  AOI22_X1 U14871 ( .A1(n12258), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13101), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14872 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14873 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14874 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11768) );
  NAND4_X1 U14875 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n11778) );
  AOI22_X1 U14876 ( .A1(n13032), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14877 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14878 ( .A1(n11789), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14879 ( .A1(n12080), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11773) );
  NAND4_X1 U14880 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11777) );
  MUX2_X1 U14881 ( .A(n12027), .B(n11779), .S(n12501), .Z(n12418) );
  NAND2_X1 U14882 ( .A1(n12418), .A2(n11780), .ZN(n11799) );
  AOI22_X1 U14883 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14884 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14885 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11767), .B1(
        n11783), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14886 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12175), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U14887 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11796) );
  AOI22_X1 U14888 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n13032), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14889 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14890 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11789), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14891 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n12080), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11791) );
  NAND4_X1 U14892 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n11795) );
  MUX2_X1 U14893 ( .A(n12003), .B(n11797), .S(n12501), .Z(n12397) );
  INV_X1 U14894 ( .A(n12397), .ZN(n11798) );
  NAND2_X1 U14895 ( .A1(n11799), .A2(n11798), .ZN(n11801) );
  AOI21_X1 U14896 ( .B1(n11802), .B2(n11801), .A(n11800), .ZN(n20042) );
  AND2_X1 U14897 ( .A1(n12173), .A2(n20055), .ZN(n11809) );
  INV_X1 U14898 ( .A(n11809), .ZN(n11803) );
  NOR2_X1 U14899 ( .A1(n16465), .A2(n11803), .ZN(n20040) );
  NAND2_X1 U14900 ( .A1(n20042), .A2(n20040), .ZN(n12511) );
  AND2_X2 U14901 ( .A1(n11837), .A2(n12957), .ZN(n11878) );
  INV_X1 U14902 ( .A(n11878), .ZN(n11804) );
  INV_X1 U14903 ( .A(n11813), .ZN(n11850) );
  NAND3_X1 U14904 ( .A1(n11804), .A2(n19347), .A3(n11850), .ZN(n11835) );
  NAND2_X1 U14905 ( .A1(n12173), .A2(n11851), .ZN(n11833) );
  NAND2_X1 U14906 ( .A1(n11833), .A2(n11815), .ZN(n11805) );
  NAND2_X1 U14907 ( .A1(n11805), .A2(n10326), .ZN(n11806) );
  NAND2_X1 U14908 ( .A1(n11806), .A2(n9948), .ZN(n11807) );
  AND2_X1 U14909 ( .A1(n11835), .A2(n11807), .ZN(n11811) );
  OAI21_X1 U14910 ( .B1(n11878), .B2(n11808), .A(n11852), .ZN(n11810) );
  NAND2_X1 U14911 ( .A1(n11810), .A2(n11809), .ZN(n11845) );
  AND2_X1 U14912 ( .A1(n11811), .A2(n11845), .ZN(n11818) );
  AND2_X2 U14913 ( .A1(n11812), .A2(n11852), .ZN(n11875) );
  NAND2_X1 U14914 ( .A1(n12193), .A2(n11851), .ZN(n11836) );
  NAND2_X1 U14915 ( .A1(n11836), .A2(n9948), .ZN(n11816) );
  NAND2_X1 U14916 ( .A1(n11874), .A2(n11816), .ZN(n11817) );
  NAND2_X1 U14917 ( .A1(n11818), .A2(n11817), .ZN(n11834) );
  AND3_X1 U14918 ( .A1(n11873), .A2(n13347), .A3(n14952), .ZN(n11819) );
  NOR2_X1 U14919 ( .A1(n11834), .A2(n11819), .ZN(n13398) );
  MUX2_X1 U14920 ( .A(n11873), .B(n11820), .S(n12173), .Z(n11821) );
  NAND3_X1 U14921 ( .A1(n11821), .A2(n13347), .A3(n20057), .ZN(n11822) );
  NAND3_X1 U14922 ( .A1(n12511), .A2(n13398), .A3(n11822), .ZN(n11823) );
  AOI21_X1 U14923 ( .B1(n20044), .B2(n11824), .A(n11823), .ZN(n11829) );
  OAI21_X1 U14924 ( .B1(n11825), .B2(n20055), .A(n11851), .ZN(n11826) );
  INV_X1 U14925 ( .A(n11826), .ZN(n11827) );
  NAND2_X1 U14926 ( .A1(n13416), .A2(n11827), .ZN(n11828) );
  OAI211_X1 U14927 ( .C1(n11830), .C2(n13416), .A(n11829), .B(n11828), .ZN(
        n11832) );
  NAND2_X1 U14928 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16478), .ZN(n19894) );
  INV_X1 U14929 ( .A(n19894), .ZN(n11831) );
  INV_X1 U14930 ( .A(n15770), .ZN(n16440) );
  NAND2_X1 U14931 ( .A1(n12502), .A2(n16440), .ZN(n13524) );
  NAND3_X1 U14932 ( .A1(n11836), .A2(n11835), .A3(n11852), .ZN(n11844) );
  NAND2_X1 U14933 ( .A1(n11844), .A2(n11839), .ZN(n11841) );
  INV_X1 U14934 ( .A(n12957), .ZN(n11853) );
  NAND2_X1 U14935 ( .A1(n11841), .A2(n11840), .ZN(n11893) );
  AND2_X1 U14936 ( .A1(n12193), .A2(n12173), .ZN(n11842) );
  NAND2_X1 U14937 ( .A1(n11842), .A2(n11848), .ZN(n11890) );
  NAND2_X1 U14938 ( .A1(n11893), .A2(n11890), .ZN(n11917) );
  NAND2_X1 U14939 ( .A1(n11917), .A2(n13351), .ZN(n11843) );
  NAND2_X1 U14940 ( .A1(n11843), .A2(n11884), .ZN(n11862) );
  INV_X1 U14941 ( .A(n12173), .ZN(n20060) );
  NAND2_X1 U14942 ( .A1(n11844), .A2(n20060), .ZN(n15753) );
  AOI21_X1 U14943 ( .B1(n15753), .B2(n11845), .A(n19341), .ZN(n11860) );
  NAND3_X1 U14944 ( .A1(n11876), .A2(n19341), .A3(n11864), .ZN(n13491) );
  OAI22_X1 U14945 ( .A1(n13351), .A2(n19347), .B1(n11815), .B2(n9948), .ZN(
        n11849) );
  INV_X1 U14946 ( .A(n11849), .ZN(n11858) );
  AND2_X1 U14947 ( .A1(n11850), .A2(n9948), .ZN(n11855) );
  MUX2_X1 U14948 ( .A(n11853), .B(n11852), .S(n11851), .Z(n11854) );
  NAND2_X1 U14949 ( .A1(n12193), .A2(n11839), .ZN(n11880) );
  NAND3_X1 U14950 ( .A1(n11855), .A2(n11854), .A3(n11880), .ZN(n11857) );
  INV_X1 U14951 ( .A(n13412), .ZN(n11856) );
  NAND3_X1 U14952 ( .A1(n11857), .A2(n11856), .A3(n11815), .ZN(n11891) );
  NAND3_X1 U14953 ( .A1(n13491), .A2(n11858), .A3(n11891), .ZN(n11859) );
  NOR2_X1 U14954 ( .A1(n11860), .A2(n11859), .ZN(n11861) );
  AND2_X1 U14955 ( .A1(n11862), .A2(n11861), .ZN(n15752) );
  INV_X1 U14956 ( .A(n11884), .ZN(n11904) );
  NAND3_X1 U14957 ( .A1(n11884), .A2(n11864), .A3(n11863), .ZN(n11865) );
  NAND2_X1 U14958 ( .A1(n15752), .A2(n11865), .ZN(n11866) );
  NAND2_X1 U14959 ( .A1(n12502), .A2(n11866), .ZN(n12163) );
  NAND2_X1 U14960 ( .A1(n13524), .A2(n12163), .ZN(n19305) );
  INV_X1 U14961 ( .A(n19305), .ZN(n15608) );
  INV_X1 U14962 ( .A(n12163), .ZN(n13529) );
  INV_X1 U14963 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15641) );
  NAND2_X1 U14964 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16380) );
  INV_X1 U14965 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15707) );
  NAND2_X1 U14966 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16406) );
  INV_X1 U14967 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12448) );
  NAND2_X1 U14968 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15739) );
  NOR3_X1 U14969 ( .A1(n15738), .A2(n12448), .A3(n15739), .ZN(n12165) );
  INV_X1 U14970 ( .A(n12165), .ZN(n11870) );
  NAND2_X1 U14971 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19304) );
  NAND2_X1 U14972 ( .A1(n13531), .A2(n19304), .ZN(n13525) );
  INV_X1 U14973 ( .A(n19304), .ZN(n11867) );
  NAND2_X1 U14974 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11867), .ZN(
        n13526) );
  NAND2_X1 U14975 ( .A1(n13529), .A2(n13526), .ZN(n13530) );
  INV_X1 U14976 ( .A(n12502), .ZN(n11869) );
  NAND2_X1 U14977 ( .A1(n19533), .A2(n20054), .ZN(n15902) );
  INV_X1 U14978 ( .A(n15902), .ZN(n11868) );
  INV_X2 U14979 ( .A(n19271), .ZN(n19150) );
  NAND2_X1 U14980 ( .A1(n11869), .A2(n19150), .ZN(n13528) );
  OAI211_X1 U14981 ( .C1(n13524), .C2(n13525), .A(n13530), .B(n13528), .ZN(
        n15737) );
  AOI21_X1 U14982 ( .B1(n19305), .B2(n11870), .A(n15737), .ZN(n15718) );
  INV_X1 U14983 ( .A(n15718), .ZN(n16411) );
  AOI21_X1 U14984 ( .B1(n19305), .B2(n16406), .A(n16411), .ZN(n15607) );
  INV_X1 U14985 ( .A(n15607), .ZN(n11871) );
  NOR2_X1 U14986 ( .A1(n15707), .A2(n11871), .ZN(n15705) );
  INV_X1 U14987 ( .A(n15705), .ZN(n16382) );
  NOR2_X1 U14988 ( .A1(n16380), .A2(n16382), .ZN(n15687) );
  NAND2_X1 U14989 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15673) );
  INV_X1 U14990 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15676) );
  NOR2_X1 U14991 ( .A1(n15673), .A2(n15676), .ZN(n12167) );
  AND2_X1 U14992 ( .A1(n15687), .A2(n12167), .ZN(n15628) );
  INV_X1 U14993 ( .A(n15737), .ZN(n11872) );
  NAND2_X1 U14994 ( .A1(n11872), .A2(n15608), .ZN(n16383) );
  NOR2_X1 U14995 ( .A1(n15628), .A2(n15688), .ZN(n15662) );
  NAND2_X1 U14996 ( .A1(n11877), .A2(n10334), .ZN(n11883) );
  NAND2_X1 U14997 ( .A1(n11878), .A2(n12173), .ZN(n11879) );
  NAND2_X1 U14998 ( .A1(n11901), .A2(n11884), .ZN(n15773) );
  NAND2_X1 U14999 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11889) );
  NOR2_X1 U15000 ( .A1(n20061), .A2(n9802), .ZN(n11887) );
  NAND2_X1 U15001 ( .A1(n11925), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11888) );
  NAND2_X1 U15002 ( .A1(n11890), .A2(n11815), .ZN(n11892) );
  NAND3_X1 U15003 ( .A1(n16465), .A2(n9948), .A3(n20060), .ZN(n11895) );
  INV_X1 U15004 ( .A(n11873), .ZN(n11894) );
  INV_X1 U15005 ( .A(n20061), .ZN(n11896) );
  NAND2_X1 U15006 ( .A1(n11931), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11899) );
  NAND2_X1 U15007 ( .A1(n20054), .A2(n16478), .ZN(n20051) );
  INV_X1 U15008 ( .A(n20051), .ZN(n16481) );
  AOI22_X1 U15009 ( .A1(n11897), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16481), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U15010 ( .A1(n11931), .A2(n11900), .ZN(n11909) );
  NAND2_X1 U15011 ( .A1(n11900), .A2(n11863), .ZN(n11903) );
  INV_X1 U15012 ( .A(n15755), .ZN(n11902) );
  NAND2_X1 U15013 ( .A1(n11903), .A2(n11902), .ZN(n11907) );
  NOR2_X1 U15014 ( .A1(n11904), .A2(n20054), .ZN(n11906) );
  NOR2_X1 U15015 ( .A1(n20051), .A2(n20036), .ZN(n11905) );
  AOI21_X1 U15016 ( .B1(n11907), .B2(n11906), .A(n11905), .ZN(n11908) );
  INV_X1 U15017 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12197) );
  INV_X1 U15018 ( .A(n12360), .ZN(n11910) );
  NAND2_X1 U15019 ( .A1(n11910), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11915) );
  NAND2_X1 U15020 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11911) );
  NAND2_X1 U15021 ( .A1(n20051), .A2(n11911), .ZN(n11912) );
  AOI21_X1 U15022 ( .B1(n11925), .B2(P2_REIP_REG_0__SCAN_IN), .A(n11912), .ZN(
        n11914) );
  NAND3_X1 U15023 ( .A1(n11915), .A2(n11914), .A3(n11913), .ZN(n11919) );
  AOI21_X1 U15024 ( .B1(n11917), .B2(n11916), .A(n20054), .ZN(n11918) );
  INV_X1 U15025 ( .A(n11921), .ZN(n11923) );
  NAND2_X1 U15026 ( .A1(n11923), .A2(n11922), .ZN(n11924) );
  INV_X1 U15027 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12396) );
  NAND2_X1 U15028 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11927) );
  NAND2_X1 U15029 ( .A1(n11925), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11926) );
  OAI211_X1 U15030 ( .C1(n12360), .C2(n12396), .A(n11927), .B(n11926), .ZN(
        n11928) );
  INV_X1 U15031 ( .A(n11928), .ZN(n11930) );
  OAI21_X1 U15032 ( .B1(n20019), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16478), 
        .ZN(n11932) );
  INV_X1 U15033 ( .A(n11946), .ZN(n11933) );
  NAND2_X1 U15034 ( .A1(n11947), .A2(n11933), .ZN(n11934) );
  INV_X1 U15035 ( .A(n11947), .ZN(n11935) );
  NAND2_X1 U15036 ( .A1(n11935), .A2(n11946), .ZN(n11936) );
  NAND2_X2 U15037 ( .A1(n11937), .A2(n11936), .ZN(n12341) );
  INV_X4 U15038 ( .A(n11939), .ZN(n12798) );
  INV_X1 U15039 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11942) );
  NAND2_X1 U15040 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U15041 ( .A1(n11925), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11940) );
  OAI211_X1 U15042 ( .C1(n12360), .C2(n11942), .A(n11941), .B(n11940), .ZN(
        n11943) );
  INV_X1 U15043 ( .A(n11943), .ZN(n11944) );
  OAI21_X2 U15044 ( .B1(n12798), .B2(n15738), .A(n11944), .ZN(n12342) );
  NOR2_X1 U15045 ( .A1(n20051), .A2(n20012), .ZN(n11945) );
  INV_X1 U15046 ( .A(n12968), .ZN(n13549) );
  OR2_X2 U15047 ( .A1(n12956), .A2(n13549), .ZN(n11965) );
  INV_X1 U15049 ( .A(n11950), .ZN(n11953) );
  INV_X1 U15050 ( .A(n11951), .ZN(n11952) );
  NAND2_X1 U15051 ( .A1(n11953), .A2(n11952), .ZN(n11955) );
  INV_X1 U15052 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11958) );
  INV_X1 U15053 ( .A(n12974), .ZN(n16418) );
  NAND2_X1 U15054 ( .A1(n16452), .A2(n16418), .ZN(n11975) );
  OAI211_X1 U15055 ( .C1(n19471), .C2(n11958), .A(n11957), .B(n20060), .ZN(
        n11962) );
  INV_X1 U15056 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11960) );
  NAND2_X1 U15057 ( .A1(n12974), .A2(n11959), .ZN(n11984) );
  INV_X1 U15058 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13112) );
  NOR2_X1 U15059 ( .A1(n11962), .A2(n11961), .ZN(n11971) );
  INV_X1 U15060 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13113) );
  INV_X1 U15061 ( .A(n11959), .ZN(n11963) );
  NAND2_X1 U15062 ( .A1(n11963), .A2(n12974), .ZN(n11986) );
  INV_X1 U15063 ( .A(n11965), .ZN(n11964) );
  NAND2_X2 U15064 ( .A1(n11964), .A2(n11956), .ZN(n12059) );
  INV_X1 U15065 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13111) );
  OAI22_X1 U15066 ( .A1(n13113), .A2(n12044), .B1(n12059), .B2(n13111), .ZN(
        n11969) );
  INV_X1 U15067 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13114) );
  OR2_X2 U15068 ( .A1(n11965), .A2(n11986), .ZN(n12054) );
  INV_X1 U15069 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11967) );
  OAI22_X1 U15070 ( .A1(n13114), .A2(n12054), .B1(n12051), .B2(n11967), .ZN(
        n11968) );
  NOR2_X1 U15071 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  NAND2_X1 U15072 ( .A1(n11971), .A2(n11970), .ZN(n12006) );
  INV_X1 U15073 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11974) );
  INV_X1 U15074 ( .A(n11986), .ZN(n11973) );
  INV_X1 U15075 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13122) );
  OAI22_X1 U15076 ( .A1(n11974), .A2(n19588), .B1(n12046), .B2(n13122), .ZN(
        n11978) );
  INV_X1 U15077 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11976) );
  INV_X1 U15078 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13120) );
  OAI22_X1 U15079 ( .A1(n11976), .A2(n12067), .B1(n12047), .B2(n13120), .ZN(
        n11977) );
  NOR2_X1 U15080 ( .A1(n11978), .A2(n11977), .ZN(n11991) );
  INV_X1 U15081 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11982) );
  INV_X1 U15082 ( .A(n11983), .ZN(n11990) );
  OR2_X2 U15083 ( .A1(n11985), .A2(n11984), .ZN(n12065) );
  INV_X1 U15084 ( .A(n12065), .ZN(n11988) );
  INV_X1 U15085 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13123) );
  NAND3_X1 U15087 ( .A1(n11991), .A2(n11990), .A3(n11989), .ZN(n12005) );
  AOI22_X1 U15088 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15089 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15090 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15091 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11993) );
  NAND4_X1 U15092 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n12002) );
  AOI22_X1 U15093 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15094 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15095 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15096 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12080), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11997) );
  NAND4_X1 U15097 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12001) );
  NAND3_X1 U15098 ( .A1(n12173), .A2(n12027), .A3(n12399), .ZN(n12031) );
  NAND2_X1 U15099 ( .A1(n12031), .A2(n12209), .ZN(n12004) );
  INV_X1 U15100 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12007) );
  INV_X1 U15101 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13177) );
  INV_X1 U15102 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13169) );
  INV_X1 U15103 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12008) );
  NOR2_X1 U15104 ( .A1(n12010), .A2(n12009), .ZN(n12024) );
  INV_X1 U15105 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13034) );
  INV_X1 U15106 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13168) );
  OAI22_X1 U15107 ( .A1(n13034), .A2(n19471), .B1(n12061), .B2(n13168), .ZN(
        n12012) );
  INV_X1 U15108 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13170) );
  INV_X1 U15109 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13179) );
  NOR2_X1 U15110 ( .A1(n12012), .A2(n12011), .ZN(n12023) );
  INV_X1 U15111 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12013) );
  INV_X1 U15112 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13178) );
  OAI22_X1 U15113 ( .A1(n12013), .A2(n12065), .B1(n12046), .B2(n13178), .ZN(
        n12015) );
  INV_X1 U15114 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13176) );
  OAI22_X1 U15115 ( .A1(n13035), .A2(n12064), .B1(n12047), .B2(n13176), .ZN(
        n12014) );
  NOR2_X1 U15116 ( .A1(n12015), .A2(n12014), .ZN(n12022) );
  INV_X1 U15117 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13167) );
  INV_X1 U15118 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12016) );
  OAI22_X1 U15119 ( .A1(n13167), .A2(n12059), .B1(n12051), .B2(n12016), .ZN(
        n12020) );
  INV_X1 U15120 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12018) );
  INV_X1 U15121 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12017) );
  OAI22_X1 U15122 ( .A1(n12018), .A2(n12058), .B1(n12050), .B2(n12017), .ZN(
        n12019) );
  NOR2_X1 U15123 ( .A1(n12020), .A2(n12019), .ZN(n12021) );
  INV_X1 U15124 ( .A(n12025), .ZN(n12218) );
  NAND2_X1 U15125 ( .A1(n12218), .A2(n12173), .ZN(n12026) );
  NAND2_X1 U15126 ( .A1(n12173), .A2(n12027), .ZN(n13384) );
  NAND2_X1 U15127 ( .A1(n13384), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13383) );
  INV_X1 U15128 ( .A(n12027), .ZN(n12195) );
  INV_X1 U15129 ( .A(n12399), .ZN(n12028) );
  XNOR2_X1 U15130 ( .A(n12195), .B(n12028), .ZN(n12029) );
  OR2_X1 U15131 ( .A1(n13383), .A2(n12029), .ZN(n12030) );
  XOR2_X1 U15132 ( .A(n12029), .B(n13383), .Z(n13390) );
  NAND2_X1 U15133 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13390), .ZN(
        n13389) );
  NAND2_X1 U15134 ( .A1(n12030), .A2(n13389), .ZN(n12032) );
  XNOR2_X1 U15135 ( .A(n13531), .B(n12032), .ZN(n13440) );
  XNOR2_X1 U15136 ( .A(n12031), .B(n12209), .ZN(n13439) );
  NAND2_X1 U15137 ( .A1(n13440), .A2(n13439), .ZN(n12034) );
  NAND2_X1 U15138 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12032), .ZN(
        n12033) );
  NAND2_X1 U15139 ( .A1(n12034), .A2(n12033), .ZN(n12035) );
  XNOR2_X1 U15140 ( .A(n12035), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14015) );
  NAND2_X1 U15141 ( .A1(n12035), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12036) );
  INV_X1 U15142 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19290) );
  NAND2_X1 U15143 ( .A1(n19274), .A2(n19290), .ZN(n12040) );
  NAND2_X1 U15144 ( .A1(n19276), .A2(n12040), .ZN(n12043) );
  INV_X1 U15145 ( .A(n19274), .ZN(n12041) );
  NAND2_X1 U15146 ( .A1(n12041), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12042) );
  INV_X1 U15147 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13221) );
  INV_X1 U15148 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13230) );
  OAI22_X1 U15149 ( .A1(n13221), .A2(n12044), .B1(n12045), .B2(n13230), .ZN(
        n12049) );
  INV_X1 U15150 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13231) );
  INV_X1 U15151 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13229) );
  OAI22_X1 U15152 ( .A1(n13231), .A2(n12046), .B1(n12047), .B2(n13229), .ZN(
        n12048) );
  NOR2_X1 U15153 ( .A1(n12049), .A2(n12048), .ZN(n12075) );
  INV_X1 U15154 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12053) );
  INV_X1 U15155 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12052) );
  OAI22_X1 U15156 ( .A1(n12053), .A2(n12050), .B1(n12051), .B2(n12052), .ZN(
        n12057) );
  INV_X1 U15157 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13222) );
  INV_X1 U15158 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13232) );
  OAI22_X1 U15159 ( .A1(n13222), .A2(n12054), .B1(n12055), .B2(n13232), .ZN(
        n12056) );
  NOR2_X1 U15160 ( .A1(n12057), .A2(n12056), .ZN(n12074) );
  INV_X1 U15161 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12060) );
  INV_X1 U15162 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13219) );
  OAI22_X1 U15163 ( .A1(n12060), .A2(n12058), .B1(n12059), .B2(n13219), .ZN(
        n12063) );
  INV_X1 U15164 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13058) );
  INV_X1 U15165 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13220) );
  OAI22_X1 U15166 ( .A1(n13058), .A2(n19471), .B1(n12061), .B2(n13220), .ZN(
        n12062) );
  NOR2_X1 U15167 ( .A1(n12063), .A2(n12062), .ZN(n12073) );
  INV_X1 U15168 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13801) );
  INV_X1 U15169 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12066) );
  OAI22_X1 U15170 ( .A1(n13801), .A2(n12064), .B1(n12065), .B2(n12066), .ZN(
        n12071) );
  INV_X1 U15171 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12069) );
  INV_X1 U15172 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12068) );
  OAI22_X1 U15173 ( .A1(n12069), .A2(n19588), .B1(n12067), .B2(n12068), .ZN(
        n12070) );
  NOR2_X1 U15174 ( .A1(n12071), .A2(n12070), .ZN(n12072) );
  NAND4_X1 U15175 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n12072), .ZN(
        n12088) );
  AOI22_X1 U15176 ( .A1(n12258), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13101), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15177 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15178 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15179 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12076) );
  NAND4_X1 U15180 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12086) );
  AOI22_X1 U15181 ( .A1(n13032), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15182 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15183 ( .A1(n11789), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15184 ( .A1(n12080), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U15185 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12085) );
  INV_X1 U15186 ( .A(n12403), .ZN(n12227) );
  NAND2_X1 U15187 ( .A1(n12227), .A2(n12173), .ZN(n12087) );
  INV_X1 U15188 ( .A(n12437), .ZN(n12089) );
  INV_X1 U15189 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15741) );
  INV_X1 U15190 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12094) );
  INV_X1 U15191 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12093) );
  OAI22_X1 U15192 ( .A1(n12094), .A2(n19588), .B1(n12067), .B2(n12093), .ZN(
        n12098) );
  INV_X1 U15193 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12096) );
  INV_X1 U15194 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12095) );
  OAI22_X1 U15195 ( .A1(n12096), .A2(n12064), .B1(n12051), .B2(n12095), .ZN(
        n12097) );
  NOR2_X1 U15196 ( .A1(n12098), .A2(n12097), .ZN(n12115) );
  INV_X1 U15197 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12100) );
  INV_X1 U15198 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12099) );
  OAI22_X1 U15199 ( .A1(n12100), .A2(n12058), .B1(n12050), .B2(n12099), .ZN(
        n12104) );
  INV_X1 U15200 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12102) );
  INV_X1 U15201 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12101) );
  OAI22_X1 U15202 ( .A1(n12102), .A2(n19471), .B1(n12055), .B2(n12101), .ZN(
        n12103) );
  NOR2_X1 U15203 ( .A1(n12104), .A2(n12103), .ZN(n12114) );
  INV_X1 U15204 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13242) );
  INV_X1 U15205 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13254) );
  OAI22_X1 U15206 ( .A1(n13242), .A2(n12044), .B1(n12045), .B2(n13254), .ZN(
        n12108) );
  INV_X1 U15207 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12106) );
  INV_X1 U15208 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12105) );
  OAI22_X1 U15209 ( .A1(n12106), .A2(n12065), .B1(n12046), .B2(n12105), .ZN(
        n12107) );
  NOR2_X1 U15210 ( .A1(n12108), .A2(n12107), .ZN(n12113) );
  INV_X1 U15211 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13241) );
  INV_X1 U15212 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12109) );
  OAI22_X1 U15213 ( .A1(n13241), .A2(n12061), .B1(n12054), .B2(n12109), .ZN(
        n12111) );
  INV_X1 U15214 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13243) );
  INV_X1 U15215 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13250) );
  OAI22_X1 U15216 ( .A1(n13243), .A2(n12059), .B1(n12047), .B2(n13250), .ZN(
        n12110) );
  NOR2_X1 U15217 ( .A1(n12111), .A2(n12110), .ZN(n12112) );
  NAND4_X1 U15218 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(
        n12127) );
  AOI22_X1 U15219 ( .A1(n12258), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13101), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15220 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15221 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15222 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12116) );
  NAND4_X1 U15223 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12125) );
  AOI22_X1 U15224 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15225 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15226 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15227 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12080), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15228 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12124) );
  NAND2_X1 U15229 ( .A1(n12404), .A2(n12173), .ZN(n12126) );
  NAND2_X1 U15230 ( .A1(n15745), .A2(n15748), .ZN(n12131) );
  NAND2_X1 U15231 ( .A1(n12131), .A2(n12130), .ZN(n12132) );
  NAND2_X1 U15232 ( .A1(n12258), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12136) );
  NAND2_X1 U15233 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12135) );
  NAND2_X1 U15234 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12134) );
  NAND2_X1 U15235 ( .A1(n11782), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12133) );
  NAND2_X1 U15236 ( .A1(n13032), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12140) );
  NAND2_X1 U15237 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12139) );
  NAND2_X1 U15238 ( .A1(n11789), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12138) );
  NAND2_X1 U15239 ( .A1(n11772), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12137) );
  NAND2_X1 U15240 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12144) );
  NAND2_X1 U15241 ( .A1(n11790), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12143) );
  NAND2_X1 U15242 ( .A1(n12080), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12142) );
  NAND2_X1 U15243 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12141) );
  NAND2_X1 U15244 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12148) );
  NAND2_X1 U15245 ( .A1(n12175), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12147) );
  NAND2_X1 U15246 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12146) );
  NAND2_X1 U15247 ( .A1(n11610), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12145) );
  NAND4_X1 U15248 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12581) );
  INV_X1 U15249 ( .A(n12581), .ZN(n12153) );
  NAND2_X1 U15250 ( .A1(n12154), .A2(n12153), .ZN(n12155) );
  NAND2_X1 U15251 ( .A1(n12160), .A2(n12155), .ZN(n12156) );
  INV_X1 U15252 ( .A(n12156), .ZN(n12157) );
  XNOR2_X1 U15253 ( .A(n12160), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15464) );
  INV_X1 U15254 ( .A(n12160), .ZN(n12161) );
  NAND2_X1 U15255 ( .A1(n12161), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12162) );
  OR2_X2 U15256 ( .A1(n16316), .A2(n15673), .ZN(n16293) );
  NOR2_X4 U15257 ( .A1(n16293), .A2(n15676), .ZN(n15664) );
  INV_X1 U15258 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15650) );
  OAI21_X1 U15259 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15608), .A(
        n15651), .ZN(n12395) );
  AND2_X1 U15260 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12505) );
  INV_X1 U15261 ( .A(n13525), .ZN(n12164) );
  OAI22_X1 U15262 ( .A1(n12164), .A2(n13524), .B1(n12163), .B2(n13526), .ZN(
        n15726) );
  NAND2_X1 U15263 ( .A1(n15726), .A2(n12165), .ZN(n16408) );
  NOR2_X1 U15264 ( .A1(n16380), .A2(n15707), .ZN(n12166) );
  NAND2_X1 U15265 ( .A1(n16393), .A2(n12166), .ZN(n16369) );
  INV_X1 U15266 ( .A(n12167), .ZN(n12168) );
  NOR2_X1 U15267 ( .A1(n16369), .A2(n12168), .ZN(n15640) );
  AOI22_X1 U15268 ( .A1(n15459), .A2(n16413), .B1(n12505), .B2(n15640), .ZN(
        n12393) );
  INV_X1 U15269 ( .A(n12170), .ZN(n12171) );
  AND2_X1 U15270 ( .A1(n15755), .A2(n12171), .ZN(n13291) );
  INV_X1 U15271 ( .A(n13291), .ZN(n16443) );
  OAI21_X1 U15272 ( .B1(n12173), .B2(n9816), .A(n16443), .ZN(n12172) );
  AOI22_X1 U15273 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15274 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15275 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15276 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12176) );
  NAND4_X1 U15277 ( .A1(n12179), .A2(n12178), .A3(n12177), .A4(n12176), .ZN(
        n12185) );
  AOI22_X1 U15278 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15279 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15280 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15281 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12080), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12180) );
  NAND4_X1 U15282 ( .A1(n12183), .A2(n12182), .A3(n12181), .A4(n12180), .ZN(
        n12184) );
  NOR2_X1 U15283 ( .A1(n12185), .A2(n12184), .ZN(n13835) );
  INV_X1 U15284 ( .A(n13835), .ZN(n12186) );
  NAND2_X1 U15285 ( .A1(n12298), .A2(n12186), .ZN(n12191) );
  NOR2_X4 U15286 ( .A1(n9802), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12835) );
  NOR2_X1 U15287 ( .A1(n11852), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12187) );
  INV_X2 U15288 ( .A(n12811), .ZN(n12821) );
  AOI22_X1 U15289 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12190) );
  INV_X4 U15290 ( .A(n12810), .ZN(n12822) );
  NAND2_X1 U15291 ( .A1(n12822), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12189) );
  AND2_X1 U15292 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12192) );
  NOR2_X1 U15293 ( .A1(n12187), .A2(n12192), .ZN(n12194) );
  INV_X1 U15294 ( .A(n12193), .ZN(n13504) );
  NAND2_X1 U15295 ( .A1(n12822), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12200) );
  INV_X1 U15296 ( .A(n11852), .ZN(n19369) );
  NAND2_X1 U15297 ( .A1(n19369), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12196) );
  OAI211_X1 U15298 ( .C1(n12173), .C2(n12197), .A(n12196), .B(n12958), .ZN(
        n12198) );
  INV_X1 U15299 ( .A(n12198), .ZN(n12199) );
  NAND2_X1 U15300 ( .A1(n12200), .A2(n12199), .ZN(n13516) );
  AOI22_X1 U15301 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n12187), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12202) );
  NAND2_X1 U15302 ( .A1(n12822), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12201) );
  AND2_X1 U15303 ( .A1(n12202), .A2(n12201), .ZN(n12205) );
  XNOR2_X1 U15304 ( .A(n13518), .B(n12205), .ZN(n13642) );
  NAND2_X1 U15305 ( .A1(n12193), .A2(n11852), .ZN(n13498) );
  MUX2_X1 U15306 ( .A(n13498), .B(n20028), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12204) );
  NAND2_X1 U15307 ( .A1(n12298), .A2(n12399), .ZN(n12203) );
  NAND2_X1 U15308 ( .A1(n12204), .A2(n12203), .ZN(n13641) );
  NAND2_X1 U15309 ( .A1(n12205), .A2(n13518), .ZN(n12206) );
  NAND2_X1 U15310 ( .A1(n13644), .A2(n12206), .ZN(n12213) );
  NAND2_X1 U15311 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12207) );
  OAI211_X1 U15312 ( .C1(n12326), .C2(n12209), .A(n12208), .B(n12207), .ZN(
        n12212) );
  XNOR2_X1 U15313 ( .A(n12213), .B(n12212), .ZN(n13533) );
  AOI22_X1 U15314 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12211) );
  NAND2_X1 U15315 ( .A1(n12822), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12210) );
  AND2_X1 U15316 ( .A1(n12211), .A2(n12210), .ZN(n13534) );
  INV_X1 U15317 ( .A(n12212), .ZN(n12214) );
  NAND2_X1 U15318 ( .A1(n12214), .A2(n12213), .ZN(n12215) );
  AOI22_X1 U15319 ( .A1(n12822), .A2(P2_REIP_REG_3__SCAN_IN), .B1(n12835), 
        .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12221) );
  NOR2_X1 U15320 ( .A1(n20012), .A2(n12958), .ZN(n12216) );
  AOI21_X1 U15321 ( .B1(n12821), .B2(P2_EAX_REG_3__SCAN_IN), .A(n12216), .ZN(
        n12217) );
  OAI21_X1 U15322 ( .B1(n12326), .B2(n12218), .A(n12217), .ZN(n12219) );
  INV_X1 U15323 ( .A(n12219), .ZN(n12220) );
  AOI22_X1 U15324 ( .A1(n12298), .A2(n12222), .B1(n12822), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15325 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12223) );
  NAND2_X1 U15326 ( .A1(n12224), .A2(n12223), .ZN(n13979) );
  INV_X1 U15327 ( .A(n13976), .ZN(n12228) );
  AOI22_X1 U15328 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U15329 ( .A1(n12822), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12225) );
  OAI211_X1 U15330 ( .C1(n12227), .C2(n12326), .A(n12226), .B(n12225), .ZN(
        n13974) );
  NAND2_X1 U15331 ( .A1(n12228), .A2(n13974), .ZN(n13978) );
  INV_X1 U15332 ( .A(n12404), .ZN(n12229) );
  NAND2_X1 U15333 ( .A1(n12298), .A2(n12229), .ZN(n12230) );
  AOI22_X1 U15334 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12232) );
  NAND2_X1 U15335 ( .A1(n12822), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12231) );
  NAND2_X1 U15336 ( .A1(n12232), .A2(n12231), .ZN(n13500) );
  AND2_X2 U15337 ( .A1(n13501), .A2(n13500), .ZN(n13503) );
  NOR2_X1 U15338 ( .A1(n13503), .A2(n12233), .ZN(n13554) );
  AOI222_X1 U15339 ( .A1(n12822), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n12835), 
        .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n12821), .C2(
        P2_EAX_REG_7__SCAN_IN), .ZN(n13553) );
  AOI22_X1 U15340 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13101), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15341 ( .A1(n11789), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15342 ( .A1(n11772), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15343 ( .A1(n13032), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12080), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12234) );
  NAND4_X1 U15344 ( .A1(n12237), .A2(n12236), .A3(n12235), .A4(n12234), .ZN(
        n12243) );
  AOI22_X1 U15345 ( .A1(n12258), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15346 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15347 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15348 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12238) );
  NAND4_X1 U15349 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n12242) );
  AOI22_X1 U15350 ( .A1(n12298), .A2(n13843), .B1(n12822), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15351 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U15352 ( .A1(n12245), .A2(n12244), .ZN(n13557) );
  AOI22_X1 U15353 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11658), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15354 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11789), .B1(
        n13032), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15355 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13033), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15356 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11772), .B1(
        n12080), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12246) );
  NAND4_X1 U15357 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12255) );
  AOI22_X1 U15358 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15359 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11783), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15360 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11610), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15361 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12250) );
  NAND4_X1 U15362 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12254) );
  AOI22_X1 U15363 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12257) );
  NAND2_X1 U15364 ( .A1(n12822), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12256) );
  OAI211_X1 U15365 ( .C1(n12996), .C2(n12326), .A(n12257), .B(n12256), .ZN(
        n13660) );
  INV_X1 U15366 ( .A(n13101), .ZN(n12285) );
  INV_X1 U15367 ( .A(n12258), .ZN(n12286) );
  OAI22_X1 U15368 ( .A1(n13167), .A2(n12285), .B1(n12286), .B2(n13177), .ZN(
        n12259) );
  INV_X1 U15369 ( .A(n12259), .ZN(n12263) );
  AOI22_X1 U15370 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15371 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15372 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12260) );
  NAND4_X1 U15373 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12269) );
  AOI22_X1 U15374 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15375 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15376 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15377 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12080), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12264) );
  NAND4_X1 U15378 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12268) );
  NAND2_X1 U15379 ( .A1(n12298), .A2(n14004), .ZN(n12272) );
  AOI22_X1 U15380 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12271) );
  NAND2_X1 U15381 ( .A1(n12822), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12270) );
  NOR2_X2 U15382 ( .A1(n15056), .A2(n15057), .ZN(n15055) );
  AOI22_X1 U15383 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15384 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15385 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15386 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12273) );
  NAND4_X1 U15387 ( .A1(n12276), .A2(n12275), .A3(n12274), .A4(n12273), .ZN(
        n12282) );
  AOI22_X1 U15388 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11789), .B1(
        n13032), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15389 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15390 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12080), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15391 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11772), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12277) );
  NAND4_X1 U15392 ( .A1(n12280), .A2(n12279), .A3(n12278), .A4(n12277), .ZN(
        n12281) );
  AOI22_X1 U15393 ( .A1(n12298), .A2(n14003), .B1(n12822), .B2(
        P2_REIP_REG_12__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15394 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12283) );
  NAND2_X1 U15395 ( .A1(n12284), .A2(n12283), .ZN(n13849) );
  NAND2_X1 U15396 ( .A1(n15055), .A2(n13849), .ZN(n13848) );
  OAI22_X1 U15397 ( .A1(n12286), .A2(n13230), .B1(n12285), .B2(n13219), .ZN(
        n12287) );
  INV_X1 U15398 ( .A(n12287), .ZN(n12291) );
  AOI22_X1 U15399 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15400 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15401 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12288) );
  NAND4_X1 U15402 ( .A1(n12291), .A2(n12290), .A3(n12289), .A4(n12288), .ZN(
        n12297) );
  AOI22_X1 U15403 ( .A1(n13032), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15404 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15405 ( .A1(n11789), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15406 ( .A1(n12080), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12292) );
  NAND4_X1 U15407 ( .A1(n12295), .A2(n12294), .A3(n12293), .A4(n12292), .ZN(
        n12296) );
  AOI22_X1 U15408 ( .A1(n12298), .A2(n14086), .B1(n12822), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U15409 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12299) );
  NOR2_X2 U15410 ( .A1(n13848), .A2(n15037), .ZN(n15678) );
  AOI22_X1 U15411 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15412 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15413 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15414 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12301) );
  NAND4_X1 U15415 ( .A1(n12304), .A2(n12303), .A3(n12302), .A4(n12301), .ZN(
        n12310) );
  AOI22_X1 U15416 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13033), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15417 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15418 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11789), .B1(
        n13032), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15419 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11772), .B1(
        n12080), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12305) );
  NAND4_X1 U15420 ( .A1(n12308), .A2(n12307), .A3(n12306), .A4(n12305), .ZN(
        n12309) );
  INV_X1 U15421 ( .A(n14088), .ZN(n12313) );
  AOI22_X1 U15422 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U15423 ( .A1(n12822), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12311) );
  OAI211_X1 U15424 ( .C1(n12313), .C2(n12326), .A(n12312), .B(n12311), .ZN(
        n15679) );
  NAND2_X1 U15425 ( .A1(n15678), .A2(n15679), .ZN(n15680) );
  AOI22_X1 U15426 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15427 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15428 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15429 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12314) );
  NAND4_X1 U15430 ( .A1(n12317), .A2(n12316), .A3(n12315), .A4(n12314), .ZN(
        n12323) );
  AOI22_X1 U15431 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15432 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15433 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15434 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12080), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12318) );
  NAND4_X1 U15435 ( .A1(n12321), .A2(n12320), .A3(n12319), .A4(n12318), .ZN(
        n12322) );
  NOR2_X1 U15436 ( .A1(n12323), .A2(n12322), .ZN(n15230) );
  AOI22_X1 U15437 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U15438 ( .A1(n12822), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12324) );
  OAI211_X1 U15439 ( .C1(n15230), .C2(n12326), .A(n12325), .B(n12324), .ZN(
        n14124) );
  INV_X1 U15440 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19942) );
  NOR2_X1 U15441 ( .A1(n12810), .A2(n19942), .ZN(n12328) );
  INV_X1 U15442 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13427) );
  OAI22_X1 U15443 ( .A1(n12813), .A2(n15650), .B1(n12811), .B2(n13427), .ZN(
        n12327) );
  OR2_X1 U15444 ( .A1(n12328), .A2(n12327), .ZN(n14125) );
  AOI22_X1 U15445 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12331) );
  NAND2_X1 U15446 ( .A1(n12822), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12330) );
  AND2_X1 U15447 ( .A1(n14129), .A2(n12332), .ZN(n12333) );
  NOR2_X1 U15448 ( .A1(n12803), .A2(n12333), .ZN(n19080) );
  AND2_X1 U15449 ( .A1(n12334), .A2(n12502), .ZN(n16412) );
  OR2_X1 U15450 ( .A1(n12798), .A2(n15641), .ZN(n12340) );
  INV_X1 U15451 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12337) );
  NAND2_X1 U15452 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U15453 ( .A1(n11925), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12335) );
  OAI211_X1 U15454 ( .C1(n12793), .C2(n12337), .A(n12336), .B(n12335), .ZN(
        n12338) );
  INV_X1 U15455 ( .A(n12338), .ZN(n12339) );
  NAND2_X1 U15456 ( .A1(n12340), .A2(n12339), .ZN(n15231) );
  INV_X1 U15457 ( .A(n12342), .ZN(n12344) );
  AOI22_X1 U15458 ( .A1(n11925), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12347) );
  NAND2_X1 U15459 ( .A1(n12795), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12346) );
  OAI211_X1 U15460 ( .C1(n12798), .C2(n19290), .A(n12347), .B(n12346), .ZN(
        n12348) );
  INV_X1 U15461 ( .A(n12348), .ZN(n13784) );
  INV_X1 U15462 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n15102) );
  OR2_X1 U15463 ( .A1(n12798), .A2(n15741), .ZN(n12350) );
  AOI22_X1 U15464 ( .A1(n11925), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12349) );
  OAI211_X1 U15465 ( .C1(n12793), .C2(n15102), .A(n12350), .B(n12349), .ZN(
        n13798) );
  OR2_X1 U15466 ( .A1(n12798), .A2(n12448), .ZN(n12355) );
  INV_X1 U15467 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13809) );
  NAND2_X1 U15468 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12352) );
  NAND2_X1 U15469 ( .A1(n11925), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12351) );
  OAI211_X1 U15470 ( .C1(n12793), .C2(n13809), .A(n12352), .B(n12351), .ZN(
        n12353) );
  INV_X1 U15471 ( .A(n12353), .ZN(n12354) );
  INV_X1 U15472 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U15473 ( .A1(n11925), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12357) );
  NAND2_X1 U15474 ( .A1(n12795), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n12356) );
  OAI211_X1 U15475 ( .C1(n12798), .C2(n15719), .A(n12357), .B(n12356), .ZN(
        n13831) );
  INV_X1 U15476 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12458) );
  OR2_X1 U15477 ( .A1(n12798), .A2(n12458), .ZN(n12363) );
  INV_X1 U15478 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n19133) );
  NAND2_X1 U15479 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12359) );
  NAND2_X1 U15480 ( .A1(n11925), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12358) );
  OAI211_X1 U15481 ( .C1(n12360), .C2(n19133), .A(n12359), .B(n12358), .ZN(
        n12361) );
  INV_X1 U15482 ( .A(n12361), .ZN(n12362) );
  INV_X1 U15483 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12366) );
  OR2_X1 U15484 ( .A1(n12798), .A2(n15707), .ZN(n12365) );
  AOI22_X1 U15485 ( .A1(n11925), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12364) );
  OAI211_X1 U15486 ( .C1(n12366), .C2(n12793), .A(n12365), .B(n12364), .ZN(
        n13836) );
  INV_X1 U15487 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16396) );
  AOI22_X1 U15488 ( .A1(n11925), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12368) );
  NAND2_X1 U15489 ( .A1(n12795), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12367) );
  OAI211_X1 U15490 ( .C1(n12798), .C2(n16396), .A(n12368), .B(n12367), .ZN(
        n12369) );
  INV_X1 U15491 ( .A(n12369), .ZN(n13911) );
  INV_X1 U15492 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16384) );
  OR2_X1 U15493 ( .A1(n12798), .A2(n16384), .ZN(n12375) );
  INV_X1 U15494 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12372) );
  NAND2_X1 U15495 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12371) );
  NAND2_X1 U15496 ( .A1(n11925), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12370) );
  OAI211_X1 U15497 ( .C1(n12793), .C2(n12372), .A(n12371), .B(n12370), .ZN(
        n12373) );
  INV_X1 U15498 ( .A(n12373), .ZN(n12374) );
  NAND2_X1 U15499 ( .A1(n12375), .A2(n12374), .ZN(n13896) );
  INV_X1 U15500 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n19122) );
  INV_X1 U15501 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16368) );
  OR2_X1 U15502 ( .A1(n12798), .A2(n16368), .ZN(n12377) );
  AOI22_X1 U15503 ( .A1(n11925), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n12376) );
  OAI211_X1 U15504 ( .C1(n19122), .C2(n12793), .A(n12377), .B(n12376), .ZN(
        n13999) );
  INV_X1 U15505 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n15040) );
  INV_X1 U15506 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16367) );
  OR2_X1 U15507 ( .A1(n12798), .A2(n16367), .ZN(n12379) );
  AOI22_X1 U15508 ( .A1(n11925), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n12378) );
  OAI211_X1 U15509 ( .C1(n15040), .C2(n12793), .A(n12379), .B(n12378), .ZN(
        n14042) );
  AOI22_X1 U15510 ( .A1(n11925), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12381) );
  NAND2_X1 U15511 ( .A1(n12795), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12380) );
  OAI211_X1 U15512 ( .C1(n12798), .C2(n15676), .A(n12381), .B(n12380), .ZN(
        n12382) );
  INV_X1 U15513 ( .A(n12382), .ZN(n14092) );
  INV_X1 U15514 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12409) );
  OR2_X1 U15515 ( .A1(n12798), .A2(n15650), .ZN(n12384) );
  AOI22_X1 U15516 ( .A1(n11925), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n12383) );
  OAI211_X1 U15517 ( .C1(n12793), .C2(n12409), .A(n12384), .B(n12383), .ZN(
        n15227) );
  INV_X1 U15518 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12387) );
  NAND2_X1 U15519 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12386) );
  NAND2_X1 U15520 ( .A1(n11925), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12385) );
  OAI211_X1 U15521 ( .C1(n12793), .C2(n12387), .A(n12386), .B(n12385), .ZN(
        n12388) );
  AOI21_X1 U15522 ( .B1(n12621), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12388), .ZN(n12389) );
  AND2_X1 U15523 ( .A1(n15226), .A2(n12389), .ZN(n12390) );
  OR2_X1 U15524 ( .A1(n15218), .A2(n12390), .ZN(n15446) );
  INV_X1 U15525 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19944) );
  OAI22_X1 U15526 ( .A1(n19308), .A2(n15446), .B1(n19944), .B2(n19150), .ZN(
        n12391) );
  AOI21_X1 U15527 ( .B1(n16387), .B2(n19080), .A(n12391), .ZN(n12392) );
  OAI21_X1 U15528 ( .B1(n12393), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12392), .ZN(n12394) );
  AOI21_X1 U15529 ( .B1(n12395), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12394), .ZN(n12504) );
  MUX2_X1 U15530 ( .A(n12397), .B(n12396), .S(n12785), .Z(n12423) );
  NOR2_X1 U15531 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n12398) );
  MUX2_X1 U15532 ( .A(n12399), .B(n12398), .S(n12785), .Z(n12424) );
  NAND2_X1 U15533 ( .A1(n12423), .A2(n12424), .ZN(n12422) );
  INV_X1 U15534 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12401) );
  MUX2_X1 U15535 ( .A(n12402), .B(n12401), .S(n12785), .Z(n12430) );
  MUX2_X1 U15536 ( .A(n12403), .B(n15102), .S(n12785), .Z(n12438) );
  MUX2_X1 U15537 ( .A(n12404), .B(P2_EBX_REG_6__SCAN_IN), .S(n12785), .Z(
        n12444) );
  INV_X1 U15538 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12405) );
  MUX2_X1 U15539 ( .A(n12581), .B(n12405), .S(n12785), .Z(n12454) );
  NAND2_X1 U15540 ( .A1(n12566), .A2(n12406), .ZN(n12463) );
  INV_X1 U15541 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13914) );
  NAND2_X1 U15542 ( .A1(n12468), .A2(n12372), .ZN(n12477) );
  NAND2_X1 U15543 ( .A1(n12566), .A2(n12477), .ZN(n12469) );
  NAND2_X1 U15544 ( .A1(n12785), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12407) );
  INV_X1 U15545 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14095) );
  NAND2_X1 U15546 ( .A1(n14095), .A2(n12337), .ZN(n12408) );
  OAI211_X1 U15547 ( .C1(n9859), .C2(P2_EBX_REG_16__SCAN_IN), .A(
        P2_EBX_REG_17__SCAN_IN), .B(n12785), .ZN(n12412) );
  NAND2_X1 U15548 ( .A1(n12409), .A2(n12387), .ZN(n12410) );
  NAND2_X1 U15549 ( .A1(n12785), .A2(n12410), .ZN(n12411) );
  INV_X1 U15550 ( .A(n12517), .ZN(n12525) );
  NAND2_X1 U15551 ( .A1(n12412), .A2(n12525), .ZN(n19077) );
  OR2_X1 U15552 ( .A1(n19077), .A2(n12153), .ZN(n12413) );
  INV_X1 U15553 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15450) );
  NAND2_X1 U15554 ( .A1(n12413), .A2(n15450), .ZN(n15395) );
  OR3_X1 U15555 ( .A1(n19077), .A2(n12153), .A3(n15450), .ZN(n12540) );
  NAND2_X1 U15556 ( .A1(n15395), .A2(n12540), .ZN(n15396) );
  INV_X1 U15557 ( .A(n12415), .ZN(n12432) );
  NAND2_X1 U15558 ( .A1(n12422), .A2(n12416), .ZN(n12417) );
  NAND2_X1 U15559 ( .A1(n12432), .A2(n12417), .ZN(n15114) );
  NAND2_X1 U15560 ( .A1(n12427), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14011) );
  INV_X1 U15561 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13552) );
  MUX2_X1 U15562 ( .A(n12418), .B(P2_EBX_REG_0__SCAN_IN), .S(n12785), .Z(
        n19177) );
  NAND2_X1 U15563 ( .A1(n19177), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13392) );
  INV_X1 U15564 ( .A(n12424), .ZN(n12420) );
  INV_X1 U15565 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n15139) );
  NAND3_X1 U15566 ( .A1(n12785), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U15567 ( .A1(n12420), .A2(n12419), .ZN(n15135) );
  NOR2_X1 U15568 ( .A1(n13392), .A2(n15135), .ZN(n12421) );
  NAND2_X1 U15569 ( .A1(n13392), .A2(n15135), .ZN(n13391) );
  OAI21_X1 U15570 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12421), .A(
        n13391), .ZN(n13443) );
  OAI21_X1 U15571 ( .B1(n12424), .B2(n12423), .A(n12422), .ZN(n15125) );
  XNOR2_X1 U15572 ( .A(n15125), .B(n13531), .ZN(n13442) );
  OR2_X1 U15573 ( .A1(n13443), .A2(n13442), .ZN(n13541) );
  INV_X1 U15574 ( .A(n15125), .ZN(n12425) );
  NAND2_X1 U15575 ( .A1(n12425), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12426) );
  AND2_X1 U15576 ( .A1(n13541), .A2(n12426), .ZN(n14013) );
  NAND2_X1 U15577 ( .A1(n14011), .A2(n14013), .ZN(n12429) );
  INV_X1 U15578 ( .A(n12427), .ZN(n12428) );
  NAND2_X1 U15579 ( .A1(n12428), .A2(n15738), .ZN(n14012) );
  INV_X1 U15580 ( .A(n12439), .ZN(n12434) );
  INV_X1 U15581 ( .A(n12430), .ZN(n12431) );
  NAND2_X1 U15582 ( .A1(n12432), .A2(n12431), .ZN(n12433) );
  NAND2_X1 U15583 ( .A1(n12434), .A2(n12433), .ZN(n19164) );
  XNOR2_X1 U15584 ( .A(n19164), .B(n19290), .ZN(n19272) );
  INV_X1 U15585 ( .A(n19164), .ZN(n12435) );
  NAND2_X1 U15586 ( .A1(n12435), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12436) );
  NAND2_X1 U15587 ( .A1(n12437), .A2(n12153), .ZN(n12440) );
  OAI21_X1 U15588 ( .B1(n12439), .B2(n12438), .A(n12445), .ZN(n15103) );
  NAND2_X1 U15589 ( .A1(n12440), .A2(n15103), .ZN(n12441) );
  XNOR2_X1 U15590 ( .A(n12441), .B(n15741), .ZN(n15734) );
  NAND2_X1 U15591 ( .A1(n15735), .A2(n15734), .ZN(n12443) );
  NAND2_X1 U15592 ( .A1(n12441), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12442) );
  AND2_X1 U15593 ( .A1(n12445), .A2(n12444), .ZN(n12446) );
  OR2_X1 U15594 ( .A1(n12446), .A2(n12456), .ZN(n19152) );
  NAND2_X1 U15595 ( .A1(n12449), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12450) );
  AND2_X1 U15596 ( .A1(n12785), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12452) );
  XNOR2_X1 U15597 ( .A(n12453), .B(n12452), .ZN(n19135) );
  OR3_X1 U15598 ( .A1(n19135), .A2(n12153), .A3(n12458), .ZN(n15469) );
  INV_X1 U15599 ( .A(n12454), .ZN(n12455) );
  XNOR2_X1 U15600 ( .A(n12456), .B(n12455), .ZN(n15090) );
  NAND2_X1 U15601 ( .A1(n15090), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15715) );
  INV_X1 U15602 ( .A(n19135), .ZN(n12457) );
  NAND2_X1 U15603 ( .A1(n12457), .A2(n12788), .ZN(n12459) );
  NAND2_X1 U15604 ( .A1(n12459), .A2(n12458), .ZN(n15470) );
  INV_X1 U15605 ( .A(n15090), .ZN(n12460) );
  NAND2_X1 U15606 ( .A1(n12460), .A2(n15719), .ZN(n15714) );
  AND2_X1 U15607 ( .A1(n15470), .A2(n15714), .ZN(n12461) );
  AND2_X1 U15608 ( .A1(n12785), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12462) );
  XNOR2_X1 U15609 ( .A(n12463), .B(n12462), .ZN(n15076) );
  NAND2_X1 U15610 ( .A1(n15076), .A2(n12788), .ZN(n12473) );
  AND2_X1 U15611 ( .A1(n12473), .A2(n15707), .ZN(n15702) );
  NAND2_X1 U15612 ( .A1(n12785), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12464) );
  OAI21_X1 U15613 ( .B1(n12465), .B2(n12464), .A(n12566), .ZN(n12466) );
  OR2_X1 U15614 ( .A1(n12468), .A2(n12466), .ZN(n15072) );
  OAI21_X1 U15615 ( .B1(n15072), .B2(n12153), .A(n16396), .ZN(n16327) );
  NAND2_X1 U15616 ( .A1(n12785), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12467) );
  OR2_X1 U15617 ( .A1(n12468), .A2(n12467), .ZN(n12471) );
  INV_X1 U15618 ( .A(n12469), .ZN(n12470) );
  AOI21_X1 U15619 ( .B1(n15052), .B2(n12788), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16313) );
  AND2_X1 U15620 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12472) );
  NAND2_X1 U15621 ( .A1(n15052), .A2(n12472), .ZN(n16311) );
  INV_X1 U15622 ( .A(n15072), .ZN(n12475) );
  AND2_X1 U15623 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12474) );
  NAND2_X1 U15624 ( .A1(n12475), .A2(n12474), .ZN(n16326) );
  AND3_X1 U15625 ( .A1(n16311), .A2(n16309), .A3(n16326), .ZN(n12476) );
  NAND3_X1 U15626 ( .A1(n12785), .A2(n12477), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n12478) );
  NAND2_X1 U15627 ( .A1(n12481), .A2(n12478), .ZN(n19121) );
  NAND2_X1 U15628 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12479) );
  NOR2_X1 U15629 ( .A1(n19121), .A2(n12479), .ZN(n15693) );
  OR2_X1 U15630 ( .A1(n19121), .A2(n12153), .ZN(n12480) );
  NAND2_X1 U15631 ( .A1(n12480), .A2(n16368), .ZN(n12523) );
  INV_X1 U15632 ( .A(n12523), .ZN(n15694) );
  XNOR2_X1 U15633 ( .A(n12481), .B(n9907), .ZN(n15045) );
  NAND2_X1 U15634 ( .A1(n15045), .A2(n12788), .ZN(n12482) );
  NAND2_X1 U15635 ( .A1(n12482), .A2(n16367), .ZN(n16289) );
  INV_X1 U15636 ( .A(n16289), .ZN(n12483) );
  OR2_X1 U15637 ( .A1(n12482), .A2(n16367), .ZN(n16290) );
  NAND2_X1 U15638 ( .A1(n12485), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12484) );
  MUX2_X1 U15639 ( .A(n12484), .B(n12485), .S(n12174), .Z(n12487) );
  INV_X1 U15640 ( .A(n12485), .ZN(n12486) );
  NAND2_X1 U15641 ( .A1(n12486), .A2(n14095), .ZN(n12492) );
  NAND2_X1 U15642 ( .A1(n12487), .A2(n12492), .ZN(n19112) );
  INV_X1 U15643 ( .A(n19112), .ZN(n12488) );
  NAND2_X1 U15644 ( .A1(n12488), .A2(n12788), .ZN(n12489) );
  NAND2_X1 U15645 ( .A1(n12489), .A2(n15676), .ZN(n15667) );
  INV_X1 U15646 ( .A(n12489), .ZN(n12490) );
  NAND2_X1 U15647 ( .A1(n12490), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15668) );
  AND2_X1 U15648 ( .A1(n12785), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12491) );
  NAND2_X1 U15649 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  NAND2_X1 U15650 ( .A1(n12493), .A2(n9859), .ZN(n19095) );
  NAND2_X1 U15651 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12494) );
  INV_X1 U15652 ( .A(n15652), .ZN(n12496) );
  OR2_X1 U15653 ( .A1(n19095), .A2(n12153), .ZN(n12495) );
  NAND2_X1 U15654 ( .A1(n12495), .A2(n15641), .ZN(n15653) );
  NAND2_X1 U15655 ( .A1(n12785), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12497) );
  MUX2_X1 U15656 ( .A(P2_EBX_REG_16__SCAN_IN), .B(n12497), .S(n9859), .Z(
        n12498) );
  AND2_X1 U15657 ( .A1(n12498), .A2(n12566), .ZN(n19085) );
  NAND2_X1 U15658 ( .A1(n19085), .A2(n12788), .ZN(n12499) );
  XNOR2_X1 U15659 ( .A(n12499), .B(n15650), .ZN(n15456) );
  AND2_X1 U15660 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12500) );
  NAND2_X1 U15661 ( .A1(n19085), .A2(n12500), .ZN(n12541) );
  XOR2_X1 U15662 ( .A(n15396), .B(n9817), .Z(n15454) );
  NOR2_X1 U15663 ( .A1(n16465), .A2(n12501), .ZN(n20039) );
  NAND2_X2 U15664 ( .A1(n12502), .A2(n20039), .ZN(n19314) );
  NAND2_X1 U15665 ( .A1(n12504), .A2(n12503), .ZN(P2_U3029) );
  AND2_X1 U15666 ( .A1(n12505), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15630) );
  AND3_X1 U15667 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12507) );
  NOR2_X1 U15668 ( .A1(n15673), .A2(n16380), .ZN(n12506) );
  NAND3_X1 U15669 ( .A1(n15630), .A2(n12507), .A3(n12506), .ZN(n12838) );
  INV_X1 U15670 ( .A(n12838), .ZN(n15609) );
  INV_X1 U15671 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15604) );
  INV_X1 U15672 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15405) );
  INV_X1 U15673 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12509) );
  INV_X1 U15674 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15555) );
  INV_X1 U15675 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15520) );
  INV_X1 U15676 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15508) );
  NAND2_X1 U15677 ( .A1(n20044), .A2(n20039), .ZN(n12512) );
  NAND2_X1 U15678 ( .A1(n12512), .A2(n12511), .ZN(n12513) );
  INV_X1 U15679 ( .A(n13349), .ZN(n12585) );
  INV_X1 U15680 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n19061) );
  INV_X1 U15681 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12514) );
  NAND2_X1 U15682 ( .A1(n19061), .A2(n12514), .ZN(n12515) );
  NAND2_X1 U15683 ( .A1(n12785), .A2(n12515), .ZN(n12516) );
  INV_X1 U15684 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n12593) );
  NAND2_X1 U15685 ( .A1(n12785), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12549) );
  NAND2_X1 U15686 ( .A1(n12785), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12518) );
  XNOR2_X1 U15687 ( .A(n12556), .B(n12518), .ZN(n16255) );
  NAND2_X1 U15688 ( .A1(n16255), .A2(n12788), .ZN(n12554) );
  INV_X1 U15689 ( .A(n12554), .ZN(n12555) );
  INV_X1 U15690 ( .A(n12519), .ZN(n12522) );
  NAND3_X1 U15691 ( .A1(n12520), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n12785), 
        .ZN(n12521) );
  NAND2_X1 U15692 ( .A1(n12522), .A2(n12521), .ZN(n15017) );
  OAI21_X1 U15693 ( .B1(n15017), .B2(n12153), .A(n15405), .ZN(n15401) );
  AND4_X1 U15694 ( .A1(n15395), .A2(n16289), .A3(n15653), .A4(n12523), .ZN(
        n12534) );
  NAND2_X1 U15695 ( .A1(n12785), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12524) );
  MUX2_X1 U15696 ( .A(n12785), .B(n12524), .S(n12525), .Z(n12526) );
  NAND2_X1 U15697 ( .A1(n12526), .A2(n12528), .ZN(n19062) );
  OR2_X1 U15698 ( .A1(n19062), .A2(n12153), .ZN(n12527) );
  INV_X1 U15699 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15629) );
  NAND2_X1 U15700 ( .A1(n12527), .A2(n15629), .ZN(n15437) );
  NAND3_X1 U15701 ( .A1(n12528), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n12785), 
        .ZN(n12530) );
  INV_X1 U15702 ( .A(n12529), .ZN(n12532) );
  NAND2_X1 U15703 ( .A1(n15018), .A2(n12788), .ZN(n12538) );
  NAND2_X1 U15704 ( .A1(n12538), .A2(n15604), .ZN(n15422) );
  NAND2_X1 U15705 ( .A1(n15437), .A2(n15422), .ZN(n15398) );
  NAND2_X1 U15706 ( .A1(n12785), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12531) );
  XNOR2_X1 U15707 ( .A(n12532), .B(n12531), .ZN(n19051) );
  AOI21_X1 U15708 ( .B1(n19051), .B2(n12788), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15413) );
  NOR2_X1 U15709 ( .A1(n15398), .A2(n15413), .ZN(n12533) );
  NAND4_X1 U15710 ( .A1(n15401), .A2(n12534), .A3(n12533), .A4(n15667), .ZN(
        n12535) );
  INV_X1 U15711 ( .A(n15017), .ZN(n12537) );
  AND2_X1 U15712 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12536) );
  NAND2_X1 U15713 ( .A1(n12537), .A2(n12536), .ZN(n15400) );
  NAND3_X1 U15714 ( .A1(n15400), .A2(n15423), .A3(n15668), .ZN(n12546) );
  NAND2_X1 U15715 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12539) );
  AND2_X1 U15716 ( .A1(n12540), .A2(n15652), .ZN(n12542) );
  NAND4_X1 U15717 ( .A1(n15436), .A2(n12542), .A3(n12541), .A4(n16290), .ZN(
        n12544) );
  AND2_X1 U15718 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12543) );
  OAI21_X2 U15719 ( .B1(n12548), .B2(n10342), .A(n12547), .ZN(n15389) );
  INV_X1 U15720 ( .A(n12549), .ZN(n12550) );
  NAND2_X1 U15721 ( .A1(n12551), .A2(n12550), .ZN(n12552) );
  NAND2_X1 U15722 ( .A1(n12556), .A2(n12552), .ZN(n15833) );
  OR2_X1 U15723 ( .A1(n15833), .A2(n12153), .ZN(n12553) );
  INV_X1 U15724 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12812) );
  NAND2_X1 U15725 ( .A1(n12553), .A2(n12812), .ZN(n15387) );
  AND2_X1 U15726 ( .A1(n12785), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12558) );
  INV_X1 U15727 ( .A(n12566), .ZN(n12557) );
  AOI21_X1 U15728 ( .B1(n12559), .B2(n12558), .A(n12557), .ZN(n12560) );
  AOI21_X1 U15729 ( .B1(n16248), .B2(n12788), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15369) );
  NAND3_X1 U15730 ( .A1(n16248), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n12788), .ZN(n15370) );
  INV_X1 U15731 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15172) );
  NAND2_X1 U15732 ( .A1(n12785), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12561) );
  OAI21_X1 U15733 ( .B1(n12562), .B2(n12561), .A(n12566), .ZN(n12563) );
  INV_X1 U15734 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15546) );
  OAI21_X1 U15735 ( .B1(n15003), .B2(n12153), .A(n15546), .ZN(n15358) );
  NAND2_X1 U15736 ( .A1(n12785), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12564) );
  OR2_X1 U15737 ( .A1(n12565), .A2(n12564), .ZN(n12567) );
  INV_X1 U15738 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U15739 ( .A1(n12612), .A2(n12565), .ZN(n14979) );
  AOI21_X1 U15740 ( .B1(n16236), .B2(n12788), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12570) );
  INV_X1 U15741 ( .A(n16236), .ZN(n12569) );
  NAND2_X1 U15742 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12568) );
  NOR2_X1 U15743 ( .A1(n12569), .A2(n12568), .ZN(n12573) );
  NOR2_X1 U15744 ( .A1(n12570), .A2(n12573), .ZN(n15353) );
  NAND2_X1 U15745 ( .A1(n12785), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12578) );
  INV_X1 U15746 ( .A(n12787), .ZN(n12572) );
  NAND2_X1 U15747 ( .A1(n12785), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12571) );
  XOR2_X1 U15748 ( .A(n12578), .B(n14981), .Z(n16219) );
  NOR2_X1 U15749 ( .A1(n16219), .A2(n12153), .ZN(n15334) );
  INV_X1 U15750 ( .A(n12573), .ZN(n12576) );
  INV_X1 U15751 ( .A(n15003), .ZN(n12575) );
  AND2_X1 U15752 ( .A1(n12581), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12574) );
  NAND2_X1 U15753 ( .A1(n12575), .A2(n12574), .ZN(n15357) );
  NAND2_X1 U15754 ( .A1(n12576), .A2(n15357), .ZN(n15329) );
  INV_X1 U15755 ( .A(n14981), .ZN(n12579) );
  NAND2_X1 U15756 ( .A1(n12785), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12580) );
  XNOR2_X1 U15757 ( .A(n12780), .B(n12580), .ZN(n14909) );
  AOI21_X1 U15758 ( .B1(n14909), .B2(n12788), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12778) );
  INV_X1 U15759 ( .A(n12778), .ZN(n12582) );
  NAND3_X1 U15760 ( .A1(n14909), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12581), .ZN(n12777) );
  NAND2_X1 U15761 ( .A1(n12582), .A2(n12777), .ZN(n12583) );
  XNOR2_X1 U15762 ( .A(n12779), .B(n12583), .ZN(n15504) );
  OR2_X1 U15763 ( .A1(n12798), .A2(n15629), .ZN(n12587) );
  AOI22_X1 U15764 ( .A1(n11925), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12586) );
  OAI211_X1 U15765 ( .C1(n12793), .C2(n19061), .A(n12587), .B(n12586), .ZN(
        n15217) );
  NAND2_X1 U15766 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12589) );
  NAND2_X1 U15767 ( .A1(n11925), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12588) );
  OAI211_X1 U15768 ( .C1(n12793), .C2(n12514), .A(n12589), .B(n12588), .ZN(
        n12590) );
  AOI21_X1 U15769 ( .B1(n12621), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12590), .ZN(n15024) );
  NAND2_X1 U15770 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12592) );
  NAND2_X1 U15771 ( .A1(n11925), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12591) );
  OAI211_X1 U15772 ( .C1(n12793), .C2(n12593), .A(n12592), .B(n12591), .ZN(
        n12594) );
  AOI21_X1 U15773 ( .B1(n12621), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12594), .ZN(n15204) );
  INV_X1 U15774 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12597) );
  NAND2_X1 U15775 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12596) );
  NAND2_X1 U15776 ( .A1(n11925), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12595) );
  OAI211_X1 U15777 ( .C1(n12793), .C2(n12597), .A(n12596), .B(n12595), .ZN(
        n12598) );
  AOI21_X1 U15778 ( .B1(n12621), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12598), .ZN(n15005) );
  INV_X1 U15779 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15832) );
  OR2_X1 U15780 ( .A1(n12798), .A2(n12812), .ZN(n12600) );
  AOI22_X1 U15781 ( .A1(n11925), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12599) );
  OAI211_X1 U15782 ( .C1(n12793), .C2(n15832), .A(n12600), .B(n12599), .ZN(
        n15194) );
  NAND2_X1 U15783 ( .A1(n15195), .A2(n15194), .ZN(n15197) );
  NAND2_X1 U15784 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12602) );
  NAND2_X1 U15785 ( .A1(n11925), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12601) );
  OAI211_X1 U15786 ( .C1(n12793), .C2(n10114), .A(n12602), .B(n12601), .ZN(
        n12603) );
  AOI21_X1 U15787 ( .B1(n12621), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12603), .ZN(n15184) );
  INV_X1 U15788 ( .A(n12604), .ZN(n15183) );
  NAND2_X1 U15789 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12606) );
  NAND2_X1 U15790 ( .A1(n11925), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12605) );
  OAI211_X1 U15791 ( .C1(n12793), .C2(n10113), .A(n12606), .B(n12605), .ZN(
        n12607) );
  AOI21_X1 U15792 ( .B1(n12621), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12607), .ZN(n15178) );
  OR2_X1 U15793 ( .A1(n12798), .A2(n15546), .ZN(n12609) );
  AOI22_X1 U15794 ( .A1(n11925), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12608) );
  OAI211_X1 U15795 ( .C1(n12793), .C2(n15172), .A(n12609), .B(n12608), .ZN(
        n14993) );
  OR2_X1 U15796 ( .A1(n12798), .A2(n10281), .ZN(n12611) );
  AOI22_X1 U15797 ( .A1(n11925), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12610) );
  OAI211_X1 U15798 ( .C1(n12793), .C2(n12612), .A(n12611), .B(n12610), .ZN(
        n15164) );
  INV_X1 U15799 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12615) );
  NAND2_X1 U15800 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12614) );
  NAND2_X1 U15801 ( .A1(n11925), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12613) );
  OAI211_X1 U15802 ( .C1(n12793), .C2(n12615), .A(n12614), .B(n12613), .ZN(
        n12616) );
  AOI21_X1 U15803 ( .B1(n12621), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12616), .ZN(n14976) );
  INV_X1 U15804 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12619) );
  NAND2_X1 U15805 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12618) );
  NAND2_X1 U15806 ( .A1(n11925), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12617) );
  OAI211_X1 U15807 ( .C1(n12793), .C2(n12619), .A(n12618), .B(n12617), .ZN(
        n12620) );
  AOI21_X1 U15808 ( .B1(n12621), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12620), .ZN(n15154) );
  INV_X1 U15809 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12624) );
  INV_X1 U15810 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15492) );
  OR2_X1 U15811 ( .A1(n12798), .A2(n15492), .ZN(n12623) );
  AOI22_X1 U15812 ( .A1(n11925), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12622) );
  OAI211_X1 U15813 ( .C1(n12793), .C2(n12624), .A(n12623), .B(n12622), .ZN(
        n12625) );
  OR2_X1 U15814 ( .A1(n9880), .A2(n12625), .ZN(n12626) );
  NAND2_X1 U15815 ( .A1(n12895), .A2(n12626), .ZN(n15499) );
  INV_X1 U15816 ( .A(n15499), .ZN(n14971) );
  INV_X1 U15817 ( .A(n16490), .ZN(n20056) );
  INV_X1 U15818 ( .A(n16485), .ZN(n12627) );
  OR2_X1 U15819 ( .A1(n20007), .A2(n15785), .ZN(n20020) );
  NAND2_X1 U15820 ( .A1(n20020), .A2(n20054), .ZN(n12629) );
  INV_X1 U15821 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14966) );
  INV_X1 U15822 ( .A(n12978), .ZN(n16479) );
  INV_X1 U15823 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20001) );
  NAND2_X1 U15824 ( .A1(n20001), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12630) );
  NAND2_X1 U15825 ( .A1(n16479), .A2(n12630), .ZN(n13386) );
  INV_X1 U15826 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15429) );
  INV_X1 U15827 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16322) );
  INV_X1 U15828 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16344) );
  NAND2_X1 U15829 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n14021), .ZN(
        n14924) );
  NAND2_X1 U15830 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n14930), .ZN(
        n14933) );
  INV_X1 U15831 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14982) );
  INV_X1 U15832 ( .A(n12947), .ZN(n12633) );
  NAND2_X1 U15833 ( .A1(n14966), .A2(n14913), .ZN(n12632) );
  NAND2_X1 U15834 ( .A1(n12633), .A2(n12632), .ZN(n14949) );
  INV_X1 U15835 ( .A(n14949), .ZN(n12634) );
  NAND2_X1 U15836 ( .A1(n19270), .A2(n12634), .ZN(n12635) );
  NAND2_X1 U15837 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19287), .ZN(n15494) );
  OAI211_X1 U15838 ( .C1(n19285), .C2(n14966), .A(n12635), .B(n15494), .ZN(
        n12636) );
  OAI21_X1 U15839 ( .B1(n15504), .B2(n19278), .A(n12637), .ZN(n12638) );
  INV_X1 U15840 ( .A(n12638), .ZN(n12639) );
  NAND2_X1 U15841 ( .A1(n20274), .A2(n20940), .ZN(n13630) );
  OR2_X1 U15842 ( .A1(n12641), .A2(n13630), .ZN(n13588) );
  NAND3_X1 U15843 ( .A1(n13580), .A2(n10428), .A3(n10470), .ZN(n13693) );
  NAND2_X1 U15844 ( .A1(n13588), .A2(n13693), .ZN(n12642) );
  NAND2_X1 U15845 ( .A1(n12642), .A2(n13678), .ZN(n12653) );
  NOR4_X1 U15846 ( .A1(n12647), .A2(n12646), .A3(n12645), .A4(n12644), .ZN(
        n12648) );
  OR2_X1 U15847 ( .A1(n12649), .A2(n12648), .ZN(n13456) );
  INV_X1 U15848 ( .A(n13456), .ZN(n13449) );
  NAND2_X1 U15849 ( .A1(n13449), .A2(n20940), .ZN(n13673) );
  NOR2_X1 U15850 ( .A1(n12643), .A2(n13673), .ZN(n13595) );
  AND4_X1 U15851 ( .A1(n10461), .A2(n14169), .A3(n14162), .A4(n10574), .ZN(
        n12650) );
  NAND2_X1 U15852 ( .A1(n12650), .A2(n13939), .ZN(n12675) );
  NOR2_X1 U15853 ( .A1(n12675), .A2(n14035), .ZN(n12651) );
  NOR2_X1 U15854 ( .A1(n13595), .A2(n12651), .ZN(n12652) );
  AND2_X1 U15855 ( .A1(n14611), .A2(n14169), .ZN(n12655) );
  NAND2_X1 U15856 ( .A1(n12855), .A2(n12655), .ZN(n12670) );
  NOR4_X1 U15857 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12659) );
  NOR4_X1 U15858 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12658) );
  NOR4_X1 U15859 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12657) );
  NOR4_X1 U15860 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12656) );
  AND4_X1 U15861 ( .A1(n12659), .A2(n12658), .A3(n12657), .A4(n12656), .ZN(
        n12664) );
  NOR4_X1 U15862 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12662) );
  NOR4_X1 U15863 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12661) );
  NOR4_X1 U15864 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12660) );
  INV_X1 U15865 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20855) );
  AND4_X1 U15866 ( .A1(n12662), .A2(n12661), .A3(n12660), .A4(n20855), .ZN(
        n12663) );
  NAND2_X1 U15867 ( .A1(n12664), .A2(n12663), .ZN(n12665) );
  INV_X1 U15868 ( .A(n14153), .ZN(n14607) );
  INV_X1 U15869 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19367) );
  NOR2_X1 U15870 ( .A1(n15981), .A2(n19367), .ZN(n12668) );
  AOI22_X1 U15871 ( .A1(n15977), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15974), .ZN(n12666) );
  INV_X1 U15872 ( .A(n12666), .ZN(n12667) );
  NOR2_X1 U15873 ( .A1(n12668), .A2(n12667), .ZN(n12669) );
  NAND2_X1 U15874 ( .A1(n12670), .A2(n12669), .ZN(P1_U2873) );
  NAND2_X1 U15875 ( .A1(n13686), .A2(n13696), .ZN(n13593) );
  NAND2_X1 U15876 ( .A1(n13593), .A2(n12676), .ZN(n12677) );
  INV_X1 U15877 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14050) );
  NAND2_X1 U15878 ( .A1(n12758), .A2(n14050), .ZN(n12683) );
  INV_X1 U15879 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12679) );
  NAND2_X1 U15880 ( .A1(n12704), .A2(n12679), .ZN(n12681) );
  NAND2_X1 U15881 ( .A1(n13709), .A2(n14050), .ZN(n12680) );
  NAND3_X1 U15882 ( .A1(n12681), .A2(n12771), .A3(n12680), .ZN(n12682) );
  NAND2_X1 U15883 ( .A1(n12683), .A2(n12682), .ZN(n12685) );
  NAND2_X1 U15884 ( .A1(n12704), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12684) );
  OAI21_X1 U15885 ( .B1(n13566), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12684), .ZN(
        n13863) );
  XNOR2_X1 U15886 ( .A(n12685), .B(n13863), .ZN(n13710) );
  NAND2_X1 U15887 ( .A1(n13710), .A2(n13709), .ZN(n13712) );
  NAND2_X1 U15888 ( .A1(n13712), .A2(n12685), .ZN(n13753) );
  MUX2_X1 U15889 ( .A(n12768), .B(n12704), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12689) );
  INV_X1 U15890 ( .A(n12704), .ZN(n12686) );
  NAND2_X1 U15891 ( .A1(n12686), .A2(n12857), .ZN(n12731) );
  NAND2_X1 U15892 ( .A1(n12857), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12687) );
  AND2_X1 U15893 ( .A1(n12731), .A2(n12687), .ZN(n12688) );
  AND2_X1 U15894 ( .A1(n12689), .A2(n12688), .ZN(n13752) );
  MUX2_X1 U15895 ( .A(n12745), .B(n12771), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12691) );
  NAND2_X1 U15896 ( .A1(n13862), .A2(n13917), .ZN(n12690) );
  NAND2_X1 U15897 ( .A1(n12691), .A2(n12690), .ZN(n13918) );
  MUX2_X1 U15898 ( .A(n12768), .B(n12704), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12694) );
  NAND2_X1 U15899 ( .A1(n12857), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12692) );
  AND2_X1 U15900 ( .A1(n12731), .A2(n12692), .ZN(n12693) );
  NAND2_X1 U15901 ( .A1(n12694), .A2(n12693), .ZN(n13925) );
  INV_X1 U15902 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20173) );
  NAND2_X1 U15903 ( .A1(n12762), .A2(n20173), .ZN(n12697) );
  NAND2_X1 U15904 ( .A1(n13709), .A2(n20173), .ZN(n12695) );
  OAI211_X1 U15905 ( .C1(n13566), .C2(n16155), .A(n12695), .B(n12704), .ZN(
        n12696) );
  NAND2_X1 U15906 ( .A1(n12697), .A2(n12696), .ZN(n14077) );
  MUX2_X1 U15907 ( .A(n12768), .B(n12704), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12700) );
  NAND2_X1 U15908 ( .A1(n12857), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12698) );
  AND2_X1 U15909 ( .A1(n12731), .A2(n12698), .ZN(n12699) );
  AND2_X1 U15910 ( .A1(n12700), .A2(n12699), .ZN(n14096) );
  INV_X1 U15911 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20168) );
  NAND2_X1 U15912 ( .A1(n12762), .A2(n20168), .ZN(n12703) );
  INV_X1 U15913 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16179) );
  NAND2_X1 U15914 ( .A1(n13709), .A2(n20168), .ZN(n12701) );
  OAI211_X1 U15915 ( .C1(n13566), .C2(n16179), .A(n12701), .B(n12704), .ZN(
        n12702) );
  MUX2_X1 U15916 ( .A(n12768), .B(n12704), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12707) );
  NAND2_X1 U15917 ( .A1(n12857), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12705) );
  AND2_X1 U15918 ( .A1(n12731), .A2(n12705), .ZN(n12706) );
  NAND2_X1 U15919 ( .A1(n12707), .A2(n12706), .ZN(n14110) );
  INV_X1 U15920 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21307) );
  NAND2_X1 U15921 ( .A1(n12762), .A2(n21307), .ZN(n12710) );
  NAND2_X1 U15922 ( .A1(n13709), .A2(n21307), .ZN(n12708) );
  OAI211_X1 U15923 ( .C1(n13566), .C2(n16152), .A(n12708), .B(n12704), .ZN(
        n12709) );
  NAND2_X1 U15924 ( .A1(n12710), .A2(n12709), .ZN(n16144) );
  INV_X1 U15925 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n21154) );
  NAND2_X1 U15926 ( .A1(n12758), .A2(n21154), .ZN(n12714) );
  INV_X1 U15927 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14781) );
  NAND2_X1 U15928 ( .A1(n12704), .A2(n14781), .ZN(n12712) );
  NAND2_X1 U15929 ( .A1(n13709), .A2(n21154), .ZN(n12711) );
  NAND3_X1 U15930 ( .A1(n12712), .A2(n12771), .A3(n12711), .ZN(n12713) );
  MUX2_X1 U15931 ( .A(n12762), .B(n13566), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12716) );
  NOR2_X1 U15932 ( .A1(n13563), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12715) );
  NOR2_X1 U15933 ( .A1(n12716), .A2(n12715), .ZN(n15959) );
  NAND2_X1 U15934 ( .A1(n15960), .A2(n15959), .ZN(n15958) );
  INV_X1 U15935 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15971) );
  NAND2_X1 U15936 ( .A1(n12758), .A2(n15971), .ZN(n12720) );
  NAND2_X1 U15937 ( .A1(n12704), .A2(n14889), .ZN(n12718) );
  NAND2_X1 U15938 ( .A1(n13709), .A2(n15971), .ZN(n12717) );
  NAND3_X1 U15939 ( .A1(n12718), .A2(n12771), .A3(n12717), .ZN(n12719) );
  INV_X1 U15940 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n21138) );
  NAND2_X1 U15941 ( .A1(n12762), .A2(n21138), .ZN(n12723) );
  NAND2_X1 U15942 ( .A1(n13709), .A2(n21138), .ZN(n12721) );
  OAI211_X1 U15943 ( .C1(n13566), .C2(n16121), .A(n12721), .B(n12704), .ZN(
        n12722) );
  NAND2_X1 U15944 ( .A1(n12723), .A2(n12722), .ZN(n14527) );
  INV_X1 U15945 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n21038) );
  NAND2_X1 U15946 ( .A1(n12758), .A2(n21038), .ZN(n12727) );
  INV_X1 U15947 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16109) );
  NAND2_X1 U15948 ( .A1(n12704), .A2(n16109), .ZN(n12725) );
  NAND2_X1 U15949 ( .A1(n13709), .A2(n21038), .ZN(n12724) );
  NAND3_X1 U15950 ( .A1(n12725), .A2(n12771), .A3(n12724), .ZN(n12726) );
  MUX2_X1 U15951 ( .A(n12745), .B(n12771), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12729) );
  NAND2_X1 U15952 ( .A1(n11278), .A2(n13862), .ZN(n12728) );
  MUX2_X1 U15953 ( .A(n12768), .B(n12704), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12733) );
  NAND2_X1 U15954 ( .A1(n12857), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12730) );
  AND2_X1 U15955 ( .A1(n12731), .A2(n12730), .ZN(n12732) );
  NAND2_X1 U15956 ( .A1(n12733), .A2(n12732), .ZN(n14509) );
  INV_X1 U15957 ( .A(n14509), .ZN(n15922) );
  MUX2_X1 U15958 ( .A(n12745), .B(n12771), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12735) );
  NAND2_X1 U15959 ( .A1(n13862), .A2(n11280), .ZN(n12734) );
  NAND2_X1 U15960 ( .A1(n12735), .A2(n12734), .ZN(n14510) );
  NOR2_X1 U15961 ( .A1(n15922), .A2(n14510), .ZN(n12736) );
  INV_X1 U15962 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21308) );
  NAND2_X1 U15963 ( .A1(n12758), .A2(n21308), .ZN(n12740) );
  NAND2_X1 U15964 ( .A1(n12704), .A2(n16085), .ZN(n12738) );
  NAND2_X1 U15965 ( .A1(n13709), .A2(n21308), .ZN(n12737) );
  NAND3_X1 U15966 ( .A1(n12738), .A2(n12771), .A3(n12737), .ZN(n12739) );
  AND2_X1 U15967 ( .A1(n12740), .A2(n12739), .ZN(n14477) );
  MUX2_X1 U15968 ( .A(n12745), .B(n12771), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12742) );
  NAND2_X1 U15969 ( .A1(n13862), .A2(n11291), .ZN(n12741) );
  NAND2_X1 U15970 ( .A1(n12742), .A2(n12741), .ZN(n14463) );
  MUX2_X1 U15971 ( .A(n12768), .B(n12704), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12744) );
  NAND2_X1 U15972 ( .A1(n12857), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12743) );
  NAND2_X1 U15973 ( .A1(n12744), .A2(n12743), .ZN(n14451) );
  MUX2_X1 U15974 ( .A(n12745), .B(n12771), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12747) );
  NAND2_X1 U15975 ( .A1(n13862), .A2(n14884), .ZN(n12746) );
  NAND2_X1 U15976 ( .A1(n12747), .A2(n12746), .ZN(n14439) );
  MUX2_X1 U15977 ( .A(n12768), .B(n12704), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12749) );
  NAND2_X1 U15978 ( .A1(n12857), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12748) );
  INV_X1 U15979 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21330) );
  NAND2_X1 U15980 ( .A1(n12762), .A2(n21330), .ZN(n12752) );
  INV_X1 U15981 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16042) );
  NAND2_X1 U15982 ( .A1(n13709), .A2(n21330), .ZN(n12750) );
  OAI211_X1 U15983 ( .C1(n13566), .C2(n16042), .A(n12750), .B(n12704), .ZN(
        n12751) );
  NAND2_X1 U15984 ( .A1(n12752), .A2(n12751), .ZN(n14410) );
  NAND2_X1 U15985 ( .A1(n12704), .A2(n14871), .ZN(n12753) );
  OAI211_X1 U15986 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n12857), .A(n12753), .B(
        n12771), .ZN(n12754) );
  OAI21_X1 U15987 ( .B1(n12768), .B2(P1_EBX_REG_24__SCAN_IN), .A(n12754), .ZN(
        n14394) );
  NAND2_X1 U15988 ( .A1(n14411), .A2(n14394), .ZN(n14396) );
  INV_X1 U15989 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21107) );
  NAND2_X1 U15990 ( .A1(n12762), .A2(n21107), .ZN(n12757) );
  NAND2_X1 U15991 ( .A1(n13709), .A2(n21107), .ZN(n12755) );
  OAI211_X1 U15992 ( .C1(n13566), .C2(n14857), .A(n12755), .B(n12704), .ZN(
        n12756) );
  NAND2_X1 U15993 ( .A1(n12757), .A2(n12756), .ZN(n14381) );
  INV_X1 U15994 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21086) );
  NAND2_X1 U15995 ( .A1(n12758), .A2(n21086), .ZN(n12761) );
  NAND2_X1 U15996 ( .A1(n12704), .A2(n16036), .ZN(n12759) );
  OAI211_X1 U15997 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n12857), .A(n12759), .B(
        n12771), .ZN(n12760) );
  INV_X1 U15998 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n21125) );
  NAND2_X1 U15999 ( .A1(n12762), .A2(n21125), .ZN(n12765) );
  INV_X1 U16000 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14855) );
  NAND2_X1 U16001 ( .A1(n13709), .A2(n21125), .ZN(n12763) );
  OAI211_X1 U16002 ( .C1(n13566), .C2(n14855), .A(n12763), .B(n12704), .ZN(
        n12764) );
  AND2_X1 U16003 ( .A1(n12765), .A2(n12764), .ZN(n14354) );
  INV_X1 U16004 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14649) );
  NAND2_X1 U16005 ( .A1(n12704), .A2(n14649), .ZN(n12766) );
  OAI211_X1 U16006 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n12857), .A(n12766), .B(
        n12771), .ZN(n12767) );
  OAI21_X1 U16007 ( .B1(n12768), .B2(P1_EBX_REG_28__SCAN_IN), .A(n12767), .ZN(
        n14344) );
  INV_X1 U16008 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n21269) );
  NAND2_X1 U16009 ( .A1(n13709), .A2(n21269), .ZN(n12769) );
  OAI21_X1 U16010 ( .B1(n13563), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12769), .ZN(n12770) );
  MUX2_X1 U16011 ( .A(n12769), .B(n12770), .S(n12771), .Z(n14330) );
  OAI22_X1 U16012 ( .A1(n14332), .A2(n12771), .B1(n12770), .B2(n9868), .ZN(
        n12774) );
  AND2_X1 U16013 ( .A1(n12857), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12772) );
  AOI21_X1 U16014 ( .B1(n13563), .B2(P1_EBX_REG_30__SCAN_IN), .A(n12772), .ZN(
        n12856) );
  INV_X1 U16015 ( .A(n12856), .ZN(n12773) );
  XNOR2_X1 U16016 ( .A(n12774), .B(n12773), .ZN(n14818) );
  INV_X1 U16017 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14319) );
  INV_X1 U16018 ( .A(n12775), .ZN(n12776) );
  OAI21_X2 U16019 ( .B1(n12779), .B2(n12778), .A(n12777), .ZN(n12892) );
  NAND2_X1 U16020 ( .A1(n12785), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12781) );
  XNOR2_X1 U16021 ( .A(n12784), .B(n12781), .ZN(n16209) );
  NAND2_X1 U16022 ( .A1(n16209), .A2(n12788), .ZN(n12782) );
  INV_X1 U16023 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12899) );
  NAND2_X1 U16024 ( .A1(n12782), .A2(n12899), .ZN(n12888) );
  NOR2_X1 U16025 ( .A1(n12782), .A2(n12899), .ZN(n12890) );
  INV_X1 U16026 ( .A(n12890), .ZN(n12783) );
  MUX2_X1 U16027 ( .A(n12787), .B(n12786), .S(n12785), .Z(n16199) );
  NAND2_X1 U16028 ( .A1(n16199), .A2(n12788), .ZN(n12789) );
  XNOR2_X1 U16029 ( .A(n12790), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12946) );
  INV_X1 U16030 ( .A(n12895), .ZN(n12794) );
  OR2_X1 U16031 ( .A1(n12798), .A2(n12899), .ZN(n12792) );
  AOI22_X1 U16032 ( .A1(n11925), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12791) );
  OAI211_X1 U16033 ( .C1(n12793), .C2(n10110), .A(n12792), .B(n12791), .ZN(
        n12894) );
  NAND2_X1 U16034 ( .A1(n12794), .A2(n12894), .ZN(n12800) );
  INV_X1 U16035 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14912) );
  AOI22_X1 U16036 ( .A1(n11925), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12797) );
  NAND2_X1 U16037 ( .A1(n12795), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12796) );
  OAI211_X1 U16038 ( .C1(n12798), .C2(n14912), .A(n12797), .B(n12796), .ZN(
        n12799) );
  INV_X1 U16039 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19946) );
  NOR2_X1 U16040 ( .A1(n12810), .A2(n19946), .ZN(n12802) );
  INV_X1 U16041 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n15319) );
  OAI22_X1 U16042 ( .A1(n12813), .A2(n15629), .B1(n12811), .B2(n15319), .ZN(
        n12801) );
  OR2_X1 U16043 ( .A1(n12802), .A2(n12801), .ZN(n15314) );
  AOI22_X1 U16044 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12805) );
  NAND2_X1 U16045 ( .A1(n12822), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U16046 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U16047 ( .A1(n12822), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U16048 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12809) );
  NAND2_X1 U16049 ( .A1(n12822), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12808) );
  NAND2_X1 U16050 ( .A1(n12809), .A2(n12808), .ZN(n15009) );
  INV_X1 U16051 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19954) );
  NOR2_X1 U16052 ( .A1(n12810), .A2(n19954), .ZN(n12815) );
  INV_X1 U16053 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15285) );
  OAI22_X1 U16054 ( .A1(n12813), .A2(n12812), .B1(n12811), .B2(n15285), .ZN(
        n12814) );
  OR2_X1 U16055 ( .A1(n12815), .A2(n12814), .ZN(n15284) );
  NAND2_X1 U16056 ( .A1(n15008), .A2(n15284), .ZN(n15283) );
  AOI22_X1 U16057 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12817) );
  NAND2_X1 U16058 ( .A1(n12822), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12816) );
  NAND2_X2 U16059 ( .A1(n15570), .A2(n10345), .ZN(n15569) );
  AOI22_X1 U16060 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12819) );
  NAND2_X1 U16061 ( .A1(n12822), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12818) );
  AND2_X1 U16062 ( .A1(n12819), .A2(n12818), .ZN(n15274) );
  INV_X1 U16063 ( .A(n15274), .ZN(n12820) );
  AOI22_X1 U16064 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12824) );
  NAND2_X1 U16065 ( .A1(n12822), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U16066 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U16067 ( .A1(n12822), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U16068 ( .A1(n12826), .A2(n12825), .ZN(n15261) );
  AOI22_X1 U16069 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U16070 ( .A1(n12822), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12827) );
  NAND2_X1 U16071 ( .A1(n12828), .A2(n12827), .ZN(n14984) );
  AND2_X2 U16072 ( .A1(n14983), .A2(n14984), .ZN(n15245) );
  AOI22_X1 U16073 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12830) );
  NAND2_X1 U16074 ( .A1(n12822), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12829) );
  NAND2_X1 U16075 ( .A1(n12830), .A2(n12829), .ZN(n15244) );
  NAND2_X2 U16076 ( .A1(n15245), .A2(n15244), .ZN(n15247) );
  AOI22_X1 U16077 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U16078 ( .A1(n12822), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12831) );
  AND2_X1 U16079 ( .A1(n12832), .A2(n12831), .ZN(n14957) );
  NOR2_X2 U16080 ( .A1(n15247), .A2(n14957), .ZN(n12896) );
  AOI22_X1 U16081 ( .A1(n12835), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n12821), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n12834) );
  NAND2_X1 U16082 ( .A1(n12822), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12833) );
  NAND2_X1 U16083 ( .A1(n12834), .A2(n12833), .ZN(n12897) );
  NAND2_X1 U16084 ( .A1(n12896), .A2(n12897), .ZN(n12837) );
  AOI222_X1 U16085 ( .A1(n12822), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12835), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n12821), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n12836) );
  XNOR2_X1 U16086 ( .A(n12837), .B(n12836), .ZN(n16204) );
  NAND2_X1 U16087 ( .A1(P2_REIP_REG_31__SCAN_IN), .A2(n19287), .ZN(n12951) );
  OAI21_X1 U16088 ( .B1(n16204), .B2(n19301), .A(n12951), .ZN(n12847) );
  NOR3_X1 U16089 ( .A1(n15508), .A2(n15520), .A3(n15492), .ZN(n12900) );
  NAND2_X1 U16090 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15527) );
  NAND2_X1 U16091 ( .A1(n16383), .A2(n15555), .ZN(n12839) );
  NAND2_X1 U16092 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15568) );
  NAND2_X1 U16093 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15594) );
  NOR3_X1 U16094 ( .A1(n15405), .A2(n12838), .A3(n15594), .ZN(n12841) );
  AOI21_X1 U16095 ( .B1(n15607), .B2(n12841), .A(n15688), .ZN(n15597) );
  AOI21_X1 U16096 ( .B1(n16383), .B2(n15568), .A(n15597), .ZN(n15556) );
  NAND2_X1 U16097 ( .A1(n12839), .A2(n15556), .ZN(n15545) );
  AOI21_X1 U16098 ( .B1(n15527), .B2(n19305), .A(n15545), .ZN(n15521) );
  OAI21_X1 U16099 ( .B1(n15608), .B2(n12900), .A(n15521), .ZN(n12904) );
  AOI21_X1 U16100 ( .B1(n12899), .B2(n19305), .A(n12904), .ZN(n12840) );
  OR2_X1 U16101 ( .A1(n12840), .A2(n14912), .ZN(n12845) );
  NAND2_X1 U16102 ( .A1(n12841), .A2(n16393), .ZN(n15585) );
  INV_X1 U16103 ( .A(n15568), .ZN(n15554) );
  NAND2_X1 U16104 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15554), .ZN(
        n12842) );
  NOR2_X1 U16105 ( .A1(n15585), .A2(n12842), .ZN(n15547) );
  INV_X1 U16106 ( .A(n15527), .ZN(n12843) );
  NAND4_X1 U16107 ( .A1(n15493), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12900), .A4(n14912), .ZN(n12844) );
  NAND2_X1 U16108 ( .A1(n12845), .A2(n12844), .ZN(n12846) );
  NOR2_X1 U16109 ( .A1(n12847), .A2(n12846), .ZN(n12848) );
  NAND2_X1 U16110 ( .A1(n10458), .A2(n20266), .ZN(n12849) );
  NOR2_X1 U16111 ( .A1(n13456), .A2(n20074), .ZN(n12850) );
  NAND2_X1 U16112 ( .A1(n13597), .A2(n12850), .ZN(n13447) );
  NOR2_X1 U16113 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20834), .ZN(n12851) );
  NAND2_X1 U16114 ( .A1(n20834), .A2(n10577), .ZN(n20935) );
  OAI21_X1 U16115 ( .B1(n20661), .B2(n20935), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n15873) );
  OAI21_X1 U16116 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n12851), .A(n15873), 
        .ZN(n12853) );
  INV_X1 U16117 ( .A(n15867), .ZN(n12852) );
  OAI21_X1 U16118 ( .B1(n12853), .B2(n12852), .A(n16162), .ZN(n12854) );
  NAND2_X1 U16119 ( .A1(n12855), .A2(n20123), .ZN(n12887) );
  MUX2_X1 U16120 ( .A(n12771), .B(n12856), .S(n14332), .Z(n12859) );
  AOI22_X1 U16121 ( .A1(n13563), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12857), .ZN(n12858) );
  OR2_X2 U16122 ( .A1(n20117), .A2(n10577), .ZN(n14036) );
  NAND2_X1 U16123 ( .A1(n20940), .A2(n21137), .ZN(n15868) );
  NAND3_X1 U16124 ( .A1(n13709), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n15868), 
        .ZN(n12860) );
  INV_X1 U16125 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20860) );
  INV_X1 U16126 ( .A(n20940), .ZN(n20846) );
  INV_X1 U16127 ( .A(n12861), .ZN(n12862) );
  NAND2_X1 U16128 ( .A1(n12862), .A2(n20837), .ZN(n20933) );
  NOR2_X1 U16129 ( .A1(n20846), .A2(n20933), .ZN(n20931) );
  INV_X1 U16130 ( .A(n20931), .ZN(n13587) );
  NAND2_X1 U16131 ( .A1(n13630), .A2(n13587), .ZN(n13676) );
  NAND2_X1 U16132 ( .A1(n13676), .A2(n21137), .ZN(n12877) );
  OR2_X1 U16133 ( .A1(n12877), .A2(n20266), .ZN(n12863) );
  OR2_X2 U16134 ( .A1(n14036), .A2(n12863), .ZN(n20148) );
  INV_X2 U16135 ( .A(n20148), .ZN(n15941) );
  NAND3_X1 U16136 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .ZN(n20147) );
  NOR2_X1 U16137 ( .A1(n21299), .A2(n20147), .ZN(n20146) );
  NAND2_X1 U16138 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n12864) );
  NOR2_X2 U16139 ( .A1(n20131), .A2(n12864), .ZN(n20112) );
  NAND2_X1 U16140 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20112), .ZN(n14114) );
  NOR2_X2 U16141 ( .A1(n20860), .A2(n14114), .ZN(n20095) );
  NAND3_X1 U16142 ( .A1(n20095), .A2(P1_REIP_REG_9__SCAN_IN), .A3(
        P1_REIP_REG_10__SCAN_IN), .ZN(n15967) );
  NAND4_X1 U16143 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n12867) );
  NOR2_X2 U16144 ( .A1(n15967), .A2(n12867), .ZN(n15921) );
  AND3_X1 U16145 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_17__SCAN_IN), .ZN(n12865) );
  AND2_X2 U16146 ( .A1(n15921), .A2(n12865), .ZN(n14431) );
  NAND3_X1 U16147 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14434) );
  NAND2_X1 U16148 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n12866) );
  NOR2_X1 U16149 ( .A1(n14434), .A2(n12866), .ZN(n14403) );
  AND2_X1 U16150 ( .A1(n14403), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n12872) );
  INV_X1 U16152 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20883) );
  INV_X1 U16153 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20879) );
  INV_X1 U16154 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21272) );
  NOR4_X2 U16155 ( .A1(n14393), .A2(n20883), .A3(n20879), .A4(n21272), .ZN(
        n14362) );
  NAND3_X1 U16156 ( .A1(n14362), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14340) );
  INV_X1 U16157 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21044) );
  INV_X1 U16158 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14626) );
  NOR4_X1 U16159 ( .A1(n14340), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21044), 
        .A4(n14626), .ZN(n12883) );
  INV_X1 U16160 ( .A(n12867), .ZN(n12870) );
  NAND2_X1 U16161 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n12869) );
  INV_X1 U16162 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21261) );
  INV_X1 U16163 ( .A(n20146), .ZN(n20116) );
  NOR4_X1 U16164 ( .A1(n20117), .A2(n20860), .A3(n21261), .A4(n20116), .ZN(
        n12868) );
  NAND3_X1 U16165 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n12868), .ZN(n14196) );
  NOR2_X1 U16166 ( .A1(n12869), .A2(n14196), .ZN(n14197) );
  NAND2_X1 U16167 ( .A1(n12870), .A2(n14197), .ZN(n14433) );
  INV_X1 U16168 ( .A(n14433), .ZN(n14491) );
  NAND3_X1 U16169 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14432) );
  INV_X1 U16170 ( .A(n14432), .ZN(n12871) );
  AND2_X1 U16171 ( .A1(n12872), .A2(n12871), .ZN(n12873) );
  NAND2_X1 U16172 ( .A1(n14491), .A2(n12873), .ZN(n14384) );
  NAND3_X1 U16173 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_25__SCAN_IN), .ZN(n12874) );
  NOR2_X1 U16174 ( .A1(n14384), .A2(n12874), .ZN(n14358) );
  NAND3_X1 U16175 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .A3(n14358), .ZN(n14333) );
  NAND2_X1 U16176 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n12876) );
  INV_X1 U16177 ( .A(n20117), .ZN(n12875) );
  OAI21_X1 U16178 ( .B1(n14333), .B2(n12876), .A(n20115), .ZN(n14317) );
  NOR2_X1 U16179 ( .A1(n14317), .A2(n21028), .ZN(n12882) );
  INV_X1 U16180 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n21166) );
  OAI22_X1 U16181 ( .A1(n20107), .A2(n21166), .B1(n12880), .B2(n20098), .ZN(
        n12881) );
  NOR3_X1 U16182 ( .A1(n12883), .A2(n12882), .A3(n12881), .ZN(n12884) );
  NAND2_X1 U16183 ( .A1(n12887), .A2(n12886), .ZN(P1_U2809) );
  INV_X1 U16184 ( .A(n12888), .ZN(n12889) );
  NOR2_X1 U16185 ( .A1(n12890), .A2(n12889), .ZN(n12891) );
  XNOR2_X1 U16186 ( .A(n12892), .B(n12891), .ZN(n12936) );
  XNOR2_X1 U16187 ( .A(n12893), .B(n12899), .ZN(n12942) );
  INV_X1 U16188 ( .A(n16211), .ZN(n12903) );
  INV_X1 U16189 ( .A(n12896), .ZN(n14959) );
  NAND2_X1 U16190 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n19287), .ZN(n12939) );
  INV_X1 U16191 ( .A(n12939), .ZN(n12898) );
  NAND3_X1 U16192 ( .A1(n15493), .A2(n12900), .A3(n12899), .ZN(n12901) );
  OAI211_X1 U16193 ( .C1(n12903), .C2(n19308), .A(n12902), .B(n12901), .ZN(
        n12907) );
  NOR2_X1 U16194 ( .A1(n12905), .A2(n12899), .ZN(n12906) );
  NOR2_X1 U16195 ( .A1(n12907), .A2(n12906), .ZN(n12908) );
  OAI21_X1 U16196 ( .B1(n12942), .B2(n19303), .A(n12908), .ZN(n12909) );
  NAND2_X1 U16197 ( .A1(n10325), .A2(n12910), .ZN(P2_U3016) );
  NOR2_X1 U16198 ( .A1(n12917), .A2(n12919), .ZN(n15879) );
  INV_X1 U16199 ( .A(n15878), .ZN(n12916) );
  INV_X1 U16200 ( .A(n12919), .ZN(n12914) );
  INV_X1 U16201 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18967) );
  AOI22_X1 U16202 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17877), .B1(
        n17779), .B2(n18967), .ZN(n12913) );
  NAND2_X1 U16203 ( .A1(n12916), .A2(n12915), .ZN(n12923) );
  INV_X1 U16204 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16507) );
  OAI22_X1 U16205 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18967), .B1(
        n12919), .B2(n12918), .ZN(n12921) );
  NAND2_X1 U16206 ( .A1(n12921), .A2(n12920), .ZN(n12922) );
  NAND2_X1 U16207 ( .A1(n12923), .A2(n12922), .ZN(n13327) );
  NAND2_X1 U16208 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16498), .ZN(
        n12924) );
  INV_X1 U16209 ( .A(n16985), .ZN(n16931) );
  INV_X1 U16210 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18935) );
  NOR2_X1 U16211 ( .A1(n18935), .A2(n16515), .ZN(n13321) );
  OAI21_X1 U16212 ( .B1(n17975), .B2(n17721), .A(n18348), .ZN(n17771) );
  OR2_X1 U16213 ( .A1(n12925), .A2(n17736), .ZN(n16503) );
  INV_X1 U16214 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16669) );
  XOR2_X1 U16215 ( .A(n16669), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12928) );
  NOR2_X1 U16216 ( .A1(n12927), .A2(n12926), .ZN(n16502) );
  OAI22_X1 U16217 ( .A1(n16503), .A2(n12928), .B1(n16502), .B2(n16669), .ZN(
        n12929) );
  AOI211_X1 U16218 ( .C1(n17828), .C2(n16931), .A(n13321), .B(n12929), .ZN(
        n12933) );
  NAND2_X1 U16219 ( .A1(n15821), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12930) );
  XNOR2_X1 U16220 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12930), .ZN(
        n13311) );
  NAND2_X1 U16221 ( .A1(n13311), .A2(n17703), .ZN(n12932) );
  NAND3_X1 U16222 ( .A1(n16508), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n17985), .ZN(n12931) );
  XOR2_X1 U16223 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12931), .Z(
        n13325) );
  NAND3_X1 U16224 ( .A1(n12933), .A2(n12932), .A3(n10335), .ZN(n12934) );
  INV_X1 U16225 ( .A(n12935), .ZN(P3_U2799) );
  INV_X1 U16226 ( .A(n12936), .ZN(n12937) );
  XNOR2_X1 U16227 ( .A(n12947), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16214) );
  NAND2_X1 U16228 ( .A1(n16355), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12938) );
  OAI211_X1 U16229 ( .C1(n16366), .C2(n16214), .A(n12939), .B(n12938), .ZN(
        n12940) );
  NAND2_X1 U16230 ( .A1(n12945), .A2(n12944), .ZN(P2_U2984) );
  INV_X1 U16231 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12948) );
  NAND2_X1 U16232 ( .A1(n16355), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12950) );
  OAI211_X1 U16233 ( .C1(n16366), .C2(n14911), .A(n12951), .B(n12950), .ZN(
        n12952) );
  OAI211_X1 U16234 ( .C1(n12955), .C2(n19278), .A(n12954), .B(n12953), .ZN(
        P2_U2983) );
  NAND2_X1 U16235 ( .A1(n12956), .A2(n12978), .ZN(n12965) );
  NAND2_X1 U16236 ( .A1(n11853), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12959) );
  NAND2_X1 U16237 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19831) );
  INV_X1 U16238 ( .A(n19831), .ZN(n12960) );
  NAND2_X1 U16239 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12960), .ZN(
        n12969) );
  INV_X1 U16240 ( .A(n12969), .ZN(n12961) );
  NAND2_X1 U16241 ( .A1(n12961), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19834) );
  OAI211_X1 U16242 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n12961), .A(
        n19834), .B(n20007), .ZN(n12962) );
  INV_X1 U16243 ( .A(n12962), .ZN(n12963) );
  AOI21_X1 U16244 ( .B1(n12979), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12963), .ZN(n12964) );
  NOR2_X1 U16245 ( .A1(n13213), .A2(n13035), .ZN(n12966) );
  NAND2_X1 U16246 ( .A1(n12991), .A2(n12966), .ZN(n13780) );
  NAND2_X1 U16247 ( .A1(n12968), .A2(n12978), .ZN(n12973) );
  NAND2_X1 U16248 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19686) );
  NAND2_X1 U16249 ( .A1(n19686), .A2(n20019), .ZN(n12970) );
  NAND2_X1 U16250 ( .A1(n12970), .A2(n12969), .ZN(n19465) );
  NOR2_X1 U16251 ( .A1(n20002), .A2(n19465), .ZN(n12971) );
  AOI21_X1 U16252 ( .B1(n12979), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12971), .ZN(n12972) );
  NAND2_X1 U16253 ( .A1(n13160), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12986) );
  AOI22_X1 U16254 ( .A1(n12979), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20007), .B2(n20036), .ZN(n12975) );
  NAND2_X1 U16255 ( .A1(n16452), .A2(n12978), .ZN(n12981) );
  NAND2_X1 U16256 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20028), .ZN(
        n19620) );
  NAND2_X1 U16257 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20036), .ZN(
        n19653) );
  NAND2_X1 U16258 ( .A1(n19620), .A2(n19653), .ZN(n19464) );
  AND2_X1 U16259 ( .A1(n20007), .A2(n19464), .ZN(n19652) );
  AOI21_X1 U16260 ( .B1(n12979), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19652), .ZN(n12980) );
  NAND2_X1 U16261 ( .A1(n12981), .A2(n12980), .ZN(n13507) );
  INV_X1 U16262 ( .A(n12982), .ZN(n15759) );
  INV_X1 U16263 ( .A(n12983), .ZN(n12984) );
  NAND2_X1 U16264 ( .A1(n15759), .A2(n12984), .ZN(n12985) );
  NAND2_X1 U16265 ( .A1(n13663), .A2(n13664), .ZN(n13662) );
  INV_X1 U16266 ( .A(n12986), .ZN(n12987) );
  NAND2_X1 U16267 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  NAND2_X1 U16268 ( .A1(n13662), .A2(n12989), .ZN(n13788) );
  NAND2_X1 U16269 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n11853), .ZN(
        n12990) );
  AND2_X1 U16270 ( .A1(n12991), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12992) );
  INV_X1 U16271 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12994) );
  NAND2_X1 U16272 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13802) );
  NOR2_X1 U16273 ( .A1(n12994), .A2(n13802), .ZN(n13842) );
  AOI22_X1 U16274 ( .A1(n12258), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13101), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U16275 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U16276 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U16277 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12998) );
  NAND4_X1 U16278 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        n13007) );
  AOI22_X1 U16279 ( .A1(n13032), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U16280 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16281 ( .A1(n11789), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U16282 ( .A1(n12080), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13002) );
  NAND4_X1 U16283 ( .A1(n13005), .A2(n13004), .A3(n13003), .A4(n13002), .ZN(
        n13006) );
  NOR2_X1 U16284 ( .A1(n13007), .A2(n13006), .ZN(n14123) );
  AOI22_X1 U16285 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U16286 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13010) );
  AOI22_X1 U16287 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13009) );
  AOI22_X1 U16288 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13008) );
  NAND4_X1 U16289 ( .A1(n13011), .A2(n13010), .A3(n13009), .A4(n13008), .ZN(
        n13017) );
  AOI22_X1 U16290 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13015) );
  AOI22_X1 U16291 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U16292 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U16293 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11790), .B1(
        n12080), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13012) );
  NAND4_X1 U16294 ( .A1(n13015), .A2(n13014), .A3(n13013), .A4(n13012), .ZN(
        n13016) );
  OR2_X1 U16295 ( .A1(n13017), .A2(n13016), .ZN(n14176) );
  AOI22_X1 U16296 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16297 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U16298 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13019) );
  AOI22_X1 U16299 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13018) );
  NAND4_X1 U16300 ( .A1(n13021), .A2(n13020), .A3(n13019), .A4(n13018), .ZN(
        n13027) );
  AOI22_X1 U16301 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U16302 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13024) );
  AOI22_X1 U16303 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13023) );
  AOI22_X1 U16304 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11790), .B1(
        n12080), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13022) );
  NAND4_X1 U16305 ( .A1(n13025), .A2(n13024), .A3(n13023), .A4(n13022), .ZN(
        n13026) );
  AOI22_X1 U16306 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U16307 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U16308 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13029) );
  AOI22_X1 U16309 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13028) );
  NAND4_X1 U16310 ( .A1(n13031), .A2(n13030), .A3(n13029), .A4(n13028), .ZN(
        n13042) );
  AOI22_X1 U16311 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U16312 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U16313 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11790), .B1(
        n12080), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13038) );
  INV_X1 U16314 ( .A(n13032), .ZN(n13060) );
  INV_X1 U16315 ( .A(n13033), .ZN(n13059) );
  OAI22_X1 U16316 ( .A1(n13035), .A2(n13060), .B1(n13059), .B2(n13034), .ZN(
        n13036) );
  INV_X1 U16317 ( .A(n13036), .ZN(n13037) );
  NAND4_X1 U16318 ( .A1(n13040), .A2(n13039), .A3(n13038), .A4(n13037), .ZN(
        n13041) );
  NOR2_X1 U16319 ( .A1(n13042), .A2(n13041), .ZN(n15212) );
  AOI22_X1 U16320 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U16321 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U16322 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U16323 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13044) );
  NAND4_X1 U16324 ( .A1(n13047), .A2(n13046), .A3(n13045), .A4(n13044), .ZN(
        n13053) );
  AOI22_X1 U16325 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13051) );
  AOI22_X1 U16326 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16327 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U16328 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11790), .B1(
        n12080), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13048) );
  NAND4_X1 U16329 ( .A1(n13051), .A2(n13050), .A3(n13049), .A4(n13048), .ZN(
        n13052) );
  NOR2_X1 U16330 ( .A1(n13053), .A2(n13052), .ZN(n15203) );
  AOI22_X1 U16331 ( .A1(n12258), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13101), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U16332 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U16333 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16334 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13054) );
  NAND4_X1 U16335 ( .A1(n13057), .A2(n13056), .A3(n13055), .A4(n13054), .ZN(
        n13067) );
  AOI22_X1 U16336 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U16337 ( .A1(n11789), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16338 ( .A1(n12080), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13063) );
  OAI22_X1 U16339 ( .A1(n13801), .A2(n13060), .B1(n13059), .B2(n13058), .ZN(
        n13061) );
  INV_X1 U16340 ( .A(n13061), .ZN(n13062) );
  NAND4_X1 U16341 ( .A1(n13065), .A2(n13064), .A3(n13063), .A4(n13062), .ZN(
        n13066) );
  OR2_X1 U16342 ( .A1(n13067), .A2(n13066), .ZN(n15200) );
  AOI22_X1 U16343 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13101), .B1(
        n12258), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16344 ( .A1(n11781), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U16345 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U16346 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13068) );
  NAND4_X1 U16347 ( .A1(n13071), .A2(n13070), .A3(n13069), .A4(n13068), .ZN(
        n13077) );
  AOI22_X1 U16348 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13032), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U16349 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13074) );
  AOI22_X1 U16350 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11789), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U16351 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11790), .B1(
        n12080), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13072) );
  NAND4_X1 U16352 ( .A1(n13075), .A2(n13074), .A3(n13073), .A4(n13072), .ZN(
        n13076) );
  NOR2_X1 U16353 ( .A1(n13077), .A2(n13076), .ZN(n15192) );
  INV_X1 U16354 ( .A(n13280), .ZN(n13252) );
  INV_X1 U16355 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13079) );
  INV_X1 U16356 ( .A(n13278), .ZN(n13251) );
  INV_X1 U16357 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13078) );
  OAI22_X1 U16358 ( .A1(n13252), .A2(n13079), .B1(n13251), .B2(n13078), .ZN(
        n13083) );
  INV_X1 U16359 ( .A(n11759), .ZN(n13255) );
  INV_X1 U16360 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13081) );
  INV_X1 U16361 ( .A(n11748), .ZN(n13253) );
  INV_X1 U16362 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13080) );
  OAI22_X1 U16363 ( .A1(n13255), .A2(n13081), .B1(n13253), .B2(n13080), .ZN(
        n13082) );
  NOR2_X1 U16364 ( .A1(n13083), .A2(n13082), .ZN(n13087) );
  AOI22_X1 U16365 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U16366 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13085) );
  XNOR2_X1 U16367 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13281) );
  NAND4_X1 U16368 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13281), .ZN(
        n13096) );
  INV_X1 U16369 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13088) );
  INV_X1 U16370 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19799) );
  OAI22_X1 U16371 ( .A1(n13252), .A2(n13088), .B1(n13251), .B2(n19799), .ZN(
        n13091) );
  INV_X1 U16372 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13089) );
  INV_X1 U16373 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19631) );
  OAI22_X1 U16374 ( .A1(n13255), .A2(n13089), .B1(n13253), .B2(n19631), .ZN(
        n13090) );
  NOR2_X1 U16375 ( .A1(n13091), .A2(n13090), .ZN(n13094) );
  INV_X1 U16376 ( .A(n13281), .ZN(n13272) );
  AOI22_X1 U16377 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16378 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13092) );
  NAND4_X1 U16379 ( .A1(n13094), .A2(n13272), .A3(n13093), .A4(n13092), .ZN(
        n13095) );
  AND2_X1 U16380 ( .A1(n13096), .A2(n13095), .ZN(n13134) );
  NAND2_X1 U16381 ( .A1(n20060), .A2(n13134), .ZN(n13108) );
  AOI22_X1 U16382 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11658), .B1(
        n11781), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16383 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13033), .B1(
        n12080), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13099) );
  AOI22_X1 U16384 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n13032), .B1(
        n11772), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U16385 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11789), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13097) );
  NAND4_X1 U16386 ( .A1(n13100), .A2(n13099), .A3(n13098), .A4(n13097), .ZN(
        n13107) );
  AOI22_X1 U16387 ( .A1(n12258), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U16388 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11767), .B1(
        n12175), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U16389 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11783), .B1(
        n11610), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U16390 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13102) );
  NAND4_X1 U16391 ( .A1(n13105), .A2(n13104), .A3(n13103), .A4(n13102), .ZN(
        n13106) );
  OR2_X1 U16392 ( .A1(n13107), .A2(n13106), .ZN(n13131) );
  XNOR2_X1 U16393 ( .A(n13108), .B(n13131), .ZN(n13137) );
  XNOR2_X1 U16394 ( .A(n13109), .B(n13137), .ZN(n15187) );
  NAND2_X1 U16395 ( .A1(n12173), .A2(n13134), .ZN(n15186) );
  OAI22_X1 U16396 ( .A1(n13255), .A2(n13112), .B1(n13251), .B2(n13111), .ZN(
        n13116) );
  OAI22_X1 U16397 ( .A1(n13252), .A2(n13114), .B1(n13253), .B2(n13113), .ZN(
        n13115) );
  NOR2_X1 U16398 ( .A1(n13116), .A2(n13115), .ZN(n13119) );
  AOI22_X1 U16399 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U16400 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13117) );
  NAND4_X1 U16401 ( .A1(n13119), .A2(n13118), .A3(n13117), .A4(n13281), .ZN(
        n13130) );
  INV_X1 U16402 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13121) );
  OAI22_X1 U16403 ( .A1(n13255), .A2(n13121), .B1(n13251), .B2(n13120), .ZN(
        n13125) );
  OAI22_X1 U16404 ( .A1(n13252), .A2(n13123), .B1(n13253), .B2(n13122), .ZN(
        n13124) );
  NOR2_X1 U16405 ( .A1(n13125), .A2(n13124), .ZN(n13128) );
  AOI22_X1 U16406 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13127) );
  AOI22_X1 U16407 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13126) );
  NAND4_X1 U16408 ( .A1(n13128), .A2(n13272), .A3(n13127), .A4(n13126), .ZN(
        n13129) );
  NAND2_X1 U16409 ( .A1(n13130), .A2(n13129), .ZN(n13138) );
  NAND2_X1 U16410 ( .A1(n13131), .A2(n13134), .ZN(n13139) );
  XOR2_X1 U16411 ( .A(n13138), .B(n13139), .Z(n13132) );
  NAND2_X1 U16412 ( .A1(n13132), .A2(n13160), .ZN(n15174) );
  INV_X1 U16413 ( .A(n13138), .ZN(n13133) );
  NAND2_X1 U16414 ( .A1(n12173), .A2(n13133), .ZN(n15177) );
  INV_X1 U16415 ( .A(n13134), .ZN(n13135) );
  NOR2_X1 U16416 ( .A1(n15177), .A2(n13135), .ZN(n13136) );
  NOR2_X1 U16417 ( .A1(n13139), .A2(n13138), .ZN(n13161) );
  INV_X1 U16418 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13141) );
  INV_X1 U16419 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13140) );
  OAI22_X1 U16420 ( .A1(n13255), .A2(n13141), .B1(n13251), .B2(n13140), .ZN(
        n13145) );
  INV_X1 U16421 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13143) );
  INV_X1 U16422 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13142) );
  OAI22_X1 U16423 ( .A1(n13252), .A2(n13143), .B1(n13253), .B2(n13142), .ZN(
        n13144) );
  NOR2_X1 U16424 ( .A1(n13145), .A2(n13144), .ZN(n13148) );
  AOI22_X1 U16425 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U16426 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13146) );
  NAND4_X1 U16427 ( .A1(n13148), .A2(n13147), .A3(n13146), .A4(n13281), .ZN(
        n13159) );
  INV_X1 U16428 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13150) );
  INV_X1 U16429 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13149) );
  OAI22_X1 U16430 ( .A1(n13255), .A2(n13150), .B1(n13251), .B2(n13149), .ZN(
        n13154) );
  INV_X1 U16431 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13152) );
  INV_X1 U16432 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13151) );
  OAI22_X1 U16433 ( .A1(n13252), .A2(n13152), .B1(n13253), .B2(n13151), .ZN(
        n13153) );
  NOR2_X1 U16434 ( .A1(n13154), .A2(n13153), .ZN(n13157) );
  AOI22_X1 U16435 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U16436 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13155) );
  NAND4_X1 U16437 ( .A1(n13157), .A2(n13272), .A3(n13156), .A4(n13155), .ZN(
        n13158) );
  NAND2_X1 U16438 ( .A1(n13161), .A2(n13162), .ZN(n13187) );
  OAI211_X1 U16439 ( .C1(n13161), .C2(n13162), .A(n13160), .B(n13187), .ZN(
        n13164) );
  INV_X1 U16440 ( .A(n13162), .ZN(n13163) );
  NOR2_X1 U16441 ( .A1(n20060), .A2(n13163), .ZN(n15170) );
  NAND2_X1 U16442 ( .A1(n15171), .A2(n15170), .ZN(n15169) );
  OAI22_X1 U16443 ( .A1(n13255), .A2(n13168), .B1(n13251), .B2(n13167), .ZN(
        n13172) );
  OAI22_X1 U16444 ( .A1(n13252), .A2(n13170), .B1(n13253), .B2(n13169), .ZN(
        n13171) );
  NOR2_X1 U16445 ( .A1(n13172), .A2(n13171), .ZN(n13175) );
  AOI22_X1 U16446 ( .A1(n13258), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13174) );
  AOI22_X1 U16447 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13173) );
  NAND4_X1 U16448 ( .A1(n13175), .A2(n13174), .A3(n13173), .A4(n13281), .ZN(
        n13186) );
  OAI22_X1 U16449 ( .A1(n13255), .A2(n13177), .B1(n13251), .B2(n13176), .ZN(
        n13181) );
  OAI22_X1 U16450 ( .A1(n13252), .A2(n13179), .B1(n13253), .B2(n13178), .ZN(
        n13180) );
  NOR2_X1 U16451 ( .A1(n13181), .A2(n13180), .ZN(n13184) );
  AOI22_X1 U16452 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13183) );
  AOI22_X1 U16453 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13182) );
  NAND4_X1 U16454 ( .A1(n13184), .A2(n13272), .A3(n13183), .A4(n13182), .ZN(
        n13185) );
  NAND2_X1 U16455 ( .A1(n13186), .A2(n13185), .ZN(n13189) );
  AOI21_X1 U16456 ( .B1(n13187), .B2(n13189), .A(n13213), .ZN(n13188) );
  OR2_X1 U16457 ( .A1(n13187), .A2(n13189), .ZN(n13214) );
  NAND2_X1 U16458 ( .A1(n13188), .A2(n13214), .ZN(n13191) );
  NOR2_X1 U16459 ( .A1(n12584), .A2(n13189), .ZN(n15163) );
  INV_X1 U16460 ( .A(n13190), .ZN(n13192) );
  INV_X1 U16461 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13194) );
  INV_X1 U16462 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13193) );
  OAI22_X1 U16463 ( .A1(n13255), .A2(n13194), .B1(n13251), .B2(n13193), .ZN(
        n13198) );
  INV_X1 U16464 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13196) );
  INV_X1 U16465 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13195) );
  OAI22_X1 U16466 ( .A1(n13252), .A2(n13196), .B1(n13253), .B2(n13195), .ZN(
        n13197) );
  NOR2_X1 U16467 ( .A1(n13198), .A2(n13197), .ZN(n13201) );
  AOI22_X1 U16468 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13200) );
  AOI22_X1 U16469 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13199) );
  NAND4_X1 U16470 ( .A1(n13201), .A2(n13200), .A3(n13199), .A4(n13281), .ZN(
        n13212) );
  INV_X1 U16471 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13203) );
  INV_X1 U16472 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13202) );
  OAI22_X1 U16473 ( .A1(n13255), .A2(n13203), .B1(n13251), .B2(n13202), .ZN(
        n13207) );
  INV_X1 U16474 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13205) );
  INV_X1 U16475 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13204) );
  OAI22_X1 U16476 ( .A1(n13252), .A2(n13205), .B1(n13253), .B2(n13204), .ZN(
        n13206) );
  NOR2_X1 U16477 ( .A1(n13207), .A2(n13206), .ZN(n13210) );
  AOI22_X1 U16478 ( .A1(n13258), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U16479 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13208) );
  NAND4_X1 U16480 ( .A1(n13210), .A2(n13272), .A3(n13209), .A4(n13208), .ZN(
        n13211) );
  NAND2_X1 U16481 ( .A1(n13212), .A2(n13211), .ZN(n13217) );
  NOR2_X1 U16482 ( .A1(n13214), .A2(n13217), .ZN(n15150) );
  AOI211_X1 U16483 ( .C1(n13217), .C2(n13214), .A(n13213), .B(n15150), .ZN(
        n13215) );
  INV_X1 U16484 ( .A(n13217), .ZN(n13218) );
  NAND2_X1 U16485 ( .A1(n12173), .A2(n13218), .ZN(n15158) );
  OAI22_X1 U16486 ( .A1(n13255), .A2(n13220), .B1(n13251), .B2(n13219), .ZN(
        n13224) );
  OAI22_X1 U16487 ( .A1(n13252), .A2(n13222), .B1(n13253), .B2(n13221), .ZN(
        n13223) );
  NOR2_X1 U16488 ( .A1(n13224), .A2(n13223), .ZN(n13228) );
  AOI22_X1 U16489 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U16490 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13226) );
  NAND4_X1 U16491 ( .A1(n13228), .A2(n13227), .A3(n13226), .A4(n13281), .ZN(
        n13239) );
  OAI22_X1 U16492 ( .A1(n13255), .A2(n13230), .B1(n13251), .B2(n13229), .ZN(
        n13234) );
  OAI22_X1 U16493 ( .A1(n13252), .A2(n13232), .B1(n13253), .B2(n13231), .ZN(
        n13233) );
  NOR2_X1 U16494 ( .A1(n13234), .A2(n13233), .ZN(n13237) );
  AOI22_X1 U16495 ( .A1(n13258), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16496 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13235) );
  NAND4_X1 U16497 ( .A1(n13237), .A2(n13272), .A3(n13236), .A4(n13235), .ZN(
        n13238) );
  AND2_X1 U16498 ( .A1(n13239), .A2(n13238), .ZN(n15153) );
  INV_X1 U16499 ( .A(n15146), .ZN(n13267) );
  AND2_X1 U16500 ( .A1(n20060), .A2(n15153), .ZN(n13240) );
  AND2_X1 U16501 ( .A1(n15150), .A2(n13240), .ZN(n13265) );
  OAI22_X1 U16502 ( .A1(n13255), .A2(n13241), .B1(n13252), .B2(n12109), .ZN(
        n13245) );
  OAI22_X1 U16503 ( .A1(n13251), .A2(n13243), .B1(n13253), .B2(n13242), .ZN(
        n13244) );
  NOR2_X1 U16504 ( .A1(n13245), .A2(n13244), .ZN(n13249) );
  AOI22_X1 U16505 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13279), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U16506 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13247) );
  NAND4_X1 U16507 ( .A1(n13249), .A2(n13248), .A3(n13247), .A4(n13281), .ZN(
        n13263) );
  OAI22_X1 U16508 ( .A1(n12101), .A2(n13252), .B1(n13251), .B2(n13250), .ZN(
        n13257) );
  OAI22_X1 U16509 ( .A1(n13255), .A2(n13254), .B1(n13253), .B2(n12105), .ZN(
        n13256) );
  NOR2_X1 U16510 ( .A1(n13257), .A2(n13256), .ZN(n13261) );
  AOI22_X1 U16511 ( .A1(n13258), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13260) );
  AOI22_X1 U16512 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13259) );
  NAND4_X1 U16513 ( .A1(n13261), .A2(n13272), .A3(n13260), .A4(n13259), .ZN(
        n13262) );
  AND2_X1 U16514 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  NAND2_X1 U16515 ( .A1(n13265), .A2(n13264), .ZN(n13268) );
  OAI21_X1 U16516 ( .B1(n13265), .B2(n13264), .A(n13268), .ZN(n15147) );
  INV_X1 U16517 ( .A(n15147), .ZN(n13266) );
  NAND2_X1 U16518 ( .A1(n13267), .A2(n13266), .ZN(n15145) );
  NAND2_X1 U16519 ( .A1(n15145), .A2(n13268), .ZN(n13290) );
  AOI22_X1 U16520 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13269), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13271) );
  AOI22_X1 U16521 ( .A1(n13275), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13270) );
  NAND2_X1 U16522 ( .A1(n13271), .A2(n13270), .ZN(n13287) );
  AOI22_X1 U16523 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U16524 ( .A1(n11759), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13273) );
  NAND3_X1 U16525 ( .A1(n13274), .A2(n13273), .A3(n13272), .ZN(n13286) );
  AOI22_X1 U16526 ( .A1(n9805), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15772), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U16527 ( .A1(n13246), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11759), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13276) );
  NAND2_X1 U16528 ( .A1(n13277), .A2(n13276), .ZN(n13285) );
  AOI22_X1 U16529 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13278), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U16530 ( .A1(n11748), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13280), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13282) );
  NAND3_X1 U16531 ( .A1(n13283), .A2(n13282), .A3(n13281), .ZN(n13284) );
  OAI22_X1 U16532 ( .A1(n13287), .A2(n13286), .B1(n13285), .B2(n13284), .ZN(
        n13288) );
  INV_X1 U16533 ( .A(n13288), .ZN(n13289) );
  XNOR2_X1 U16534 ( .A(n13290), .B(n13289), .ZN(n14314) );
  NAND2_X1 U16535 ( .A1(n16444), .A2(n13291), .ZN(n13400) );
  NAND2_X1 U16536 ( .A1(n13400), .A2(n11865), .ZN(n13292) );
  NAND2_X1 U16537 ( .A1(n16211), .A2(n15235), .ZN(n13294) );
  NAND2_X1 U16538 ( .A1(n15221), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13293) );
  OAI21_X1 U16539 ( .B1(n14314), .B2(n15237), .A(n10348), .ZN(P2_U2857) );
  NAND2_X2 U16540 ( .A1(n18936), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18939) );
  OAI21_X1 U16541 ( .B1(n9803), .B2(n16646), .A(n19006), .ZN(n13295) );
  NAND2_X1 U16542 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19009) );
  OAI21_X1 U16543 ( .B1(n13296), .B2(n13295), .A(n19009), .ZN(n16628) );
  NOR2_X1 U16544 ( .A1(n13297), .A2(n16628), .ZN(n13304) );
  INV_X1 U16545 ( .A(n13298), .ZN(n13309) );
  OAI21_X1 U16546 ( .B1(n13309), .B2(n13300), .A(n13299), .ZN(n13302) );
  NAND2_X1 U16547 ( .A1(n13302), .A2(n13301), .ZN(n15812) );
  OAI21_X1 U16548 ( .B1(n13305), .B2(n13762), .A(n18772), .ZN(n13306) );
  NAND2_X1 U16549 ( .A1(n18776), .A2(n13310), .ZN(n16518) );
  NAND2_X1 U16550 ( .A1(n9829), .A2(n18293), .ZN(n18302) );
  NAND2_X1 U16551 ( .A1(n18776), .A2(n18293), .ZN(n18300) );
  NOR2_X1 U16552 ( .A1(n13310), .A2(n18300), .ZN(n18150) );
  NOR2_X1 U16553 ( .A1(n13312), .A2(n16507), .ZN(n13316) );
  NAND2_X1 U16554 ( .A1(n18293), .A2(n18235), .ZN(n18282) );
  AOI21_X1 U16555 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18208) );
  INV_X1 U16556 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18258) );
  NOR3_X1 U16557 ( .A1(n18258), .A2(n18251), .A3(n18246), .ZN(n18233) );
  NAND2_X1 U16558 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18233), .ZN(
        n18211) );
  NOR2_X1 U16559 ( .A1(n18210), .A2(n18211), .ZN(n18213) );
  NAND2_X1 U16560 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18213), .ZN(
        n18087) );
  NOR2_X1 U16561 ( .A1(n18208), .A2(n18087), .ZN(n18110) );
  NAND2_X1 U16562 ( .A1(n16506), .A2(n18110), .ZN(n18047) );
  OAI21_X1 U16563 ( .B1(n13313), .B2(n18047), .A(n10076), .ZN(n17987) );
  NAND2_X1 U16564 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18268) );
  NOR2_X1 U16565 ( .A1(n18087), .A2(n18268), .ZN(n18109) );
  NAND2_X1 U16566 ( .A1(n16506), .A2(n18109), .ZN(n13317) );
  INV_X1 U16567 ( .A(n13317), .ZN(n18090) );
  NAND2_X1 U16568 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18090), .ZN(
        n18111) );
  NAND2_X1 U16569 ( .A1(n13318), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16513) );
  OAI21_X1 U16570 ( .B1(n18111), .B2(n16513), .A(n18814), .ZN(n13315) );
  OAI21_X1 U16571 ( .B1(n13313), .B2(n13317), .A(n18796), .ZN(n13314) );
  NAND4_X1 U16572 ( .A1(n18236), .A2(n17987), .A3(n13315), .A4(n13314), .ZN(
        n16520) );
  NAND2_X1 U16573 ( .A1(n16515), .A2(n16520), .ZN(n15820) );
  OAI21_X1 U16574 ( .B1(n13316), .B2(n18282), .A(n15820), .ZN(n13322) );
  AOI21_X1 U16575 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18814), .A(
        n18796), .ZN(n18269) );
  OAI22_X1 U16576 ( .A1(n18809), .A2(n18047), .B1(n13317), .B2(n18269), .ZN(
        n18011) );
  NAND4_X1 U16577 ( .A1(n13319), .A2(n13318), .A3(n18293), .A4(n18011), .ZN(
        n15826) );
  NOR4_X1 U16578 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15827), .A3(
        n16507), .A4(n15826), .ZN(n13320) );
  AOI211_X1 U16579 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n13322), .A(
        n13321), .B(n13320), .ZN(n13323) );
  AOI21_X1 U16580 ( .B1(n13327), .B2(n18194), .A(n13326), .ZN(n13328) );
  INV_X1 U16581 ( .A(n13328), .ZN(P3_U2831) );
  NOR2_X1 U16582 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13330) );
  NOR4_X1 U16583 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13329) );
  NAND4_X1 U16584 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13330), .A4(n13329), .ZN(n13343) );
  NOR4_X1 U16585 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        n21289), .A4(n21130), .ZN(n13332) );
  NOR4_X1 U16586 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13331)
         );
  NAND3_X1 U16587 ( .A1(n14609), .A2(n13332), .A3(n13331), .ZN(U214) );
  NOR4_X1 U16588 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13336) );
  NOR4_X1 U16589 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13335) );
  NOR4_X1 U16590 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13334) );
  NOR4_X1 U16591 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13333) );
  NAND4_X1 U16592 ( .A1(n13336), .A2(n13335), .A3(n13334), .A4(n13333), .ZN(
        n13341) );
  NOR4_X1 U16593 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13339) );
  NOR4_X1 U16594 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13338) );
  NOR4_X1 U16595 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13337) );
  NAND4_X1 U16596 ( .A1(n13339), .A2(n13338), .A3(n13337), .A4(n19918), .ZN(
        n13340) );
  NOR2_X1 U16597 ( .A1(n19316), .A2(n13343), .ZN(n16533) );
  NAND2_X1 U16598 ( .A1(n16533), .A2(U214), .ZN(U212) );
  INV_X1 U16599 ( .A(n11874), .ZN(n13414) );
  NAND2_X1 U16600 ( .A1(n14963), .A2(n13414), .ZN(n15132) );
  INV_X1 U16601 ( .A(n15132), .ZN(n19189) );
  INV_X1 U16602 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20070) );
  INV_X1 U16603 ( .A(n13344), .ZN(n13345) );
  INV_X1 U16604 ( .A(n14955), .ZN(n13346) );
  NAND2_X1 U16605 ( .A1(n20007), .A2(n16478), .ZN(n19026) );
  OAI211_X1 U16606 ( .C1(n19189), .C2(n20070), .A(n13346), .B(n19026), .ZN(
        P2_U2814) );
  INV_X1 U16607 ( .A(n13347), .ZN(n16438) );
  NOR2_X1 U16608 ( .A1(n13495), .A2(n14952), .ZN(n13348) );
  NAND2_X1 U16609 ( .A1(n13397), .A2(n13348), .ZN(n16470) );
  AND2_X1 U16610 ( .A1(n16470), .A2(n13493), .ZN(n20038) );
  OAI21_X1 U16611 ( .B1(n13350), .B2(n20038), .A(n13349), .ZN(P2_U2819) );
  INV_X1 U16612 ( .A(n13351), .ZN(n13355) );
  INV_X1 U16613 ( .A(n20052), .ZN(n13354) );
  INV_X1 U16614 ( .A(n19026), .ZN(n13352) );
  OAI21_X1 U16615 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n13352), .A(n13354), 
        .ZN(n13353) );
  OAI21_X1 U16616 ( .B1(n13355), .B2(n13354), .A(n13353), .ZN(P2_U3612) );
  INV_X1 U16617 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13359) );
  AND2_X1 U16618 ( .A1(n14955), .A2(n20057), .ZN(n13356) );
  OR2_X1 U16619 ( .A1(n19266), .A2(n13356), .ZN(n13360) );
  AND2_X1 U16620 ( .A1(n13356), .A2(n12584), .ZN(n19261) );
  INV_X1 U16621 ( .A(n19261), .ZN(n13358) );
  AOI22_X1 U16622 ( .A1(n19318), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19316), .ZN(n14009) );
  INV_X1 U16623 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13357) );
  OAI222_X1 U16624 ( .A1(n13359), .A2(n13360), .B1(n13358), .B2(n14009), .C1(
        n13357), .C2(n13490), .ZN(P2_U2982) );
  AOI22_X1 U16625 ( .A1(n19263), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n19266), .ZN(n13361) );
  AOI22_X1 U16626 ( .A1(n19318), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19316), .ZN(n19332) );
  INV_X1 U16627 ( .A(n19332), .ZN(n14177) );
  NAND2_X1 U16628 ( .A1(n19261), .A2(n14177), .ZN(n13482) );
  NAND2_X1 U16629 ( .A1(n13361), .A2(n13482), .ZN(P2_U2953) );
  AOI22_X1 U16630 ( .A1(n19263), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n19266), .ZN(n13362) );
  OAI22_X1 U16631 ( .A1(n19316), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19318), .ZN(n19371) );
  INV_X1 U16632 ( .A(n19371), .ZN(n16265) );
  NAND2_X1 U16633 ( .A1(n19261), .A2(n16265), .ZN(n13462) );
  NAND2_X1 U16634 ( .A1(n13362), .A2(n13462), .ZN(P2_U2959) );
  AOI22_X1 U16635 ( .A1(n19263), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n19266), .ZN(n13363) );
  AOI22_X1 U16636 ( .A1(n19318), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19316), .ZN(n19342) );
  INV_X1 U16637 ( .A(n19342), .ZN(n15307) );
  NAND2_X1 U16638 ( .A1(n19261), .A2(n15307), .ZN(n13468) );
  NAND2_X1 U16639 ( .A1(n13363), .A2(n13468), .ZN(P2_U2955) );
  AOI22_X1 U16640 ( .A1(n19263), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U16641 ( .A1(n19318), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19316), .ZN(n19336) );
  INV_X1 U16642 ( .A(n19336), .ZN(n15317) );
  NAND2_X1 U16643 ( .A1(n19261), .A2(n15317), .ZN(n13466) );
  NAND2_X1 U16644 ( .A1(n13364), .A2(n13466), .ZN(P2_U2954) );
  AOI22_X1 U16645 ( .A1(n19263), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19266), .ZN(n13365) );
  AOI22_X1 U16646 ( .A1(n19318), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19316), .ZN(n13850) );
  INV_X1 U16647 ( .A(n13850), .ZN(n15248) );
  NAND2_X1 U16648 ( .A1(n19261), .A2(n15248), .ZN(n13474) );
  NAND2_X1 U16649 ( .A1(n13365), .A2(n13474), .ZN(P2_U2979) );
  AOI22_X1 U16650 ( .A1(n19263), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n19266), .ZN(n13368) );
  INV_X1 U16651 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16565) );
  OR2_X1 U16652 ( .A1(n19316), .A2(n16565), .ZN(n13367) );
  NAND2_X1 U16653 ( .A1(n19316), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13366) );
  NAND2_X1 U16654 ( .A1(n13367), .A2(n13366), .ZN(n15279) );
  NAND2_X1 U16655 ( .A1(n19261), .A2(n15279), .ZN(n13464) );
  NAND2_X1 U16656 ( .A1(n13368), .A2(n13464), .ZN(P2_U2960) );
  AOI22_X1 U16657 ( .A1(n19263), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n19266), .ZN(n13371) );
  INV_X1 U16658 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16561) );
  OR2_X1 U16659 ( .A1(n19316), .A2(n16561), .ZN(n13370) );
  NAND2_X1 U16660 ( .A1(n19316), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13369) );
  NAND2_X1 U16661 ( .A1(n13370), .A2(n13369), .ZN(n15266) );
  NAND2_X1 U16662 ( .A1(n19261), .A2(n15266), .ZN(n13476) );
  NAND2_X1 U16663 ( .A1(n13371), .A2(n13476), .ZN(P2_U2962) );
  AOI22_X1 U16664 ( .A1(n19263), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13372) );
  AOI22_X1 U16665 ( .A1(n19318), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19316), .ZN(n19323) );
  INV_X1 U16666 ( .A(n19323), .ZN(n14133) );
  NAND2_X1 U16667 ( .A1(n19261), .A2(n14133), .ZN(n13470) );
  NAND2_X1 U16668 ( .A1(n13372), .A2(n13470), .ZN(P2_U2952) );
  AOI22_X1 U16669 ( .A1(n19263), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n19266), .ZN(n13373) );
  AOI22_X1 U16670 ( .A1(n19318), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19316), .ZN(n19353) );
  INV_X1 U16671 ( .A(n19353), .ZN(n15291) );
  NAND2_X1 U16672 ( .A1(n19261), .A2(n15291), .ZN(n13472) );
  NAND2_X1 U16673 ( .A1(n13373), .A2(n13472), .ZN(P2_U2957) );
  AOI22_X1 U16674 ( .A1(n19263), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13375) );
  AOI22_X1 U16675 ( .A1(n19318), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19316), .ZN(n19359) );
  INV_X1 U16676 ( .A(n19359), .ZN(n13374) );
  NAND2_X1 U16677 ( .A1(n19261), .A2(n13374), .ZN(n13480) );
  NAND2_X1 U16678 ( .A1(n13375), .A2(n13480), .ZN(P2_U2958) );
  AOI22_X1 U16679 ( .A1(n19263), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U16680 ( .A1(n19318), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19316), .ZN(n19348) );
  INV_X1 U16681 ( .A(n19348), .ZN(n15301) );
  NAND2_X1 U16682 ( .A1(n19261), .A2(n15301), .ZN(n13478) );
  NAND2_X1 U16683 ( .A1(n13376), .A2(n13478), .ZN(P2_U2956) );
  INV_X1 U16684 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19239) );
  NAND2_X1 U16685 ( .A1(n19263), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13379) );
  INV_X1 U16686 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16563) );
  OR2_X1 U16687 ( .A1(n19316), .A2(n16563), .ZN(n13378) );
  NAND2_X1 U16688 ( .A1(n19316), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13377) );
  NAND2_X1 U16689 ( .A1(n13378), .A2(n13377), .ZN(n19212) );
  NAND2_X1 U16690 ( .A1(n19261), .A2(n19212), .ZN(n13380) );
  OAI211_X1 U16691 ( .C1(n19239), .C2(n13490), .A(n13379), .B(n13380), .ZN(
        P2_U2976) );
  INV_X1 U16692 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U16693 ( .A1(n19263), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13381) );
  OAI211_X1 U16694 ( .C1(n13434), .C2(n13490), .A(n13381), .B(n13380), .ZN(
        P2_U2961) );
  OAI21_X1 U16695 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19177), .A(
        n13392), .ZN(n13382) );
  INV_X1 U16696 ( .A(n13382), .ZN(n16421) );
  OAI21_X1 U16697 ( .B1(n13384), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13383), .ZN(n16424) );
  NAND2_X1 U16698 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(n19287), .ZN(n16422) );
  OAI21_X1 U16699 ( .B1(n19277), .B2(n16424), .A(n16422), .ZN(n13385) );
  AOI21_X1 U16700 ( .B1(n16361), .B2(n16421), .A(n13385), .ZN(n13388) );
  OAI21_X1 U16701 ( .B1(n16355), .B2(n13386), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13387) );
  OAI211_X1 U16702 ( .C1(n19317), .C2(n16418), .A(n13388), .B(n13387), .ZN(
        P2_U3014) );
  INV_X1 U16703 ( .A(n16452), .ZN(n19307) );
  OAI21_X1 U16704 ( .B1(n13390), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13389), .ZN(n19302) );
  NAND2_X1 U16705 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19287), .ZN(n19312) );
  OAI21_X1 U16706 ( .B1(n19277), .B2(n19302), .A(n19312), .ZN(n13395) );
  OAI21_X1 U16707 ( .B1(n13392), .B2(n15135), .A(n13391), .ZN(n13393) );
  XNOR2_X1 U16708 ( .A(n13393), .B(n15783), .ZN(n19315) );
  OAI22_X1 U16709 ( .A1(n19315), .A2(n19278), .B1(n16366), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13394) );
  AOI211_X1 U16710 ( .C1(n16355), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13395), .B(n13394), .ZN(n13396) );
  OAI21_X1 U16711 ( .B1(n19307), .B2(n19317), .A(n13396), .ZN(P2_U3013) );
  OR2_X1 U16712 ( .A1(n16444), .A2(n15770), .ZN(n13492) );
  NAND2_X1 U16713 ( .A1(n13397), .A2(n13495), .ZN(n13399) );
  AND2_X1 U16714 ( .A1(n13399), .A2(n13398), .ZN(n13401) );
  AND3_X1 U16715 ( .A1(n13492), .A2(n13401), .A3(n13400), .ZN(n13406) );
  INV_X1 U16716 ( .A(n13416), .ZN(n13404) );
  NOR2_X1 U16717 ( .A1(n11874), .A2(n13402), .ZN(n13403) );
  NAND2_X1 U16718 ( .A1(n13404), .A2(n13403), .ZN(n13405) );
  NAND2_X1 U16719 ( .A1(n13406), .A2(n13405), .ZN(n16474) );
  NAND2_X1 U16720 ( .A1(n16474), .A2(n13493), .ZN(n13408) );
  NAND2_X1 U16721 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16485), .ZN(n16497) );
  INV_X1 U16722 ( .A(n16497), .ZN(n15905) );
  AOI22_X1 U16723 ( .A1(n15905), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n20054), .ZN(n13407) );
  NAND2_X1 U16724 ( .A1(n13408), .A2(n13407), .ZN(n19999) );
  INV_X1 U16725 ( .A(n15785), .ZN(n20004) );
  AND2_X1 U16726 ( .A1(n13410), .A2(n13409), .ZN(n13411) );
  NAND2_X1 U16727 ( .A1(n13412), .A2(n13411), .ZN(n16462) );
  OR3_X1 U16728 ( .A1(n19996), .A2(n20004), .A3(n16462), .ZN(n13413) );
  OAI21_X1 U16729 ( .B1(n16473), .B2(n19999), .A(n13413), .ZN(P2_U3595) );
  INV_X1 U16730 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13420) );
  NAND2_X1 U16731 ( .A1(n13414), .A2(n13493), .ZN(n13415) );
  NAND2_X1 U16732 ( .A1(n16485), .A2(n20054), .ZN(n13418) );
  INV_X2 U16733 ( .A(n13418), .ZN(n19227) );
  AOI22_X1 U16734 ( .A1(n19227), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13419) );
  OAI21_X1 U16735 ( .B1(n13420), .B2(n19219), .A(n13419), .ZN(P2_U2931) );
  INV_X1 U16736 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13422) );
  AOI22_X1 U16737 ( .A1(n19227), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13421) );
  OAI21_X1 U16738 ( .B1(n13422), .B2(n19219), .A(n13421), .ZN(P2_U2928) );
  AOI22_X1 U16739 ( .A1(n19227), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13423) );
  OAI21_X1 U16740 ( .B1(n15319), .B2(n19219), .A(n13423), .ZN(P2_U2933) );
  INV_X1 U16741 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U16742 ( .A1(n19227), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13424) );
  OAI21_X1 U16743 ( .B1(n13425), .B2(n19219), .A(n13424), .ZN(P2_U2932) );
  AOI22_X1 U16744 ( .A1(n19227), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13426) );
  OAI21_X1 U16745 ( .B1(n13427), .B2(n19219), .A(n13426), .ZN(P2_U2935) );
  INV_X1 U16746 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14179) );
  AOI22_X1 U16747 ( .A1(n19227), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13428) );
  OAI21_X1 U16748 ( .B1(n14179), .B2(n19219), .A(n13428), .ZN(P2_U2934) );
  AOI22_X1 U16749 ( .A1(n19227), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13429) );
  OAI21_X1 U16750 ( .B1(n15285), .B2(n19219), .A(n13429), .ZN(P2_U2929) );
  INV_X1 U16751 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U16752 ( .A1(n19227), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13430) );
  OAI21_X1 U16753 ( .B1(n13431), .B2(n19219), .A(n13430), .ZN(P2_U2930) );
  INV_X1 U16754 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15263) );
  AOI22_X1 U16755 ( .A1(n19227), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13432) );
  OAI21_X1 U16756 ( .B1(n15263), .B2(n19219), .A(n13432), .ZN(P2_U2925) );
  AOI22_X1 U16757 ( .A1(n19227), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13433) );
  OAI21_X1 U16758 ( .B1(n13434), .B2(n19219), .A(n13433), .ZN(P2_U2926) );
  INV_X1 U16759 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15277) );
  AOI22_X1 U16760 ( .A1(n19227), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13435) );
  OAI21_X1 U16761 ( .B1(n15277), .B2(n19219), .A(n13435), .ZN(P2_U2927) );
  INV_X1 U16762 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U16763 ( .A1(n19227), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13436) );
  OAI21_X1 U16764 ( .B1(n13487), .B2(n19219), .A(n13436), .ZN(P2_U2924) );
  INV_X1 U16765 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U16766 ( .A1(n19227), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13437) );
  OAI21_X1 U16767 ( .B1(n13438), .B2(n19219), .A(n13437), .ZN(P2_U2923) );
  AOI21_X1 U16768 ( .B1(n15136), .B2(n15126), .A(n14021), .ZN(n15121) );
  XNOR2_X1 U16769 ( .A(n13440), .B(n13439), .ZN(n13543) );
  INV_X1 U16770 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19917) );
  NAND2_X1 U16771 ( .A1(n19287), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U16772 ( .A1(n16355), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13441) );
  OAI211_X1 U16773 ( .C1(n13543), .C2(n19277), .A(n13539), .B(n13441), .ZN(
        n13445) );
  NAND2_X1 U16774 ( .A1(n13443), .A2(n13442), .ZN(n13540) );
  AND3_X1 U16775 ( .A1(n13541), .A2(n16361), .A3(n13540), .ZN(n13444) );
  AOI211_X1 U16776 ( .C1(n19270), .C2(n15121), .A(n13445), .B(n13444), .ZN(
        n13446) );
  OAI21_X1 U16777 ( .B1(n13549), .B2(n19317), .A(n13446), .ZN(P2_U3012) );
  INV_X1 U16778 ( .A(n13447), .ZN(n13448) );
  INV_X1 U16779 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21302) );
  NAND2_X1 U16780 ( .A1(n20698), .A2(n20834), .ZN(n20077) );
  OAI211_X1 U16781 ( .C1(n13448), .C2(n21302), .A(n13651), .B(n20077), .ZN(
        P1_U2801) );
  NAND2_X1 U16782 ( .A1(n13597), .A2(n13449), .ZN(n13450) );
  NAND2_X1 U16783 ( .A1(n12641), .A2(n13450), .ZN(n13452) );
  NAND2_X1 U16784 ( .A1(n13686), .A2(n14035), .ZN(n13451) );
  NAND2_X1 U16785 ( .A1(n13452), .A2(n13451), .ZN(n20075) );
  NAND2_X1 U16786 ( .A1(n13453), .A2(n20940), .ZN(n20929) );
  INV_X1 U16787 ( .A(n14028), .ZN(n20934) );
  OAI21_X1 U16788 ( .B1(n20929), .B2(n20934), .A(n13587), .ZN(n13454) );
  NOR2_X1 U16789 ( .A1(n20075), .A2(n13454), .ZN(n15857) );
  OR2_X1 U16790 ( .A1(n15857), .A2(n20074), .ZN(n13459) );
  INV_X1 U16791 ( .A(n13459), .ZN(n20081) );
  INV_X1 U16792 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13461) );
  NAND3_X1 U16793 ( .A1(n12641), .A2(n15859), .A3(n13693), .ZN(n13455) );
  NAND2_X1 U16794 ( .A1(n13455), .A2(n13686), .ZN(n13458) );
  AOI22_X1 U16795 ( .A1(n13678), .A2(n13696), .B1(n13597), .B2(n13456), .ZN(
        n13457) );
  AND2_X1 U16796 ( .A1(n13458), .A2(n13457), .ZN(n15860) );
  OR2_X1 U16797 ( .A1(n13459), .A2(n15860), .ZN(n13460) );
  OAI21_X1 U16798 ( .B1(n20081), .B2(n13461), .A(n13460), .ZN(P1_U3484) );
  AOI22_X1 U16799 ( .A1(n19263), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13463) );
  NAND2_X1 U16800 ( .A1(n13463), .A2(n13462), .ZN(P2_U2974) );
  AOI22_X1 U16801 ( .A1(n19263), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13465) );
  NAND2_X1 U16802 ( .A1(n13465), .A2(n13464), .ZN(P2_U2975) );
  AOI22_X1 U16803 ( .A1(n19263), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13467) );
  NAND2_X1 U16804 ( .A1(n13467), .A2(n13466), .ZN(P2_U2969) );
  AOI22_X1 U16805 ( .A1(n19263), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U16806 ( .A1(n13469), .A2(n13468), .ZN(P2_U2970) );
  AOI22_X1 U16807 ( .A1(n19263), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13471) );
  NAND2_X1 U16808 ( .A1(n13471), .A2(n13470), .ZN(P2_U2967) );
  AOI22_X1 U16809 ( .A1(n19263), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13473) );
  NAND2_X1 U16810 ( .A1(n13473), .A2(n13472), .ZN(P2_U2972) );
  AOI22_X1 U16811 ( .A1(n19263), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19266), .ZN(n13475) );
  NAND2_X1 U16812 ( .A1(n13475), .A2(n13474), .ZN(P2_U2964) );
  AOI22_X1 U16813 ( .A1(n19263), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n19266), .ZN(n13477) );
  NAND2_X1 U16814 ( .A1(n13477), .A2(n13476), .ZN(P2_U2977) );
  AOI22_X1 U16815 ( .A1(n19263), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13479) );
  NAND2_X1 U16816 ( .A1(n13479), .A2(n13478), .ZN(P2_U2971) );
  AOI22_X1 U16817 ( .A1(n19263), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13481) );
  NAND2_X1 U16818 ( .A1(n13481), .A2(n13480), .ZN(P2_U2973) );
  AOI22_X1 U16819 ( .A1(n19263), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13483) );
  NAND2_X1 U16820 ( .A1(n13483), .A2(n13482), .ZN(P2_U2968) );
  NAND2_X1 U16821 ( .A1(n19263), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13486) );
  INV_X1 U16822 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16559) );
  OR2_X1 U16823 ( .A1(n19316), .A2(n16559), .ZN(n13485) );
  NAND2_X1 U16824 ( .A1(n19316), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13484) );
  NAND2_X1 U16825 ( .A1(n13485), .A2(n13484), .ZN(n19209) );
  NAND2_X1 U16826 ( .A1(n19261), .A2(n19209), .ZN(n13488) );
  OAI211_X1 U16827 ( .C1(n13487), .C2(n13490), .A(n13486), .B(n13488), .ZN(
        P2_U2963) );
  INV_X1 U16828 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19235) );
  NAND2_X1 U16829 ( .A1(n19263), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13489) );
  OAI211_X1 U16830 ( .C1(n19235), .C2(n13490), .A(n13489), .B(n13488), .ZN(
        P2_U2978) );
  INV_X1 U16831 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n13505) );
  NAND2_X1 U16832 ( .A1(n13492), .A2(n13491), .ZN(n13494) );
  NAND2_X1 U16833 ( .A1(n13494), .A2(n13493), .ZN(n13497) );
  NAND2_X1 U16834 ( .A1(n20052), .A2(n13495), .ZN(n13496) );
  INV_X1 U16835 ( .A(n13498), .ZN(n13499) );
  NOR2_X1 U16836 ( .A1(n13501), .A2(n13500), .ZN(n13502) );
  OR2_X1 U16837 ( .A1(n13503), .A2(n13502), .ZN(n19158) );
  OAI222_X1 U16838 ( .A1(n13505), .A2(n19217), .B1(n14010), .B2(n19359), .C1(
        n19158), .C2(n19206), .ZN(P2_U2913) );
  NAND2_X1 U16839 ( .A1(n13508), .A2(n13507), .ZN(n13509) );
  MUX2_X1 U16840 ( .A(n15139), .B(n19307), .S(n15235), .Z(n13510) );
  OAI21_X1 U16841 ( .B1(n19994), .B2(n15237), .A(n13510), .ZN(P2_U2886) );
  INV_X1 U16842 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13512) );
  AND2_X1 U16843 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12958), .ZN(n13511) );
  OAI211_X1 U16844 ( .C1(n12173), .C2(n13512), .A(n12957), .B(n13511), .ZN(
        n13513) );
  INV_X1 U16845 ( .A(n13513), .ZN(n13514) );
  AOI21_X1 U16846 ( .B1(n20031), .B2(n16268), .A(n19198), .ZN(n13523) );
  OR2_X1 U16847 ( .A1(n13516), .A2(n13515), .ZN(n13517) );
  NAND2_X1 U16848 ( .A1(n13518), .A2(n13517), .ZN(n19178) );
  NOR2_X1 U16849 ( .A1(n14010), .A2(n19323), .ZN(n13521) );
  INV_X1 U16850 ( .A(n19178), .ZN(n13519) );
  NOR3_X1 U16851 ( .A1(n20031), .A2(n13519), .A3(n15327), .ZN(n13520) );
  AOI211_X1 U16852 ( .C1(P2_EAX_REG_0__SCAN_IN), .C2(n19203), .A(n13521), .B(
        n13520), .ZN(n13522) );
  OAI21_X1 U16853 ( .B1(n13523), .B2(n19178), .A(n13522), .ZN(P2_U2919) );
  AOI21_X1 U16854 ( .B1(n13526), .B2(n13525), .A(n13524), .ZN(n13527) );
  INV_X1 U16855 ( .A(n13527), .ZN(n13548) );
  INV_X1 U16856 ( .A(n13528), .ZN(n19311) );
  AOI21_X1 U16857 ( .B1(n13529), .B2(n19304), .A(n19311), .ZN(n13532) );
  OAI22_X1 U16858 ( .A1(n13532), .A2(n13531), .B1(n19304), .B2(n13530), .ZN(
        n13546) );
  INV_X1 U16859 ( .A(n13533), .ZN(n13536) );
  INV_X1 U16860 ( .A(n13534), .ZN(n13535) );
  NAND2_X1 U16861 ( .A1(n13536), .A2(n13535), .ZN(n13538) );
  OAI21_X1 U16862 ( .B1(n19301), .B2(n15127), .A(n13539), .ZN(n13545) );
  NAND3_X1 U16863 ( .A1(n13541), .A2(n19296), .A3(n13540), .ZN(n13542) );
  OAI21_X1 U16864 ( .B1(n13543), .B2(n19303), .A(n13542), .ZN(n13544) );
  NOR3_X1 U16865 ( .A1(n13546), .A2(n13545), .A3(n13544), .ZN(n13547) );
  OAI211_X1 U16866 ( .C1(n19308), .C2(n13549), .A(n13548), .B(n13547), .ZN(
        P2_U3044) );
  NAND2_X1 U16867 ( .A1(n19586), .A2(n15224), .ZN(n13551) );
  NAND2_X1 U16868 ( .A1(n12974), .A2(n15235), .ZN(n13550) );
  OAI211_X1 U16869 ( .C1(n15235), .C2(n13552), .A(n13551), .B(n13550), .ZN(
        P2_U2887) );
  INV_X1 U16870 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n13556) );
  AOI21_X1 U16871 ( .B1(n13554), .B2(n13553), .A(n9889), .ZN(n13555) );
  INV_X1 U16872 ( .A(n13555), .ZN(n15720) );
  OAI222_X1 U16873 ( .A1(n13556), .A2(n19217), .B1(n14010), .B2(n19371), .C1(
        n15720), .C2(n19206), .ZN(P2_U2912) );
  INV_X1 U16874 ( .A(n15279), .ZN(n13558) );
  OAI21_X1 U16875 ( .B1(n13557), .B2(n9889), .A(n15079), .ZN(n19146) );
  INV_X1 U16876 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19241) );
  OAI222_X1 U16877 ( .A1(n14010), .A2(n13558), .B1(n19146), .B2(n19206), .C1(
        n19217), .C2(n19241), .ZN(P2_U2911) );
  NAND2_X1 U16878 ( .A1(n13597), .A2(n20274), .ZN(n13948) );
  OAI21_X1 U16879 ( .B1(n10458), .B2(n14028), .A(n13560), .ZN(n13561) );
  AOI21_X1 U16880 ( .B1(n13563), .B2(n13562), .A(n13561), .ZN(n13570) );
  OR2_X1 U16881 ( .A1(n13564), .A2(n13939), .ZN(n13565) );
  NAND2_X1 U16882 ( .A1(n11230), .A2(n10469), .ZN(n13684) );
  NAND2_X1 U16883 ( .A1(n13568), .A2(n13567), .ZN(n13598) );
  NAND4_X1 U16884 ( .A1(n13571), .A2(n13570), .A3(n13569), .A4(n13598), .ZN(
        n13702) );
  INV_X1 U16885 ( .A(n13702), .ZN(n13577) );
  INV_X1 U16886 ( .A(n13698), .ZN(n13574) );
  NAND2_X1 U16887 ( .A1(n13574), .A2(n13573), .ZN(n13575) );
  NOR2_X1 U16888 ( .A1(n13572), .A2(n13575), .ZN(n13576) );
  NAND3_X1 U16889 ( .A1(n13577), .A2(n13576), .A3(n12643), .ZN(n13935) );
  NAND2_X1 U16890 ( .A1(n20731), .A2(n13935), .ZN(n13582) );
  INV_X1 U16891 ( .A(n13578), .ZN(n13579) );
  INV_X1 U16892 ( .A(n13612), .ZN(n13611) );
  NAND3_X1 U16893 ( .A1(n13580), .A2(n13579), .A3(n13611), .ZN(n13581) );
  OAI211_X1 U16894 ( .C1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n13948), .A(
        n13582), .B(n13581), .ZN(n15847) );
  INV_X1 U16895 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13583) );
  AOI22_X1 U16896 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n12679), .B2(n13583), .ZN(
        n13620) );
  INV_X1 U16897 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20265) );
  NOR2_X1 U16898 ( .A1(n20834), .A2(n20265), .ZN(n13621) );
  INV_X1 U16899 ( .A(n13621), .ZN(n13584) );
  NOR2_X1 U16900 ( .A1(n13620), .A2(n13584), .ZN(n13586) );
  INV_X1 U16901 ( .A(n20905), .ZN(n15875) );
  NOR3_X1 U16902 ( .A1(n13578), .A2(n13612), .A3(n15875), .ZN(n13585) );
  AOI211_X1 U16903 ( .C1(n15847), .C2(n20906), .A(n13586), .B(n13585), .ZN(
        n13607) );
  NAND2_X1 U16904 ( .A1(n13588), .A2(n13587), .ZN(n13591) );
  INV_X1 U16905 ( .A(n13572), .ZN(n13589) );
  NAND2_X1 U16906 ( .A1(n13948), .A2(n13589), .ZN(n13590) );
  INV_X1 U16907 ( .A(n13693), .ZN(n13610) );
  AOI21_X1 U16908 ( .B1(n13591), .B2(n13590), .A(n13610), .ZN(n13592) );
  OR2_X1 U16909 ( .A1(n13592), .A2(n13686), .ZN(n13602) );
  OAI21_X1 U16910 ( .B1(n14028), .B2(n20281), .A(n13593), .ZN(n13594) );
  OR2_X1 U16911 ( .A1(n13595), .A2(n13594), .ZN(n13600) );
  OR2_X1 U16912 ( .A1(n13597), .A2(n13596), .ZN(n13599) );
  NAND2_X1 U16913 ( .A1(n13599), .A2(n13598), .ZN(n13683) );
  NOR2_X1 U16914 ( .A1(n13600), .A2(n13683), .ZN(n13601) );
  NAND2_X1 U16915 ( .A1(n15846), .A2(n13690), .ZN(n13605) );
  INV_X1 U16916 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21151) );
  NAND2_X1 U16917 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n16190) );
  OR2_X1 U16918 ( .A1(n20936), .A2(n16190), .ZN(n16195) );
  NOR2_X1 U16919 ( .A1(n21151), .A2(n16195), .ZN(n13603) );
  NOR2_X1 U16920 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20661), .ZN(n16194) );
  NOR2_X1 U16921 ( .A1(n13603), .A2(n16194), .ZN(n13604) );
  NAND2_X1 U16922 ( .A1(n20909), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13606) );
  OAI21_X1 U16923 ( .B1(n13607), .B2(n20909), .A(n13606), .ZN(P1_U3473) );
  INV_X1 U16924 ( .A(n13948), .ZN(n13616) );
  XNOR2_X1 U16925 ( .A(n13940), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13615) );
  NOR2_X1 U16926 ( .A1(n13610), .A2(n13696), .ZN(n13946) );
  INV_X1 U16927 ( .A(n13946), .ZN(n13614) );
  NAND2_X1 U16928 ( .A1(n13611), .A2(n10009), .ZN(n13944) );
  NAND2_X1 U16929 ( .A1(n13612), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13936) );
  AND2_X1 U16930 ( .A1(n13944), .A2(n13936), .ZN(n13619) );
  INV_X1 U16931 ( .A(n13619), .ZN(n13613) );
  AOI22_X1 U16932 ( .A1(n13616), .A2(n13615), .B1(n13614), .B2(n13613), .ZN(
        n13618) );
  NAND3_X1 U16933 ( .A1(n13951), .A2(n13939), .A3(n13619), .ZN(n13617) );
  OAI211_X1 U16934 ( .C1(n13609), .C2(n13951), .A(n13618), .B(n13617), .ZN(
        n13934) );
  AOI222_X1 U16935 ( .A1(n13934), .A2(n20906), .B1(n13621), .B2(n13620), .C1(
        n20905), .C2(n13619), .ZN(n13623) );
  NAND2_X1 U16936 ( .A1(n20909), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13622) );
  OAI21_X1 U16937 ( .B1(n13623), .B2(n20909), .A(n13622), .ZN(P1_U3472) );
  INV_X1 U16938 ( .A(n10591), .ZN(n13987) );
  OAI22_X1 U16939 ( .A1(n13987), .A2(n13951), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13624), .ZN(n15845) );
  OAI22_X1 U16940 ( .A1(n20834), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15875), .ZN(n13625) );
  AOI21_X1 U16941 ( .B1(n15845), .B2(n20906), .A(n13625), .ZN(n13627) );
  NOR2_X1 U16942 ( .A1(n13948), .A2(n10323), .ZN(n15844) );
  AOI22_X1 U16943 ( .A1(n20909), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20906), .B2(n15844), .ZN(n13626) );
  OAI21_X1 U16944 ( .B1(n13627), .B2(n20909), .A(n13626), .ZN(P1_U3474) );
  OAI21_X4 U16945 ( .B1(n13629), .B2(n20940), .A(n13628), .ZN(n20223) );
  INV_X1 U16946 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21292) );
  INV_X1 U16947 ( .A(DATAI_14_), .ZN(n21059) );
  NAND2_X1 U16948 ( .A1(n14607), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13631) );
  OAI21_X1 U16949 ( .B1(n14609), .B2(n21059), .A(n13631), .ZN(n20247) );
  AOI22_X1 U16950 ( .A1(n20248), .A2(n20247), .B1(n20223), .B2(
        P1_UWORD_REG_14__SCAN_IN), .ZN(n13632) );
  OAI21_X1 U16951 ( .B1(n20212), .B2(n21292), .A(n13632), .ZN(P1_U2951) );
  INV_X1 U16952 ( .A(DATAI_12_), .ZN(n21057) );
  NAND2_X1 U16953 ( .A1(n14607), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13633) );
  OAI21_X1 U16954 ( .B1(n14609), .B2(n21057), .A(n13633), .ZN(n20241) );
  AOI22_X1 U16955 ( .A1(n20248), .A2(n20241), .B1(n20223), .B2(
        P1_UWORD_REG_12__SCAN_IN), .ZN(n13634) );
  OAI21_X1 U16956 ( .B1(n20212), .B2(n11076), .A(n13634), .ZN(P1_U2949) );
  INV_X1 U16957 ( .A(n20909), .ZN(n13640) );
  INV_X1 U16958 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13639) );
  INV_X1 U16959 ( .A(n20411), .ZN(n20652) );
  OR2_X1 U16960 ( .A1(n13635), .A2(n20652), .ZN(n13636) );
  XNOR2_X1 U16961 ( .A(n13636), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20145) );
  INV_X1 U16962 ( .A(n12643), .ZN(n13637) );
  NAND4_X1 U16963 ( .A1(n20145), .A2(n20906), .A3(n13637), .A4(n13640), .ZN(
        n13638) );
  OAI21_X1 U16964 ( .B1(n13640), .B2(n13639), .A(n13638), .ZN(P1_U3468) );
  NOR2_X1 U16965 ( .A1(n20031), .A2(n19178), .ZN(n13646) );
  NAND2_X1 U16966 ( .A1(n13642), .A2(n13641), .ZN(n13643) );
  NAND2_X1 U16967 ( .A1(n13644), .A2(n13643), .ZN(n20026) );
  INV_X1 U16968 ( .A(n20026), .ZN(n19300) );
  NAND2_X1 U16969 ( .A1(n19994), .A2(n19300), .ZN(n13819) );
  OAI21_X1 U16970 ( .B1(n19994), .B2(n19300), .A(n13819), .ZN(n13645) );
  NOR2_X1 U16971 ( .A1(n13645), .A2(n13646), .ZN(n13821) );
  AOI21_X1 U16972 ( .B1(n13646), .B2(n13645), .A(n13821), .ZN(n13649) );
  AOI22_X1 U16973 ( .A1(n19198), .A2(n20026), .B1(n19203), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13648) );
  NAND2_X1 U16974 ( .A1(n19213), .A2(n14177), .ZN(n13647) );
  OAI211_X1 U16975 ( .C1(n13649), .C2(n15327), .A(n13648), .B(n13647), .ZN(
        P2_U2918) );
  OAI22_X1 U16976 ( .A1(n13651), .A2(n20274), .B1(n13948), .B2(n13650), .ZN(
        n13653) );
  INV_X1 U16977 ( .A(n20933), .ZN(n13652) );
  NOR2_X1 U16978 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16190), .ZN(n13869) );
  NOR2_X4 U16979 ( .A1(n20180), .A2(n20941), .ZN(n20195) );
  AOI22_X1 U16980 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20195), .B1(n13869), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13654) );
  OAI21_X1 U16981 ( .B1(n21292), .B2(n13880), .A(n13654), .ZN(P1_U2906) );
  AOI22_X1 U16982 ( .A1(n13869), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13655) );
  OAI21_X1 U16983 ( .B1(n10976), .B2(n13880), .A(n13655), .ZN(P1_U2913) );
  AOI22_X1 U16984 ( .A1(n13869), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13656) );
  OAI21_X1 U16985 ( .B1(n10995), .B2(n13880), .A(n13656), .ZN(P1_U2912) );
  AOI22_X1 U16986 ( .A1(n13869), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13657) );
  OAI21_X1 U16987 ( .B1(n11076), .B2(n13880), .A(n13657), .ZN(P1_U2908) );
  AOI22_X1 U16988 ( .A1(n13869), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13658) );
  OAI21_X1 U16989 ( .B1(n11100), .B2(n13880), .A(n13658), .ZN(P1_U2907) );
  AOI22_X1 U16990 ( .A1(n13869), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13659) );
  OAI21_X1 U16991 ( .B1(n11017), .B2(n13880), .A(n13659), .ZN(P1_U2911) );
  XNOR2_X1 U16992 ( .A(n13660), .B(n9888), .ZN(n16399) );
  AOI22_X1 U16993 ( .A1(n19213), .A2(n15266), .B1(n19203), .B2(
        P2_EAX_REG_10__SCAN_IN), .ZN(n13661) );
  OAI21_X1 U16994 ( .B1(n19206), .B2(n16399), .A(n13661), .ZN(P2_U2909) );
  MUX2_X1 U16995 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n15764), .S(n15235), .Z(
        n13666) );
  AOI21_X1 U16996 ( .B1(n19466), .B2(n15224), .A(n13666), .ZN(n13667) );
  INV_X1 U16997 ( .A(n13667), .ZN(P2_U2885) );
  INV_X1 U16998 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20197) );
  INV_X1 U16999 ( .A(DATAI_8_), .ZN(n21172) );
  NAND2_X1 U17000 ( .A1(n14607), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13668) );
  OAI21_X1 U17001 ( .B1(n14609), .B2(n21172), .A(n13668), .ZN(n14564) );
  NAND2_X1 U17002 ( .A1(n20248), .A2(n14564), .ZN(n13670) );
  NAND2_X1 U17003 ( .A1(n20223), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13669) );
  OAI211_X1 U17004 ( .C1(n20212), .C2(n20197), .A(n13670), .B(n13669), .ZN(
        P1_U2960) );
  NAND2_X1 U17005 ( .A1(n20223), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13671) );
  OAI211_X1 U17006 ( .C1(n20212), .C2(n10995), .A(n13671), .B(n13670), .ZN(
        P1_U2945) );
  XNOR2_X1 U17007 ( .A(n13672), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13747) );
  NAND2_X1 U17008 ( .A1(n20274), .A2(n20933), .ZN(n13675) );
  INV_X1 U17009 ( .A(n13673), .ZN(n13674) );
  NAND2_X1 U17010 ( .A1(n13675), .A2(n13674), .ZN(n13682) );
  NAND2_X1 U17011 ( .A1(n13572), .A2(n13676), .ZN(n13677) );
  NAND2_X1 U17012 ( .A1(n13679), .A2(n13678), .ZN(n13681) );
  MUX2_X1 U17013 ( .A(n13682), .B(n13681), .S(n13680), .Z(n13689) );
  INV_X1 U17014 ( .A(n13683), .ZN(n13688) );
  INV_X1 U17015 ( .A(n13684), .ZN(n13685) );
  NAND2_X1 U17016 ( .A1(n13686), .A2(n13685), .ZN(n13687) );
  NAND3_X1 U17017 ( .A1(n13689), .A2(n13688), .A3(n13687), .ZN(n13691) );
  OAI211_X1 U17018 ( .C1(n14162), .C2(n13705), .A(n15859), .B(n13693), .ZN(
        n13694) );
  NOR2_X1 U17019 ( .A1(n13692), .A2(n13694), .ZN(n13695) );
  NAND2_X1 U17020 ( .A1(n13714), .A2(n16162), .ZN(n20263) );
  INV_X1 U17021 ( .A(n13696), .ZN(n13697) );
  NAND2_X1 U17022 ( .A1(n13698), .A2(n20266), .ZN(n13700) );
  NAND2_X1 U17023 ( .A1(n13700), .A2(n13699), .ZN(n13701) );
  NOR2_X1 U17024 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  NAND2_X1 U17025 ( .A1(n15888), .A2(n16070), .ZN(n13713) );
  NAND2_X1 U17026 ( .A1(n20265), .A2(n13713), .ZN(n20256) );
  AOI21_X1 U17027 ( .B1(n20263), .B2(n20256), .A(n12679), .ZN(n13704) );
  INV_X1 U17028 ( .A(n13704), .ZN(n13718) );
  OAI22_X1 U17029 ( .A1(n12641), .A2(n20274), .B1(n13706), .B2(n13705), .ZN(
        n13707) );
  INV_X1 U17030 ( .A(n13707), .ZN(n13708) );
  OR2_X1 U17031 ( .A1(n13710), .A2(n13709), .ZN(n13711) );
  NAND2_X1 U17032 ( .A1(n13712), .A2(n13711), .ZN(n14047) );
  INV_X1 U17033 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21275) );
  NOR2_X1 U17034 ( .A1(n16162), .A2(n21275), .ZN(n13743) );
  INV_X1 U17035 ( .A(n13713), .ZN(n13715) );
  NAND2_X1 U17036 ( .A1(n20265), .A2(n20264), .ZN(n13750) );
  AND3_X1 U17037 ( .A1(n16160), .A2(n13750), .A3(n12679), .ZN(n13716) );
  AOI211_X1 U17038 ( .C1(n16173), .C2(n14047), .A(n13743), .B(n13716), .ZN(
        n13717) );
  OAI211_X1 U17039 ( .C1(n13747), .C2(n16182), .A(n13718), .B(n13717), .ZN(
        P1_U3030) );
  INV_X1 U17040 ( .A(n13719), .ZN(n13722) );
  OAI21_X1 U17041 ( .B1(n13722), .B2(n13721), .A(n13720), .ZN(n14038) );
  OR2_X1 U17042 ( .A1(n13723), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13724) );
  AND2_X1 U17043 ( .A1(n13725), .A2(n13724), .ZN(n20261) );
  OAI21_X1 U17044 ( .B1(n16015), .B2(n13726), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13728) );
  INV_X1 U17045 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13727) );
  OR2_X1 U17046 ( .A1(n16162), .A2(n13727), .ZN(n20255) );
  NAND2_X1 U17047 ( .A1(n13728), .A2(n20255), .ZN(n13729) );
  AOI21_X1 U17048 ( .B1(n20261), .B2(n11296), .A(n13729), .ZN(n13730) );
  OAI21_X1 U17049 ( .B1(n14038), .B2(n13814), .A(n13730), .ZN(P1_U2999) );
  INV_X1 U17050 ( .A(DATAI_13_), .ZN(n13732) );
  NAND2_X1 U17051 ( .A1(n14607), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13731) );
  OAI21_X1 U17052 ( .B1(n14609), .B2(n13732), .A(n13731), .ZN(n20244) );
  AOI22_X1 U17053 ( .A1(n20248), .A2(n20244), .B1(n20223), .B2(
        P1_UWORD_REG_13__SCAN_IN), .ZN(n13733) );
  OAI21_X1 U17054 ( .B1(n20212), .B2(n11100), .A(n13733), .ZN(P1_U2950) );
  INV_X1 U17055 ( .A(DATAI_9_), .ZN(n13735) );
  NAND2_X1 U17056 ( .A1(n14607), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13734) );
  OAI21_X1 U17057 ( .B1(n14609), .B2(n13735), .A(n13734), .ZN(n20232) );
  AOI22_X1 U17058 ( .A1(n20248), .A2(n20232), .B1(n20223), .B2(
        P1_UWORD_REG_9__SCAN_IN), .ZN(n13736) );
  OAI21_X1 U17059 ( .B1(n20212), .B2(n11017), .A(n13736), .ZN(P1_U2946) );
  INV_X1 U17060 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n21105) );
  INV_X1 U17061 ( .A(DATAI_11_), .ZN(n21052) );
  NAND2_X1 U17062 ( .A1(n14607), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13737) );
  OAI21_X1 U17063 ( .B1(n14609), .B2(n21052), .A(n13737), .ZN(n20238) );
  AOI22_X1 U17064 ( .A1(n20248), .A2(n20238), .B1(n20223), .B2(
        P1_UWORD_REG_11__SCAN_IN), .ZN(n13738) );
  OAI21_X1 U17065 ( .B1(n20212), .B2(n21105), .A(n13738), .ZN(P1_U2948) );
  INV_X1 U17066 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21258) );
  INV_X1 U17067 ( .A(DATAI_10_), .ZN(n21253) );
  NAND2_X1 U17068 ( .A1(n14607), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13739) );
  OAI21_X1 U17069 ( .B1(n14609), .B2(n21253), .A(n13739), .ZN(n20235) );
  AOI22_X1 U17070 ( .A1(n20248), .A2(n20235), .B1(n20223), .B2(
        P1_UWORD_REG_10__SCAN_IN), .ZN(n13740) );
  OAI21_X1 U17071 ( .B1(n20212), .B2(n21258), .A(n13740), .ZN(P1_U2947) );
  OAI21_X1 U17072 ( .B1(n13742), .B2(n13741), .A(n13812), .ZN(n14054) );
  INV_X1 U17073 ( .A(n14054), .ZN(n13992) );
  AOI21_X1 U17074 ( .B1(n16015), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13743), .ZN(n13744) );
  OAI21_X1 U17075 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16022), .A(
        n13744), .ZN(n13745) );
  AOI21_X1 U17076 ( .B1(n13992), .B2(n16025), .A(n13745), .ZN(n13746) );
  OAI21_X1 U17077 ( .B1(n13747), .B2(n20080), .A(n13746), .ZN(P1_U2998) );
  XNOR2_X1 U17078 ( .A(n13749), .B(n13748), .ZN(n13818) );
  NAND2_X1 U17079 ( .A1(n16070), .A2(n20264), .ZN(n15891) );
  NAND2_X1 U17080 ( .A1(n15891), .A2(n13750), .ZN(n14896) );
  NOR2_X1 U17081 ( .A1(n12679), .A2(n14896), .ZN(n13759) );
  INV_X1 U17082 ( .A(n15891), .ZN(n16158) );
  OAI21_X1 U17083 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16070), .A(
        n20263), .ZN(n14800) );
  INV_X1 U17084 ( .A(n14800), .ZN(n15887) );
  NAND3_X1 U17085 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n14803), .ZN(n13751) );
  OAI211_X1 U17086 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n16158), .A(
        n15887), .B(n13751), .ZN(n13758) );
  NAND2_X1 U17087 ( .A1(n13753), .A2(n13752), .ZN(n13754) );
  NAND2_X1 U17088 ( .A1(n13919), .A2(n13754), .ZN(n14304) );
  INV_X2 U17089 ( .A(n16162), .ZN(n16174) );
  NAND2_X1 U17090 ( .A1(n16174), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13756) );
  AOI21_X1 U17091 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14080) );
  NAND2_X1 U17092 ( .A1(n14803), .A2(n14080), .ZN(n13755) );
  OAI211_X1 U17093 ( .C1(n20258), .C2(n14304), .A(n13756), .B(n13755), .ZN(
        n13757) );
  AOI221_X1 U17094 ( .B1(n13759), .B2(n11216), .C1(n13758), .C2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n13757), .ZN(n13760) );
  OAI21_X1 U17095 ( .B1(n16182), .B2(n13818), .A(n13760), .ZN(P1_U3029) );
  NOR3_X1 U17096 ( .A1(n17393), .A2(n13762), .A3(n13761), .ZN(n13763) );
  NOR4_X4 U17097 ( .A1(n19008), .A2(n18314), .A3(n15907), .A4(n18846), .ZN(
        n17344) );
  INV_X1 U17098 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17002) );
  NAND2_X1 U17099 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17332) );
  NOR2_X1 U17100 ( .A1(n17002), .A2(n17332), .ZN(n17325) );
  NAND3_X1 U17101 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17325), .ZN(n13775) );
  NAND3_X1 U17102 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17322), .ZN(n17315) );
  INV_X1 U17103 ( .A(n17315), .ZN(n17313) );
  NAND2_X1 U17104 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17313), .ZN(n17269) );
  AOI22_X1 U17105 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11392), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13774) );
  AOI22_X1 U17106 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13766) );
  AOI22_X1 U17107 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13765) );
  OAI211_X1 U17108 ( .C1(n13764), .C2(n18317), .A(n13766), .B(n13765), .ZN(
        n13772) );
  AOI22_X1 U17109 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13770) );
  AOI22_X1 U17110 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13769) );
  AOI22_X1 U17111 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13768) );
  NAND2_X1 U17112 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13767) );
  NAND4_X1 U17113 ( .A1(n13770), .A2(n13769), .A3(n13768), .A4(n13767), .ZN(
        n13771) );
  AOI211_X1 U17114 ( .C1(n9810), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n13772), .B(n13771), .ZN(n13773) );
  OAI211_X1 U17115 ( .C1(n15798), .C2(n17203), .A(n13774), .B(n13773), .ZN(
        n17465) );
  OAI222_X1 U17116 ( .A1(n17341), .A2(P3_EBX_REG_8__SCAN_IN), .B1(n17341), 
        .B2(n17269), .C1(n17324), .C2(n17465), .ZN(n13779) );
  NAND3_X1 U17117 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n14210) );
  INV_X1 U17118 ( .A(n14210), .ZN(n13777) );
  INV_X1 U17119 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n13776) );
  NAND2_X1 U17120 ( .A1(n18350), .A2(n17344), .ZN(n17338) );
  NAND3_X1 U17121 ( .A1(n13777), .A2(n13776), .A3(n17328), .ZN(n13778) );
  NAND2_X1 U17122 ( .A1(n13779), .A2(n13778), .ZN(P3_U2695) );
  NAND2_X1 U17123 ( .A1(n13780), .A2(n10336), .ZN(n13782) );
  INV_X1 U17124 ( .A(n13781), .ZN(n13803) );
  OAI21_X1 U17125 ( .B1(n13783), .B2(n13782), .A(n13803), .ZN(n13994) );
  AOI21_X1 U17126 ( .B1(n13785), .B2(n13784), .A(n13797), .ZN(n19281) );
  INV_X1 U17127 ( .A(n19281), .ZN(n19292) );
  NOR2_X1 U17128 ( .A1(n19292), .A2(n15221), .ZN(n13786) );
  AOI21_X1 U17129 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n15221), .A(n13786), .ZN(
        n13787) );
  OAI21_X1 U17130 ( .B1(n13994), .B2(n15237), .A(n13787), .ZN(P2_U2883) );
  INV_X1 U17131 ( .A(n19987), .ZN(n20009) );
  INV_X1 U17132 ( .A(n10039), .ZN(n16425) );
  MUX2_X1 U17133 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n16425), .S(n15235), .Z(
        n13790) );
  AOI21_X1 U17134 ( .B1(n20009), .B2(n15224), .A(n13790), .ZN(n13791) );
  INV_X1 U17135 ( .A(n13791), .ZN(P2_U2884) );
  NAND2_X1 U17136 ( .A1(n13795), .A2(n13792), .ZN(n13793) );
  INV_X1 U17137 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20211) );
  INV_X1 U17138 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16584) );
  NAND2_X1 U17139 ( .A1(n14607), .A2(n16584), .ZN(n13794) );
  OAI21_X1 U17140 ( .B1(n14609), .B2(DATAI_0_), .A(n13794), .ZN(n20267) );
  OAI222_X1 U17141 ( .A1(n14624), .A2(n14038), .B1(n14611), .B2(n20211), .C1(
        n20267), .C2(n14610), .ZN(P1_U2904) );
  XOR2_X1 U17142 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13803), .Z(n13800)
         );
  OAI21_X1 U17143 ( .B1(n13798), .B2(n13797), .A(n13805), .ZN(n16356) );
  MUX2_X1 U17144 ( .A(n15102), .B(n16356), .S(n15235), .Z(n13799) );
  OAI21_X1 U17145 ( .B1(n13800), .B2(n15237), .A(n13799), .ZN(P2_U2882) );
  NOR2_X1 U17146 ( .A1(n13803), .A2(n13801), .ZN(n13804) );
  OR2_X1 U17147 ( .A1(n13803), .A2(n13802), .ZN(n13829) );
  OAI211_X1 U17148 ( .C1(n13804), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15224), .B(n13829), .ZN(n13808) );
  AOI21_X1 U17149 ( .B1(n13806), .B2(n13805), .A(n13830), .ZN(n19155) );
  NAND2_X1 U17150 ( .A1(n19155), .A2(n15235), .ZN(n13807) );
  OAI211_X1 U17151 ( .C1(n15235), .C2(n13809), .A(n13808), .B(n13807), .ZN(
        P2_U2881) );
  INV_X1 U17152 ( .A(n13810), .ZN(n13811) );
  AOI21_X1 U17153 ( .B1(n13813), .B2(n13812), .A(n13811), .ZN(n14296) );
  INV_X1 U17154 ( .A(n13814), .ZN(n16001) );
  AOI22_X1 U17155 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13815) );
  OAI21_X1 U17156 ( .B1(n14297), .B2(n16022), .A(n13815), .ZN(n13816) );
  AOI21_X1 U17157 ( .B1(n14296), .B2(n16001), .A(n13816), .ZN(n13817) );
  OAI21_X1 U17158 ( .B1(n20080), .B2(n13818), .A(n13817), .ZN(P1_U2997) );
  INV_X1 U17159 ( .A(n13819), .ZN(n13820) );
  NOR2_X1 U17160 ( .A1(n13821), .A2(n13820), .ZN(n13823) );
  NAND2_X1 U17161 ( .A1(n20015), .A2(n15127), .ZN(n13887) );
  OAI21_X1 U17162 ( .B1(n20015), .B2(n15127), .A(n13887), .ZN(n13822) );
  NOR2_X1 U17163 ( .A1(n13823), .A2(n13822), .ZN(n13889) );
  AOI21_X1 U17164 ( .B1(n13823), .B2(n13822), .A(n13889), .ZN(n13826) );
  INV_X1 U17165 ( .A(n15127), .ZN(n20017) );
  AOI22_X1 U17166 ( .A1(n20017), .A2(n19198), .B1(n19203), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13825) );
  NAND2_X1 U17167 ( .A1(n19213), .A2(n15317), .ZN(n13824) );
  OAI211_X1 U17168 ( .C1(n13826), .C2(n15327), .A(n13825), .B(n13824), .ZN(
        P2_U2917) );
  INV_X1 U17169 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20208) );
  INV_X1 U17170 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16579) );
  NAND2_X1 U17171 ( .A1(n14609), .A2(n16579), .ZN(n13827) );
  OAI21_X1 U17172 ( .B1(n14609), .B2(DATAI_1_), .A(n13827), .ZN(n20276) );
  OAI222_X1 U17173 ( .A1(n14054), .A2(n14624), .B1(n14611), .B2(n20208), .C1(
        n20276), .C2(n14610), .ZN(P1_U2903) );
  INV_X1 U17174 ( .A(n14296), .ZN(n13865) );
  INV_X1 U17175 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20206) );
  INV_X1 U17176 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16577) );
  NAND2_X1 U17177 ( .A1(n14609), .A2(n16577), .ZN(n13828) );
  OAI21_X1 U17178 ( .B1(n14609), .B2(DATAI_2_), .A(n13828), .ZN(n20283) );
  OAI222_X1 U17179 ( .A1(n13865), .A2(n14624), .B1(n14611), .B2(n20206), .C1(
        n20283), .C2(n14610), .ZN(P1_U2902) );
  XOR2_X1 U17180 ( .A(n13829), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13833)
         );
  OAI21_X1 U17181 ( .B1(n13831), .B2(n13830), .A(n13840), .ZN(n16354) );
  MUX2_X1 U17182 ( .A(n12405), .B(n16354), .S(n15235), .Z(n13832) );
  OAI21_X1 U17183 ( .B1(n13833), .B2(n15237), .A(n13832), .ZN(P2_U2880) );
  XNOR2_X1 U17184 ( .A(n13834), .B(n13835), .ZN(n13838) );
  OAI21_X1 U17185 ( .B1(n13836), .B2(n13839), .A(n13910), .ZN(n16338) );
  MUX2_X1 U17186 ( .A(n12366), .B(n16338), .S(n15235), .Z(n13837) );
  OAI21_X1 U17187 ( .B1(n13838), .B2(n15237), .A(n13837), .ZN(P2_U2878) );
  AOI21_X1 U17188 ( .B1(n13841), .B2(n13840), .A(n13839), .ZN(n19142) );
  INV_X1 U17189 ( .A(n19142), .ZN(n13847) );
  AND2_X1 U17190 ( .A1(n13781), .A2(n13842), .ZN(n13844) );
  OAI211_X1 U17191 ( .C1(n13844), .C2(n13843), .A(n13834), .B(n15224), .ZN(
        n13846) );
  NAND2_X1 U17192 ( .A1(n15221), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13845) );
  OAI211_X1 U17193 ( .C1(n13847), .C2(n15221), .A(n13846), .B(n13845), .ZN(
        P2_U2879) );
  OAI21_X1 U17194 ( .B1(n13849), .B2(n15055), .A(n13848), .ZN(n19132) );
  INV_X1 U17195 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19233) );
  OAI222_X1 U17196 ( .A1(n14010), .A2(n13850), .B1(n19132), .B2(n19206), .C1(
        n19217), .C2(n19233), .ZN(P2_U2907) );
  XNOR2_X1 U17197 ( .A(n13852), .B(n13851), .ZN(n13924) );
  OR2_X1 U17198 ( .A1(n13855), .A2(n13854), .ZN(n13856) );
  AND2_X1 U17199 ( .A1(n13853), .A2(n13856), .ZN(n20177) );
  INV_X1 U17200 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14063) );
  NOR2_X1 U17201 ( .A1(n16162), .A2(n14063), .ZN(n13921) );
  AOI21_X1 U17202 ( .B1(n16015), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13921), .ZN(n13857) );
  OAI21_X1 U17203 ( .B1(n14067), .B2(n16022), .A(n13857), .ZN(n13858) );
  AOI21_X1 U17204 ( .B1(n20177), .B2(n16001), .A(n13858), .ZN(n13859) );
  OAI21_X1 U17205 ( .B1(n13924), .B2(n20080), .A(n13859), .ZN(P1_U2996) );
  INV_X1 U17206 ( .A(n20177), .ZN(n14072) );
  NAND2_X1 U17207 ( .A1(n14153), .A2(DATAI_3_), .ZN(n13861) );
  NAND2_X1 U17208 ( .A1(n14609), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13860) );
  INV_X1 U17209 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20204) );
  OAI222_X1 U17210 ( .A1(n14624), .A2(n14072), .B1(n20288), .B2(n14610), .C1(
        n14611), .C2(n20204), .ZN(P1_U2901) );
  NAND2_X1 U17211 ( .A1(n13862), .A2(n20265), .ZN(n13864) );
  NAND2_X1 U17212 ( .A1(n13864), .A2(n13863), .ZN(n20257) );
  INV_X1 U17213 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n21141) );
  OAI222_X1 U17214 ( .A1(n20257), .A2(n14521), .B1(n21141), .B2(n20179), .C1(
        n14038), .C2(n14532), .ZN(P1_U2872) );
  INV_X1 U17215 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n21290) );
  OAI222_X1 U17216 ( .A1(n14304), .A2(n14521), .B1(n20179), .B2(n21290), .C1(
        n13865), .C2(n14532), .ZN(P1_U2870) );
  INV_X1 U17217 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21167) );
  AOI22_X1 U17218 ( .A1(n13869), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13866) );
  OAI21_X1 U17219 ( .B1(n21167), .B2(n13880), .A(n13866), .ZN(P1_U2915) );
  AOI22_X1 U17220 ( .A1(n13869), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13867) );
  OAI21_X1 U17221 ( .B1(n21258), .B2(n13880), .A(n13867), .ZN(P1_U2910) );
  INV_X1 U17222 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n21274) );
  AOI22_X1 U17223 ( .A1(n13869), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13868) );
  OAI21_X1 U17224 ( .B1(n21274), .B2(n13880), .A(n13868), .ZN(P1_U2914) );
  AOI22_X1 U17225 ( .A1(n13869), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13870) );
  OAI21_X1 U17226 ( .B1(n21105), .B2(n13880), .A(n13870), .ZN(P1_U2909) );
  INV_X1 U17227 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U17228 ( .A1(n20941), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13871) );
  OAI21_X1 U17229 ( .B1(n13872), .B2(n13880), .A(n13871), .ZN(P1_U2917) );
  INV_X1 U17230 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U17231 ( .A1(n20941), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13873) );
  OAI21_X1 U17232 ( .B1(n13874), .B2(n13880), .A(n13873), .ZN(P1_U2919) );
  INV_X1 U17233 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U17234 ( .A1(n20941), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13875) );
  OAI21_X1 U17235 ( .B1(n13876), .B2(n13880), .A(n13875), .ZN(P1_U2918) );
  INV_X1 U17236 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13878) );
  AOI22_X1 U17237 ( .A1(n20941), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13877) );
  OAI21_X1 U17238 ( .B1(n13878), .B2(n13880), .A(n13877), .ZN(P1_U2920) );
  AOI22_X1 U17239 ( .A1(n20941), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13879) );
  OAI21_X1 U17240 ( .B1(n10916), .B2(n13880), .A(n13879), .ZN(P1_U2916) );
  NAND2_X1 U17241 ( .A1(n13853), .A2(n13882), .ZN(n13883) );
  AND2_X1 U17242 ( .A1(n13881), .A2(n13883), .ZN(n20158) );
  NAND2_X1 U17243 ( .A1(n14153), .A2(DATAI_4_), .ZN(n13885) );
  NAND2_X1 U17244 ( .A1(n14609), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13884) );
  AND2_X1 U17245 ( .A1(n13885), .A2(n13884), .ZN(n20227) );
  INV_X1 U17246 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20202) );
  OAI222_X1 U17247 ( .A1(n13927), .A2(n14624), .B1(n20227), .B2(n14610), .C1(
        n20202), .C2(n14611), .ZN(P1_U2900) );
  XNOR2_X1 U17248 ( .A(n13886), .B(n9908), .ZN(n20008) );
  XOR2_X1 U17249 ( .A(n20008), .B(n19987), .Z(n13891) );
  INV_X1 U17250 ( .A(n13887), .ZN(n13888) );
  NOR2_X1 U17251 ( .A1(n13889), .A2(n13888), .ZN(n13890) );
  NOR2_X1 U17252 ( .A1(n13890), .A2(n13891), .ZN(n13982) );
  AOI21_X1 U17253 ( .B1(n13891), .B2(n13890), .A(n13982), .ZN(n13894) );
  AOI22_X1 U17254 ( .A1(n19213), .A2(n15307), .B1(n19203), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n13893) );
  NAND2_X1 U17255 ( .A1(n19198), .A2(n20008), .ZN(n13892) );
  OAI211_X1 U17256 ( .C1(n13894), .C2(n15327), .A(n13893), .B(n13892), .ZN(
        P2_U2916) );
  XNOR2_X1 U17257 ( .A(n13895), .B(n14004), .ZN(n13900) );
  NOR2_X1 U17258 ( .A1(n13896), .A2(n13909), .ZN(n13897) );
  NOR2_X1 U17259 ( .A1(n14000), .A2(n13897), .ZN(n16388) );
  NOR2_X1 U17260 ( .A1(n15235), .A2(n12372), .ZN(n13898) );
  AOI21_X1 U17261 ( .B1(n16388), .B2(n15235), .A(n13898), .ZN(n13899) );
  OAI21_X1 U17262 ( .B1(n13900), .B2(n15237), .A(n13899), .ZN(P2_U2876) );
  XNOR2_X1 U17263 ( .A(n13901), .B(n13902), .ZN(n13933) );
  INV_X1 U17264 ( .A(n13903), .ZN(n20141) );
  NOR2_X1 U17265 ( .A1(n16162), .A2(n21299), .ZN(n13929) );
  AOI21_X1 U17266 ( .B1(n16015), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13929), .ZN(n13904) );
  OAI21_X1 U17267 ( .B1(n20141), .B2(n16022), .A(n13904), .ZN(n13905) );
  AOI21_X1 U17268 ( .B1(n20158), .B2(n16025), .A(n13905), .ZN(n13906) );
  OAI21_X1 U17269 ( .B1(n13933), .B2(n20080), .A(n13906), .ZN(P1_U2995) );
  INV_X1 U17270 ( .A(n13895), .ZN(n13907) );
  OAI211_X1 U17271 ( .C1(n9911), .C2(n13908), .A(n13907), .B(n15224), .ZN(
        n13913) );
  AOI21_X1 U17272 ( .B1(n13911), .B2(n13910), .A(n13909), .ZN(n16398) );
  NAND2_X1 U17273 ( .A1(n16398), .A2(n15235), .ZN(n13912) );
  OAI211_X1 U17274 ( .C1(n15235), .C2(n13914), .A(n13913), .B(n13912), .ZN(
        P2_U2877) );
  NOR2_X1 U17275 ( .A1(n11216), .A2(n12679), .ZN(n13915) );
  OAI21_X1 U17276 ( .B1(n13915), .B2(n16158), .A(n15887), .ZN(n16137) );
  AOI21_X1 U17277 ( .B1(n14803), .B2(n14080), .A(n16137), .ZN(n13916) );
  INV_X1 U17278 ( .A(n13916), .ZN(n13930) );
  NOR3_X1 U17279 ( .A1(n11216), .A2(n12679), .A3(n14896), .ZN(n16154) );
  NOR2_X1 U17280 ( .A1(n14803), .A2(n16154), .ZN(n16141) );
  NOR2_X1 U17281 ( .A1(n14080), .A2(n16141), .ZN(n14898) );
  AOI22_X1 U17282 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13930), .B1(
        n14898), .B2(n13917), .ZN(n13923) );
  AND2_X1 U17283 ( .A1(n13919), .A2(n13918), .ZN(n13920) );
  NOR2_X1 U17284 ( .A1(n9922), .A2(n13920), .ZN(n20174) );
  AOI21_X1 U17285 ( .B1(n16173), .B2(n20174), .A(n13921), .ZN(n13922) );
  OAI211_X1 U17286 ( .C1(n16182), .C2(n13924), .A(n13923), .B(n13922), .ZN(
        P1_U3028) );
  OR2_X1 U17287 ( .A1(n9922), .A2(n13925), .ZN(n13926) );
  NAND2_X1 U17288 ( .A1(n14078), .A2(n13926), .ZN(n20154) );
  INV_X1 U17289 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21095) );
  OAI222_X1 U17290 ( .A1(n20154), .A2(n14521), .B1(n20179), .B2(n21095), .C1(
        n13927), .C2(n14532), .ZN(P1_U2868) );
  NAND2_X1 U17291 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14897) );
  OAI211_X1 U17292 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n14898), .B(n14897), .ZN(n13932) );
  NOR2_X1 U17293 ( .A1(n20258), .A2(n20154), .ZN(n13928) );
  AOI211_X1 U17294 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n13930), .A(
        n13929), .B(n13928), .ZN(n13931) );
  OAI211_X1 U17295 ( .C1(n16182), .C2(n13933), .A(n13932), .B(n13931), .ZN(
        P1_U3027) );
  NOR2_X1 U17296 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20834), .ZN(n13955) );
  MUX2_X1 U17297 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13934), .S(
        n15846), .Z(n15852) );
  AOI22_X1 U17298 ( .A1(n13955), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20834), .B2(n15852), .ZN(n13958) );
  NAND2_X1 U17299 ( .A1(n20913), .A2(n13935), .ZN(n13953) );
  NAND2_X1 U17300 ( .A1(n13936), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13937) );
  NAND2_X1 U17301 ( .A1(n13938), .A2(n13937), .ZN(n20904) );
  AND2_X1 U17302 ( .A1(n13939), .A2(n20904), .ZN(n13950) );
  MUX2_X1 U17303 ( .A(n13941), .B(n9823), .S(n13940), .Z(n13943) );
  OR2_X1 U17304 ( .A1(n13943), .A2(n13942), .ZN(n13947) );
  XNOR2_X1 U17305 ( .A(n13944), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13945) );
  OAI22_X1 U17306 ( .A1(n13948), .A2(n13947), .B1(n13946), .B2(n13945), .ZN(
        n13949) );
  AOI21_X1 U17307 ( .B1(n13951), .B2(n13950), .A(n13949), .ZN(n13952) );
  NAND2_X1 U17308 ( .A1(n13953), .A2(n13952), .ZN(n20907) );
  NOR2_X1 U17309 ( .A1(n15846), .A2(n10010), .ZN(n13954) );
  AOI21_X1 U17310 ( .B1(n20907), .B2(n15846), .A(n13954), .ZN(n15853) );
  INV_X1 U17311 ( .A(n15853), .ZN(n13956) );
  AOI22_X1 U17312 ( .A1(n13956), .A2(n20834), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13955), .ZN(n13957) );
  NOR2_X1 U17313 ( .A1(n15856), .A2(n13578), .ZN(n13986) );
  NAND2_X1 U17314 ( .A1(n15846), .A2(n20834), .ZN(n13959) );
  NOR2_X1 U17315 ( .A1(n13959), .A2(n12643), .ZN(n13962) );
  NAND2_X1 U17316 ( .A1(n13959), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13960) );
  NOR2_X1 U17317 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13960), .ZN(n13961) );
  AOI21_X1 U17318 ( .B1(n20145), .B2(n13962), .A(n13961), .ZN(n15861) );
  INV_X1 U17319 ( .A(n15861), .ZN(n13985) );
  NOR3_X1 U17320 ( .A1(n13986), .A2(P1_FLUSH_REG_SCAN_IN), .A3(n13985), .ZN(
        n13964) );
  NAND2_X1 U17321 ( .A1(n20339), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20623) );
  XOR2_X1 U17322 ( .A(n20623), .B(n11217), .Z(n13965) );
  NAND2_X1 U17323 ( .A1(n20661), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20914) );
  INV_X1 U17324 ( .A(n20914), .ZN(n14907) );
  OAI22_X1 U17325 ( .A1(n13965), .A2(n20920), .B1(n13609), .B2(n14907), .ZN(
        n13966) );
  NAND2_X1 U17326 ( .A1(n20923), .A2(n13966), .ZN(n13967) );
  OAI21_X1 U17327 ( .B1(n20923), .B2(n11143), .A(n13967), .ZN(P1_U3476) );
  NAND2_X1 U17328 ( .A1(n13881), .A2(n13969), .ZN(n13970) );
  AND2_X1 U17329 ( .A1(n13968), .A2(n13970), .ZN(n20171) );
  INV_X1 U17330 ( .A(n20171), .ZN(n13973) );
  NAND2_X1 U17331 ( .A1(n14153), .A2(DATAI_5_), .ZN(n13972) );
  NAND2_X1 U17332 ( .A1(n14609), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13971) );
  AND2_X1 U17333 ( .A1(n13972), .A2(n13971), .ZN(n20295) );
  OAI222_X1 U17334 ( .A1(n14624), .A2(n13973), .B1(n20295), .B2(n14610), .C1(
        n14611), .C2(n10675), .ZN(P1_U2899) );
  INV_X1 U17335 ( .A(n13974), .ZN(n13975) );
  NAND2_X1 U17336 ( .A1(n13976), .A2(n13975), .ZN(n13977) );
  NAND2_X1 U17337 ( .A1(n13978), .A2(n13977), .ZN(n15736) );
  NOR2_X1 U17338 ( .A1(n20009), .A2(n20008), .ZN(n13981) );
  XOR2_X1 U17339 ( .A(n13980), .B(n13979), .Z(n19167) );
  INV_X1 U17340 ( .A(n19167), .ZN(n19293) );
  OAI21_X1 U17341 ( .B1(n13982), .B2(n13981), .A(n19293), .ZN(n13995) );
  INV_X1 U17342 ( .A(n13994), .ZN(n19169) );
  NAND3_X1 U17343 ( .A1(n13995), .A2(n16268), .A3(n19169), .ZN(n13984) );
  AOI22_X1 U17344 ( .A1(n19213), .A2(n15291), .B1(n19203), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n13983) );
  OAI211_X1 U17345 ( .C1(n19206), .C2(n15736), .A(n13984), .B(n13983), .ZN(
        P2_U2914) );
  NOR3_X1 U17346 ( .A1(n13986), .A2(n16190), .A3(n13985), .ZN(n15866) );
  OAI22_X1 U17347 ( .A1(n20338), .A2(n20920), .B1(n13987), .B2(n14907), .ZN(
        n13988) );
  OAI21_X1 U17348 ( .B1(n15866), .B2(n13988), .A(n20923), .ZN(n13989) );
  OAI21_X1 U17349 ( .B1(n20923), .B2(n20696), .A(n13989), .ZN(P1_U3478) );
  INV_X1 U17350 ( .A(n14047), .ZN(n13990) );
  OAI22_X1 U17351 ( .A1(n14521), .A2(n13990), .B1(n14050), .B2(n20179), .ZN(
        n13991) );
  AOI21_X1 U17352 ( .B1(n13992), .B2(n20176), .A(n13991), .ZN(n13993) );
  INV_X1 U17353 ( .A(n13993), .ZN(P1_U2871) );
  XNOR2_X1 U17354 ( .A(n13995), .B(n13994), .ZN(n13996) );
  NAND2_X1 U17355 ( .A1(n13996), .A2(n16268), .ZN(n13998) );
  AOI22_X1 U17356 ( .A1(n19213), .A2(n15301), .B1(n19203), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13997) );
  OAI211_X1 U17357 ( .C1(n19293), .C2(n15310), .A(n13998), .B(n13997), .ZN(
        P2_U2915) );
  NOR2_X1 U17358 ( .A1(n14000), .A2(n13999), .ZN(n14001) );
  OR2_X1 U17359 ( .A1(n14043), .A2(n14001), .ZN(n16301) );
  AOI21_X1 U17360 ( .B1(n13895), .B2(n14004), .A(n14003), .ZN(n14005) );
  OR3_X1 U17361 ( .A1(n14002), .A2(n14005), .A3(n15237), .ZN(n14007) );
  NAND2_X1 U17362 ( .A1(n15221), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14006) );
  OAI211_X1 U17363 ( .C1(n16301), .C2(n15221), .A(n14007), .B(n14006), .ZN(
        P2_U2875) );
  XNOR2_X1 U17364 ( .A(n14124), .B(n14008), .ZN(n19110) );
  OAI222_X1 U17365 ( .A1(n19110), .A2(n19206), .B1(n14010), .B2(n14009), .C1(
        n19217), .C2(n13357), .ZN(P2_U2904) );
  NAND2_X1 U17366 ( .A1(n14012), .A2(n9815), .ZN(n14014) );
  XNOR2_X1 U17367 ( .A(n14014), .B(n14013), .ZN(n14027) );
  XOR2_X1 U17368 ( .A(n12414), .B(n14015), .Z(n14025) );
  MUX2_X1 U17369 ( .A(n15737), .B(n15726), .S(n15738), .Z(n14019) );
  INV_X1 U17370 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19919) );
  NOR2_X1 U17371 ( .A1(n19919), .A2(n19150), .ZN(n14016) );
  AOI21_X1 U17372 ( .B1(n16387), .B2(n20008), .A(n14016), .ZN(n14017) );
  OAI21_X1 U17373 ( .B1(n10039), .B2(n19308), .A(n14017), .ZN(n14018) );
  AOI211_X1 U17374 ( .C1(n14025), .C2(n16413), .A(n14019), .B(n14018), .ZN(
        n14020) );
  OAI21_X1 U17375 ( .B1(n14027), .B2(n19314), .A(n14020), .ZN(P2_U3043) );
  OAI21_X1 U17376 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14021), .A(
        n14924), .ZN(n15110) );
  NAND2_X1 U17377 ( .A1(n16425), .A2(n19282), .ZN(n14023) );
  AOI22_X1 U17378 ( .A1(n16355), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n19287), .B2(P2_REIP_REG_3__SCAN_IN), .ZN(n14022) );
  OAI211_X1 U17379 ( .C1(n15110), .C2(n16366), .A(n14023), .B(n14022), .ZN(
        n14024) );
  AOI21_X1 U17380 ( .B1(n14025), .B2(n16350), .A(n14024), .ZN(n14026) );
  OAI21_X1 U17381 ( .B1(n14027), .B2(n19278), .A(n14026), .ZN(P2_U3011) );
  NOR2_X1 U17382 ( .A1(n14036), .A2(n14028), .ZN(n20144) );
  OAI22_X1 U17383 ( .A1(n21141), .A2(n20107), .B1(n20155), .B2(n20257), .ZN(
        n14029) );
  INV_X1 U17384 ( .A(n14029), .ZN(n14034) );
  OAI21_X1 U17385 ( .B1(n20127), .B2(n20139), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14033) );
  OAI211_X1 U17386 ( .C1(n20106), .C2(n13727), .A(n14034), .B(n14033), .ZN(
        n14040) );
  NOR2_X1 U17387 ( .A1(n14036), .A2(n14035), .ZN(n14037) );
  OR2_X1 U17388 ( .A1(n20123), .A2(n14037), .ZN(n20157) );
  NOR2_X1 U17389 ( .A1(n14038), .A2(n14071), .ZN(n14039) );
  AOI211_X1 U17390 ( .C1(n20144), .C2(n10591), .A(n14040), .B(n14039), .ZN(
        n14041) );
  INV_X1 U17391 ( .A(n14041), .ZN(P1_U2840) );
  XNOR2_X1 U17392 ( .A(n14002), .B(n14086), .ZN(n14046) );
  OR2_X1 U17393 ( .A1(n14043), .A2(n14042), .ZN(n14044) );
  NAND2_X1 U17394 ( .A1(n14044), .A2(n14091), .ZN(n16376) );
  MUX2_X1 U17395 ( .A(n16376), .B(n15040), .S(n15221), .Z(n14045) );
  OAI21_X1 U17396 ( .B1(n14046), .B2(n15237), .A(n14045), .ZN(P2_U2874) );
  NOR2_X1 U17397 ( .A1(n20142), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14052) );
  AOI22_X1 U17398 ( .A1(n15941), .A2(n21275), .B1(n20130), .B2(n14047), .ZN(
        n14049) );
  AOI22_X1 U17399 ( .A1(n20139), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20117), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14048) );
  OAI211_X1 U17400 ( .C1(n14050), .C2(n20107), .A(n14049), .B(n14048), .ZN(
        n14051) );
  AOI211_X1 U17401 ( .C1(n20144), .C2(n20731), .A(n14052), .B(n14051), .ZN(
        n14053) );
  OAI21_X1 U17402 ( .B1(n14054), .B2(n14071), .A(n14053), .ZN(P1_U2839) );
  XNOR2_X1 U17403 ( .A(n14055), .B(n14056), .ZN(n16183) );
  AOI21_X1 U17404 ( .B1(n14059), .B2(n13968), .A(n14058), .ZN(n20124) );
  INV_X1 U17405 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21255) );
  NOR2_X1 U17406 ( .A1(n16162), .A2(n21255), .ZN(n16186) );
  AOI21_X1 U17407 ( .B1(n16015), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16186), .ZN(n14060) );
  OAI21_X1 U17408 ( .B1(n20120), .B2(n16022), .A(n14060), .ZN(n14061) );
  AOI21_X1 U17409 ( .B1(n20124), .B2(n16025), .A(n14061), .ZN(n14062) );
  OAI21_X1 U17410 ( .B1(n20080), .B2(n16183), .A(n14062), .ZN(P1_U2993) );
  INV_X1 U17411 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n21284) );
  NAND4_X1 U17412 ( .A1(n15941), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .A4(n14063), .ZN(n14065) );
  AOI21_X1 U17413 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .A(n20148), .ZN(n14299) );
  OR2_X1 U17414 ( .A1(n20117), .A2(n14299), .ZN(n14300) );
  AOI22_X1 U17415 ( .A1(n20139), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n14300), .ZN(n14064) );
  OAI211_X1 U17416 ( .C1(n21284), .C2(n20107), .A(n14065), .B(n14064), .ZN(
        n14069) );
  INV_X1 U17417 ( .A(n20174), .ZN(n14066) );
  OAI22_X1 U17418 ( .A1(n20142), .A2(n14067), .B1(n20155), .B2(n14066), .ZN(
        n14068) );
  OAI21_X1 U17419 ( .B1(n14072), .B2(n14071), .A(n14070), .ZN(P1_U2837) );
  INV_X1 U17420 ( .A(n20124), .ZN(n14099) );
  NAND2_X1 U17421 ( .A1(n14153), .A2(DATAI_6_), .ZN(n14074) );
  NAND2_X1 U17422 ( .A1(n14609), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14073) );
  AND2_X1 U17423 ( .A1(n14074), .A2(n14073), .ZN(n20303) );
  OAI222_X1 U17424 ( .A1(n14624), .A2(n14099), .B1(n20303), .B2(n14610), .C1(
        n14611), .C2(n10696), .ZN(P1_U2898) );
  XOR2_X1 U17425 ( .A(n14075), .B(n14076), .Z(n16026) );
  NAND2_X1 U17426 ( .A1(n14078), .A2(n14077), .ZN(n14079) );
  NAND2_X1 U17427 ( .A1(n14097), .A2(n14079), .ZN(n20169) );
  NOR3_X1 U17428 ( .A1(n11216), .A2(n12679), .A3(n14897), .ZN(n16159) );
  NOR3_X1 U17429 ( .A1(n14897), .A2(n16155), .A3(n14080), .ZN(n16135) );
  INV_X1 U17430 ( .A(n16135), .ZN(n14791) );
  AOI21_X1 U17431 ( .B1(n14803), .B2(n14791), .A(n14800), .ZN(n16157) );
  OAI21_X1 U17432 ( .B1(n16159), .B2(n16158), .A(n16157), .ZN(n14082) );
  NOR2_X1 U17433 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14897), .ZN(
        n14081) );
  AOI22_X1 U17434 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14082), .B1(
        n14898), .B2(n14081), .ZN(n14083) );
  NAND2_X1 U17435 ( .A1(n16174), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16027) );
  OAI211_X1 U17436 ( .C1(n20258), .C2(n20169), .A(n14083), .B(n16027), .ZN(
        n14084) );
  AOI21_X1 U17437 ( .B1(n20260), .B2(n16026), .A(n14084), .ZN(n14085) );
  INV_X1 U17438 ( .A(n14085), .ZN(P1_U3026) );
  AND2_X1 U17439 ( .A1(n14002), .A2(n14086), .ZN(n14089) );
  OAI211_X1 U17440 ( .C1(n14089), .C2(n14088), .A(n15224), .B(n14087), .ZN(
        n14094) );
  AOI21_X1 U17441 ( .B1(n14092), .B2(n14091), .A(n14090), .ZN(n19117) );
  NAND2_X1 U17442 ( .A1(n19117), .A2(n15235), .ZN(n14093) );
  OAI211_X1 U17443 ( .C1(n15235), .C2(n14095), .A(n14094), .B(n14093), .ZN(
        P2_U2873) );
  AND2_X1 U17444 ( .A1(n14097), .A2(n14096), .ZN(n14098) );
  OR2_X1 U17445 ( .A1(n14098), .A2(n16170), .ZN(n20119) );
  INV_X1 U17446 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14100) );
  OAI222_X1 U17447 ( .A1(n20119), .A2(n14521), .B1(n20179), .B2(n14100), .C1(
        n14099), .C2(n14532), .ZN(P1_U2866) );
  OR2_X1 U17448 ( .A1(n14058), .A2(n14102), .ZN(n14103) );
  AND2_X1 U17449 ( .A1(n14101), .A2(n14103), .ZN(n20166) );
  INV_X1 U17450 ( .A(n20166), .ZN(n14106) );
  NAND2_X1 U17451 ( .A1(n14153), .A2(DATAI_7_), .ZN(n14105) );
  NAND2_X1 U17452 ( .A1(n14609), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14104) );
  AND2_X1 U17453 ( .A1(n14105), .A2(n14104), .ZN(n20231) );
  OAI222_X1 U17454 ( .A1(n14624), .A2(n14106), .B1(n20231), .B2(n14610), .C1(
        n14611), .C2(n10706), .ZN(P1_U2897) );
  AOI21_X1 U17455 ( .B1(n14108), .B2(n14101), .A(n14107), .ZN(n14144) );
  INV_X1 U17456 ( .A(n14144), .ZN(n14119) );
  AOI22_X1 U17457 ( .A1(n14622), .A2(n14564), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15974), .ZN(n14109) );
  OAI21_X1 U17458 ( .B1(n14119), .B2(n14624), .A(n14109), .ZN(P1_U2896) );
  OAI21_X1 U17459 ( .B1(n16172), .B2(n14110), .A(n16145), .ZN(n16163) );
  INV_X1 U17460 ( .A(n16163), .ZN(n14117) );
  OR2_X1 U17461 ( .A1(n20117), .A2(n20077), .ZN(n20134) );
  AOI21_X1 U17462 ( .B1(n20139), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20138), .ZN(n14112) );
  NAND2_X1 U17463 ( .A1(n20152), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n14111) );
  OAI211_X1 U17464 ( .C1(n20142), .C2(n14142), .A(n14112), .B(n14111), .ZN(
        n14116) );
  NAND2_X1 U17465 ( .A1(n20115), .A2(n14196), .ZN(n14113) );
  AOI21_X1 U17466 ( .B1(n20860), .B2(n14114), .A(n14113), .ZN(n14115) );
  AOI211_X1 U17467 ( .C1(n14117), .C2(n20130), .A(n14116), .B(n14115), .ZN(
        n14118) );
  OAI21_X1 U17468 ( .B1(n14119), .B2(n20099), .A(n14118), .ZN(P1_U2832) );
  INV_X1 U17469 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21271) );
  OAI222_X1 U17470 ( .A1(n14119), .A2(n14532), .B1(n20179), .B2(n21271), .C1(
        n16163), .C2(n14521), .ZN(P1_U2864) );
  AOI21_X1 U17471 ( .B1(n14123), .B2(n14120), .A(n14122), .ZN(n15225) );
  NAND2_X1 U17472 ( .A1(n14124), .A2(n14008), .ZN(n14127) );
  INV_X1 U17473 ( .A(n14125), .ZN(n14126) );
  NAND2_X1 U17474 ( .A1(n14127), .A2(n14126), .ZN(n14128) );
  NAND2_X1 U17475 ( .A1(n14129), .A2(n14128), .ZN(n19094) );
  NOR2_X1 U17476 ( .A1(n19369), .A2(n12957), .ZN(n14130) );
  AOI22_X1 U17477 ( .A1(n19200), .A2(BUF1_REG_16__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n14135) );
  AOI22_X1 U17478 ( .A1(n16266), .A2(n14133), .B1(n19203), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14134) );
  OAI211_X1 U17479 ( .C1(n15310), .C2(n19094), .A(n14135), .B(n14134), .ZN(
        n14136) );
  AOI21_X1 U17480 ( .B1(n15225), .B2(n16268), .A(n14136), .ZN(n14137) );
  INV_X1 U17481 ( .A(n14137), .ZN(P2_U2903) );
  XOR2_X1 U17482 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14139), .Z(
        n14140) );
  XNOR2_X1 U17483 ( .A(n9819), .B(n14140), .ZN(n16161) );
  AOI22_X1 U17484 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14141) );
  OAI21_X1 U17485 ( .B1(n14142), .B2(n16022), .A(n14141), .ZN(n14143) );
  AOI21_X1 U17486 ( .B1(n14144), .B2(n16025), .A(n14143), .ZN(n14145) );
  OAI21_X1 U17487 ( .B1(n20080), .B2(n16161), .A(n14145), .ZN(P1_U2991) );
  AND2_X1 U17488 ( .A1(n10317), .A2(n14146), .ZN(n14148) );
  OR2_X1 U17489 ( .A1(n14148), .A2(n14147), .ZN(n20163) );
  AOI22_X1 U17490 ( .A1(n14622), .A2(n20232), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15974), .ZN(n14149) );
  OAI21_X1 U17491 ( .B1(n20163), .B2(n14624), .A(n14149), .ZN(P1_U2895) );
  INV_X1 U17492 ( .A(n11217), .ZN(n20521) );
  NOR3_X1 U17493 ( .A1(n20334), .A2(n20828), .A3(n20920), .ZN(n14151) );
  AND2_X1 U17494 ( .A1(n20698), .A2(n21137), .ZN(n20915) );
  NOR2_X1 U17495 ( .A1(n14151), .A2(n20915), .ZN(n14154) );
  INV_X1 U17496 ( .A(n13609), .ZN(n14152) );
  OR2_X1 U17497 ( .A1(n20913), .A2(n14152), .ZN(n20380) );
  OR2_X1 U17498 ( .A1(n20380), .A2(n20731), .ZN(n14159) );
  NAND2_X1 U17499 ( .A1(n20523), .A2(n20578), .ZN(n20413) );
  NOR2_X1 U17500 ( .A1(n14155), .A2(n10577), .ZN(n20580) );
  INV_X1 U17501 ( .A(n20580), .ZN(n20525) );
  OAI22_X1 U17502 ( .A1(n14154), .A2(n14159), .B1(n20413), .B2(n20525), .ZN(
        n20307) );
  INV_X1 U17503 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16537) );
  INV_X1 U17504 ( .A(DATAI_28_), .ZN(n21286) );
  INV_X1 U17505 ( .A(n14609), .ZN(n14153) );
  OAI22_X1 U17506 ( .A1(n16537), .A2(n20306), .B1(n21286), .B2(n20304), .ZN(
        n20750) );
  INV_X1 U17507 ( .A(n20750), .ZN(n20810) );
  INV_X1 U17508 ( .A(n14154), .ZN(n14160) );
  INV_X1 U17509 ( .A(n14155), .ZN(n14156) );
  NOR2_X1 U17510 ( .A1(n14156), .A2(n10577), .ZN(n20654) );
  INV_X1 U17511 ( .A(n20584), .ZN(n20343) );
  INV_X1 U17512 ( .A(n20413), .ZN(n14157) );
  NAND3_X1 U17513 ( .A1(n20617), .A2(n11143), .A3(n20655), .ZN(n20314) );
  NOR2_X1 U17514 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20314), .ZN(
        n20294) );
  OAI22_X1 U17515 ( .A1(n14157), .A2(n10577), .B1(n20294), .B2(n20661), .ZN(
        n14158) );
  AOI211_X2 U17516 ( .C1(n14160), .C2(n14159), .A(n20343), .B(n14158), .ZN(
        n20311) );
  INV_X1 U17517 ( .A(n20311), .ZN(n14168) );
  NAND2_X1 U17518 ( .A1(n14168), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14164) );
  INV_X1 U17519 ( .A(DATAI_20_), .ZN(n21032) );
  INV_X1 U17520 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19346) );
  OAI22_X2 U17521 ( .A1(n21032), .A2(n20304), .B1(n19346), .B2(n20306), .ZN(
        n20807) );
  NOR2_X2 U17522 ( .A1(n20273), .A2(n14162), .ZN(n20805) );
  AOI22_X1 U17523 ( .A1(n20334), .A2(n20807), .B1(n20294), .B2(n20805), .ZN(
        n14163) );
  OAI211_X1 U17524 ( .C1(n20803), .C2(n20810), .A(n14164), .B(n14163), .ZN(
        n14165) );
  AOI21_X1 U17525 ( .B1(n20806), .B2(n20307), .A(n14165), .ZN(n14166) );
  INV_X1 U17526 ( .A(n14166), .ZN(P1_U3037) );
  INV_X1 U17527 ( .A(DATAI_31_), .ZN(n14167) );
  OAI22_X1 U17528 ( .A1(n14167), .A2(n20304), .B1(n19367), .B2(n20306), .ZN(
        n20764) );
  INV_X1 U17529 ( .A(n20764), .ZN(n20833) );
  NAND2_X1 U17530 ( .A1(n14168), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14171) );
  INV_X1 U17531 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n19363) );
  INV_X1 U17532 ( .A(DATAI_23_), .ZN(n21021) );
  NOR2_X2 U17533 ( .A1(n20273), .A2(n14169), .ZN(n20824) );
  AOI22_X1 U17534 ( .A1(n20334), .A2(n20827), .B1(n20294), .B2(n20824), .ZN(
        n14170) );
  OAI211_X1 U17535 ( .C1(n20803), .C2(n20833), .A(n14171), .B(n14170), .ZN(
        n14172) );
  AOI21_X1 U17536 ( .B1(n20826), .B2(n20307), .A(n14172), .ZN(n14173) );
  INV_X1 U17537 ( .A(n14173), .ZN(P1_U3040) );
  INV_X1 U17538 ( .A(n14174), .ZN(n14175) );
  OAI21_X1 U17539 ( .B1(n14122), .B2(n14176), .A(n14175), .ZN(n15223) );
  NAND2_X1 U17540 ( .A1(n16266), .A2(n14177), .ZN(n14178) );
  OAI21_X1 U17541 ( .B1(n14179), .B2(n19217), .A(n14178), .ZN(n14182) );
  INV_X1 U17542 ( .A(n19200), .ZN(n15323) );
  INV_X1 U17543 ( .A(n19197), .ZN(n15321) );
  INV_X1 U17544 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14180) );
  OAI22_X1 U17545 ( .A1(n15323), .A2(n20277), .B1(n15321), .B2(n14180), .ZN(
        n14181) );
  AOI211_X1 U17546 ( .C1(n19198), .C2(n19080), .A(n14182), .B(n14181), .ZN(
        n14183) );
  OAI21_X1 U17547 ( .B1(n15223), .B2(n15327), .A(n14183), .ZN(P2_U2902) );
  XOR2_X1 U17548 ( .A(n14184), .B(n14147), .Z(n14787) );
  AND2_X1 U17549 ( .A1(n16147), .A2(n14185), .ZN(n14186) );
  OR2_X1 U17550 ( .A1(n15960), .A2(n14186), .ZN(n14198) );
  OAI22_X1 U17551 ( .A1(n14198), .A2(n14521), .B1(n21154), .B2(n20179), .ZN(
        n14187) );
  AOI21_X1 U17552 ( .B1(n14787), .B2(n20176), .A(n14187), .ZN(n14188) );
  INV_X1 U17553 ( .A(n14188), .ZN(P1_U2862) );
  XNOR2_X1 U17554 ( .A(n14729), .B(n16152), .ZN(n14189) );
  XNOR2_X1 U17555 ( .A(n14190), .B(n14189), .ZN(n16149) );
  NAND2_X1 U17556 ( .A1(n16149), .A2(n11296), .ZN(n14194) );
  INV_X1 U17557 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14191) );
  OAI22_X1 U17558 ( .A1(n16029), .A2(n20097), .B1(n16162), .B2(n14191), .ZN(
        n14192) );
  AOI21_X1 U17559 ( .B1(n16024), .B2(n20096), .A(n14192), .ZN(n14193) );
  OAI211_X1 U17560 ( .C1(n13814), .C2(n20163), .A(n14194), .B(n14193), .ZN(
        P1_U2990) );
  INV_X1 U17561 ( .A(n14787), .ZN(n14204) );
  AOI22_X1 U17562 ( .A1(n14622), .A2(n20235), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15974), .ZN(n14195) );
  OAI21_X1 U17563 ( .B1(n14204), .B2(n14624), .A(n14195), .ZN(P1_U2894) );
  AOI21_X1 U17564 ( .B1(n20115), .B2(n14196), .A(n14191), .ZN(n20105) );
  NOR2_X1 U17565 ( .A1(n14197), .A2(n20106), .ZN(n15964) );
  OAI21_X1 U17566 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n20105), .A(n15964), 
        .ZN(n14203) );
  INV_X1 U17567 ( .A(n14198), .ZN(n16138) );
  NOR2_X1 U17568 ( .A1(n20107), .A2(n21154), .ZN(n14199) );
  AOI211_X1 U17569 ( .C1(n20139), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20138), .B(n14199), .ZN(n14200) );
  OAI21_X1 U17570 ( .B1(n14785), .B2(n20142), .A(n14200), .ZN(n14201) );
  AOI21_X1 U17571 ( .B1(n16138), .B2(n20130), .A(n14201), .ZN(n14202) );
  OAI211_X1 U17572 ( .C1(n14204), .C2(n20099), .A(n14203), .B(n14202), .ZN(
        P1_U2830) );
  NAND3_X1 U17573 ( .A1(n15818), .A2(n17307), .A3(n18783), .ZN(n18304) );
  NOR2_X1 U17574 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18304), .ZN(n14205) );
  NAND2_X1 U17575 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .ZN(n18856) );
  INV_X1 U17576 ( .A(n18856), .ZN(n18857) );
  NAND2_X1 U17577 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18857), .ZN(n18952) );
  OAI21_X1 U17578 ( .B1(n14205), .B2(n18952), .A(n18356), .ZN(n18310) );
  INV_X1 U17579 ( .A(n18310), .ZN(n14207) );
  NOR2_X1 U17580 ( .A1(n18966), .A2(n19007), .ZN(n18855) );
  INV_X1 U17581 ( .A(n18855), .ZN(n17944) );
  AOI22_X1 U17582 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n14206), .B2(n17944), .ZN(n15807) );
  NOR2_X1 U17583 ( .A1(n14207), .A2(n15807), .ZN(n14209) );
  NOR2_X1 U17584 ( .A1(n18954), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18355) );
  OR2_X1 U17585 ( .A1(n18355), .A2(n14207), .ZN(n15805) );
  OR2_X1 U17586 ( .A1(n18613), .A2(n15805), .ZN(n14208) );
  MUX2_X1 U17587 ( .A(n14209), .B(n14208), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AND2_X1 U17588 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17073) );
  INV_X1 U17589 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17035) );
  INV_X1 U17590 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16753) );
  INV_X1 U17591 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16778) );
  INV_X1 U17592 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17176) );
  INV_X1 U17593 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17206) );
  INV_X1 U17594 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17225) );
  INV_X1 U17595 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16648) );
  NOR2_X1 U17596 ( .A1(n16648), .A2(n14210), .ZN(n14211) );
  AND4_X1 U17597 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(n14211), .ZN(n15803) );
  NAND3_X1 U17598 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n15803), .ZN(n15802) );
  INV_X1 U17599 ( .A(n15802), .ZN(n14212) );
  NOR2_X1 U17600 ( .A1(n17393), .A2(n17032), .ZN(n17141) );
  NAND2_X1 U17601 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17141), .ZN(n17129) );
  NAND2_X1 U17602 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17098), .ZN(n17092) );
  NAND2_X1 U17603 ( .A1(n17324), .A2(n17079), .ZN(n17077) );
  OAI21_X1 U17604 ( .B1(n17073), .B2(n17338), .A(n17077), .ZN(n17074) );
  AOI22_X1 U17605 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14213) );
  OAI21_X1 U17606 ( .B1(n11340), .B2(n18340), .A(n14213), .ZN(n14223) );
  AOI22_X1 U17607 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14220) );
  OAI22_X1 U17608 ( .A1(n17307), .A2(n17120), .B1(n11489), .B2(n17114), .ZN(
        n14218) );
  AOI22_X1 U17609 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11331), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14216) );
  AOI22_X1 U17610 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14215) );
  AOI22_X1 U17611 ( .A1(n17276), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14214) );
  NAND3_X1 U17612 ( .A1(n14216), .A2(n14215), .A3(n14214), .ZN(n14217) );
  AOI211_X1 U17613 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n14218), .B(n14217), .ZN(n14219) );
  OAI211_X1 U17614 ( .C1(n17172), .C2(n14221), .A(n14220), .B(n14219), .ZN(
        n14222) );
  AOI211_X1 U17615 ( .C1(n17228), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n14223), .B(n14222), .ZN(n14292) );
  AOI22_X1 U17616 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14224) );
  OAI21_X1 U17617 ( .B1(n17145), .B2(n17258), .A(n14224), .ZN(n14233) );
  AOI22_X1 U17618 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11378), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14231) );
  AOI22_X1 U17619 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14225) );
  OAI21_X1 U17620 ( .B1(n13764), .B2(n18385), .A(n14225), .ZN(n14229) );
  AOI22_X1 U17621 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U17622 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14226) );
  OAI211_X1 U17623 ( .C1(n11489), .C2(n17146), .A(n14227), .B(n14226), .ZN(
        n14228) );
  AOI211_X1 U17624 ( .C1(n17276), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n14229), .B(n14228), .ZN(n14230) );
  OAI211_X1 U17625 ( .C1(n10327), .C2(n18737), .A(n14231), .B(n14230), .ZN(
        n14232) );
  AOI211_X1 U17626 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n14233), .B(n14232), .ZN(n17080) );
  AOI22_X1 U17627 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14234) );
  OAI21_X1 U17628 ( .B1(n15798), .B2(n18568), .A(n14234), .ZN(n14245) );
  AOI22_X1 U17629 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14242) );
  INV_X1 U17630 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14236) );
  AOI22_X1 U17631 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11378), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14235) );
  OAI21_X1 U17632 ( .B1(n17296), .B2(n14236), .A(n14235), .ZN(n14240) );
  AOI22_X1 U17633 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14238) );
  AOI22_X1 U17634 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14237) );
  OAI211_X1 U17635 ( .C1(n11489), .C2(n17301), .A(n14238), .B(n14237), .ZN(
        n14239) );
  AOI211_X1 U17636 ( .C1(n9810), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n14240), .B(n14239), .ZN(n14241) );
  OAI211_X1 U17637 ( .C1(n17172), .C2(n14243), .A(n14242), .B(n14241), .ZN(
        n14244) );
  AOI211_X1 U17638 ( .C1(n11331), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n14245), .B(n14244), .ZN(n17089) );
  AOI22_X1 U17639 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14256) );
  AOI22_X1 U17640 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14247) );
  AOI22_X1 U17641 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14246) );
  OAI211_X1 U17642 ( .C1(n17296), .C2(n14248), .A(n14247), .B(n14246), .ZN(
        n14254) );
  AOI22_X1 U17643 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14252) );
  AOI22_X1 U17644 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14251) );
  AOI22_X1 U17645 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U17646 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n14249) );
  NAND4_X1 U17647 ( .A1(n14252), .A2(n14251), .A3(n14250), .A4(n14249), .ZN(
        n14253) );
  AOI211_X1 U17648 ( .C1(n9809), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n14254), .B(n14253), .ZN(n14255) );
  OAI211_X1 U17649 ( .C1(n17219), .C2(n17203), .A(n14256), .B(n14255), .ZN(
        n17094) );
  AOI22_X1 U17650 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9810), .B1(
        n17243), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14267) );
  AOI22_X1 U17651 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17292), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n15791), .ZN(n14257) );
  OAI21_X1 U17652 ( .B1(n9858), .B2(n14258), .A(n14257), .ZN(n14265) );
  OAI22_X1 U17653 ( .A1(n17057), .A2(n17145), .B1(n17307), .B2(n18354), .ZN(
        n14259) );
  AOI21_X1 U17654 ( .B1(n17298), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n14259), .ZN(n14263) );
  AOI22_X1 U17655 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14262) );
  AOI22_X1 U17656 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17297), .ZN(n14261) );
  AOI22_X1 U17657 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n9804), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14260) );
  NAND4_X1 U17658 ( .A1(n14263), .A2(n14262), .A3(n14261), .A4(n14260), .ZN(
        n14264) );
  AOI211_X1 U17659 ( .C1(n9808), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n14265), .B(n14264), .ZN(n14266) );
  OAI211_X1 U17660 ( .C1(n11489), .C2(n18397), .A(n14267), .B(n14266), .ZN(
        n17095) );
  NAND2_X1 U17661 ( .A1(n17094), .A2(n17095), .ZN(n17093) );
  NOR2_X1 U17662 ( .A1(n17089), .A2(n17093), .ZN(n17086) );
  AOI22_X1 U17663 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11378), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14278) );
  AOI22_X1 U17664 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14268) );
  OAI21_X1 U17665 ( .B1(n10327), .B2(n18730), .A(n14268), .ZN(n14276) );
  AOI22_X1 U17666 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9809), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14273) );
  INV_X1 U17667 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U17668 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14270) );
  AOI22_X1 U17669 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14269) );
  OAI211_X1 U17670 ( .C1(n17296), .C2(n17275), .A(n14270), .B(n14269), .ZN(
        n14271) );
  AOI21_X1 U17671 ( .B1(n9810), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(n14271), .ZN(n14272) );
  OAI211_X1 U17672 ( .C1(n17172), .C2(n14274), .A(n14273), .B(n14272), .ZN(
        n14275) );
  AOI211_X1 U17673 ( .C1(n11331), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n14276), .B(n14275), .ZN(n14277) );
  OAI211_X1 U17674 ( .C1(n11450), .C2(n14279), .A(n14278), .B(n14277), .ZN(
        n17085) );
  NAND2_X1 U17675 ( .A1(n17086), .A2(n17085), .ZN(n17084) );
  NOR2_X1 U17676 ( .A1(n17080), .A2(n17084), .ZN(n17367) );
  AOI22_X1 U17677 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14290) );
  INV_X1 U17678 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U17679 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14281) );
  AOI22_X1 U17680 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14280) );
  OAI211_X1 U17681 ( .C1(n11489), .C2(n17248), .A(n14281), .B(n14280), .ZN(
        n14288) );
  AOI22_X1 U17682 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14286) );
  AOI22_X1 U17683 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14285) );
  AOI22_X1 U17684 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14284) );
  NAND2_X1 U17685 ( .A1(n9804), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14283) );
  NAND4_X1 U17686 ( .A1(n14286), .A2(n14285), .A3(n14284), .A4(n14283), .ZN(
        n14287) );
  AOI211_X1 U17687 ( .C1(n17276), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n14288), .B(n14287), .ZN(n14289) );
  OAI211_X1 U17688 ( .C1(n17172), .C2(n14291), .A(n14290), .B(n14289), .ZN(
        n17366) );
  NAND2_X1 U17689 ( .A1(n17367), .A2(n17366), .ZN(n17365) );
  NOR2_X1 U17690 ( .A1(n14292), .A2(n17365), .ZN(n17071) );
  AOI21_X1 U17691 ( .B1(n14292), .B2(n17365), .A(n17071), .ZN(n17360) );
  AOI22_X1 U17692 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17074), .B1(n17341), 
        .B2(n17360), .ZN(n14295) );
  INV_X1 U17693 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14293) );
  INV_X1 U17694 ( .A(n17079), .ZN(n17082) );
  NAND3_X1 U17695 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14293), .A3(n17082), 
        .ZN(n14294) );
  NAND2_X1 U17696 ( .A1(n14295), .A2(n14294), .ZN(P3_U2675) );
  INV_X1 U17697 ( .A(n20144), .ZN(n14309) );
  NAND2_X1 U17698 ( .A1(n14296), .A2(n20157), .ZN(n14308) );
  INV_X1 U17699 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14303) );
  INV_X1 U17700 ( .A(n14297), .ZN(n14298) );
  NAND2_X1 U17701 ( .A1(n20127), .A2(n14298), .ZN(n14302) );
  AOI22_X1 U17702 ( .A1(n14300), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n14299), .ZN(n14301) );
  OAI211_X1 U17703 ( .C1(n20098), .C2(n14303), .A(n14302), .B(n14301), .ZN(
        n14306) );
  OAI22_X1 U17704 ( .A1(n21290), .A2(n20107), .B1(n20155), .B2(n14304), .ZN(
        n14305) );
  NOR2_X1 U17705 ( .A1(n14306), .A2(n14305), .ZN(n14307) );
  OAI211_X1 U17706 ( .C1(n14309), .C2(n13609), .A(n14308), .B(n14307), .ZN(
        P1_U2838) );
  INV_X1 U17707 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14535) );
  MUX2_X1 U17708 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n19316), .Z(n19260) );
  AOI22_X1 U17709 ( .A1(n16266), .A2(n19260), .B1(n19203), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14311) );
  NAND2_X1 U17710 ( .A1(n19197), .A2(BUF2_REG_30__SCAN_IN), .ZN(n14310) );
  OAI211_X1 U17711 ( .C1(n15323), .C2(n14535), .A(n14311), .B(n14310), .ZN(
        n14312) );
  AOI21_X1 U17712 ( .B1(n16210), .B2(n19198), .A(n14312), .ZN(n14313) );
  OAI21_X1 U17713 ( .B1(n14314), .B2(n15327), .A(n14313), .ZN(P2_U2889) );
  INV_X1 U17714 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21256) );
  NAND2_X1 U17715 ( .A1(n20077), .A2(n21256), .ZN(n14316) );
  MUX2_X1 U17716 ( .A(n14316), .B(n14315), .S(n20938), .Z(P1_U3487) );
  INV_X1 U17717 ( .A(n14317), .ZN(n14325) );
  OAI21_X1 U17718 ( .B1(n14340), .B2(n21044), .A(n14626), .ZN(n14324) );
  INV_X1 U17719 ( .A(n14627), .ZN(n14321) );
  OAI22_X1 U17720 ( .A1(n20107), .A2(n14319), .B1(n14318), .B2(n20098), .ZN(
        n14320) );
  AOI21_X1 U17721 ( .B1(n14321), .B2(n20127), .A(n14320), .ZN(n14322) );
  OAI21_X1 U17722 ( .B1(n14818), .B2(n20155), .A(n14322), .ZN(n14323) );
  AOI21_X1 U17723 ( .B1(n14325), .B2(n14324), .A(n14323), .ZN(n14326) );
  OAI21_X1 U17724 ( .B1(n14634), .B2(n20099), .A(n14326), .ZN(P1_U2810) );
  NAND2_X1 U17725 ( .A1(n14638), .A2(n20123), .ZN(n14339) );
  AND2_X1 U17726 ( .A1(n9868), .A2(n14330), .ZN(n14331) );
  INV_X1 U17727 ( .A(n14832), .ZN(n14337) );
  NAND2_X1 U17728 ( .A1(n20115), .A2(n14333), .ZN(n14348) );
  OAI22_X1 U17729 ( .A1(n20107), .A2(n21269), .B1(n14639), .B2(n20098), .ZN(
        n14334) );
  AOI21_X1 U17730 ( .B1(n14641), .B2(n20127), .A(n14334), .ZN(n14335) );
  OAI21_X1 U17731 ( .B1(n21044), .B2(n14348), .A(n14335), .ZN(n14336) );
  AOI21_X1 U17732 ( .B1(n14337), .B2(n20130), .A(n14336), .ZN(n14338) );
  OAI211_X1 U17733 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14340), .A(n14339), 
        .B(n14338), .ZN(P1_U2811) );
  INV_X1 U17734 ( .A(n14655), .ZN(n14548) );
  OR2_X1 U17735 ( .A1(n14356), .A2(n14344), .ZN(n14345) );
  AND2_X1 U17736 ( .A1(n9868), .A2(n14345), .ZN(n14500) );
  INV_X1 U17737 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21268) );
  INV_X1 U17738 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n21153) );
  OAI22_X1 U17739 ( .A1(n20107), .A2(n21153), .B1(n14653), .B2(n20098), .ZN(
        n14346) );
  AOI21_X1 U17740 ( .B1(n14651), .B2(n20127), .A(n14346), .ZN(n14347) );
  OAI21_X1 U17741 ( .B1(n21268), .B2(n14348), .A(n14347), .ZN(n14349) );
  AOI21_X1 U17742 ( .B1(n14500), .B2(n20130), .A(n14349), .ZN(n14351) );
  NAND3_X1 U17743 ( .A1(n14362), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n21268), 
        .ZN(n14350) );
  OAI211_X1 U17744 ( .C1(n14548), .C2(n20099), .A(n14351), .B(n14350), .ZN(
        P1_U2812) );
  OAI21_X1 U17745 ( .B1(n14352), .B2(n14353), .A(n14341), .ZN(n14667) );
  INV_X1 U17746 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21103) );
  NOR2_X1 U17747 ( .A1(n14369), .A2(n14354), .ZN(n14355) );
  OR2_X1 U17748 ( .A1(n14356), .A2(n14355), .ZN(n14850) );
  OAI22_X1 U17749 ( .A1(n20107), .A2(n21125), .B1(n14657), .B2(n20098), .ZN(
        n14357) );
  AOI21_X1 U17750 ( .B1(n14659), .B2(n20127), .A(n14357), .ZN(n14360) );
  NOR2_X1 U17751 ( .A1(n14358), .A2(n20106), .ZN(n14371) );
  NAND2_X1 U17752 ( .A1(n14371), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14359) );
  OAI211_X1 U17753 ( .C1(n14850), .C2(n20155), .A(n14360), .B(n14359), .ZN(
        n14361) );
  AOI21_X1 U17754 ( .B1(n14362), .B2(n21103), .A(n14361), .ZN(n14363) );
  OAI21_X1 U17755 ( .B1(n14667), .B2(n20099), .A(n14363), .ZN(P1_U2813) );
  INV_X1 U17756 ( .A(n14352), .ZN(n14366) );
  AND2_X1 U17757 ( .A1(n9857), .A2(n14368), .ZN(n14370) );
  OR2_X1 U17758 ( .A1(n14370), .A2(n14369), .ZN(n16040) );
  INV_X1 U17759 ( .A(n16040), .ZN(n14376) );
  NAND2_X1 U17760 ( .A1(n14371), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14373) );
  AOI22_X1 U17761 ( .A1(n20152), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20139), .ZN(n14372) );
  OAI211_X1 U17762 ( .C1(n20142), .C2(n14668), .A(n14373), .B(n14372), .ZN(
        n14375) );
  NOR4_X1 U17763 ( .A1(n14393), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n20883), 
        .A4(n20879), .ZN(n14374) );
  AOI211_X1 U17764 ( .C1(n14376), .C2(n20130), .A(n14375), .B(n14374), .ZN(
        n14377) );
  OAI21_X1 U17765 ( .B1(n14675), .B2(n20099), .A(n14377), .ZN(P1_U2814) );
  AOI21_X1 U17766 ( .B1(n14379), .B2(n14378), .A(n14365), .ZN(n14685) );
  XNOR2_X1 U17767 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14380) );
  NOR2_X1 U17768 ( .A1(n14393), .A2(n14380), .ZN(n14388) );
  NAND2_X1 U17769 ( .A1(n14396), .A2(n14381), .ZN(n14382) );
  NAND2_X1 U17770 ( .A1(n9857), .A2(n14382), .ZN(n14860) );
  OAI22_X1 U17771 ( .A1(n20107), .A2(n21107), .B1(n14683), .B2(n20098), .ZN(
        n14383) );
  AOI21_X1 U17772 ( .B1(n14681), .B2(n20127), .A(n14383), .ZN(n14386) );
  NAND2_X1 U17773 ( .A1(n14384), .A2(n20115), .ZN(n14417) );
  OR2_X1 U17774 ( .A1(n14417), .A2(n20883), .ZN(n14385) );
  OAI211_X1 U17775 ( .C1(n14860), .C2(n20155), .A(n14386), .B(n14385), .ZN(
        n14387) );
  AOI211_X1 U17776 ( .C1(n14685), .C2(n20123), .A(n14388), .B(n14387), .ZN(
        n14389) );
  INV_X1 U17777 ( .A(n14389), .ZN(P1_U2815) );
  INV_X1 U17778 ( .A(n14378), .ZN(n14391) );
  AOI21_X1 U17779 ( .B1(n14392), .B2(n14390), .A(n14391), .ZN(n14691) );
  INV_X1 U17780 ( .A(n14691), .ZN(n14570) );
  INV_X1 U17781 ( .A(n14393), .ZN(n14401) );
  OR2_X1 U17782 ( .A1(n14411), .A2(n14394), .ZN(n14395) );
  NAND2_X1 U17783 ( .A1(n14396), .A2(n14395), .ZN(n14874) );
  INV_X1 U17784 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21293) );
  OAI22_X1 U17785 ( .A1(n20107), .A2(n21293), .B1(n14692), .B2(n20098), .ZN(
        n14397) );
  AOI21_X1 U17786 ( .B1(n14694), .B2(n20127), .A(n14397), .ZN(n14399) );
  OR2_X1 U17787 ( .A1(n14417), .A2(n20879), .ZN(n14398) );
  OAI211_X1 U17788 ( .C1(n14874), .C2(n20155), .A(n14399), .B(n14398), .ZN(
        n14400) );
  AOI21_X1 U17789 ( .B1(n14401), .B2(n20879), .A(n14400), .ZN(n14402) );
  OAI21_X1 U17790 ( .B1(n14570), .B2(n20099), .A(n14402), .ZN(P1_U2816) );
  AOI21_X1 U17791 ( .B1(n14431), .B2(n14403), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14418) );
  INV_X1 U17792 ( .A(n14405), .ZN(n14407) );
  INV_X1 U17793 ( .A(n14390), .ZN(n14406) );
  NAND2_X1 U17794 ( .A1(n14702), .A2(n20123), .ZN(n14416) );
  OAI22_X1 U17795 ( .A1(n20107), .A2(n21330), .B1(n14409), .B2(n20098), .ZN(
        n14414) );
  AND2_X1 U17796 ( .A1(n14425), .A2(n14410), .ZN(n14412) );
  OR2_X1 U17797 ( .A1(n14412), .A2(n14411), .ZN(n16048) );
  NOR2_X1 U17798 ( .A1(n16048), .A2(n20155), .ZN(n14413) );
  AOI211_X1 U17799 ( .C1(n20127), .C2(n14698), .A(n14414), .B(n14413), .ZN(
        n14415) );
  OAI211_X1 U17800 ( .C1(n14418), .C2(n14417), .A(n14416), .B(n14415), .ZN(
        P1_U2817) );
  INV_X1 U17801 ( .A(n14419), .ZN(n14420) );
  AOI21_X1 U17802 ( .B1(n14420), .B2(n14438), .A(n14421), .ZN(n14422) );
  NOR2_X1 U17803 ( .A1(n14422), .A2(n14405), .ZN(n14710) );
  INV_X1 U17804 ( .A(n14710), .ZN(n14502) );
  NAND2_X1 U17805 ( .A1(n14441), .A2(n14423), .ZN(n14424) );
  NAND2_X1 U17806 ( .A1(n14425), .A2(n14424), .ZN(n16059) );
  INV_X1 U17807 ( .A(n16059), .ZN(n14429) );
  AOI22_X1 U17808 ( .A1(n20152), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20139), .ZN(n14426) );
  OAI21_X1 U17809 ( .B1(n20142), .B2(n14708), .A(n14426), .ZN(n14428) );
  INV_X1 U17810 ( .A(n14431), .ZN(n14487) );
  INV_X1 U17811 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21018) );
  NOR4_X1 U17812 ( .A1(n14487), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n14434), 
        .A4(n21018), .ZN(n14427) );
  AOI211_X1 U17813 ( .C1(n14429), .C2(n20130), .A(n14428), .B(n14427), .ZN(
        n14437) );
  NOR2_X1 U17814 ( .A1(n14434), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14430) );
  AND2_X1 U17815 ( .A1(n14431), .A2(n14430), .ZN(n14447) );
  OAI21_X1 U17816 ( .B1(n14433), .B2(n14432), .A(n20115), .ZN(n15919) );
  NAND2_X1 U17817 ( .A1(n20115), .A2(n14434), .ZN(n14435) );
  NAND2_X1 U17818 ( .A1(n15919), .A2(n14435), .ZN(n14456) );
  OAI21_X1 U17819 ( .B1(n14447), .B2(n14456), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14436) );
  OAI211_X1 U17820 ( .C1(n14502), .C2(n20099), .A(n14437), .B(n14436), .ZN(
        P1_U2818) );
  XNOR2_X1 U17821 ( .A(n14420), .B(n14438), .ZN(n14719) );
  NAND2_X1 U17822 ( .A1(n14453), .A2(n14439), .ZN(n14440) );
  NAND2_X1 U17823 ( .A1(n14441), .A2(n14440), .ZN(n14879) );
  INV_X1 U17824 ( .A(n14716), .ZN(n14444) );
  INV_X1 U17825 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n21164) );
  OAI22_X1 U17826 ( .A1(n20107), .A2(n21164), .B1(n14442), .B2(n20098), .ZN(
        n14443) );
  AOI21_X1 U17827 ( .B1(n14444), .B2(n20127), .A(n14443), .ZN(n14445) );
  OAI21_X1 U17828 ( .B1(n14879), .B2(n20155), .A(n14445), .ZN(n14446) );
  AOI21_X1 U17829 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n14456), .A(n14446), 
        .ZN(n14449) );
  INV_X1 U17830 ( .A(n14447), .ZN(n14448) );
  OAI211_X1 U17831 ( .C1(n14719), .C2(n20099), .A(n14449), .B(n14448), .ZN(
        P1_U2819) );
  INV_X1 U17832 ( .A(n9875), .ZN(n14461) );
  AOI21_X1 U17833 ( .B1(n14450), .B2(n14461), .A(n14420), .ZN(n14585) );
  INV_X1 U17834 ( .A(n14585), .ZN(n14724) );
  INV_X1 U17835 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n21082) );
  OAI22_X1 U17836 ( .A1(n20107), .A2(n21082), .B1(n14723), .B2(n20098), .ZN(
        n14455) );
  OR2_X1 U17837 ( .A1(n14465), .A2(n14451), .ZN(n14452) );
  NAND2_X1 U17838 ( .A1(n14453), .A2(n14452), .ZN(n15896) );
  NOR2_X1 U17839 ( .A1(n15896), .A2(n20155), .ZN(n14454) );
  AOI211_X1 U17840 ( .C1(n20127), .C2(n14727), .A(n14455), .B(n14454), .ZN(
        n14459) );
  INV_X1 U17841 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21041) );
  INV_X1 U17842 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21039) );
  NOR3_X1 U17843 ( .A1(n14487), .A2(n21041), .A3(n21039), .ZN(n14457) );
  OAI21_X1 U17844 ( .B1(n14457), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14456), 
        .ZN(n14458) );
  OAI211_X1 U17845 ( .C1(n14724), .C2(n20099), .A(n14459), .B(n14458), .ZN(
        P1_U2820) );
  INV_X1 U17846 ( .A(n14460), .ZN(n14462) );
  OAI21_X1 U17847 ( .B1(n9837), .B2(n14462), .A(n14461), .ZN(n14733) );
  INV_X1 U17848 ( .A(n15919), .ZN(n14484) );
  AND2_X1 U17849 ( .A1(n9832), .A2(n14463), .ZN(n14464) );
  NOR2_X1 U17850 ( .A1(n14465), .A2(n14464), .ZN(n16061) );
  INV_X1 U17851 ( .A(n16061), .ZN(n14469) );
  NAND2_X1 U17852 ( .A1(n20152), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n14466) );
  OAI211_X1 U17853 ( .C1(n20098), .C2(n14732), .A(n14466), .B(n20134), .ZN(
        n14467) );
  AOI21_X1 U17854 ( .B1(n14736), .B2(n20127), .A(n14467), .ZN(n14468) );
  OAI21_X1 U17855 ( .B1(n14469), .B2(n20155), .A(n14468), .ZN(n14472) );
  XNOR2_X1 U17856 ( .A(P1_REIP_REG_19__SCAN_IN), .B(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14470) );
  NOR2_X1 U17857 ( .A1(n14487), .A2(n14470), .ZN(n14471) );
  AOI211_X1 U17858 ( .C1(n14484), .C2(P1_REIP_REG_19__SCAN_IN), .A(n14472), 
        .B(n14471), .ZN(n14473) );
  OAI21_X1 U17859 ( .B1(n14733), .B2(n20099), .A(n14473), .ZN(P1_U2821) );
  INV_X1 U17860 ( .A(n14474), .ZN(n14476) );
  NAND2_X1 U17861 ( .A1(n14745), .A2(n20123), .ZN(n14486) );
  NAND2_X1 U17862 ( .A1(n9909), .A2(n14477), .ZN(n14478) );
  NAND2_X1 U17863 ( .A1(n9832), .A2(n14478), .ZN(n16079) );
  INV_X1 U17864 ( .A(n14743), .ZN(n14481) );
  NAND2_X1 U17865 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n20139), .ZN(
        n14479) );
  OAI211_X1 U17866 ( .C1(n20107), .C2(n21308), .A(n14479), .B(n20134), .ZN(
        n14480) );
  AOI21_X1 U17867 ( .B1(n14481), .B2(n20127), .A(n14480), .ZN(n14482) );
  OAI21_X1 U17868 ( .B1(n16079), .B2(n20155), .A(n14482), .ZN(n14483) );
  AOI21_X1 U17869 ( .B1(n14484), .B2(P1_REIP_REG_18__SCAN_IN), .A(n14483), 
        .ZN(n14485) );
  OAI211_X1 U17870 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n14487), .A(n14486), 
        .B(n14485), .ZN(P1_U2822) );
  OAI21_X1 U17871 ( .B1(n10835), .B2(n10834), .A(n14490), .ZN(n14763) );
  INV_X1 U17872 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21122) );
  NOR2_X1 U17873 ( .A1(n14491), .A2(n20106), .ZN(n15936) );
  AOI22_X1 U17874 ( .A1(n15936), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n20152), 
        .B2(P1_EBX_REG_15__SCAN_IN), .ZN(n14492) );
  OAI211_X1 U17875 ( .C1(n20098), .C2(n14493), .A(n14492), .B(n20134), .ZN(
        n14494) );
  AOI21_X1 U17876 ( .B1(n15921), .B2(n21122), .A(n14494), .ZN(n14499) );
  NOR2_X1 U17877 ( .A1(n14519), .A2(n14495), .ZN(n14496) );
  OR2_X1 U17878 ( .A1(n15923), .A2(n14496), .ZN(n16101) );
  OAI22_X1 U17879 ( .A1(n16101), .A2(n20155), .B1(n14765), .B2(n20142), .ZN(
        n14497) );
  INV_X1 U17880 ( .A(n14497), .ZN(n14498) );
  OAI211_X1 U17881 ( .C1(n14763), .C2(n20099), .A(n14499), .B(n14498), .ZN(
        P1_U2825) );
  OAI22_X1 U17882 ( .A1(n14790), .A2(n14521), .B1(n20179), .B2(n21166), .ZN(
        P1_U2841) );
  INV_X1 U17883 ( .A(n14638), .ZN(n14543) );
  OAI222_X1 U17884 ( .A1(n14532), .A2(n14543), .B1(n21269), .B2(n20179), .C1(
        n14832), .C2(n14521), .ZN(P1_U2843) );
  INV_X1 U17885 ( .A(n14500), .ZN(n14841) );
  OAI222_X1 U17886 ( .A1(n14841), .A2(n14521), .B1(n21153), .B2(n20179), .C1(
        n14548), .C2(n14532), .ZN(P1_U2844) );
  OAI222_X1 U17887 ( .A1(n14532), .A2(n14667), .B1(n21125), .B2(n20179), .C1(
        n14850), .C2(n14521), .ZN(P1_U2845) );
  OAI222_X1 U17888 ( .A1(n16040), .A2(n14521), .B1(n21086), .B2(n20179), .C1(
        n14675), .C2(n14532), .ZN(P1_U2846) );
  INV_X1 U17889 ( .A(n14685), .ZN(n14563) );
  OAI222_X1 U17890 ( .A1(n14532), .A2(n14563), .B1(n21107), .B2(n20179), .C1(
        n14860), .C2(n14521), .ZN(P1_U2847) );
  OAI222_X1 U17891 ( .A1(n14532), .A2(n14570), .B1(n21293), .B2(n20179), .C1(
        n14874), .C2(n14521), .ZN(P1_U2848) );
  INV_X1 U17892 ( .A(n14702), .ZN(n14501) );
  OAI222_X1 U17893 ( .A1(n16048), .A2(n14521), .B1(n21330), .B2(n20179), .C1(
        n14501), .C2(n14532), .ZN(P1_U2849) );
  INV_X1 U17894 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n21287) );
  OAI222_X1 U17895 ( .A1(n16059), .A2(n14521), .B1(n21287), .B2(n20179), .C1(
        n14502), .C2(n14532), .ZN(P1_U2850) );
  OAI222_X1 U17896 ( .A1(n14879), .A2(n14521), .B1(n21164), .B2(n20179), .C1(
        n14532), .C2(n14719), .ZN(P1_U2851) );
  OAI222_X1 U17897 ( .A1(n14724), .A2(n14532), .B1(n21082), .B2(n20179), .C1(
        n15896), .C2(n14521), .ZN(P1_U2852) );
  AOI22_X1 U17898 ( .A1(n16061), .A2(n20175), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14530), .ZN(n14503) );
  OAI21_X1 U17899 ( .B1(n14733), .B2(n14532), .A(n14503), .ZN(P1_U2853) );
  OAI22_X1 U17900 ( .A1(n16079), .A2(n14521), .B1(n21308), .B2(n20179), .ZN(
        n14504) );
  AOI21_X1 U17901 ( .B1(n14745), .B2(n20176), .A(n14504), .ZN(n14505) );
  INV_X1 U17902 ( .A(n14505), .ZN(P1_U2854) );
  AND2_X1 U17903 ( .A1(n14506), .A2(n14507), .ZN(n14508) );
  OR2_X1 U17904 ( .A1(n14508), .A2(n14475), .ZN(n15915) );
  INV_X1 U17905 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14513) );
  NAND2_X1 U17906 ( .A1(n15923), .A2(n14509), .ZN(n14511) );
  NAND2_X1 U17907 ( .A1(n14511), .A2(n14510), .ZN(n14512) );
  NAND2_X1 U17908 ( .A1(n14512), .A2(n9909), .ZN(n16087) );
  OAI222_X1 U17909 ( .A1(n15915), .A2(n14532), .B1(n14513), .B2(n20179), .C1(
        n14521), .C2(n16087), .ZN(P1_U2855) );
  INV_X1 U17910 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14514) );
  OAI222_X1 U17911 ( .A1(n16101), .A2(n14521), .B1(n14514), .B2(n20179), .C1(
        n14763), .C2(n14532), .ZN(P1_U2857) );
  OR2_X1 U17912 ( .A1(n14515), .A2(n14516), .ZN(n14517) );
  AND2_X1 U17913 ( .A1(n14488), .A2(n14517), .ZN(n15997) );
  AND2_X1 U17914 ( .A1(n14528), .A2(n14518), .ZN(n14520) );
  OR2_X1 U17915 ( .A1(n14520), .A2(n14519), .ZN(n16116) );
  OAI22_X1 U17916 ( .A1(n16116), .A2(n14521), .B1(n21038), .B2(n20179), .ZN(
        n14522) );
  AOI21_X1 U17917 ( .B1(n15997), .B2(n20176), .A(n14522), .ZN(n14523) );
  INV_X1 U17918 ( .A(n14523), .ZN(P1_U2858) );
  AOI21_X1 U17919 ( .B1(n14525), .B2(n14524), .A(n14515), .ZN(n14526) );
  INV_X1 U17920 ( .A(n14526), .ZN(n15944) );
  OAI21_X1 U17921 ( .B1(n15958), .B2(n14903), .A(n14527), .ZN(n14529) );
  AND2_X1 U17922 ( .A1(n14529), .A2(n14528), .ZN(n16117) );
  AOI22_X1 U17923 ( .A1(n16117), .A2(n20175), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14530), .ZN(n14531) );
  OAI21_X1 U17924 ( .B1(n15944), .B2(n14532), .A(n14531), .ZN(P1_U2859) );
  NAND2_X1 U17925 ( .A1(n15977), .A2(DATAI_30_), .ZN(n14534) );
  AOI22_X1 U17926 ( .A1(n15976), .A2(n20247), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n15974), .ZN(n14533) );
  OAI211_X1 U17927 ( .C1(n15981), .C2(n14535), .A(n14534), .B(n14533), .ZN(
        n14536) );
  INV_X1 U17928 ( .A(n14536), .ZN(n14537) );
  OAI21_X1 U17929 ( .B1(n14634), .B2(n14624), .A(n14537), .ZN(P1_U2874) );
  INV_X1 U17930 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14540) );
  NAND2_X1 U17931 ( .A1(n15977), .A2(DATAI_29_), .ZN(n14539) );
  AOI22_X1 U17932 ( .A1(n15976), .A2(n20244), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15974), .ZN(n14538) );
  OAI211_X1 U17933 ( .C1(n15981), .C2(n14540), .A(n14539), .B(n14538), .ZN(
        n14541) );
  INV_X1 U17934 ( .A(n14541), .ZN(n14542) );
  OAI21_X1 U17935 ( .B1(n14543), .B2(n14624), .A(n14542), .ZN(P1_U2875) );
  NAND2_X1 U17936 ( .A1(n15977), .A2(DATAI_28_), .ZN(n14545) );
  AOI22_X1 U17937 ( .A1(n15976), .A2(n20241), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n15974), .ZN(n14544) );
  OAI211_X1 U17938 ( .C1(n15981), .C2(n16537), .A(n14545), .B(n14544), .ZN(
        n14546) );
  INV_X1 U17939 ( .A(n14546), .ZN(n14547) );
  OAI21_X1 U17940 ( .B1(n14548), .B2(n14624), .A(n14547), .ZN(P1_U2876) );
  INV_X1 U17941 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n14551) );
  NAND2_X1 U17942 ( .A1(n15977), .A2(DATAI_27_), .ZN(n14550) );
  AOI22_X1 U17943 ( .A1(n15976), .A2(n20238), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15974), .ZN(n14549) );
  OAI211_X1 U17944 ( .C1(n15981), .C2(n14551), .A(n14550), .B(n14549), .ZN(
        n14552) );
  INV_X1 U17945 ( .A(n14552), .ZN(n14553) );
  OAI21_X1 U17946 ( .B1(n14667), .B2(n14624), .A(n14553), .ZN(P1_U2877) );
  INV_X1 U17947 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n15260) );
  NAND2_X1 U17948 ( .A1(n15977), .A2(DATAI_26_), .ZN(n14555) );
  AOI22_X1 U17949 ( .A1(n15976), .A2(n20235), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n15974), .ZN(n14554) );
  OAI211_X1 U17950 ( .C1(n15981), .C2(n15260), .A(n14555), .B(n14554), .ZN(
        n14556) );
  INV_X1 U17951 ( .A(n14556), .ZN(n14557) );
  OAI21_X1 U17952 ( .B1(n14675), .B2(n14624), .A(n14557), .ZN(P1_U2878) );
  INV_X1 U17953 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14560) );
  NAND2_X1 U17954 ( .A1(n15977), .A2(DATAI_25_), .ZN(n14559) );
  AOI22_X1 U17955 ( .A1(n15976), .A2(n20232), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n15974), .ZN(n14558) );
  OAI211_X1 U17956 ( .C1(n14560), .C2(n15981), .A(n14559), .B(n14558), .ZN(
        n14561) );
  INV_X1 U17957 ( .A(n14561), .ZN(n14562) );
  OAI21_X1 U17958 ( .B1(n14563), .B2(n14624), .A(n14562), .ZN(P1_U2879) );
  INV_X1 U17959 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14567) );
  NAND2_X1 U17960 ( .A1(n15977), .A2(DATAI_24_), .ZN(n14566) );
  AOI22_X1 U17961 ( .A1(n15976), .A2(n14564), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n15974), .ZN(n14565) );
  OAI211_X1 U17962 ( .C1(n14567), .C2(n15981), .A(n14566), .B(n14565), .ZN(
        n14568) );
  INV_X1 U17963 ( .A(n14568), .ZN(n14569) );
  OAI21_X1 U17964 ( .B1(n14570), .B2(n14624), .A(n14569), .ZN(P1_U2880) );
  NAND2_X1 U17965 ( .A1(n14702), .A2(n15978), .ZN(n14574) );
  NAND2_X1 U17966 ( .A1(n15974), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n14571) );
  OAI21_X1 U17967 ( .B1(n14597), .B2(n20231), .A(n14571), .ZN(n14572) );
  AOI21_X1 U17968 ( .B1(n15977), .B2(DATAI_23_), .A(n14572), .ZN(n14573) );
  OAI211_X1 U17969 ( .C1(n15981), .C2(n19363), .A(n14574), .B(n14573), .ZN(
        P1_U2881) );
  INV_X1 U17970 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14579) );
  NAND2_X1 U17971 ( .A1(n14710), .A2(n15978), .ZN(n14578) );
  NAND2_X1 U17972 ( .A1(n15974), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n14575) );
  OAI21_X1 U17973 ( .B1(n14597), .B2(n20303), .A(n14575), .ZN(n14576) );
  AOI21_X1 U17974 ( .B1(n15977), .B2(DATAI_22_), .A(n14576), .ZN(n14577) );
  OAI211_X1 U17975 ( .C1(n15981), .C2(n14579), .A(n14578), .B(n14577), .ZN(
        P1_U2882) );
  INV_X1 U17976 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20296) );
  NAND2_X1 U17977 ( .A1(n15977), .A2(DATAI_21_), .ZN(n14582) );
  INV_X1 U17978 ( .A(n20295), .ZN(n14580) );
  AOI22_X1 U17979 ( .A1(n15976), .A2(n14580), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n15974), .ZN(n14581) );
  OAI211_X1 U17980 ( .C1(n20296), .C2(n15981), .A(n14582), .B(n14581), .ZN(
        n14583) );
  INV_X1 U17981 ( .A(n14583), .ZN(n14584) );
  OAI21_X1 U17982 ( .B1(n14719), .B2(n14624), .A(n14584), .ZN(P1_U2883) );
  NAND2_X1 U17983 ( .A1(n14585), .A2(n15978), .ZN(n14589) );
  NAND2_X1 U17984 ( .A1(n15974), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n14586) );
  OAI21_X1 U17985 ( .B1(n14597), .B2(n20227), .A(n14586), .ZN(n14587) );
  AOI21_X1 U17986 ( .B1(n15977), .B2(DATAI_20_), .A(n14587), .ZN(n14588) );
  OAI211_X1 U17987 ( .C1(n15981), .C2(n19346), .A(n14589), .B(n14588), .ZN(
        P1_U2884) );
  INV_X1 U17988 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14593) );
  NAND2_X1 U17989 ( .A1(n15977), .A2(DATAI_19_), .ZN(n14592) );
  INV_X1 U17990 ( .A(n20288), .ZN(n14590) );
  AOI22_X1 U17991 ( .A1(n15976), .A2(n14590), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15974), .ZN(n14591) );
  OAI211_X1 U17992 ( .C1(n14593), .C2(n15981), .A(n14592), .B(n14591), .ZN(
        n14594) );
  INV_X1 U17993 ( .A(n14594), .ZN(n14595) );
  OAI21_X1 U17994 ( .B1(n14733), .B2(n14624), .A(n14595), .ZN(P1_U2885) );
  INV_X1 U17995 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n15322) );
  NAND2_X1 U17996 ( .A1(n14745), .A2(n15978), .ZN(n14600) );
  NAND2_X1 U17997 ( .A1(n15974), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n14596) );
  OAI21_X1 U17998 ( .B1(n14597), .B2(n20283), .A(n14596), .ZN(n14598) );
  AOI21_X1 U17999 ( .B1(n15977), .B2(DATAI_18_), .A(n14598), .ZN(n14599) );
  OAI211_X1 U18000 ( .C1(n15981), .C2(n15322), .A(n14600), .B(n14599), .ZN(
        P1_U2886) );
  NAND2_X1 U18001 ( .A1(n15977), .A2(DATAI_17_), .ZN(n14603) );
  INV_X1 U18002 ( .A(n20276), .ZN(n14601) );
  AOI22_X1 U18003 ( .A1(n15976), .A2(n14601), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n15974), .ZN(n14602) );
  OAI211_X1 U18004 ( .C1(n20277), .C2(n15981), .A(n14603), .B(n14602), .ZN(
        n14604) );
  INV_X1 U18005 ( .A(n14604), .ZN(n14605) );
  OAI21_X1 U18006 ( .B1(n15915), .B2(n14624), .A(n14605), .ZN(P1_U2887) );
  INV_X1 U18007 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20182) );
  INV_X1 U18008 ( .A(DATAI_15_), .ZN(n14606) );
  NOR2_X1 U18009 ( .A1(n14607), .A2(n14606), .ZN(n14608) );
  AOI21_X1 U18010 ( .B1(n14609), .B2(BUF1_REG_15__SCAN_IN), .A(n14608), .ZN(
        n20254) );
  OAI222_X1 U18011 ( .A1(n14763), .A2(n14624), .B1(n14611), .B2(n20182), .C1(
        n14610), .C2(n20254), .ZN(P1_U2889) );
  INV_X1 U18012 ( .A(n15997), .ZN(n14613) );
  AOI22_X1 U18013 ( .A1(n14622), .A2(n20247), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15974), .ZN(n14612) );
  OAI21_X1 U18014 ( .B1(n14613), .B2(n14624), .A(n14612), .ZN(P1_U2890) );
  AOI22_X1 U18015 ( .A1(n14622), .A2(n20244), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15974), .ZN(n14614) );
  OAI21_X1 U18016 ( .B1(n15944), .B2(n14624), .A(n14614), .ZN(P1_U2891) );
  OAI21_X1 U18017 ( .B1(n14615), .B2(n14616), .A(n14524), .ZN(n15950) );
  AOI22_X1 U18018 ( .A1(n14622), .A2(n20241), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15974), .ZN(n14617) );
  OAI21_X1 U18019 ( .B1(n15950), .B2(n14624), .A(n14617), .ZN(P1_U2892) );
  INV_X1 U18020 ( .A(n14619), .ZN(n14620) );
  AOI21_X1 U18021 ( .B1(n14621), .B2(n14618), .A(n14620), .ZN(n16011) );
  INV_X1 U18022 ( .A(n16011), .ZN(n14625) );
  AOI22_X1 U18023 ( .A1(n14622), .A2(n20238), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15974), .ZN(n14623) );
  OAI21_X1 U18024 ( .B1(n14625), .B2(n14624), .A(n14623), .ZN(P1_U2893) );
  NOR2_X1 U18025 ( .A1(n16162), .A2(n14626), .ZN(n14819) );
  NOR2_X1 U18026 ( .A1(n16022), .A2(n14627), .ZN(n14628) );
  AOI211_X1 U18027 ( .C1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n16015), .A(
        n14819), .B(n14628), .ZN(n14633) );
  XNOR2_X1 U18028 ( .A(n14631), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14817) );
  NAND2_X1 U18029 ( .A1(n14817), .A2(n11296), .ZN(n14632) );
  OAI211_X1 U18030 ( .C1(n14634), .C2(n13814), .A(n14633), .B(n14632), .ZN(
        P1_U2969) );
  MUX2_X1 U18031 ( .A(n14751), .B(n14636), .S(n14635), .Z(n14637) );
  INV_X1 U18032 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14828) );
  XNOR2_X1 U18033 ( .A(n14637), .B(n14828), .ZN(n14837) );
  NAND2_X1 U18034 ( .A1(n14638), .A2(n16025), .ZN(n14643) );
  NOR2_X1 U18035 ( .A1(n16162), .A2(n21044), .ZN(n14830) );
  NOR2_X1 U18036 ( .A1(n16029), .A2(n14639), .ZN(n14640) );
  AOI211_X1 U18037 ( .C1(n14641), .C2(n16024), .A(n14830), .B(n14640), .ZN(
        n14642) );
  OAI211_X1 U18038 ( .C1(n20080), .C2(n14837), .A(n14643), .B(n14642), .ZN(
        P1_U2970) );
  NOR3_X1 U18039 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14644) );
  NAND4_X1 U18040 ( .A1(n14751), .A2(n14644), .A3(n14871), .A4(n16042), .ZN(
        n14648) );
  NAND3_X1 U18041 ( .A1(n14729), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14647) );
  INV_X1 U18042 ( .A(n14645), .ZN(n14687) );
  AOI21_X1 U18043 ( .B1(n14729), .B2(n14805), .A(n14687), .ZN(n14646) );
  MUX2_X1 U18044 ( .A(n14648), .B(n14647), .S(n14646), .Z(n14650) );
  XNOR2_X1 U18045 ( .A(n14650), .B(n14649), .ZN(n14846) );
  NAND2_X1 U18046 ( .A1(n16024), .A2(n14651), .ZN(n14652) );
  NAND2_X1 U18047 ( .A1(n16174), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14840) );
  OAI211_X1 U18048 ( .C1(n16029), .C2(n14653), .A(n14652), .B(n14840), .ZN(
        n14654) );
  AOI21_X1 U18049 ( .B1(n14655), .B2(n16025), .A(n14654), .ZN(n14656) );
  OAI21_X1 U18050 ( .B1(n14846), .B2(n20080), .A(n14656), .ZN(P1_U2971) );
  NAND2_X1 U18051 ( .A1(n16174), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14849) );
  OAI21_X1 U18052 ( .B1(n16029), .B2(n14657), .A(n14849), .ZN(n14658) );
  AOI21_X1 U18053 ( .B1(n16024), .B2(n14659), .A(n14658), .ZN(n14666) );
  NAND2_X1 U18054 ( .A1(n14661), .A2(n9972), .ZN(n14663) );
  MUX2_X1 U18055 ( .A(n14663), .B(n14662), .S(n14751), .Z(n14664) );
  XNOR2_X1 U18056 ( .A(n14664), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14847) );
  NAND2_X1 U18057 ( .A1(n14847), .A2(n11296), .ZN(n14665) );
  OAI211_X1 U18058 ( .C1(n14667), .C2(n13814), .A(n14666), .B(n14665), .ZN(
        P1_U2972) );
  NOR2_X1 U18059 ( .A1(n16162), .A2(n21272), .ZN(n16034) );
  NOR2_X1 U18060 ( .A1(n16022), .A2(n14668), .ZN(n14669) );
  AOI211_X1 U18061 ( .C1(n16015), .C2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16034), .B(n14669), .ZN(n14674) );
  OAI21_X1 U18062 ( .B1(n14687), .B2(n14805), .A(n14729), .ZN(n14670) );
  NAND2_X1 U18063 ( .A1(n14671), .A2(n14670), .ZN(n14672) );
  XNOR2_X1 U18064 ( .A(n14672), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16035) );
  NAND2_X1 U18065 ( .A1(n16035), .A2(n11296), .ZN(n14673) );
  OAI211_X1 U18066 ( .C1(n14675), .C2(n13814), .A(n14674), .B(n14673), .ZN(
        P1_U2973) );
  MUX2_X1 U18067 ( .A(n14871), .B(n14676), .S(n14751), .Z(n14679) );
  NAND2_X1 U18068 ( .A1(n14677), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14688) );
  AND2_X1 U18069 ( .A1(n14688), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14678) );
  NOR2_X1 U18070 ( .A1(n14679), .A2(n14678), .ZN(n14680) );
  XNOR2_X1 U18071 ( .A(n14680), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14863) );
  NAND2_X1 U18072 ( .A1(n16024), .A2(n14681), .ZN(n14682) );
  NAND2_X1 U18073 ( .A1(n16174), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14859) );
  OAI211_X1 U18074 ( .C1(n16029), .C2(n14683), .A(n14682), .B(n14859), .ZN(
        n14684) );
  AOI21_X1 U18075 ( .B1(n14685), .B2(n16025), .A(n14684), .ZN(n14686) );
  OAI21_X1 U18076 ( .B1(n20080), .B2(n14863), .A(n14686), .ZN(P1_U2974) );
  NAND2_X1 U18077 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  MUX2_X1 U18078 ( .A(n14689), .B(n14688), .S(n14729), .Z(n14690) );
  NAND2_X1 U18079 ( .A1(n14691), .A2(n16025), .ZN(n14696) );
  NOR2_X1 U18080 ( .A1(n16162), .A2(n20879), .ZN(n14870) );
  NOR2_X1 U18081 ( .A1(n16029), .A2(n14692), .ZN(n14693) );
  AOI211_X1 U18082 ( .C1(n16024), .C2(n14694), .A(n14870), .B(n14693), .ZN(
        n14695) );
  OAI211_X1 U18083 ( .C1(n14864), .C2(n20080), .A(n14696), .B(n14695), .ZN(
        P1_U2975) );
  XNOR2_X1 U18084 ( .A(n14729), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14697) );
  XNOR2_X1 U18085 ( .A(n14645), .B(n14697), .ZN(n16044) );
  INV_X1 U18086 ( .A(n14698), .ZN(n14700) );
  AOI22_X1 U18087 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14699) );
  OAI21_X1 U18088 ( .B1(n14700), .B2(n16022), .A(n14699), .ZN(n14701) );
  AOI21_X1 U18089 ( .B1(n14702), .B2(n16025), .A(n14701), .ZN(n14703) );
  OAI21_X1 U18090 ( .B1(n16044), .B2(n20080), .A(n14703), .ZN(P1_U2976) );
  NAND2_X1 U18091 ( .A1(n14705), .A2(n14704), .ZN(n14706) );
  XOR2_X1 U18092 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14706), .Z(
        n16051) );
  AOI22_X1 U18093 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14707) );
  OAI21_X1 U18094 ( .B1(n14708), .B2(n16022), .A(n14707), .ZN(n14709) );
  AOI21_X1 U18095 ( .B1(n14710), .B2(n16025), .A(n14709), .ZN(n14711) );
  OAI21_X1 U18096 ( .B1(n20080), .B2(n16051), .A(n14711), .ZN(P1_U2977) );
  NAND3_X1 U18097 ( .A1(n14751), .A2(n11291), .A3(n16085), .ZN(n14712) );
  NOR2_X1 U18098 ( .A1(n14739), .A2(n14712), .ZN(n14720) );
  NOR2_X1 U18099 ( .A1(n14751), .A2(n14866), .ZN(n14713) );
  AOI22_X1 U18100 ( .A1(n14720), .A2(n14794), .B1(n14738), .B2(n14713), .ZN(
        n14714) );
  XNOR2_X1 U18101 ( .A(n14714), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14878) );
  NOR2_X1 U18102 ( .A1(n16162), .A2(n21018), .ZN(n14881) );
  AOI21_X1 U18103 ( .B1(n16015), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14881), .ZN(n14715) );
  OAI21_X1 U18104 ( .B1(n14716), .B2(n16022), .A(n14715), .ZN(n14717) );
  AOI21_X1 U18105 ( .B1(n14878), .B2(n11296), .A(n14717), .ZN(n14718) );
  OAI21_X1 U18106 ( .B1(n14719), .B2(n13814), .A(n14718), .ZN(P1_U2978) );
  AND3_X1 U18107 ( .A1(n14738), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14729), .ZN(n14721) );
  NOR2_X1 U18108 ( .A1(n14721), .A2(n14720), .ZN(n14722) );
  XNOR2_X1 U18109 ( .A(n14722), .B(n14794), .ZN(n15895) );
  INV_X1 U18110 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21131) );
  OAI22_X1 U18111 ( .A1(n16029), .A2(n14723), .B1(n16162), .B2(n21131), .ZN(
        n14726) );
  NOR2_X1 U18112 ( .A1(n14724), .A2(n13814), .ZN(n14725) );
  AOI211_X1 U18113 ( .C1(n16024), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        n14728) );
  OAI21_X1 U18114 ( .B1(n15895), .B2(n20080), .A(n14728), .ZN(P1_U2979) );
  NOR2_X1 U18115 ( .A1(n14729), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14730) );
  MUX2_X1 U18116 ( .A(n14730), .B(n14729), .S(n14738), .Z(n14731) );
  XNOR2_X1 U18117 ( .A(n14731), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16060) );
  OAI22_X1 U18118 ( .A1(n16029), .A2(n14732), .B1(n16162), .B2(n21041), .ZN(
        n14735) );
  NOR2_X1 U18119 ( .A1(n14733), .A2(n13814), .ZN(n14734) );
  AOI211_X1 U18120 ( .C1(n16024), .C2(n14736), .A(n14735), .B(n14734), .ZN(
        n14737) );
  OAI21_X1 U18121 ( .B1(n20080), .B2(n16060), .A(n14737), .ZN(P1_U2980) );
  OAI21_X1 U18122 ( .B1(n14740), .B2(n14739), .A(n9974), .ZN(n16080) );
  NOR2_X1 U18123 ( .A1(n16162), .A2(n21039), .ZN(n16083) );
  INV_X1 U18124 ( .A(n16083), .ZN(n14742) );
  NAND2_X1 U18125 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14741) );
  OAI211_X1 U18126 ( .C1(n16022), .C2(n14743), .A(n14742), .B(n14741), .ZN(
        n14744) );
  AOI21_X1 U18127 ( .B1(n14745), .B2(n16025), .A(n14744), .ZN(n14746) );
  OAI21_X1 U18128 ( .B1(n20080), .B2(n16080), .A(n14746), .ZN(P1_U2981) );
  AOI21_X1 U18129 ( .B1(n14729), .B2(n16109), .A(n15993), .ZN(n14750) );
  AND2_X1 U18130 ( .A1(n14751), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14759) );
  INV_X1 U18131 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14755) );
  OAI22_X1 U18132 ( .A1(n16029), .A2(n15912), .B1(n16162), .B2(n14755), .ZN(
        n14757) );
  NOR2_X1 U18133 ( .A1(n15915), .A2(n13814), .ZN(n14756) );
  AOI211_X1 U18134 ( .C1(n16024), .C2(n15914), .A(n14757), .B(n14756), .ZN(
        n14758) );
  OAI21_X1 U18135 ( .B1(n16086), .B2(n20080), .A(n14758), .ZN(P1_U2982) );
  INV_X1 U18136 ( .A(n14759), .ZN(n14760) );
  NAND2_X1 U18137 ( .A1(n14760), .A2(n15984), .ZN(n14761) );
  AOI22_X1 U18138 ( .A1(n9820), .A2(n15984), .B1(n14762), .B2(n14761), .ZN(
        n16103) );
  INV_X1 U18139 ( .A(n14763), .ZN(n14767) );
  AOI22_X1 U18140 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14764) );
  OAI21_X1 U18141 ( .B1(n14765), .B2(n16022), .A(n14764), .ZN(n14766) );
  AOI21_X1 U18142 ( .B1(n14767), .B2(n16025), .A(n14766), .ZN(n14768) );
  OAI21_X1 U18143 ( .B1(n16103), .B2(n20080), .A(n14768), .ZN(P1_U2984) );
  AND2_X1 U18144 ( .A1(n16006), .A2(n14769), .ZN(n14886) );
  OAI21_X1 U18145 ( .B1(n14886), .B2(n14770), .A(n14888), .ZN(n14772) );
  XNOR2_X1 U18146 ( .A(n14772), .B(n14771), .ZN(n16118) );
  INV_X1 U18147 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14773) );
  OAI22_X1 U18148 ( .A1(n16029), .A2(n14774), .B1(n16162), .B2(n14773), .ZN(
        n14776) );
  NOR2_X1 U18149 ( .A1(n15944), .A2(n13814), .ZN(n14775) );
  AOI211_X1 U18150 ( .C1(n16024), .C2(n15947), .A(n14776), .B(n14775), .ZN(
        n14777) );
  OAI21_X1 U18151 ( .B1(n20080), .B2(n16118), .A(n14777), .ZN(P1_U2986) );
  NAND2_X1 U18152 ( .A1(n14780), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14779) );
  XNOR2_X1 U18153 ( .A(n14747), .B(n14781), .ZN(n14778) );
  MUX2_X1 U18154 ( .A(n14779), .B(n14778), .S(n14729), .Z(n14783) );
  INV_X1 U18155 ( .A(n14780), .ZN(n14782) );
  NAND3_X1 U18156 ( .A1(n14782), .A2(n14751), .A3(n14781), .ZN(n16007) );
  NAND2_X1 U18157 ( .A1(n14783), .A2(n16007), .ZN(n16139) );
  INV_X1 U18158 ( .A(n16139), .ZN(n14789) );
  AOI22_X1 U18159 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14784) );
  OAI21_X1 U18160 ( .B1(n14785), .B2(n16022), .A(n14784), .ZN(n14786) );
  AOI21_X1 U18161 ( .B1(n14787), .B2(n16025), .A(n14786), .ZN(n14788) );
  OAI21_X1 U18162 ( .B1(n14789), .B2(n20080), .A(n14788), .ZN(P1_U2989) );
  INV_X1 U18163 ( .A(n14790), .ZN(n14799) );
  NAND3_X1 U18164 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16078) );
  NAND2_X1 U18165 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16159), .ZN(
        n14892) );
  INV_X1 U18166 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16009) );
  INV_X1 U18167 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16168) );
  NOR3_X1 U18168 ( .A1(n16168), .A2(n16179), .A3(n16165), .ZN(n16136) );
  NAND3_X1 U18169 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16136), .ZN(n14893) );
  NOR2_X1 U18170 ( .A1(n16009), .A2(n14893), .ZN(n14901) );
  NAND2_X1 U18171 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14901), .ZN(
        n14792) );
  NOR2_X1 U18172 ( .A1(n14892), .A2(n14792), .ZN(n16071) );
  NAND2_X1 U18173 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16071), .ZN(
        n14793) );
  NOR2_X1 U18174 ( .A1(n14792), .A2(n14791), .ZN(n16113) );
  NAND2_X1 U18175 ( .A1(n14803), .A2(n16113), .ZN(n16077) );
  OAI21_X1 U18176 ( .B1(n16070), .B2(n14793), .A(n16077), .ZN(n16119) );
  NAND2_X1 U18177 ( .A1(n15889), .A2(n16119), .ZN(n15893) );
  INV_X1 U18178 ( .A(n16071), .ZN(n16128) );
  NOR2_X1 U18179 ( .A1(n16128), .A2(n14896), .ZN(n16075) );
  NAND2_X1 U18180 ( .A1(n15889), .A2(n16075), .ZN(n14869) );
  NAND2_X1 U18181 ( .A1(n15893), .A2(n14869), .ZN(n16065) );
  NAND2_X1 U18182 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16065), .ZN(
        n15901) );
  INV_X1 U18183 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16053) );
  NOR2_X1 U18184 ( .A1(n14884), .A2(n16053), .ZN(n16052) );
  AND3_X1 U18185 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n16052), .ZN(n14795) );
  AND2_X1 U18186 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14807) );
  NAND2_X1 U18187 ( .A1(n16037), .A2(n14807), .ZN(n14848) );
  NAND2_X1 U18188 ( .A1(n14838), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14796) );
  OR2_X1 U18189 ( .A1(n14848), .A2(n14796), .ZN(n14822) );
  INV_X1 U18190 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14821) );
  NOR3_X1 U18191 ( .A1(n14822), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14821), .ZN(n14797) );
  AOI211_X1 U18192 ( .C1(n14799), .C2(n16173), .A(n14798), .B(n14797), .ZN(
        n14815) );
  OAI211_X1 U18193 ( .C1(n16071), .C2(n16158), .A(n16113), .B(n15889), .ZN(
        n14801) );
  AOI221_X1 U18194 ( .B1(n14801), .B2(n16160), .C1(n14866), .C2(n16160), .A(
        n14800), .ZN(n16049) );
  INV_X1 U18195 ( .A(n16052), .ZN(n14865) );
  NAND2_X1 U18196 ( .A1(n16160), .A2(n14865), .ZN(n14802) );
  AND2_X1 U18197 ( .A1(n16049), .A2(n14802), .ZN(n16043) );
  NAND2_X1 U18198 ( .A1(n14803), .A2(n16042), .ZN(n14804) );
  NAND2_X1 U18199 ( .A1(n16160), .A2(n14805), .ZN(n14806) );
  NAND2_X1 U18200 ( .A1(n14868), .A2(n14806), .ZN(n16031) );
  INV_X1 U18201 ( .A(n14807), .ZN(n14808) );
  OR2_X1 U18202 ( .A1(n16031), .A2(n14808), .ZN(n14809) );
  INV_X1 U18203 ( .A(n16160), .ZN(n16074) );
  NAND2_X1 U18204 ( .A1(n14868), .A2(n16074), .ZN(n14813) );
  NAND2_X1 U18205 ( .A1(n14809), .A2(n14813), .ZN(n14856) );
  INV_X1 U18206 ( .A(n14838), .ZN(n14810) );
  NAND2_X1 U18207 ( .A1(n14813), .A2(n14810), .ZN(n14811) );
  NAND2_X1 U18208 ( .A1(n14856), .A2(n14811), .ZN(n14835) );
  AND2_X1 U18209 ( .A1(n16160), .A2(n14828), .ZN(n14812) );
  NAND3_X1 U18210 ( .A1(n14824), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14813), .ZN(n14814) );
  OAI211_X1 U18211 ( .C1(n14816), .C2(n16182), .A(n14815), .B(n14814), .ZN(
        P1_U3000) );
  INV_X1 U18212 ( .A(n14817), .ZN(n14827) );
  INV_X1 U18213 ( .A(n14818), .ZN(n14820) );
  AOI21_X1 U18214 ( .B1(n14820), .B2(n16173), .A(n14819), .ZN(n14826) );
  NAND2_X1 U18215 ( .A1(n14822), .A2(n14821), .ZN(n14823) );
  NAND2_X1 U18216 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  OAI211_X1 U18217 ( .C1(n14827), .C2(n16182), .A(n14826), .B(n14825), .ZN(
        P1_U3001) );
  NAND2_X1 U18218 ( .A1(n14838), .A2(n14828), .ZN(n14829) );
  NOR2_X1 U18219 ( .A1(n14848), .A2(n14829), .ZN(n14834) );
  INV_X1 U18220 ( .A(n14830), .ZN(n14831) );
  OAI21_X1 U18221 ( .B1(n14832), .B2(n20258), .A(n14831), .ZN(n14833) );
  AOI211_X1 U18222 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14835), .A(
        n14834), .B(n14833), .ZN(n14836) );
  OAI21_X1 U18223 ( .B1(n14837), .B2(n16182), .A(n14836), .ZN(P1_U3002) );
  INV_X1 U18224 ( .A(n14856), .ZN(n14844) );
  NOR3_X1 U18225 ( .A1(n14848), .A2(n14839), .A3(n14838), .ZN(n14843) );
  OAI21_X1 U18226 ( .B1(n14841), .B2(n20258), .A(n14840), .ZN(n14842) );
  AOI211_X1 U18227 ( .C1(n14844), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14843), .B(n14842), .ZN(n14845) );
  OAI21_X1 U18228 ( .B1(n14846), .B2(n16182), .A(n14845), .ZN(P1_U3003) );
  NAND2_X1 U18229 ( .A1(n14847), .A2(n20260), .ZN(n14854) );
  INV_X1 U18230 ( .A(n14848), .ZN(n14852) );
  OAI21_X1 U18231 ( .B1(n14850), .B2(n20258), .A(n14849), .ZN(n14851) );
  AOI21_X1 U18232 ( .B1(n14852), .B2(n14855), .A(n14851), .ZN(n14853) );
  OAI211_X1 U18233 ( .C1(n14856), .C2(n14855), .A(n14854), .B(n14853), .ZN(
        P1_U3004) );
  NAND2_X1 U18234 ( .A1(n16037), .A2(n14857), .ZN(n14858) );
  OAI211_X1 U18235 ( .C1(n14860), .C2(n20258), .A(n14859), .B(n14858), .ZN(
        n14861) );
  AOI21_X1 U18236 ( .B1(n16031), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14861), .ZN(n14862) );
  OAI21_X1 U18237 ( .B1(n14863), .B2(n16182), .A(n14862), .ZN(P1_U3006) );
  NOR2_X1 U18238 ( .A1(n14864), .A2(n16182), .ZN(n14877) );
  NOR3_X1 U18239 ( .A1(n14866), .A2(n14865), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16041) );
  INV_X1 U18240 ( .A(n16041), .ZN(n14867) );
  AOI221_X1 U18241 ( .B1(n14869), .B2(n14868), .C1(n14867), .C2(n14868), .A(
        n14871), .ZN(n14876) );
  INV_X1 U18242 ( .A(n14870), .ZN(n14873) );
  NAND4_X1 U18243 ( .A1(n16055), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n16052), .A4(n14871), .ZN(n14872) );
  OAI211_X1 U18244 ( .C1(n14874), .C2(n20258), .A(n14873), .B(n14872), .ZN(
        n14875) );
  OR3_X1 U18245 ( .A1(n14877), .A2(n14876), .A3(n14875), .ZN(P1_U3007) );
  NAND2_X1 U18246 ( .A1(n14878), .A2(n20260), .ZN(n14883) );
  NOR2_X1 U18247 ( .A1(n14879), .A2(n20258), .ZN(n14880) );
  AOI211_X1 U18248 ( .C1(n16055), .C2(n14884), .A(n14881), .B(n14880), .ZN(
        n14882) );
  OAI211_X1 U18249 ( .C1(n16049), .C2(n14884), .A(n14883), .B(n14882), .ZN(
        P1_U3010) );
  INV_X1 U18250 ( .A(n14885), .ZN(n14887) );
  AOI21_X1 U18251 ( .B1(n14751), .B2(n14887), .A(n14886), .ZN(n14891) );
  OAI21_X1 U18252 ( .B1(n14889), .B2(n14729), .A(n14888), .ZN(n14890) );
  XNOR2_X1 U18253 ( .A(n14891), .B(n14890), .ZN(n16005) );
  OR2_X1 U18254 ( .A1(n14893), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16134) );
  OAI21_X1 U18255 ( .B1(n14893), .B2(n14892), .A(n15891), .ZN(n14894) );
  OAI211_X1 U18256 ( .C1(n14901), .C2(n15888), .A(n16157), .B(n14894), .ZN(
        n16130) );
  INV_X1 U18257 ( .A(n16130), .ZN(n14895) );
  OAI21_X1 U18258 ( .B1(n14896), .B2(n16134), .A(n14895), .ZN(n14902) );
  INV_X1 U18259 ( .A(n14897), .ZN(n14899) );
  NAND3_X1 U18260 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14899), .A3(
        n14898), .ZN(n16181) );
  NOR2_X1 U18261 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16181), .ZN(
        n14900) );
  AOI22_X1 U18262 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14902), .B1(
        n14901), .B2(n14900), .ZN(n14905) );
  XOR2_X1 U18263 ( .A(n14903), .B(n15958), .Z(n15969) );
  AOI22_X1 U18264 ( .A1(n15969), .A2(n16173), .B1(n16174), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14904) );
  OAI211_X1 U18265 ( .C1(n16005), .C2(n16182), .A(n14905), .B(n14904), .ZN(
        P1_U3019) );
  OAI211_X1 U18266 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20339), .A(n20623), 
        .B(n20698), .ZN(n14906) );
  OAI21_X1 U18267 ( .B1(n13559), .B2(n14907), .A(n14906), .ZN(n14908) );
  MUX2_X1 U18268 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14908), .S(
        n20923), .Z(P1_U3477) );
  INV_X1 U18269 ( .A(n14909), .ZN(n14974) );
  NAND2_X1 U18270 ( .A1(n20052), .A2(n11863), .ZN(n14951) );
  INV_X1 U18271 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16201) );
  NAND2_X1 U18272 ( .A1(n20057), .A2(n20001), .ZN(n14953) );
  INV_X1 U18273 ( .A(n14953), .ZN(n14910) );
  OAI21_X1 U18274 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n14914), .A(
        n14913), .ZN(n16226) );
  INV_X1 U18275 ( .A(n14947), .ZN(n14915) );
  OAI21_X1 U18276 ( .B1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n14915), .A(
        n10182), .ZN(n15347) );
  INV_X1 U18277 ( .A(n14916), .ZN(n14944) );
  INV_X1 U18278 ( .A(n14919), .ZN(n14917) );
  NAND2_X1 U18279 ( .A1(n14917), .A2(n16243), .ZN(n14918) );
  NAND2_X1 U18280 ( .A1(n14944), .A2(n14918), .ZN(n16251) );
  AOI21_X1 U18281 ( .B1(n14942), .B2(n10178), .A(n14919), .ZN(n15380) );
  INV_X1 U18282 ( .A(n15380), .ZN(n16260) );
  INV_X1 U18283 ( .A(n14922), .ZN(n14921) );
  INV_X1 U18284 ( .A(n14943), .ZN(n14920) );
  OAI21_X1 U18285 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n14921), .A(
        n14920), .ZN(n15406) );
  OAI21_X1 U18286 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n14939), .A(
        n14922), .ZN(n19053) );
  INV_X1 U18287 ( .A(n19053), .ZN(n19050) );
  OAI21_X1 U18288 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n9885), .A(
        n14938), .ZN(n15443) );
  INV_X1 U18289 ( .A(n15443), .ZN(n19066) );
  OAI21_X1 U18290 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14934), .A(
        n14937), .ZN(n19089) );
  OAI21_X1 U18291 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n14932), .A(
        n14935), .ZN(n16287) );
  INV_X1 U18292 ( .A(n16287), .ZN(n19116) );
  OAI21_X1 U18293 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n14930), .A(
        n14933), .ZN(n16307) );
  INV_X1 U18294 ( .A(n16307), .ZN(n19127) );
  OAI21_X1 U18295 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9886), .A(
        n14931), .ZN(n16334) );
  INV_X1 U18296 ( .A(n16334), .ZN(n15063) );
  OAI21_X1 U18297 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n14923), .A(
        n14929), .ZN(n15473) );
  INV_X1 U18298 ( .A(n15473), .ZN(n19141) );
  AOI21_X1 U18299 ( .B1(n19151), .B2(n14925), .A(n14928), .ZN(n19149) );
  AOI21_X1 U18300 ( .B1(n19286), .B2(n14924), .A(n14926), .ZN(n19269) );
  AOI22_X1 U18301 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20054), .ZN(n15757) );
  AOI22_X1 U18302 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n15136), .B2(n20054), .ZN(
        n15134) );
  NAND2_X1 U18303 ( .A1(n15757), .A2(n15134), .ZN(n15133) );
  NOR2_X1 U18304 ( .A1(n15121), .A2(n15133), .ZN(n15109) );
  NAND2_X1 U18305 ( .A1(n15109), .A2(n15110), .ZN(n19170) );
  NOR2_X1 U18306 ( .A1(n19269), .A2(n19170), .ZN(n15097) );
  OAI21_X1 U18307 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n14926), .A(
        n14925), .ZN(n16365) );
  NAND2_X1 U18308 ( .A1(n15097), .A2(n16365), .ZN(n19147) );
  NOR2_X1 U18309 ( .A1(n19149), .A2(n19147), .ZN(n15086) );
  OAI21_X1 U18310 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14928), .A(
        n14927), .ZN(n16345) );
  NAND2_X1 U18311 ( .A1(n15086), .A2(n16345), .ZN(n19139) );
  NOR2_X1 U18312 ( .A1(n19141), .A2(n19139), .ZN(n15073) );
  AOI21_X1 U18313 ( .B1(n16344), .B2(n14929), .A(n9886), .ZN(n16335) );
  INV_X1 U18314 ( .A(n16335), .ZN(n15074) );
  NAND2_X1 U18315 ( .A1(n15073), .A2(n15074), .ZN(n15061) );
  NOR2_X1 U18316 ( .A1(n15063), .A2(n15061), .ZN(n15048) );
  AOI21_X1 U18317 ( .B1(n16322), .B2(n14931), .A(n14930), .ZN(n16308) );
  INV_X1 U18318 ( .A(n16308), .ZN(n15049) );
  NAND2_X1 U18319 ( .A1(n15048), .A2(n15049), .ZN(n19125) );
  NOR2_X1 U18320 ( .A1(n19127), .A2(n19125), .ZN(n15036) );
  AOI21_X1 U18321 ( .B1(n16300), .B2(n14933), .A(n14932), .ZN(n16288) );
  INV_X1 U18322 ( .A(n16288), .ZN(n15035) );
  NAND2_X1 U18323 ( .A1(n15036), .A2(n15035), .ZN(n19114) );
  NOR2_X1 U18324 ( .A1(n19116), .A2(n19114), .ZN(n19107) );
  AOI21_X1 U18325 ( .B1(n16281), .B2(n14935), .A(n14934), .ZN(n16273) );
  INV_X1 U18326 ( .A(n16273), .ZN(n19106) );
  NAND2_X1 U18327 ( .A1(n19107), .A2(n19106), .ZN(n19104) );
  INV_X1 U18328 ( .A(n19104), .ZN(n14936) );
  NAND2_X1 U18329 ( .A1(n19089), .A2(n14936), .ZN(n19074) );
  AOI21_X1 U18330 ( .B1(n15447), .B2(n14937), .A(n9885), .ZN(n19075) );
  OR2_X1 U18331 ( .A1(n19074), .A2(n19075), .ZN(n19065) );
  NOR2_X1 U18332 ( .A1(n19066), .A2(n19065), .ZN(n15020) );
  NAND2_X1 U18333 ( .A1(n14938), .A2(n15429), .ZN(n14941) );
  INV_X1 U18334 ( .A(n14939), .ZN(n14940) );
  NAND2_X1 U18335 ( .A1(n14941), .A2(n14940), .ZN(n15433) );
  NAND2_X1 U18336 ( .A1(n15020), .A2(n15433), .ZN(n19049) );
  OAI21_X1 U18337 ( .B1(n19050), .B2(n19049), .A(n15019), .ZN(n19048) );
  NAND2_X1 U18338 ( .A1(n15406), .A2(n19048), .ZN(n15004) );
  NAND2_X1 U18339 ( .A1(n15019), .A2(n15004), .ZN(n15838) );
  OAI21_X1 U18340 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n14943), .A(
        n14942), .ZN(n15839) );
  NAND2_X1 U18341 ( .A1(n9807), .A2(n15837), .ZN(n16259) );
  NAND2_X1 U18342 ( .A1(n16260), .A2(n16259), .ZN(n16258) );
  NAND2_X1 U18343 ( .A1(n9807), .A2(n16258), .ZN(n16250) );
  NAND2_X1 U18344 ( .A1(n16251), .A2(n16250), .ZN(n16249) );
  NAND2_X1 U18345 ( .A1(n9807), .A2(n16249), .ZN(n14992) );
  INV_X1 U18346 ( .A(n14948), .ZN(n14946) );
  INV_X1 U18347 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15363) );
  NAND2_X1 U18348 ( .A1(n14944), .A2(n15363), .ZN(n14945) );
  NAND2_X1 U18349 ( .A1(n14946), .A2(n14945), .ZN(n15362) );
  NAND2_X1 U18350 ( .A1(n9807), .A2(n14991), .ZN(n16238) );
  OAI21_X1 U18351 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n14948), .A(
        n14947), .ZN(n16239) );
  NAND2_X1 U18352 ( .A1(n9807), .A2(n16237), .ZN(n14978) );
  NAND2_X1 U18353 ( .A1(n15347), .A2(n14978), .ZN(n14977) );
  NAND2_X1 U18354 ( .A1(n9807), .A2(n14977), .ZN(n16225) );
  NAND2_X1 U18355 ( .A1(n16226), .A2(n16225), .ZN(n16224) );
  NAND2_X1 U18356 ( .A1(n9807), .A2(n16224), .ZN(n14950) );
  NOR3_X1 U18357 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n16478), .A3(n15902), 
        .ZN(n15122) );
  OAI211_X1 U18358 ( .C1(n14950), .C2(n14949), .A(n19190), .B(n16198), .ZN(
        n14973) );
  INV_X1 U18359 ( .A(n20057), .ZN(n19897) );
  NAND2_X1 U18360 ( .A1(n20001), .A2(n14952), .ZN(n14960) );
  NAND2_X1 U18361 ( .A1(n19266), .A2(n14960), .ZN(n16200) );
  AND2_X1 U18362 ( .A1(n16201), .A2(n14953), .ZN(n14954) );
  NAND2_X1 U18363 ( .A1(n14955), .A2(n14954), .ZN(n14956) );
  NAND2_X1 U18364 ( .A1(n15247), .A2(n14957), .ZN(n14958) );
  INV_X1 U18365 ( .A(n14960), .ZN(n14961) );
  AND3_X1 U18366 ( .A1(n12173), .A2(n14961), .A3(n20055), .ZN(n14962) );
  AND2_X1 U18367 ( .A1(n11873), .A2(n14962), .ZN(n16482) );
  NAND2_X1 U18368 ( .A1(n15496), .A2(n19168), .ZN(n14969) );
  NAND2_X1 U18369 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19533), .ZN(n19887) );
  NOR2_X1 U18370 ( .A1(n19894), .A2(n19887), .ZN(n16489) );
  NAND2_X1 U18371 ( .A1(n19150), .A2(n19891), .ZN(n14964) );
  OR2_X1 U18372 ( .A1(n16489), .A2(n14964), .ZN(n14965) );
  NOR2_X2 U18373 ( .A1(n19166), .A2(n12958), .ZN(n19193) );
  INV_X1 U18374 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19968) );
  OAI22_X1 U18375 ( .A1(n14966), .A2(n19163), .B1(n19968), .B2(n19181), .ZN(
        n14967) );
  INV_X1 U18376 ( .A(n14967), .ZN(n14968) );
  OAI211_X1 U18377 ( .C1(n12624), .C2(n19134), .A(n14969), .B(n14968), .ZN(
        n14970) );
  AOI21_X1 U18378 ( .B1(n14971), .B2(n19188), .A(n14970), .ZN(n14972) );
  OAI211_X1 U18379 ( .C1(n14974), .C2(n19186), .A(n14973), .B(n14972), .ZN(
        P2_U2826) );
  OAI211_X1 U18380 ( .C1(n14978), .C2(n15347), .A(n19190), .B(n14977), .ZN(
        n14990) );
  NAND3_X1 U18381 ( .A1(n12785), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n14979), 
        .ZN(n14980) );
  NAND2_X1 U18382 ( .A1(n14981), .A2(n14980), .ZN(n15330) );
  INV_X1 U18383 ( .A(n15330), .ZN(n14988) );
  INV_X1 U18384 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19965) );
  OAI22_X1 U18385 ( .A1(n14982), .A2(n19163), .B1(n19965), .B2(n19181), .ZN(
        n14987) );
  NOR2_X1 U18386 ( .A1(n14983), .A2(n14984), .ZN(n14985) );
  OR2_X1 U18387 ( .A1(n15245), .A2(n14985), .ZN(n15516) );
  OAI22_X1 U18388 ( .A1(n15516), .A2(n19179), .B1(n12615), .B2(n19134), .ZN(
        n14986) );
  AOI211_X1 U18389 ( .C1(n19102), .C2(n14988), .A(n14987), .B(n14986), .ZN(
        n14989) );
  OAI211_X1 U18390 ( .C1(n15514), .C2(n19157), .A(n14990), .B(n14989), .ZN(
        P2_U2828) );
  OAI211_X1 U18391 ( .C1(n14992), .C2(n15362), .A(n19190), .B(n14991), .ZN(
        n15002) );
  NOR2_X1 U18392 ( .A1(n15179), .A2(n14993), .ZN(n14994) );
  OR2_X1 U18393 ( .A1(n15165), .A2(n14994), .ZN(n15543) );
  INV_X1 U18394 ( .A(n15543), .ZN(n15000) );
  INV_X1 U18395 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19960) );
  OAI22_X1 U18396 ( .A1(n15363), .A2(n19163), .B1(n19960), .B2(n19181), .ZN(
        n14999) );
  AND2_X1 U18397 ( .A1(n15276), .A2(n14995), .ZN(n14996) );
  NOR2_X1 U18398 ( .A1(n9834), .A2(n14996), .ZN(n15540) );
  INV_X1 U18399 ( .A(n15540), .ZN(n14997) );
  OAI22_X1 U18400 ( .A1(n14997), .A2(n19179), .B1(n19134), .B2(n15172), .ZN(
        n14998) );
  AOI211_X1 U18401 ( .C1(n15000), .C2(n19188), .A(n14999), .B(n14998), .ZN(
        n15001) );
  OAI211_X1 U18402 ( .C1(n19186), .C2(n15003), .A(n15002), .B(n15001), .ZN(
        P2_U2830) );
  OAI211_X1 U18403 ( .C1(n19048), .C2(n15406), .A(n19190), .B(n15004), .ZN(
        n15016) );
  INV_X1 U18404 ( .A(n15195), .ZN(n15007) );
  NAND2_X1 U18405 ( .A1(n15207), .A2(n15005), .ZN(n15006) );
  NAND2_X1 U18406 ( .A1(n15007), .A2(n15006), .ZN(n15409) );
  INV_X1 U18407 ( .A(n15409), .ZN(n15591) );
  NOR2_X1 U18408 ( .A1(n15299), .A2(n15009), .ZN(n15010) );
  OR2_X1 U18409 ( .A1(n15008), .A2(n15010), .ZN(n15593) );
  INV_X1 U18410 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19952) );
  OAI22_X1 U18411 ( .A1(n15011), .A2(n19163), .B1(n19952), .B2(n19181), .ZN(
        n15012) );
  AOI21_X1 U18412 ( .B1(n19183), .B2(P2_EBX_REG_21__SCAN_IN), .A(n15012), .ZN(
        n15013) );
  OAI21_X1 U18413 ( .B1(n15593), .B2(n19179), .A(n15013), .ZN(n15014) );
  AOI21_X1 U18414 ( .B1(n15591), .B2(n19188), .A(n15014), .ZN(n15015) );
  OAI211_X1 U18415 ( .C1(n19186), .C2(n15017), .A(n15016), .B(n15015), .ZN(
        P2_U2834) );
  INV_X1 U18416 ( .A(n15018), .ZN(n15034) );
  NOR2_X1 U18417 ( .A1(n15758), .A2(n15020), .ZN(n15021) );
  XNOR2_X1 U18418 ( .A(n15021), .B(n15433), .ZN(n15022) );
  NAND2_X1 U18419 ( .A1(n15022), .A2(n19190), .ZN(n15033) );
  NAND2_X1 U18420 ( .A1(n15023), .A2(n15024), .ZN(n15025) );
  NAND2_X1 U18421 ( .A1(n15316), .A2(n15026), .ZN(n15027) );
  NAND2_X1 U18422 ( .A1(n15298), .A2(n15027), .ZN(n15620) );
  NAND2_X1 U18423 ( .A1(n19166), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15028) );
  OAI211_X1 U18424 ( .C1(n15429), .C2(n19163), .A(n15028), .B(n19150), .ZN(
        n15029) );
  AOI21_X1 U18425 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19183), .A(n15029), .ZN(
        n15030) );
  OAI21_X1 U18426 ( .B1(n15620), .B2(n19179), .A(n15030), .ZN(n15031) );
  AOI21_X1 U18427 ( .B1(n15617), .B2(n19188), .A(n15031), .ZN(n15032) );
  OAI211_X1 U18428 ( .C1(n19186), .C2(n15034), .A(n15033), .B(n15032), .ZN(
        P2_U2836) );
  NAND2_X1 U18429 ( .A1(n19190), .A2(n15019), .ZN(n16208) );
  INV_X1 U18430 ( .A(n16208), .ZN(n19105) );
  OAI211_X1 U18431 ( .C1(n15036), .C2(n15035), .A(n19105), .B(n19114), .ZN(
        n15047) );
  NAND2_X1 U18432 ( .A1(n15758), .A2(n19190), .ZN(n19100) );
  INV_X1 U18433 ( .A(n19100), .ZN(n19192) );
  AOI21_X1 U18434 ( .B1(n15037), .B2(n13848), .A(n15678), .ZN(n19207) );
  INV_X1 U18435 ( .A(n19207), .ZN(n15039) );
  AOI22_X1 U18436 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19193), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19166), .ZN(n15038) );
  OAI211_X1 U18437 ( .C1(n15039), .C2(n19179), .A(n15038), .B(n19150), .ZN(
        n15042) );
  NOR2_X1 U18438 ( .A1(n19134), .A2(n15040), .ZN(n15041) );
  AOI211_X1 U18439 ( .C1(n16288), .C2(n19192), .A(n15042), .B(n15041), .ZN(
        n15043) );
  OAI21_X1 U18440 ( .B1(n16376), .B2(n19157), .A(n15043), .ZN(n15044) );
  AOI21_X1 U18441 ( .B1(n15045), .B2(n19102), .A(n15044), .ZN(n15046) );
  NAND2_X1 U18442 ( .A1(n15047), .A2(n15046), .ZN(P2_U2842) );
  NOR2_X1 U18443 ( .A1(n15758), .A2(n15048), .ZN(n15050) );
  XNOR2_X1 U18444 ( .A(n15050), .B(n15049), .ZN(n15051) );
  NAND2_X1 U18445 ( .A1(n15051), .A2(n15122), .ZN(n15060) );
  INV_X1 U18446 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19932) );
  AOI22_X1 U18447 ( .A1(n15052), .A2(n19102), .B1(P2_EBX_REG_11__SCAN_IN), 
        .B2(n19183), .ZN(n15053) );
  OAI211_X1 U18448 ( .C1(n19932), .C2(n19181), .A(n15053), .B(n19150), .ZN(
        n15054) );
  AOI21_X1 U18449 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19193), .A(
        n15054), .ZN(n15059) );
  AOI21_X1 U18450 ( .B1(n15057), .B2(n15056), .A(n15055), .ZN(n19210) );
  AOI22_X1 U18451 ( .A1(n16388), .A2(n19188), .B1(n19168), .B2(n19210), .ZN(
        n15058) );
  NAND3_X1 U18452 ( .A1(n15060), .A2(n15059), .A3(n15058), .ZN(P2_U2844) );
  NAND2_X1 U18453 ( .A1(n9807), .A2(n15061), .ZN(n15062) );
  XNOR2_X1 U18454 ( .A(n15063), .B(n15062), .ZN(n15064) );
  NAND2_X1 U18455 ( .A1(n15064), .A2(n19190), .ZN(n15071) );
  INV_X1 U18456 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n15068) );
  INV_X1 U18457 ( .A(n16399), .ZN(n15065) );
  AOI22_X1 U18458 ( .A1(n19183), .A2(P2_EBX_REG_10__SCAN_IN), .B1(n19168), 
        .B2(n15065), .ZN(n15067) );
  AOI21_X1 U18459 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19193), .A(
        n19287), .ZN(n15066) );
  OAI211_X1 U18460 ( .C1(n15068), .C2(n19181), .A(n15067), .B(n15066), .ZN(
        n15069) );
  AOI21_X1 U18461 ( .B1(n16398), .B2(n19188), .A(n15069), .ZN(n15070) );
  OAI211_X1 U18462 ( .C1(n19186), .C2(n15072), .A(n15071), .B(n15070), .ZN(
        P2_U2845) );
  NOR2_X1 U18463 ( .A1(n15758), .A2(n15073), .ZN(n15075) );
  XNOR2_X1 U18464 ( .A(n15075), .B(n15074), .ZN(n15084) );
  INV_X1 U18465 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19929) );
  AOI22_X1 U18466 ( .A1(n15076), .A2(n19102), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19183), .ZN(n15077) );
  OAI211_X1 U18467 ( .C1(n19929), .C2(n19181), .A(n15077), .B(n19150), .ZN(
        n15078) );
  AOI21_X1 U18468 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19193), .A(
        n15078), .ZN(n15082) );
  AOI21_X1 U18469 ( .B1(n15080), .B2(n15079), .A(n9888), .ZN(n19214) );
  NAND2_X1 U18470 ( .A1(n19214), .A2(n19168), .ZN(n15081) );
  OAI211_X1 U18471 ( .C1(n19157), .C2(n16338), .A(n15082), .B(n15081), .ZN(
        n15083) );
  AOI21_X1 U18472 ( .B1(n15084), .B2(n19190), .A(n15083), .ZN(n15085) );
  INV_X1 U18473 ( .A(n15085), .ZN(P2_U2846) );
  NOR2_X1 U18474 ( .A1(n15758), .A2(n15086), .ZN(n15087) );
  XNOR2_X1 U18475 ( .A(n15087), .B(n16345), .ZN(n15088) );
  NAND2_X1 U18476 ( .A1(n15088), .A2(n19190), .ZN(n15096) );
  INV_X1 U18477 ( .A(n16354), .ZN(n15094) );
  INV_X1 U18478 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n15089) );
  OAI21_X1 U18479 ( .B1(n19181), .B2(n15089), .A(n19150), .ZN(n15093) );
  INV_X1 U18480 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16346) );
  AOI22_X1 U18481 ( .A1(n15090), .A2(n19102), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19183), .ZN(n15091) );
  OAI21_X1 U18482 ( .B1(n16346), .B2(n19163), .A(n15091), .ZN(n15092) );
  AOI211_X1 U18483 ( .C1(n15094), .C2(n19188), .A(n15093), .B(n15092), .ZN(
        n15095) );
  OAI211_X1 U18484 ( .C1(n15720), .C2(n19179), .A(n15096), .B(n15095), .ZN(
        P2_U2848) );
  NOR2_X1 U18485 ( .A1(n15758), .A2(n15097), .ZN(n15098) );
  XNOR2_X1 U18486 ( .A(n15098), .B(n16365), .ZN(n15099) );
  NAND2_X1 U18487 ( .A1(n15099), .A2(n19190), .ZN(n15108) );
  INV_X1 U18488 ( .A(n16356), .ZN(n15106) );
  INV_X1 U18489 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19922) );
  OAI21_X1 U18490 ( .B1(n19922), .B2(n19181), .A(n19150), .ZN(n15100) );
  AOI21_X1 U18491 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19193), .A(
        n15100), .ZN(n15101) );
  OAI21_X1 U18492 ( .B1(n19134), .B2(n15102), .A(n15101), .ZN(n15105) );
  NOR2_X1 U18493 ( .A1(n15103), .A2(n19186), .ZN(n15104) );
  AOI211_X1 U18494 ( .C1(n15106), .C2(n19188), .A(n15105), .B(n15104), .ZN(
        n15107) );
  OAI211_X1 U18495 ( .C1(n15736), .C2(n19179), .A(n15108), .B(n15107), .ZN(
        P2_U2850) );
  NOR2_X1 U18496 ( .A1(n15758), .A2(n15109), .ZN(n15111) );
  XNOR2_X1 U18497 ( .A(n15111), .B(n15110), .ZN(n15112) );
  NAND2_X1 U18498 ( .A1(n15112), .A2(n15122), .ZN(n15119) );
  AOI22_X1 U18499 ( .A1(n19183), .A2(P2_EBX_REG_3__SCAN_IN), .B1(n19168), .B2(
        n20008), .ZN(n15113) );
  OAI21_X1 U18500 ( .B1(n15114), .B2(n19186), .A(n15113), .ZN(n15117) );
  INV_X1 U18501 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15115) );
  OAI22_X1 U18502 ( .A1(n15115), .A2(n19163), .B1(n19919), .B2(n19181), .ZN(
        n15116) );
  AOI211_X1 U18503 ( .C1(n19188), .C2(n16425), .A(n15117), .B(n15116), .ZN(
        n15118) );
  OAI211_X1 U18504 ( .C1(n19987), .C2(n15132), .A(n15119), .B(n15118), .ZN(
        P2_U2852) );
  NAND2_X1 U18505 ( .A1(n9807), .A2(n15133), .ZN(n15120) );
  XNOR2_X1 U18506 ( .A(n15121), .B(n15120), .ZN(n15123) );
  NAND2_X1 U18507 ( .A1(n15123), .A2(n15122), .ZN(n15131) );
  AOI22_X1 U18508 ( .A1(n19166), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n19183), .ZN(n15124) );
  OAI21_X1 U18509 ( .B1(n15125), .B2(n19186), .A(n15124), .ZN(n15129) );
  OAI22_X1 U18510 ( .A1(n15127), .A2(n19179), .B1(n15126), .B2(n19163), .ZN(
        n15128) );
  AOI211_X1 U18511 ( .C1(n19188), .C2(n15764), .A(n15129), .B(n15128), .ZN(
        n15130) );
  OAI211_X1 U18512 ( .C1(n15132), .C2(n20015), .A(n15131), .B(n15130), .ZN(
        P2_U2853) );
  OAI211_X1 U18513 ( .C1(n15757), .C2(n15134), .A(n15019), .B(n15133), .ZN(
        n15782) );
  NOR2_X1 U18514 ( .A1(n19186), .A2(n15135), .ZN(n15141) );
  AOI22_X1 U18515 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19193), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19166), .ZN(n15138) );
  NAND2_X1 U18516 ( .A1(n19192), .A2(n15136), .ZN(n15137) );
  OAI211_X1 U18517 ( .C1(n19134), .C2(n15139), .A(n15138), .B(n15137), .ZN(
        n15140) );
  AOI211_X1 U18518 ( .C1(n19168), .C2(n20026), .A(n15141), .B(n15140), .ZN(
        n15142) );
  OAI21_X1 U18519 ( .B1(n19307), .B2(n19157), .A(n15142), .ZN(n15143) );
  AOI21_X1 U18520 ( .B1(n20022), .B2(n19189), .A(n15143), .ZN(n15144) );
  OAI21_X1 U18521 ( .B1(n15782), .B2(n19891), .A(n15144), .ZN(P2_U2854) );
  MUX2_X1 U18522 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16205), .S(n15235), .Z(
        P2_U2856) );
  NAND2_X1 U18523 ( .A1(n15146), .A2(n15147), .ZN(n15239) );
  NAND3_X1 U18524 ( .A1(n15145), .A2(n15239), .A3(n15224), .ZN(n15149) );
  NAND2_X1 U18525 ( .A1(n15221), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15148) );
  OAI211_X1 U18526 ( .C1(n15221), .C2(n15499), .A(n15149), .B(n15148), .ZN(
        P2_U2858) );
  NOR2_X1 U18527 ( .A1(n15151), .A2(n15150), .ZN(n15152) );
  XOR2_X1 U18528 ( .A(n15153), .B(n15152), .Z(n15253) );
  AND2_X1 U18529 ( .A1(n9876), .A2(n15154), .ZN(n15155) );
  OR2_X1 U18530 ( .A1(n15155), .A2(n9880), .ZN(n16222) );
  NOR2_X1 U18531 ( .A1(n16222), .A2(n15221), .ZN(n15156) );
  AOI21_X1 U18532 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15221), .A(n15156), .ZN(
        n15157) );
  OAI21_X1 U18533 ( .B1(n15253), .B2(n15237), .A(n15157), .ZN(P2_U2859) );
  NAND2_X1 U18534 ( .A1(n15221), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15160) );
  OAI21_X1 U18535 ( .B1(n15161), .B2(n15163), .A(n15162), .ZN(n15268) );
  OR2_X1 U18536 ( .A1(n15165), .A2(n15164), .ZN(n15166) );
  NAND2_X1 U18537 ( .A1(n14975), .A2(n15166), .ZN(n16234) );
  NOR2_X1 U18538 ( .A1(n16234), .A2(n15221), .ZN(n15167) );
  AOI21_X1 U18539 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15221), .A(n15167), .ZN(
        n15168) );
  OAI21_X1 U18540 ( .B1(n15268), .B2(n15237), .A(n15168), .ZN(P2_U2861) );
  OAI21_X1 U18541 ( .B1(n15171), .B2(n15170), .A(n15169), .ZN(n15269) );
  MUX2_X1 U18542 ( .A(n15543), .B(n15172), .S(n15221), .Z(n15173) );
  OAI21_X1 U18543 ( .B1(n15269), .B2(n15237), .A(n15173), .ZN(P2_U2862) );
  AOI21_X1 U18544 ( .B1(n15175), .B2(n15174), .A(n9901), .ZN(n15176) );
  XOR2_X1 U18545 ( .A(n15177), .B(n15176), .Z(n15282) );
  AND2_X1 U18546 ( .A1(n15183), .A2(n15178), .ZN(n15180) );
  OR2_X1 U18547 ( .A1(n15180), .A2(n15179), .ZN(n16246) );
  NOR2_X1 U18548 ( .A1(n16246), .A2(n15221), .ZN(n15181) );
  AOI21_X1 U18549 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15221), .A(n15181), .ZN(
        n15182) );
  OAI21_X1 U18550 ( .B1(n15282), .B2(n15237), .A(n15182), .ZN(P2_U2863) );
  AOI21_X1 U18551 ( .B1(n15184), .B2(n15197), .A(n12604), .ZN(n16257) );
  INV_X1 U18552 ( .A(n16257), .ZN(n15190) );
  AOI21_X1 U18553 ( .B1(n15187), .B2(n15186), .A(n15185), .ZN(n16269) );
  NAND2_X1 U18554 ( .A1(n16269), .A2(n15224), .ZN(n15189) );
  NAND2_X1 U18555 ( .A1(n15221), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15188) );
  OAI211_X1 U18556 ( .C1(n15190), .C2(n15221), .A(n15189), .B(n15188), .ZN(
        P2_U2864) );
  AOI21_X1 U18557 ( .B1(n15192), .B2(n15191), .A(n13109), .ZN(n15193) );
  INV_X1 U18558 ( .A(n15193), .ZN(n15290) );
  OR2_X1 U18559 ( .A1(n15195), .A2(n15194), .ZN(n15196) );
  AND2_X1 U18560 ( .A1(n15197), .A2(n15196), .ZN(n15836) );
  INV_X1 U18561 ( .A(n15836), .ZN(n15391) );
  MUX2_X1 U18562 ( .A(n15391), .B(n15832), .S(n15221), .Z(n15198) );
  OAI21_X1 U18563 ( .B1(n15290), .B2(n15237), .A(n15198), .ZN(P2_U2865) );
  OAI21_X1 U18564 ( .B1(n15199), .B2(n15200), .A(n15191), .ZN(n15296) );
  MUX2_X1 U18565 ( .A(n12597), .B(n15409), .S(n15235), .Z(n15201) );
  OAI21_X1 U18566 ( .B1(n15296), .B2(n15237), .A(n15201), .ZN(P2_U2866) );
  AOI21_X1 U18567 ( .B1(n15203), .B2(n15202), .A(n15199), .ZN(n15305) );
  NAND2_X1 U18568 ( .A1(n15305), .A2(n15224), .ZN(n15209) );
  NAND2_X1 U18569 ( .A1(n15205), .A2(n15204), .ZN(n15206) );
  NAND2_X1 U18570 ( .A1(n19057), .A2(n15235), .ZN(n15208) );
  OAI211_X1 U18571 ( .C1(n15235), .C2(n12593), .A(n15209), .B(n15208), .ZN(
        P2_U2867) );
  INV_X1 U18572 ( .A(n15617), .ZN(n15215) );
  INV_X1 U18573 ( .A(n15202), .ZN(n15211) );
  AOI21_X1 U18574 ( .B1(n15212), .B2(n15210), .A(n15211), .ZN(n15312) );
  NAND2_X1 U18575 ( .A1(n15312), .A2(n15224), .ZN(n15214) );
  NAND2_X1 U18576 ( .A1(n15221), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15213) );
  OAI211_X1 U18577 ( .C1(n15215), .C2(n15221), .A(n15214), .B(n15213), .ZN(
        P2_U2868) );
  OAI21_X1 U18578 ( .B1(n14174), .B2(n15216), .A(n15210), .ZN(n15328) );
  OAI21_X1 U18579 ( .B1(n15218), .B2(n15217), .A(n15023), .ZN(n19067) );
  MUX2_X1 U18580 ( .A(n19061), .B(n19067), .S(n15235), .Z(n15219) );
  OAI21_X1 U18581 ( .B1(n15328), .B2(n15237), .A(n15219), .ZN(P2_U2869) );
  NOR2_X1 U18582 ( .A1(n15446), .A2(n15221), .ZN(n15220) );
  AOI21_X1 U18583 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15221), .A(n15220), .ZN(
        n15222) );
  OAI21_X1 U18584 ( .B1(n15223), .B2(n15237), .A(n15222), .ZN(P2_U2870) );
  NAND2_X1 U18585 ( .A1(n15225), .A2(n15224), .ZN(n15229) );
  OAI21_X1 U18586 ( .B1(n15233), .B2(n15227), .A(n15226), .ZN(n15643) );
  INV_X1 U18587 ( .A(n15643), .ZN(n19090) );
  NAND2_X1 U18588 ( .A1(n19090), .A2(n15235), .ZN(n15228) );
  OAI211_X1 U18589 ( .C1(n15235), .C2(n12409), .A(n15229), .B(n15228), .ZN(
        P2_U2871) );
  XNOR2_X1 U18590 ( .A(n14087), .B(n15230), .ZN(n15238) );
  NOR2_X1 U18591 ( .A1(n15231), .A2(n14090), .ZN(n15232) );
  NOR2_X1 U18592 ( .A1(n15233), .A2(n15232), .ZN(n19098) );
  NOR2_X1 U18593 ( .A1(n15235), .A2(n12337), .ZN(n15234) );
  AOI21_X1 U18594 ( .B1(n19098), .B2(n15235), .A(n15234), .ZN(n15236) );
  OAI21_X1 U18595 ( .B1(n15238), .B2(n15237), .A(n15236), .ZN(P2_U2872) );
  NAND3_X1 U18596 ( .A1(n15145), .A2(n15239), .A3(n16268), .ZN(n15243) );
  MUX2_X1 U18597 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n19316), .Z(n19258) );
  AOI22_X1 U18598 ( .A1(n16266), .A2(n19258), .B1(n19203), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15242) );
  AOI22_X1 U18599 ( .A1(n19200), .A2(BUF1_REG_29__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15241) );
  NAND2_X1 U18600 ( .A1(n15496), .A2(n19198), .ZN(n15240) );
  NAND4_X1 U18601 ( .A1(n15243), .A2(n15242), .A3(n15241), .A4(n15240), .ZN(
        P2_U2890) );
  OR2_X1 U18602 ( .A1(n15245), .A2(n15244), .ZN(n15246) );
  AOI22_X1 U18603 ( .A1(n16266), .A2(n15248), .B1(n19203), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15250) );
  AOI22_X1 U18604 ( .A1(n19200), .A2(BUF1_REG_28__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15249) );
  OAI211_X1 U18605 ( .C1(n16221), .C2(n15310), .A(n15250), .B(n15249), .ZN(
        n15251) );
  INV_X1 U18606 ( .A(n15251), .ZN(n15252) );
  OAI21_X1 U18607 ( .B1(n15253), .B2(n15327), .A(n15252), .ZN(P2_U2891) );
  AOI22_X1 U18608 ( .A1(n16266), .A2(n19209), .B1(n19203), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15255) );
  AOI22_X1 U18609 ( .A1(n19200), .A2(BUF1_REG_27__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15254) );
  OAI211_X1 U18610 ( .C1(n15516), .C2(n15310), .A(n15255), .B(n15254), .ZN(
        n15256) );
  AOI21_X1 U18611 ( .B1(n15257), .B2(n16268), .A(n15256), .ZN(n15258) );
  INV_X1 U18612 ( .A(n15258), .ZN(P2_U2892) );
  INV_X1 U18613 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n15259) );
  OAI22_X1 U18614 ( .A1(n15323), .A2(n15260), .B1(n15321), .B2(n15259), .ZN(
        n15265) );
  NOR2_X1 U18615 ( .A1(n9834), .A2(n15261), .ZN(n15262) );
  OR2_X1 U18616 ( .A1(n14983), .A2(n15262), .ZN(n16242) );
  OAI22_X1 U18617 ( .A1(n16242), .A2(n15310), .B1(n19217), .B2(n15263), .ZN(
        n15264) );
  AOI211_X1 U18618 ( .C1(n16266), .C2(n15266), .A(n15265), .B(n15264), .ZN(
        n15267) );
  OAI21_X1 U18619 ( .B1(n15268), .B2(n15327), .A(n15267), .ZN(P2_U2893) );
  OR2_X1 U18620 ( .A1(n15269), .A2(n15327), .ZN(n15273) );
  AOI22_X1 U18621 ( .A1(n16266), .A2(n19212), .B1(n19203), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15272) );
  AOI22_X1 U18622 ( .A1(n19200), .A2(BUF1_REG_25__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15271) );
  NAND2_X1 U18623 ( .A1(n15540), .A2(n19198), .ZN(n15270) );
  NAND4_X1 U18624 ( .A1(n15273), .A2(n15272), .A3(n15271), .A4(n15270), .ZN(
        P2_U2894) );
  NAND2_X1 U18625 ( .A1(n15569), .A2(n15274), .ZN(n15275) );
  NAND2_X1 U18626 ( .A1(n15276), .A2(n15275), .ZN(n16254) );
  OAI22_X1 U18627 ( .A1(n16254), .A2(n15310), .B1(n19217), .B2(n15277), .ZN(
        n15278) );
  AOI21_X1 U18628 ( .B1(n16266), .B2(n15279), .A(n15278), .ZN(n15281) );
  AOI22_X1 U18629 ( .A1(n19200), .A2(BUF1_REG_24__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15280) );
  OAI211_X1 U18630 ( .C1(n15282), .C2(n15327), .A(n15281), .B(n15280), .ZN(
        P2_U2895) );
  OAI21_X1 U18631 ( .B1(n15008), .B2(n15284), .A(n15283), .ZN(n15580) );
  INV_X1 U18632 ( .A(n15580), .ZN(n15835) );
  INV_X1 U18633 ( .A(n16266), .ZN(n15286) );
  OAI22_X1 U18634 ( .A1(n15286), .A2(n19359), .B1(n15285), .B2(n19217), .ZN(
        n15287) );
  AOI21_X1 U18635 ( .B1(n19198), .B2(n15835), .A(n15287), .ZN(n15289) );
  AOI22_X1 U18636 ( .A1(n19200), .A2(BUF1_REG_22__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n15288) );
  OAI211_X1 U18637 ( .C1(n15290), .C2(n15327), .A(n15289), .B(n15288), .ZN(
        P2_U2897) );
  AOI22_X1 U18638 ( .A1(n19200), .A2(BUF1_REG_21__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15293) );
  AOI22_X1 U18639 ( .A1(n16266), .A2(n15291), .B1(n19203), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15292) );
  OAI211_X1 U18640 ( .C1(n15310), .C2(n15593), .A(n15293), .B(n15292), .ZN(
        n15294) );
  INV_X1 U18641 ( .A(n15294), .ZN(n15295) );
  OAI21_X1 U18642 ( .B1(n15296), .B2(n15327), .A(n15295), .ZN(P2_U2898) );
  AND2_X1 U18643 ( .A1(n15298), .A2(n15297), .ZN(n15300) );
  OR2_X1 U18644 ( .A1(n15300), .A2(n15299), .ZN(n19060) );
  AOI22_X1 U18645 ( .A1(n19200), .A2(BUF1_REG_20__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n15303) );
  AOI22_X1 U18646 ( .A1(n16266), .A2(n15301), .B1(n19203), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15302) );
  OAI211_X1 U18647 ( .C1(n15310), .C2(n19060), .A(n15303), .B(n15302), .ZN(
        n15304) );
  AOI21_X1 U18648 ( .B1(n15305), .B2(n16268), .A(n15304), .ZN(n15306) );
  INV_X1 U18649 ( .A(n15306), .ZN(P2_U2899) );
  AOI22_X1 U18650 ( .A1(n19200), .A2(BUF1_REG_19__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15309) );
  AOI22_X1 U18651 ( .A1(n16266), .A2(n15307), .B1(n19203), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15308) );
  OAI211_X1 U18652 ( .C1(n15310), .C2(n15620), .A(n15309), .B(n15308), .ZN(
        n15311) );
  AOI21_X1 U18653 ( .B1(n15312), .B2(n16268), .A(n15311), .ZN(n15313) );
  INV_X1 U18654 ( .A(n15313), .ZN(P2_U2900) );
  OR2_X1 U18655 ( .A1(n12803), .A2(n15314), .ZN(n15315) );
  NAND2_X1 U18656 ( .A1(n15316), .A2(n15315), .ZN(n19072) );
  INV_X1 U18657 ( .A(n19072), .ZN(n15632) );
  NAND2_X1 U18658 ( .A1(n16266), .A2(n15317), .ZN(n15318) );
  OAI21_X1 U18659 ( .B1(n15319), .B2(n19217), .A(n15318), .ZN(n15325) );
  INV_X1 U18660 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n15320) );
  OAI22_X1 U18661 ( .A1(n15323), .A2(n15322), .B1(n15321), .B2(n15320), .ZN(
        n15324) );
  AOI211_X1 U18662 ( .C1(n19198), .C2(n15632), .A(n15325), .B(n15324), .ZN(
        n15326) );
  OAI21_X1 U18663 ( .B1(n15328), .B2(n15327), .A(n15326), .ZN(P2_U2901) );
  NOR2_X1 U18664 ( .A1(n15330), .A2(n12153), .ZN(n15333) );
  XNOR2_X1 U18665 ( .A(n15331), .B(n15333), .ZN(n15343) );
  INV_X1 U18666 ( .A(n15331), .ZN(n15332) );
  AOI22_X1 U18667 ( .A1(n15343), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n15333), .B2(n15332), .ZN(n15336) );
  XNOR2_X1 U18668 ( .A(n15334), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15335) );
  XNOR2_X1 U18669 ( .A(n15336), .B(n15335), .ZN(n15513) );
  AND2_X1 U18670 ( .A1(n15337), .A2(n15508), .ZN(n15338) );
  NOR2_X1 U18671 ( .A1(n12510), .A2(n15338), .ZN(n15511) );
  INV_X1 U18672 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19966) );
  NOR2_X1 U18673 ( .A1(n19966), .A2(n19150), .ZN(n15505) );
  NOR2_X1 U18674 ( .A1(n16366), .A2(n16226), .ZN(n15339) );
  AOI211_X1 U18675 ( .C1(n16355), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15505), .B(n15339), .ZN(n15340) );
  OAI21_X1 U18676 ( .B1(n16222), .B2(n19317), .A(n15340), .ZN(n15341) );
  AOI21_X1 U18677 ( .B1(n15511), .B2(n16350), .A(n15341), .ZN(n15342) );
  OAI21_X1 U18678 ( .B1(n15513), .B2(n19278), .A(n15342), .ZN(P2_U2986) );
  XNOR2_X1 U18679 ( .A(n15343), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15526) );
  INV_X1 U18680 ( .A(n15337), .ZN(n15345) );
  AOI21_X1 U18681 ( .B1(n15520), .B2(n15344), .A(n15345), .ZN(n15524) );
  NOR2_X1 U18682 ( .A1(n15514), .A2(n19317), .ZN(n15349) );
  NAND2_X1 U18683 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n19287), .ZN(n15515) );
  NAND2_X1 U18684 ( .A1(n16355), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15346) );
  OAI211_X1 U18685 ( .C1(n16366), .C2(n15347), .A(n15515), .B(n15346), .ZN(
        n15348) );
  AOI211_X1 U18686 ( .C1(n15524), .C2(n16350), .A(n15349), .B(n15348), .ZN(
        n15350) );
  OAI21_X1 U18687 ( .B1(n15526), .B2(n19278), .A(n15350), .ZN(P2_U2987) );
  INV_X1 U18688 ( .A(n15357), .ZN(n15351) );
  AOI21_X1 U18689 ( .B1(n15359), .B2(n15358), .A(n15351), .ZN(n15352) );
  XOR2_X1 U18690 ( .A(n15353), .B(n15352), .Z(n15539) );
  INV_X1 U18691 ( .A(n16234), .ZN(n15531) );
  NAND2_X1 U18692 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19287), .ZN(n15529) );
  NAND2_X1 U18693 ( .A1(n16355), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15354) );
  OAI211_X1 U18694 ( .C1(n16366), .C2(n16239), .A(n15529), .B(n15354), .ZN(
        n15356) );
  NAND2_X1 U18695 ( .A1(n15358), .A2(n15357), .ZN(n15360) );
  XOR2_X1 U18696 ( .A(n15360), .B(n15359), .Z(n15553) );
  INV_X1 U18697 ( .A(n9877), .ZN(n15361) );
  AOI21_X1 U18698 ( .B1(n15546), .B2(n15361), .A(n15355), .ZN(n15551) );
  INV_X1 U18699 ( .A(n15362), .ZN(n15365) );
  NAND2_X1 U18700 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19287), .ZN(n15542) );
  OAI21_X1 U18701 ( .B1(n19285), .B2(n15363), .A(n15542), .ZN(n15364) );
  AOI21_X1 U18702 ( .B1(n19270), .B2(n15365), .A(n15364), .ZN(n15366) );
  OAI21_X1 U18703 ( .B1(n15543), .B2(n19317), .A(n15366), .ZN(n15367) );
  AOI21_X1 U18704 ( .B1(n15551), .B2(n16350), .A(n15367), .ZN(n15368) );
  OAI21_X1 U18705 ( .B1(n15553), .B2(n19278), .A(n15368), .ZN(P2_U2989) );
  INV_X1 U18706 ( .A(n15369), .ZN(n15371) );
  NAND2_X1 U18707 ( .A1(n15371), .A2(n15370), .ZN(n15372) );
  XNOR2_X1 U18708 ( .A(n15373), .B(n15372), .ZN(n15567) );
  AOI21_X1 U18709 ( .B1(n15555), .B2(n9835), .A(n9877), .ZN(n15565) );
  NOR2_X1 U18710 ( .A1(n16246), .A2(n19317), .ZN(n15376) );
  NAND2_X1 U18711 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19287), .ZN(n15559) );
  NAND2_X1 U18712 ( .A1(n16355), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15374) );
  OAI211_X1 U18713 ( .C1(n16366), .C2(n16251), .A(n15559), .B(n15374), .ZN(
        n15375) );
  AOI211_X1 U18714 ( .C1(n15565), .C2(n16350), .A(n15376), .B(n15375), .ZN(
        n15377) );
  OAI21_X1 U18715 ( .B1(n15567), .B2(n19278), .A(n15377), .ZN(P2_U2990) );
  INV_X1 U18716 ( .A(n15378), .ZN(n15379) );
  OAI21_X1 U18717 ( .B1(n15379), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n9835), .ZN(n15579) );
  NAND2_X1 U18718 ( .A1(n19270), .A2(n15380), .ZN(n15381) );
  NAND2_X1 U18719 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19287), .ZN(n15571) );
  OAI211_X1 U18720 ( .C1(n19285), .C2(n10178), .A(n15381), .B(n15571), .ZN(
        n15384) );
  NOR3_X1 U18721 ( .A1(n15382), .A2(n15575), .A3(n19278), .ZN(n15383) );
  AOI211_X1 U18722 ( .C1(n19282), .C2(n16257), .A(n15384), .B(n15383), .ZN(
        n15385) );
  OAI21_X1 U18723 ( .B1(n19277), .B2(n15579), .A(n15385), .ZN(P2_U2991) );
  OAI21_X1 U18724 ( .B1(n15386), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15378), .ZN(n15589) );
  NAND2_X1 U18725 ( .A1(n9893), .A2(n15387), .ZN(n15388) );
  XNOR2_X1 U18726 ( .A(n15389), .B(n15388), .ZN(n15587) );
  OAI22_X1 U18727 ( .A1(n19954), .A2(n19150), .B1(n16366), .B2(n15839), .ZN(
        n15393) );
  INV_X1 U18728 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15390) );
  OAI22_X1 U18729 ( .A1(n15391), .A2(n19317), .B1(n15390), .B2(n19285), .ZN(
        n15392) );
  AOI211_X1 U18730 ( .C1(n15587), .C2(n16361), .A(n15393), .B(n15392), .ZN(
        n15394) );
  OAI21_X1 U18731 ( .B1(n19277), .B2(n15589), .A(n15394), .ZN(P2_U2992) );
  INV_X1 U18732 ( .A(n15413), .ZN(n15399) );
  AOI21_X1 U18733 ( .B1(n15415), .B2(n15399), .A(n15412), .ZN(n15403) );
  NAND2_X1 U18734 ( .A1(n15401), .A2(n15400), .ZN(n15402) );
  XNOR2_X1 U18735 ( .A(n15403), .B(n15402), .ZN(n15601) );
  AOI21_X1 U18736 ( .B1(n15405), .B2(n15404), .A(n15386), .ZN(n15598) );
  NOR2_X1 U18737 ( .A1(n19952), .A2(n19150), .ZN(n15590) );
  NOR2_X1 U18738 ( .A1(n16366), .A2(n15406), .ZN(n15407) );
  AOI211_X1 U18739 ( .C1(n16355), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15590), .B(n15407), .ZN(n15408) );
  OAI21_X1 U18740 ( .B1(n15409), .B2(n19317), .A(n15408), .ZN(n15410) );
  AOI21_X1 U18741 ( .B1(n15598), .B2(n16350), .A(n15410), .ZN(n15411) );
  OAI21_X1 U18742 ( .B1(n15601), .B2(n19278), .A(n15411), .ZN(P2_U2993) );
  NOR2_X1 U18743 ( .A1(n15413), .A2(n15412), .ZN(n15414) );
  XNOR2_X1 U18744 ( .A(n15415), .B(n15414), .ZN(n15616) );
  INV_X1 U18745 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19950) );
  NOR2_X1 U18746 ( .A1(n19950), .A2(n19150), .ZN(n15602) );
  AOI21_X1 U18747 ( .B1(n16355), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15602), .ZN(n15416) );
  OAI21_X1 U18748 ( .B1(n16366), .B2(n19053), .A(n15416), .ZN(n15420) );
  INV_X1 U18749 ( .A(n15417), .ZN(n15418) );
  OAI21_X1 U18750 ( .B1(n15418), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15404), .ZN(n15613) );
  NOR2_X1 U18751 ( .A1(n15613), .A2(n19277), .ZN(n15419) );
  AOI211_X1 U18752 ( .C1(n19282), .C2(n19057), .A(n15420), .B(n15419), .ZN(
        n15421) );
  OAI21_X1 U18753 ( .B1(n15616), .B2(n19278), .A(n15421), .ZN(P2_U2994) );
  NAND2_X1 U18754 ( .A1(n15423), .A2(n15422), .ZN(n15427) );
  INV_X1 U18755 ( .A(n15437), .ZN(n15424) );
  NOR2_X1 U18756 ( .A1(n15425), .A2(n15424), .ZN(n15426) );
  XOR2_X1 U18757 ( .A(n15427), .B(n15426), .Z(n15627) );
  NAND2_X1 U18758 ( .A1(n15428), .A2(n15604), .ZN(n15624) );
  NAND3_X1 U18759 ( .A1(n15417), .A2(n16350), .A3(n15624), .ZN(n15432) );
  NAND2_X1 U18760 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n19287), .ZN(n15618) );
  OAI21_X1 U18761 ( .B1(n19285), .B2(n15429), .A(n15618), .ZN(n15430) );
  AOI21_X1 U18762 ( .B1(n15617), .B2(n19282), .A(n15430), .ZN(n15431) );
  OAI211_X1 U18763 ( .C1(n16366), .C2(n15433), .A(n15432), .B(n15431), .ZN(
        n15434) );
  INV_X1 U18764 ( .A(n15434), .ZN(n15435) );
  OAI21_X1 U18765 ( .B1(n15627), .B2(n19278), .A(n15435), .ZN(P2_U2995) );
  NAND2_X1 U18766 ( .A1(n15437), .A2(n15436), .ZN(n15438) );
  XNOR2_X1 U18767 ( .A(n15439), .B(n15438), .ZN(n15639) );
  INV_X1 U18768 ( .A(n15428), .ZN(n15440) );
  NOR2_X1 U18769 ( .A1(n9869), .A2(n15440), .ZN(n15637) );
  NOR2_X1 U18770 ( .A1(n19946), .A2(n19150), .ZN(n15631) );
  NOR2_X1 U18771 ( .A1(n19067), .A2(n19317), .ZN(n15441) );
  AOI211_X1 U18772 ( .C1(n16355), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15631), .B(n15441), .ZN(n15442) );
  OAI21_X1 U18773 ( .B1(n15443), .B2(n16366), .A(n15442), .ZN(n15444) );
  AOI21_X1 U18774 ( .B1(n15637), .B2(n16350), .A(n15444), .ZN(n15445) );
  OAI21_X1 U18775 ( .B1(n15639), .B2(n19278), .A(n15445), .ZN(P2_U2996) );
  INV_X1 U18776 ( .A(n15446), .ZN(n19081) );
  NOR2_X1 U18777 ( .A1(n19944), .A2(n19150), .ZN(n15449) );
  INV_X1 U18778 ( .A(n19075), .ZN(n19084) );
  OAI22_X1 U18779 ( .A1(n15447), .A2(n19285), .B1(n16366), .B2(n19084), .ZN(
        n15448) );
  AOI211_X1 U18780 ( .C1(n19282), .C2(n19081), .A(n15449), .B(n15448), .ZN(
        n15453) );
  XNOR2_X1 U18781 ( .A(n15459), .B(n15450), .ZN(n15451) );
  NAND2_X1 U18782 ( .A1(n15451), .A2(n16350), .ZN(n15452) );
  OAI211_X1 U18783 ( .C1(n15454), .C2(n19278), .A(n15453), .B(n15452), .ZN(
        P2_U2997) );
  XOR2_X1 U18784 ( .A(n15456), .B(n15455), .Z(n15647) );
  INV_X1 U18785 ( .A(n15647), .ZN(n15462) );
  NOR2_X1 U18786 ( .A1(n19942), .A2(n19150), .ZN(n15458) );
  OAI22_X1 U18787 ( .A1(n10181), .A2(n19285), .B1(n16366), .B2(n19089), .ZN(
        n15457) );
  AOI211_X1 U18788 ( .C1(n19282), .C2(n19090), .A(n15458), .B(n15457), .ZN(
        n15461) );
  INV_X1 U18789 ( .A(n15642), .ZN(n16274) );
  OAI211_X1 U18790 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16274), .A(
        n10151), .B(n16350), .ZN(n15460) );
  OAI211_X1 U18791 ( .C1(n15462), .C2(n19278), .A(n15461), .B(n15460), .ZN(
        P2_U2998) );
  OAI21_X1 U18792 ( .B1(n15465), .B2(n15464), .A(n15463), .ZN(n15466) );
  INV_X1 U18793 ( .A(n15466), .ZN(n16414) );
  NAND2_X1 U18794 ( .A1(n15467), .A2(n15714), .ZN(n15468) );
  NAND2_X1 U18795 ( .A1(n15468), .A2(n15715), .ZN(n15472) );
  AND2_X1 U18796 ( .A1(n15470), .A2(n15469), .ZN(n15471) );
  XNOR2_X1 U18797 ( .A(n15472), .B(n15471), .ZN(n16417) );
  AOI22_X1 U18798 ( .A1(n19282), .A2(n19142), .B1(n16355), .B2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15476) );
  INV_X1 U18799 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19927) );
  OAI22_X1 U18800 ( .A1(n19927), .A2(n19150), .B1(n16366), .B2(n15473), .ZN(
        n15474) );
  INV_X1 U18801 ( .A(n15474), .ZN(n15475) );
  OAI211_X1 U18802 ( .C1(n16417), .C2(n19278), .A(n15476), .B(n15475), .ZN(
        n15477) );
  AOI21_X1 U18803 ( .B1(n16414), .B2(n16350), .A(n15477), .ZN(n15478) );
  INV_X1 U18804 ( .A(n15478), .ZN(P2_U3006) );
  OAI21_X1 U18805 ( .B1(n15480), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15479), .ZN(n15725) );
  XOR2_X1 U18806 ( .A(n15482), .B(n15481), .Z(n15724) );
  NAND2_X1 U18807 ( .A1(n15724), .A2(n16361), .ZN(n15487) );
  INV_X1 U18808 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19924) );
  OAI22_X1 U18809 ( .A1(n19151), .A2(n19285), .B1(n19924), .B2(n19150), .ZN(
        n15485) );
  INV_X1 U18810 ( .A(n19149), .ZN(n15483) );
  NOR2_X1 U18811 ( .A1(n16366), .A2(n15483), .ZN(n15484) );
  AOI211_X1 U18812 ( .C1(n19155), .C2(n19282), .A(n15485), .B(n15484), .ZN(
        n15486) );
  OAI211_X1 U18813 ( .C1(n19277), .C2(n15725), .A(n15487), .B(n15486), .ZN(
        P2_U3008) );
  INV_X1 U18814 ( .A(n15488), .ZN(n15502) );
  INV_X1 U18815 ( .A(n15493), .ZN(n15489) );
  NOR2_X1 U18816 ( .A1(n15489), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15523) );
  INV_X1 U18817 ( .A(n15521), .ZN(n15490) );
  NOR2_X1 U18818 ( .A1(n15523), .A2(n15490), .ZN(n15509) );
  AND2_X1 U18819 ( .A1(n15508), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15491) );
  NAND2_X1 U18820 ( .A1(n15493), .A2(n15491), .ZN(n15507) );
  AOI21_X1 U18821 ( .B1(n15509), .B2(n15507), .A(n15492), .ZN(n15501) );
  NAND4_X1 U18822 ( .A1(n15493), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A4(n15492), .ZN(n15498) );
  INV_X1 U18823 ( .A(n15494), .ZN(n15495) );
  AOI21_X1 U18824 ( .B1(n15496), .B2(n16387), .A(n15495), .ZN(n15497) );
  OAI211_X1 U18825 ( .C1(n19308), .C2(n15499), .A(n15498), .B(n15497), .ZN(
        n15500) );
  OAI21_X1 U18826 ( .B1(n15504), .B2(n19314), .A(n15503), .ZN(P2_U3017) );
  INV_X1 U18827 ( .A(n16222), .ZN(n15506) );
  AOI21_X1 U18828 ( .B1(n15511), .B2(n16413), .A(n15510), .ZN(n15512) );
  OAI21_X1 U18829 ( .B1(n15513), .B2(n19314), .A(n15512), .ZN(P2_U3018) );
  INV_X1 U18830 ( .A(n15514), .ZN(n15518) );
  OAI21_X1 U18831 ( .B1(n15516), .B2(n19301), .A(n15515), .ZN(n15517) );
  AOI21_X1 U18832 ( .B1(n15518), .B2(n16412), .A(n15517), .ZN(n15519) );
  OAI21_X1 U18833 ( .B1(n15521), .B2(n15520), .A(n15519), .ZN(n15522) );
  AOI211_X1 U18834 ( .C1(n15524), .C2(n16413), .A(n15523), .B(n15522), .ZN(
        n15525) );
  OAI21_X1 U18835 ( .B1(n15526), .B2(n19314), .A(n15525), .ZN(P2_U3019) );
  OAI21_X1 U18836 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n15527), .ZN(n15528) );
  INV_X1 U18837 ( .A(n15528), .ZN(n15537) );
  NAND2_X1 U18838 ( .A1(n15545), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15533) );
  OAI21_X1 U18839 ( .B1(n16242), .B2(n19301), .A(n15529), .ZN(n15530) );
  AOI21_X1 U18840 ( .B1(n15531), .B2(n16412), .A(n15530), .ZN(n15532) );
  NAND2_X1 U18841 ( .A1(n15533), .A2(n15532), .ZN(n15536) );
  NOR2_X1 U18842 ( .A1(n15534), .A2(n19303), .ZN(n15535) );
  AOI211_X1 U18843 ( .C1(n15547), .C2(n15537), .A(n15536), .B(n15535), .ZN(
        n15538) );
  OAI21_X1 U18844 ( .B1(n15539), .B2(n19314), .A(n15538), .ZN(P2_U3020) );
  NAND2_X1 U18845 ( .A1(n15540), .A2(n16387), .ZN(n15541) );
  OAI211_X1 U18846 ( .C1(n15543), .C2(n19308), .A(n15542), .B(n15541), .ZN(
        n15544) );
  AOI21_X1 U18847 ( .B1(n15545), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15544), .ZN(n15549) );
  NAND2_X1 U18848 ( .A1(n15547), .A2(n15546), .ZN(n15548) );
  NAND2_X1 U18849 ( .A1(n15549), .A2(n15548), .ZN(n15550) );
  AOI21_X1 U18850 ( .B1(n15551), .B2(n16413), .A(n15550), .ZN(n15552) );
  OAI21_X1 U18851 ( .B1(n15553), .B2(n19314), .A(n15552), .ZN(P2_U3021) );
  NAND2_X1 U18852 ( .A1(n15555), .A2(n15554), .ZN(n15563) );
  INV_X1 U18853 ( .A(n16246), .ZN(n15561) );
  INV_X1 U18854 ( .A(n15556), .ZN(n15557) );
  NAND2_X1 U18855 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15557), .ZN(
        n15558) );
  OAI211_X1 U18856 ( .C1(n16254), .C2(n19301), .A(n15559), .B(n15558), .ZN(
        n15560) );
  AOI21_X1 U18857 ( .B1(n15561), .B2(n16412), .A(n15560), .ZN(n15562) );
  OAI21_X1 U18858 ( .B1(n15585), .B2(n15563), .A(n15562), .ZN(n15564) );
  AOI21_X1 U18859 ( .B1(n15565), .B2(n16413), .A(n15564), .ZN(n15566) );
  OAI21_X1 U18860 ( .B1(n15567), .B2(n19314), .A(n15566), .ZN(P2_U3022) );
  OAI21_X1 U18861 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n15568), .ZN(n15574) );
  INV_X1 U18862 ( .A(n15283), .ZN(n15570) );
  OAI21_X1 U18863 ( .B1(n15570), .B2(n10345), .A(n15569), .ZN(n16256) );
  OAI21_X1 U18864 ( .B1(n16256), .B2(n19301), .A(n15571), .ZN(n15572) );
  AOI21_X1 U18865 ( .B1(n16257), .B2(n16412), .A(n15572), .ZN(n15573) );
  OAI21_X1 U18866 ( .B1(n15585), .B2(n15574), .A(n15573), .ZN(n15577) );
  NOR3_X1 U18867 ( .A1(n15382), .A2(n15575), .A3(n19314), .ZN(n15576) );
  AOI211_X1 U18868 ( .C1(n15597), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15577), .B(n15576), .ZN(n15578) );
  OAI21_X1 U18869 ( .B1(n19303), .B2(n15579), .A(n15578), .ZN(P2_U3023) );
  NAND2_X1 U18870 ( .A1(n15597), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15584) );
  NOR2_X1 U18871 ( .A1(n19954), .A2(n19150), .ZN(n15582) );
  NOR2_X1 U18872 ( .A1(n19301), .A2(n15580), .ZN(n15581) );
  AOI211_X1 U18873 ( .C1(n15836), .C2(n16412), .A(n15582), .B(n15581), .ZN(
        n15583) );
  OAI211_X1 U18874 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15585), .A(
        n15584), .B(n15583), .ZN(n15586) );
  AOI21_X1 U18875 ( .B1(n15587), .B2(n19296), .A(n15586), .ZN(n15588) );
  OAI21_X1 U18876 ( .B1(n19303), .B2(n15589), .A(n15588), .ZN(P2_U3024) );
  AOI21_X1 U18877 ( .B1(n15591), .B2(n16412), .A(n15590), .ZN(n15592) );
  OAI21_X1 U18878 ( .B1(n19301), .B2(n15593), .A(n15592), .ZN(n15596) );
  NAND2_X1 U18879 ( .A1(n16393), .A2(n15609), .ZN(n15610) );
  NOR3_X1 U18880 ( .A1(n15610), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15594), .ZN(n15595) );
  AOI211_X1 U18881 ( .C1(n15597), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15596), .B(n15595), .ZN(n15600) );
  NAND2_X1 U18882 ( .A1(n15598), .A2(n16413), .ZN(n15599) );
  OAI211_X1 U18883 ( .C1(n15601), .C2(n19314), .A(n15600), .B(n15599), .ZN(
        P2_U3025) );
  INV_X1 U18884 ( .A(n15602), .ZN(n15603) );
  OAI21_X1 U18885 ( .B1(n19301), .B2(n19060), .A(n15603), .ZN(n15606) );
  NOR3_X1 U18886 ( .A1(n15610), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15604), .ZN(n15605) );
  AOI211_X1 U18887 ( .C1(n19057), .C2(n16412), .A(n15606), .B(n15605), .ZN(
        n15612) );
  OAI21_X1 U18888 ( .B1(n15609), .B2(n15608), .A(n15607), .ZN(n15623) );
  NOR2_X1 U18889 ( .A1(n15610), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15621) );
  OAI21_X1 U18890 ( .B1(n15623), .B2(n15621), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15611) );
  OAI211_X1 U18891 ( .C1(n15613), .C2(n19303), .A(n15612), .B(n15611), .ZN(
        n15614) );
  INV_X1 U18892 ( .A(n15614), .ZN(n15615) );
  OAI21_X1 U18893 ( .B1(n15616), .B2(n19314), .A(n15615), .ZN(P2_U3026) );
  NAND2_X1 U18894 ( .A1(n15617), .A2(n16412), .ZN(n15619) );
  OAI211_X1 U18895 ( .C1(n19301), .C2(n15620), .A(n15619), .B(n15618), .ZN(
        n15622) );
  AOI211_X1 U18896 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15623), .A(
        n15622), .B(n15621), .ZN(n15626) );
  NAND3_X1 U18897 ( .A1(n15417), .A2(n16413), .A3(n15624), .ZN(n15625) );
  OAI211_X1 U18898 ( .C1(n15627), .C2(n19314), .A(n15626), .B(n15625), .ZN(
        P2_U3027) );
  AOI211_X1 U18899 ( .C1(n15628), .C2(n15630), .A(n15688), .B(n15629), .ZN(
        n15636) );
  NAND3_X1 U18900 ( .A1(n15640), .A2(n15630), .A3(n15629), .ZN(n15634) );
  AOI21_X1 U18901 ( .B1(n16387), .B2(n15632), .A(n15631), .ZN(n15633) );
  OAI211_X1 U18902 ( .C1(n19067), .C2(n19308), .A(n15634), .B(n15633), .ZN(
        n15635) );
  AOI211_X1 U18903 ( .C1(n15637), .C2(n16413), .A(n15636), .B(n15635), .ZN(
        n15638) );
  OAI21_X1 U18904 ( .B1(n15639), .B2(n19314), .A(n15638), .ZN(P2_U3028) );
  INV_X1 U18905 ( .A(n15640), .ZN(n15659) );
  OAI22_X1 U18906 ( .A1(n15642), .A2(n19303), .B1(n15641), .B2(n15659), .ZN(
        n15646) );
  NOR2_X1 U18907 ( .A1(n19308), .A2(n15643), .ZN(n15645) );
  OAI22_X1 U18908 ( .A1(n19301), .A2(n19094), .B1(n19942), .B2(n19150), .ZN(
        n15644) );
  AOI211_X1 U18909 ( .C1(n15646), .C2(n15650), .A(n15645), .B(n15644), .ZN(
        n15649) );
  NAND2_X1 U18910 ( .A1(n15647), .A2(n19296), .ZN(n15648) );
  OAI211_X1 U18911 ( .C1(n15651), .C2(n15650), .A(n15649), .B(n15648), .ZN(
        P2_U3030) );
  NAND2_X1 U18912 ( .A1(n15653), .A2(n15652), .ZN(n15655) );
  XOR2_X1 U18913 ( .A(n15655), .B(n15654), .Z(n16276) );
  INV_X1 U18914 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19940) );
  NOR2_X1 U18915 ( .A1(n19940), .A2(n19150), .ZN(n15657) );
  NOR2_X1 U18916 ( .A1(n19301), .A2(n19110), .ZN(n15656) );
  AOI211_X1 U18917 ( .C1(n19098), .C2(n16412), .A(n15657), .B(n15656), .ZN(
        n15658) );
  OAI21_X1 U18918 ( .B1(n15659), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15658), .ZN(n15661) );
  NOR2_X1 U18919 ( .A1(n15664), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16275) );
  NOR3_X1 U18920 ( .A1(n16275), .A2(n16274), .A3(n19303), .ZN(n15660) );
  AOI211_X1 U18921 ( .C1(n15662), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15661), .B(n15660), .ZN(n15663) );
  OAI21_X1 U18922 ( .B1(n16276), .B2(n19314), .A(n15663), .ZN(P2_U3031) );
  INV_X1 U18923 ( .A(n16293), .ZN(n15666) );
  INV_X1 U18924 ( .A(n15664), .ZN(n15665) );
  OAI21_X1 U18925 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15666), .A(
        n15665), .ZN(n16282) );
  INV_X1 U18926 ( .A(n15668), .ZN(n15671) );
  AND2_X1 U18927 ( .A1(n15668), .A2(n15667), .ZN(n15670) );
  OAI22_X1 U18928 ( .A1(n15672), .A2(n15671), .B1(n15670), .B2(n15669), .ZN(
        n16283) );
  NOR2_X1 U18929 ( .A1(n15673), .A2(n16369), .ZN(n15677) );
  INV_X1 U18930 ( .A(n15673), .ZN(n15674) );
  OAI22_X1 U18931 ( .A1(n15687), .A2(n15688), .B1(n15674), .B2(n16369), .ZN(
        n16371) );
  INV_X1 U18932 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19938) );
  NOR2_X1 U18933 ( .A1(n19938), .A2(n19150), .ZN(n15675) );
  AOI221_X1 U18934 ( .B1(n15677), .B2(n15676), .C1(n16371), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n15675), .ZN(n15684) );
  OR2_X1 U18935 ( .A1(n15679), .A2(n15678), .ZN(n15681) );
  NAND2_X1 U18936 ( .A1(n15681), .A2(n15680), .ZN(n19205) );
  INV_X1 U18937 ( .A(n19205), .ZN(n15682) );
  AOI22_X1 U18938 ( .A1(n16387), .A2(n15682), .B1(n16412), .B2(n19117), .ZN(
        n15683) );
  OAI211_X1 U18939 ( .C1(n16283), .C2(n19314), .A(n15684), .B(n15683), .ZN(
        n15685) );
  INV_X1 U18940 ( .A(n15685), .ZN(n15686) );
  OAI21_X1 U18941 ( .B1(n19303), .B2(n16282), .A(n15686), .ZN(P2_U3032) );
  XNOR2_X1 U18942 ( .A(n16316), .B(n16368), .ZN(n16303) );
  INV_X1 U18943 ( .A(n16369), .ZN(n15699) );
  NOR2_X1 U18944 ( .A1(n15688), .A2(n15687), .ZN(n15691) );
  INV_X1 U18945 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19934) );
  NOR2_X1 U18946 ( .A1(n19934), .A2(n19150), .ZN(n15690) );
  NOR2_X1 U18947 ( .A1(n19308), .A2(n16301), .ZN(n15689) );
  AOI211_X1 U18948 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15691), .A(
        n15690), .B(n15689), .ZN(n15692) );
  OAI21_X1 U18949 ( .B1(n19301), .B2(n19132), .A(n15692), .ZN(n15698) );
  NOR2_X1 U18950 ( .A1(n15694), .A2(n15693), .ZN(n15695) );
  XNOR2_X1 U18951 ( .A(n15696), .B(n15695), .ZN(n16302) );
  NOR2_X1 U18952 ( .A1(n16302), .A2(n19314), .ZN(n15697) );
  AOI211_X1 U18953 ( .C1(n15699), .C2(n16368), .A(n15698), .B(n15697), .ZN(
        n15700) );
  OAI21_X1 U18954 ( .B1(n19303), .B2(n16303), .A(n15700), .ZN(P2_U3034) );
  NAND2_X1 U18955 ( .A1(n16325), .A2(n16309), .ZN(n15704) );
  INV_X1 U18956 ( .A(n16309), .ZN(n16324) );
  OAI21_X1 U18957 ( .B1(n15702), .B2(n16324), .A(n15701), .ZN(n15703) );
  NAND2_X1 U18958 ( .A1(n15704), .A2(n15703), .ZN(n16339) );
  NOR2_X1 U18959 ( .A1(n12508), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16337) );
  INV_X1 U18960 ( .A(n16323), .ZN(n16336) );
  OR3_X1 U18961 ( .A1(n16337), .A2(n16336), .A3(n19303), .ZN(n15711) );
  OAI22_X1 U18962 ( .A1(n19308), .A2(n16338), .B1(n19929), .B2(n19150), .ZN(
        n15709) );
  INV_X1 U18963 ( .A(n16393), .ZN(n15706) );
  AOI21_X1 U18964 ( .B1(n15707), .B2(n15706), .A(n15705), .ZN(n15708) );
  AOI211_X1 U18965 ( .C1(n16387), .C2(n19214), .A(n15709), .B(n15708), .ZN(
        n15710) );
  OAI211_X1 U18966 ( .C1(n16339), .C2(n19314), .A(n15711), .B(n15710), .ZN(
        P2_U3037) );
  OAI21_X1 U18967 ( .B1(n15712), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15713), .ZN(n16348) );
  NAND2_X1 U18968 ( .A1(n15715), .A2(n15714), .ZN(n15716) );
  XNOR2_X1 U18969 ( .A(n15467), .B(n15716), .ZN(n16349) );
  NAND2_X1 U18970 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19287), .ZN(n15717) );
  OAI221_X1 U18971 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16408), .C1(
        n15719), .C2(n15718), .A(n15717), .ZN(n15722) );
  OAI22_X1 U18972 ( .A1(n15720), .A2(n19301), .B1(n19308), .B2(n16354), .ZN(
        n15721) );
  AOI211_X1 U18973 ( .C1(n16349), .C2(n19296), .A(n15722), .B(n15721), .ZN(
        n15723) );
  OAI21_X1 U18974 ( .B1(n16348), .B2(n19303), .A(n15723), .ZN(P2_U3039) );
  INV_X1 U18975 ( .A(n15724), .ZN(n15733) );
  INV_X1 U18976 ( .A(n15725), .ZN(n15731) );
  NAND2_X1 U18977 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15726), .ZN(
        n19291) );
  NOR2_X1 U18978 ( .A1(n15739), .A2(n19291), .ZN(n15727) );
  MUX2_X1 U18979 ( .A(n15727), .B(n16411), .S(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n15730) );
  AOI22_X1 U18980 ( .A1(n16412), .A2(n19155), .B1(n19287), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n15728) );
  OAI21_X1 U18981 ( .B1(n19158), .B2(n19301), .A(n15728), .ZN(n15729) );
  AOI211_X1 U18982 ( .C1(n15731), .C2(n16413), .A(n15730), .B(n15729), .ZN(
        n15732) );
  OAI21_X1 U18983 ( .B1(n15733), .B2(n19314), .A(n15732), .ZN(P2_U3040) );
  XOR2_X1 U18984 ( .A(n15735), .B(n15734), .Z(n16362) );
  INV_X1 U18985 ( .A(n16362), .ZN(n15751) );
  INV_X1 U18986 ( .A(n15736), .ZN(n15744) );
  OAI22_X1 U18987 ( .A1(n19308), .A2(n16356), .B1(n19922), .B2(n19150), .ZN(
        n15743) );
  AOI21_X1 U18988 ( .B1(n15738), .B2(n19305), .A(n15737), .ZN(n19289) );
  OAI21_X1 U18989 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n15739), .ZN(n15740) );
  OAI22_X1 U18990 ( .A1(n19289), .A2(n15741), .B1(n19291), .B2(n15740), .ZN(
        n15742) );
  AOI211_X1 U18991 ( .C1(n16387), .C2(n15744), .A(n15743), .B(n15742), .ZN(
        n15750) );
  NOR2_X1 U18992 ( .A1(n10042), .A2(n15745), .ZN(n16358) );
  AOI21_X1 U18993 ( .B1(n15748), .B2(n15747), .A(n15746), .ZN(n16357) );
  OR3_X1 U18994 ( .A1(n16358), .A2(n16357), .A3(n19303), .ZN(n15749) );
  OAI211_X1 U18995 ( .C1(n15751), .C2(n19314), .A(n15750), .B(n15749), .ZN(
        P2_U3041) );
  INV_X1 U18996 ( .A(n15753), .ZN(n15754) );
  NOR2_X1 U18997 ( .A1(n15755), .A2(n15754), .ZN(n16447) );
  INV_X1 U18998 ( .A(n16447), .ZN(n15756) );
  AOI22_X1 U18999 ( .A1(n12974), .A2(n16451), .B1(n15761), .B2(n15756), .ZN(
        n16454) );
  INV_X1 U19000 ( .A(n16454), .ZN(n15760) );
  INV_X1 U19001 ( .A(n19995), .ZN(n16491) );
  NOR2_X1 U19002 ( .A1(n15758), .A2(n15757), .ZN(n19191) );
  AOI21_X1 U19003 ( .B1(n15758), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19191), .ZN(n15784) );
  AOI222_X1 U19004 ( .A1(n15760), .A2(n15785), .B1(n15759), .B2(n16491), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15784), .ZN(n15763) );
  AOI21_X1 U19005 ( .B1(n15785), .B2(n11897), .A(n19996), .ZN(n15762) );
  OAI22_X1 U19006 ( .A1(n15763), .A2(n19996), .B1(n15762), .B2(n15761), .ZN(
        P2_U3601) );
  NAND2_X1 U19007 ( .A1(n15764), .A2(n16451), .ZN(n15781) );
  INV_X1 U19008 ( .A(n15766), .ZN(n15767) );
  NAND2_X1 U19009 ( .A1(n11897), .A2(n15767), .ZN(n16426) );
  INV_X1 U19010 ( .A(n15768), .ZN(n16450) );
  NAND2_X1 U19011 ( .A1(n16450), .A2(n15769), .ZN(n16430) );
  INV_X1 U19012 ( .A(n16430), .ZN(n15771) );
  NAND2_X1 U19013 ( .A1(n16443), .A2(n15770), .ZN(n16431) );
  OAI21_X1 U19014 ( .B1(n15772), .B2(n15771), .A(n16431), .ZN(n15778) );
  NAND2_X1 U19015 ( .A1(n15773), .A2(n11865), .ZN(n15775) );
  NAND2_X1 U19016 ( .A1(n15775), .A2(n9811), .ZN(n16427) );
  INV_X1 U19017 ( .A(n16427), .ZN(n15776) );
  NAND2_X1 U19018 ( .A1(n15776), .A2(n16430), .ZN(n15777) );
  OAI211_X1 U19019 ( .C1(n15765), .C2(n16426), .A(n15778), .B(n15777), .ZN(
        n15779) );
  INV_X1 U19020 ( .A(n15779), .ZN(n15780) );
  NAND2_X1 U19021 ( .A1(n15781), .A2(n15780), .ZN(n16436) );
  OAI21_X1 U19022 ( .B1(n9807), .B2(n15783), .A(n15782), .ZN(n19991) );
  NOR2_X1 U19023 ( .A1(n15784), .A2(n16478), .ZN(n19990) );
  AOI222_X1 U19024 ( .A1(n16436), .A2(n15785), .B1(n19991), .B2(n19990), .C1(
        n16491), .C2(n19466), .ZN(n15787) );
  NAND2_X1 U19025 ( .A1(n19996), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15786) );
  OAI21_X1 U19026 ( .B1(n15787), .B2(n19996), .A(n15786), .ZN(P2_U3599) );
  INV_X1 U19027 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15789) );
  AOI22_X1 U19028 ( .A1(n11300), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15788) );
  OAI21_X1 U19029 ( .B1(n17219), .B2(n15789), .A(n15788), .ZN(n15800) );
  AOI22_X1 U19030 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15797) );
  AOI22_X1 U19031 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15790) );
  OAI21_X1 U19032 ( .B1(n10328), .B2(n17114), .A(n15790), .ZN(n15795) );
  AOI22_X1 U19033 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15793) );
  AOI22_X1 U19034 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15792) );
  OAI211_X1 U19035 ( .C1(n11489), .C2(n17120), .A(n15793), .B(n15792), .ZN(
        n15794) );
  AOI211_X1 U19036 ( .C1(n9804), .C2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n15795), .B(n15794), .ZN(n15796) );
  OAI211_X1 U19037 ( .C1(n15798), .C2(n17116), .A(n15797), .B(n15796), .ZN(
        n15799) );
  AOI211_X1 U19038 ( .C1(n11331), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15800), .B(n15799), .ZN(n17443) );
  INV_X1 U19039 ( .A(n17328), .ZN(n15801) );
  NOR2_X1 U19040 ( .A1(n15802), .A2(n15801), .ZN(n17227) );
  NAND2_X1 U19041 ( .A1(n15803), .A2(n17328), .ZN(n17256) );
  INV_X1 U19042 ( .A(n17256), .ZN(n17272) );
  AOI22_X1 U19043 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17336), .B1(
        P3_EBX_REG_12__SCAN_IN), .B2(n17272), .ZN(n15804) );
  OAI22_X1 U19044 ( .A1(n17443), .A2(n17324), .B1(n17227), .B2(n15804), .ZN(
        P3_U2690) );
  NAND2_X1 U19045 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18492) );
  NOR2_X1 U19046 ( .A1(n19003), .A2(n18855), .ZN(n15806) );
  AOI221_X1 U19047 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18492), .C1(n15806), 
        .C2(n18492), .A(n15805), .ZN(n18309) );
  NOR2_X1 U19048 ( .A1(n15807), .A2(n18821), .ZN(n15808) );
  OAI21_X1 U19049 ( .B1(n15808), .B2(n18613), .A(n18310), .ZN(n18307) );
  AOI22_X1 U19050 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18309), .B1(
        n18307), .B2(n18826), .ZN(P3_U2865) );
  NAND2_X1 U19051 ( .A1(n18779), .A2(n19009), .ZN(n15815) );
  OR2_X1 U19052 ( .A1(n16646), .A2(n17541), .ZN(n18839) );
  AOI211_X1 U19053 ( .C1(n15813), .C2(n18772), .A(n15909), .B(n15812), .ZN(
        n15814) );
  NOR2_X1 U19054 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18954), .ZN(n18313) );
  INV_X1 U19055 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18305) );
  NOR2_X1 U19056 ( .A1(n18305), .A2(n18952), .ZN(n15816) );
  INV_X1 U19057 ( .A(n18988), .ZN(n18985) );
  INV_X1 U19058 ( .A(n18956), .ZN(n18983) );
  AOI21_X1 U19059 ( .B1(n15818), .B2(n18783), .A(n15817), .ZN(n18836) );
  NAND3_X1 U19060 ( .A1(n18985), .A2(n18983), .A3(n18836), .ZN(n15819) );
  OAI21_X1 U19061 ( .B1(n18985), .B2(n18783), .A(n15819), .ZN(P3_U3284) );
  NOR2_X1 U19062 ( .A1(n10076), .A2(n18796), .ZN(n18190) );
  NOR2_X1 U19063 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18190), .ZN(
        n16521) );
  INV_X1 U19064 ( .A(n16521), .ZN(n15824) );
  INV_X1 U19065 ( .A(n18150), .ZN(n18218) );
  OAI21_X1 U19066 ( .B1(n15821), .B2(n18218), .A(n15820), .ZN(n15822) );
  AOI21_X1 U19067 ( .B1(n18277), .B2(n15823), .A(n15822), .ZN(n15880) );
  OAI221_X1 U19068 ( .B1(n18282), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C1(n18282), .C2(n15824), .A(n15880), .ZN(n15828) );
  NAND2_X1 U19069 ( .A1(n18150), .A2(n16524), .ZN(n15825) );
  OAI211_X1 U19070 ( .C1(n18302), .C2(n16522), .A(n15826), .B(n15825), .ZN(
        n15882) );
  AOI22_X1 U19071 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15828), .B1(
        n15882), .B2(n15827), .ZN(n15830) );
  OAI211_X1 U19072 ( .C1(n15831), .C2(n18223), .A(n15830), .B(n15829), .ZN(
        P3_U2833) );
  AOI22_X1 U19073 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19193), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19166), .ZN(n15843) );
  OAI22_X1 U19074 ( .A1(n15833), .A2(n19186), .B1(n19134), .B2(n15832), .ZN(
        n15834) );
  INV_X1 U19075 ( .A(n15834), .ZN(n15842) );
  AOI22_X1 U19076 ( .A1(n15836), .A2(n19188), .B1(n15835), .B2(n19168), .ZN(
        n15841) );
  OAI211_X1 U19077 ( .C1(n15839), .C2(n15838), .A(n19190), .B(n15837), .ZN(
        n15840) );
  NAND4_X1 U19078 ( .A1(n15843), .A2(n15842), .A3(n15841), .A4(n15840), .ZN(
        P2_U2833) );
  NOR3_X1 U19079 ( .A1(n15845), .A2(n15844), .A3(n20696), .ZN(n15850) );
  INV_X1 U19080 ( .A(n15850), .ZN(n15848) );
  OAI211_X1 U19081 ( .C1(n15848), .C2(n20655), .A(n15847), .B(n15846), .ZN(
        n15849) );
  OAI21_X1 U19082 ( .B1(n15850), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15849), .ZN(n15851) );
  AOI222_X1 U19083 ( .A1(n11143), .A2(n15852), .B1(n11143), .B2(n15851), .C1(
        n15852), .C2(n15851), .ZN(n15854) );
  AND2_X1 U19084 ( .A1(n15854), .A2(n15853), .ZN(n15855) );
  OAI22_X1 U19085 ( .A1(n15855), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n15854), .B2(n15853), .ZN(n15864) );
  INV_X1 U19086 ( .A(n15856), .ZN(n15863) );
  OAI21_X1 U19087 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15857), .ZN(n15858) );
  NAND4_X1 U19088 ( .A1(n15861), .A2(n15860), .A3(n15859), .A4(n15858), .ZN(
        n15862) );
  AOI211_X1 U19089 ( .C1(n15864), .C2(n11147), .A(n15863), .B(n15862), .ZN(
        n15865) );
  INV_X1 U19090 ( .A(n15865), .ZN(n15872) );
  AOI21_X1 U19091 ( .B1(n15871), .B2(n15872), .A(n15866), .ZN(n15877) );
  NOR2_X1 U19092 ( .A1(n20940), .A2(n15867), .ZN(n15870) );
  OR4_X1 U19093 ( .A1(n12641), .A2(n20274), .A3(n20933), .A4(n15868), .ZN(
        n15869) );
  OAI21_X1 U19094 ( .B1(n15871), .B2(n15870), .A(n15869), .ZN(n16192) );
  AOI221_X1 U19095 ( .B1(n20936), .B2(n20834), .C1(n15872), .C2(n20834), .A(
        n16192), .ZN(n15874) );
  AOI211_X1 U19096 ( .C1(n20846), .C2(n10577), .A(n15874), .B(n15873), .ZN(
        n16189) );
  INV_X1 U19097 ( .A(n15874), .ZN(n16197) );
  OAI21_X1 U19098 ( .B1(n15875), .B2(n20935), .A(n16197), .ZN(n15876) );
  AOI22_X1 U19099 ( .A1(n15877), .A2(n16189), .B1(n20936), .B2(n15876), .ZN(
        P1_U3161) );
  AOI21_X1 U19100 ( .B1(n15879), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15878), .ZN(n16511) );
  OAI21_X1 U19101 ( .B1(n16508), .B2(n18282), .A(n15880), .ZN(n15881) );
  AOI22_X1 U19102 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15881), .B1(
        n18296), .B2(P3_REIP_REG_30__SCAN_IN), .ZN(n15884) );
  NAND3_X1 U19103 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16507), .A3(
        n15882), .ZN(n15883) );
  OAI211_X1 U19104 ( .C1(n16511), .C2(n18223), .A(n15884), .B(n15883), .ZN(
        P3_U2832) );
  INV_X1 U19105 ( .A(HOLD), .ZN(n20842) );
  NAND2_X1 U19106 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20852), .ZN(n20845) );
  INV_X1 U19107 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20840) );
  NOR2_X1 U19108 ( .A1(n20837), .A2(n20840), .ZN(n15885) );
  AND2_X1 U19109 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20846), .ZN(n20843) );
  AOI221_X1 U19110 ( .B1(n20842), .B2(n15885), .C1(n20852), .C2(n15885), .A(
        n20843), .ZN(n15886) );
  OAI211_X1 U19111 ( .C1(n20842), .C2(n20845), .A(n15886), .B(n20933), .ZN(
        P1_U3195) );
  AND2_X1 U19112 ( .A1(n20195), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NAND2_X1 U19113 ( .A1(n16071), .A2(n15889), .ZN(n15892) );
  OAI21_X1 U19114 ( .B1(n16113), .B2(n15888), .A(n15887), .ZN(n16073) );
  OAI22_X1 U19115 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n20264), .B1(
        n15889), .B2(n15888), .ZN(n15890) );
  AOI211_X1 U19116 ( .C1(n15892), .C2(n15891), .A(n16073), .B(n15890), .ZN(
        n16063) );
  OAI21_X1 U19117 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15893), .A(
        n16063), .ZN(n15894) );
  AOI22_X1 U19118 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15894), .B1(
        n16174), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15900) );
  INV_X1 U19119 ( .A(n15895), .ZN(n15898) );
  INV_X1 U19120 ( .A(n15896), .ZN(n15897) );
  AOI22_X1 U19121 ( .A1(n15898), .A2(n20260), .B1(n16173), .B2(n15897), .ZN(
        n15899) );
  OAI211_X1 U19122 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15901), .A(
        n15900), .B(n15899), .ZN(P1_U3011) );
  NOR3_X1 U19123 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20054), .A3(n20057), 
        .ZN(n16487) );
  OAI22_X1 U19124 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n15902), .B1(
        P2_STATE2_REG_2__SCAN_IN), .B2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15903)
         );
  NOR3_X1 U19125 ( .A1(n16487), .A2(n15905), .A3(n15903), .ZN(P2_U3178) );
  INV_X1 U19126 ( .A(n20044), .ZN(n15904) );
  AOI221_X1 U19127 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15905), .C1(n15904), .C2(
        n15905), .A(n19836), .ZN(n20034) );
  INV_X1 U19128 ( .A(n20034), .ZN(n20035) );
  NOR2_X1 U19129 ( .A1(n15906), .A2(n20035), .ZN(P2_U3047) );
  NAND2_X1 U19130 ( .A1(n18350), .A2(n15911), .ZN(n17486) );
  INV_X1 U19131 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17574) );
  AOI22_X1 U19132 ( .A1(n17498), .A2(BUF2_REG_0__SCAN_IN), .B1(n17497), .B2(
        n17978), .ZN(n15910) );
  OAI221_X1 U19133 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17486), .C1(n17574), 
        .C2(n15911), .A(n15910), .ZN(P3_U2735) );
  INV_X1 U19134 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21042) );
  NOR2_X1 U19135 ( .A1(n21042), .A2(n21122), .ZN(n15932) );
  AOI21_X1 U19136 ( .B1(n15921), .B2(n15932), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n15920) );
  OAI22_X1 U19137 ( .A1(n20107), .A2(n14513), .B1(n15912), .B2(n20098), .ZN(
        n15913) );
  AOI211_X1 U19138 ( .C1(n20127), .C2(n15914), .A(n20138), .B(n15913), .ZN(
        n15918) );
  OAI22_X1 U19139 ( .A1(n15915), .A2(n20099), .B1(n20155), .B2(n16087), .ZN(
        n15916) );
  INV_X1 U19140 ( .A(n15916), .ZN(n15917) );
  OAI211_X1 U19141 ( .C1(n15920), .C2(n15919), .A(n15918), .B(n15917), .ZN(
        P1_U2823) );
  OAI21_X1 U19142 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15921), .ZN(n15931) );
  XNOR2_X1 U19143 ( .A(n15923), .B(n15922), .ZN(n16095) );
  AOI22_X1 U19144 ( .A1(n15936), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n20130), 
        .B2(n16095), .ZN(n15930) );
  INV_X1 U19145 ( .A(n14506), .ZN(n15924) );
  AOI21_X1 U19146 ( .B1(n15925), .B2(n14490), .A(n15924), .ZN(n15988) );
  AOI21_X1 U19147 ( .B1(n20139), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20138), .ZN(n15927) );
  NAND2_X1 U19148 ( .A1(n20152), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n15926) );
  OAI211_X1 U19149 ( .C1(n20142), .C2(n15991), .A(n15927), .B(n15926), .ZN(
        n15928) );
  AOI21_X1 U19150 ( .B1(n15988), .B2(n20123), .A(n15928), .ZN(n15929) );
  OAI211_X1 U19151 ( .C1(n15932), .C2(n15931), .A(n15930), .B(n15929), .ZN(
        P1_U2824) );
  INV_X1 U19152 ( .A(n15996), .ZN(n15933) );
  OAI22_X1 U19153 ( .A1(n16116), .A2(n20155), .B1(n20142), .B2(n15933), .ZN(
        n15934) );
  INV_X1 U19154 ( .A(n15934), .ZN(n15939) );
  AOI22_X1 U19155 ( .A1(n20152), .A2(P1_EBX_REG_14__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n20139), .ZN(n15938) );
  INV_X1 U19156 ( .A(n15967), .ZN(n15949) );
  NAND3_X1 U19157 ( .A1(n15949), .A2(P1_REIP_REG_12__SCAN_IN), .A3(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15943) );
  INV_X1 U19158 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21300) );
  OAI21_X1 U19159 ( .B1(n14773), .B2(n15943), .A(n21300), .ZN(n15935) );
  AOI22_X1 U19160 ( .A1(n15997), .A2(n20123), .B1(n15936), .B2(n15935), .ZN(
        n15937) );
  NAND4_X1 U19161 ( .A1(n15939), .A2(n15938), .A3(n15937), .A4(n20134), .ZN(
        P1_U2826) );
  NAND2_X1 U19162 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15940) );
  AOI21_X1 U19163 ( .B1(n15941), .B2(n15940), .A(n15964), .ZN(n15957) );
  AOI22_X1 U19164 ( .A1(n16117), .A2(n20130), .B1(n20152), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15942) );
  OAI211_X1 U19165 ( .C1(n20098), .C2(n14774), .A(n15942), .B(n20134), .ZN(
        n15946) );
  OAI22_X1 U19166 ( .A1(n15944), .A2(n20099), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n15943), .ZN(n15945) );
  AOI211_X1 U19167 ( .C1(n15947), .C2(n20127), .A(n15946), .B(n15945), .ZN(
        n15948) );
  OAI21_X1 U19168 ( .B1(n15957), .B2(n14773), .A(n15948), .ZN(P1_U2827) );
  AOI21_X1 U19169 ( .B1(n15949), .B2(P1_REIP_REG_11__SCAN_IN), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15956) );
  AOI22_X1 U19170 ( .A1(n15969), .A2(n20130), .B1(n20127), .B2(n16000), .ZN(
        n15955) );
  INV_X1 U19171 ( .A(n15950), .ZN(n16002) );
  NOR2_X1 U19172 ( .A1(n20107), .A2(n15971), .ZN(n15953) );
  OAI21_X1 U19173 ( .B1(n20098), .B2(n15951), .A(n20134), .ZN(n15952) );
  AOI211_X1 U19174 ( .C1(n16002), .C2(n20123), .A(n15953), .B(n15952), .ZN(
        n15954) );
  OAI211_X1 U19175 ( .C1(n15957), .C2(n15956), .A(n15955), .B(n15954), .ZN(
        P1_U2828) );
  OAI21_X1 U19176 ( .B1(n15960), .B2(n15959), .A(n15958), .ZN(n15961) );
  INV_X1 U19177 ( .A(n15961), .ZN(n16129) );
  AOI22_X1 U19178 ( .A1(n16129), .A2(n20130), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n20152), .ZN(n15962) );
  OAI21_X1 U19179 ( .B1(n16014), .B2(n20142), .A(n15962), .ZN(n15963) );
  AOI211_X1 U19180 ( .C1(n20139), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20138), .B(n15963), .ZN(n15966) );
  AOI22_X1 U19181 ( .A1(n16011), .A2(n20123), .B1(n15964), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15965) );
  OAI211_X1 U19182 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15967), .A(n15966), 
        .B(n15965), .ZN(P1_U2829) );
  INV_X1 U19183 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21170) );
  AOI22_X1 U19184 ( .A1(n15988), .A2(n20176), .B1(n20175), .B2(n16095), .ZN(
        n15968) );
  OAI21_X1 U19185 ( .B1(n20179), .B2(n21170), .A(n15968), .ZN(P1_U2856) );
  AOI22_X1 U19186 ( .A1(n16002), .A2(n20176), .B1(n20175), .B2(n15969), .ZN(
        n15970) );
  OAI21_X1 U19187 ( .B1(n20179), .B2(n15971), .A(n15970), .ZN(P1_U2860) );
  INV_X1 U19188 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15973) );
  AOI22_X1 U19189 ( .A1(n16011), .A2(n20176), .B1(n20175), .B2(n16129), .ZN(
        n15972) );
  OAI21_X1 U19190 ( .B1(n20179), .B2(n15973), .A(n15972), .ZN(P1_U2861) );
  INV_X1 U19191 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20268) );
  INV_X1 U19192 ( .A(n20267), .ZN(n15975) );
  AOI22_X1 U19193 ( .A1(n15976), .A2(n15975), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15974), .ZN(n15980) );
  AOI22_X1 U19194 ( .A1(n15988), .A2(n15978), .B1(n15977), .B2(DATAI_16_), 
        .ZN(n15979) );
  OAI211_X1 U19195 ( .C1(n15981), .C2(n20268), .A(n15980), .B(n15979), .ZN(
        P1_U2888) );
  AOI22_X1 U19196 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15990) );
  INV_X1 U19197 ( .A(n9820), .ZN(n15985) );
  AOI21_X1 U19198 ( .B1(n15985), .B2(n15984), .A(n15983), .ZN(n15987) );
  NOR2_X1 U19199 ( .A1(n15987), .A2(n15986), .ZN(n16096) );
  AOI22_X1 U19200 ( .A1(n16096), .A2(n11296), .B1(n15988), .B2(n16025), .ZN(
        n15989) );
  OAI211_X1 U19201 ( .C1(n16022), .C2(n15991), .A(n15990), .B(n15989), .ZN(
        P1_U2983) );
  NAND2_X1 U19202 ( .A1(n9821), .A2(n15992), .ZN(n15995) );
  XNOR2_X1 U19203 ( .A(n14729), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15994) );
  XNOR2_X1 U19204 ( .A(n15995), .B(n15994), .ZN(n16110) );
  AOI22_X1 U19205 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15999) );
  AOI22_X1 U19206 ( .A1(n15997), .A2(n16025), .B1(n16024), .B2(n15996), .ZN(
        n15998) );
  OAI211_X1 U19207 ( .C1(n16110), .C2(n20080), .A(n15999), .B(n15998), .ZN(
        P1_U2985) );
  AOI22_X1 U19208 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16004) );
  AOI22_X1 U19209 ( .A1(n16002), .A2(n16001), .B1(n16024), .B2(n16000), .ZN(
        n16003) );
  OAI211_X1 U19210 ( .C1(n16005), .C2(n20080), .A(n16004), .B(n16003), .ZN(
        P1_U2987) );
  AOI22_X1 U19211 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16013) );
  NAND3_X1 U19212 ( .A1(n16006), .A2(n14729), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16008) );
  NAND2_X1 U19213 ( .A1(n16008), .A2(n16007), .ZN(n16010) );
  XNOR2_X1 U19214 ( .A(n16010), .B(n16009), .ZN(n16131) );
  AOI22_X1 U19215 ( .A1(n16025), .A2(n16011), .B1(n16131), .B2(n11296), .ZN(
        n16012) );
  OAI211_X1 U19216 ( .C1(n16022), .C2(n16014), .A(n16013), .B(n16012), .ZN(
        P1_U2988) );
  AOI22_X1 U19217 ( .A1(n16015), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16174), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16021) );
  NAND2_X1 U19218 ( .A1(n16018), .A2(n16017), .ZN(n16019) );
  XNOR2_X1 U19219 ( .A(n16016), .B(n16019), .ZN(n16176) );
  AOI22_X1 U19220 ( .A1(n16176), .A2(n11296), .B1(n16025), .B2(n20166), .ZN(
        n16020) );
  OAI211_X1 U19221 ( .C1(n16022), .C2(n20110), .A(n16021), .B(n16020), .ZN(
        P1_U2992) );
  INV_X1 U19222 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16030) );
  INV_X1 U19223 ( .A(n16023), .ZN(n20128) );
  AOI222_X1 U19224 ( .A1(n16026), .A2(n11296), .B1(n16025), .B2(n20171), .C1(
        n20128), .C2(n16024), .ZN(n16028) );
  OAI211_X1 U19225 ( .C1(n16030), .C2(n16029), .A(n16028), .B(n16027), .ZN(
        P1_U2994) );
  INV_X1 U19226 ( .A(n16031), .ZN(n16032) );
  NOR2_X1 U19227 ( .A1(n16032), .A2(n16036), .ZN(n16033) );
  AOI211_X1 U19228 ( .C1(n16035), .C2(n20260), .A(n16034), .B(n16033), .ZN(
        n16039) );
  NAND3_X1 U19229 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n16037), .A3(
        n16036), .ZN(n16038) );
  OAI211_X1 U19230 ( .C1(n16040), .C2(n20258), .A(n16039), .B(n16038), .ZN(
        P1_U3005) );
  AOI22_X1 U19231 ( .A1(n16174), .A2(P1_REIP_REG_23__SCAN_IN), .B1(n16041), 
        .B2(n16065), .ZN(n16047) );
  OAI22_X1 U19232 ( .A1(n16044), .A2(n16182), .B1(n16043), .B2(n16042), .ZN(
        n16045) );
  INV_X1 U19233 ( .A(n16045), .ZN(n16046) );
  OAI211_X1 U19234 ( .C1(n20258), .C2(n16048), .A(n16047), .B(n16046), .ZN(
        P1_U3008) );
  INV_X1 U19235 ( .A(n16049), .ZN(n16050) );
  AOI22_X1 U19236 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16050), .B1(
        n16174), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16058) );
  INV_X1 U19237 ( .A(n16051), .ZN(n16056) );
  AOI21_X1 U19238 ( .B1(n14884), .B2(n16053), .A(n16052), .ZN(n16054) );
  AOI22_X1 U19239 ( .A1(n16056), .A2(n20260), .B1(n16055), .B2(n16054), .ZN(
        n16057) );
  OAI211_X1 U19240 ( .C1(n20258), .C2(n16059), .A(n16058), .B(n16057), .ZN(
        P1_U3009) );
  INV_X1 U19241 ( .A(n16060), .ZN(n16062) );
  AOI22_X1 U19242 ( .A1(n16062), .A2(n20260), .B1(n16173), .B2(n16061), .ZN(
        n16068) );
  INV_X1 U19243 ( .A(n16063), .ZN(n16066) );
  NOR2_X1 U19244 ( .A1(n16162), .A2(n21041), .ZN(n16064) );
  AOI221_X1 U19245 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16066), 
        .C1(n11291), .C2(n16065), .A(n16064), .ZN(n16067) );
  NAND2_X1 U19246 ( .A1(n16068), .A2(n16067), .ZN(P1_U3012) );
  INV_X1 U19247 ( .A(n20264), .ZN(n16069) );
  OAI21_X1 U19248 ( .B1(n16121), .B2(n16128), .A(n16069), .ZN(n16127) );
  OAI21_X1 U19249 ( .B1(n16071), .B2(n16070), .A(n16127), .ZN(n16072) );
  AOI211_X1 U19250 ( .C1(n16121), .C2(n16119), .A(n16073), .B(n16072), .ZN(
        n16120) );
  OAI21_X1 U19251 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16074), .A(
        n16120), .ZN(n16104) );
  AOI21_X1 U19252 ( .B1(n16160), .B2(n16078), .A(n16104), .ZN(n16093) );
  INV_X1 U19253 ( .A(n16075), .ZN(n16076) );
  AOI211_X1 U19254 ( .C1(n16077), .C2(n16076), .A(n16109), .B(n16121), .ZN(
        n16094) );
  INV_X1 U19255 ( .A(n16094), .ZN(n16108) );
  NOR3_X1 U19256 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16078), .A3(
        n16108), .ZN(n16082) );
  OAI22_X1 U19257 ( .A1(n16080), .A2(n16182), .B1(n20258), .B2(n16079), .ZN(
        n16081) );
  NOR3_X1 U19258 ( .A1(n16083), .A2(n16082), .A3(n16081), .ZN(n16084) );
  OAI21_X1 U19259 ( .B1(n16093), .B2(n16085), .A(n16084), .ZN(P1_U3013) );
  AND2_X1 U19260 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16100) );
  AOI21_X1 U19261 ( .B1(n16100), .B2(n16094), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16092) );
  INV_X1 U19262 ( .A(n16086), .ZN(n16089) );
  INV_X1 U19263 ( .A(n16087), .ZN(n16088) );
  NAND2_X1 U19264 ( .A1(n16174), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16090) );
  OAI211_X1 U19265 ( .C1(n16093), .C2(n16092), .A(n16091), .B(n16090), .ZN(
        P1_U3014) );
  OAI21_X1 U19266 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16094), .ZN(n16099) );
  AOI22_X1 U19267 ( .A1(n16174), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n16173), 
        .B2(n16095), .ZN(n16098) );
  AOI22_X1 U19268 ( .A1(n16096), .A2(n20260), .B1(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16104), .ZN(n16097) );
  OAI211_X1 U19269 ( .C1(n16100), .C2(n16099), .A(n16098), .B(n16097), .ZN(
        P1_U3015) );
  INV_X1 U19270 ( .A(n16101), .ZN(n16102) );
  AOI22_X1 U19271 ( .A1(n16174), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n16173), 
        .B2(n16102), .ZN(n16107) );
  INV_X1 U19272 ( .A(n16103), .ZN(n16105) );
  AOI22_X1 U19273 ( .A1(n16105), .A2(n20260), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16104), .ZN(n16106) );
  OAI211_X1 U19274 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16108), .A(
        n16107), .B(n16106), .ZN(P1_U3016) );
  NOR3_X1 U19275 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16141), .A3(
        n16121), .ZN(n16112) );
  OAI22_X1 U19276 ( .A1(n16110), .A2(n16182), .B1(n16120), .B2(n16109), .ZN(
        n16111) );
  AOI21_X1 U19277 ( .B1(n16113), .B2(n16112), .A(n16111), .ZN(n16115) );
  NAND2_X1 U19278 ( .A1(n16174), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16114) );
  OAI211_X1 U19279 ( .C1(n20258), .C2(n16116), .A(n16115), .B(n16114), .ZN(
        P1_U3017) );
  AOI22_X1 U19280 ( .A1(n16174), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n16173), 
        .B2(n16117), .ZN(n16126) );
  INV_X1 U19281 ( .A(n16118), .ZN(n16124) );
  INV_X1 U19282 ( .A(n16119), .ZN(n16122) );
  AOI21_X1 U19283 ( .B1(n16122), .B2(n16121), .A(n16120), .ZN(n16123) );
  AOI21_X1 U19284 ( .B1(n16124), .B2(n20260), .A(n16123), .ZN(n16125) );
  OAI211_X1 U19285 ( .C1(n16128), .C2(n16127), .A(n16126), .B(n16125), .ZN(
        P1_U3018) );
  AOI22_X1 U19286 ( .A1(n16174), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n16173), 
        .B2(n16129), .ZN(n16133) );
  AOI22_X1 U19287 ( .A1(n16131), .A2(n20260), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16130), .ZN(n16132) );
  OAI211_X1 U19288 ( .C1(n16181), .C2(n16134), .A(n16133), .B(n16132), .ZN(
        P1_U3020) );
  NAND2_X1 U19289 ( .A1(n16136), .A2(n16135), .ZN(n16140) );
  AOI21_X1 U19290 ( .B1(n16160), .B2(n16140), .A(n16137), .ZN(n16153) );
  AOI222_X1 U19291 ( .A1(n16139), .A2(n20260), .B1(n16173), .B2(n16138), .C1(
        P1_REIP_REG_10__SCAN_IN), .C2(n16174), .ZN(n16143) );
  NOR2_X1 U19292 ( .A1(n16141), .A2(n16140), .ZN(n16148) );
  OAI221_X1 U19293 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14781), .C2(n16152), .A(
        n16148), .ZN(n16142) );
  OAI211_X1 U19294 ( .C1(n16153), .C2(n14781), .A(n16143), .B(n16142), .ZN(
        P1_U3021) );
  NAND2_X1 U19295 ( .A1(n16145), .A2(n16144), .ZN(n16146) );
  AND2_X1 U19296 ( .A1(n16147), .A2(n16146), .ZN(n20161) );
  AOI22_X1 U19297 ( .A1(n16174), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n16173), 
        .B2(n20161), .ZN(n16151) );
  AOI22_X1 U19298 ( .A1(n16149), .A2(n20260), .B1(n16148), .B2(n16152), .ZN(
        n16150) );
  OAI211_X1 U19299 ( .C1(n16153), .C2(n16152), .A(n16151), .B(n16150), .ZN(
        P1_U3022) );
  NAND2_X1 U19300 ( .A1(n16155), .A2(n16154), .ZN(n16156) );
  OAI211_X1 U19301 ( .C1(n16159), .C2(n16158), .A(n16157), .B(n16156), .ZN(
        n16185) );
  AOI21_X1 U19302 ( .B1(n16165), .B2(n16160), .A(n16185), .ZN(n16180) );
  OAI222_X1 U19303 ( .A1(n16163), .A2(n20258), .B1(n16162), .B2(n20860), .C1(
        n16182), .C2(n16161), .ZN(n16164) );
  INV_X1 U19304 ( .A(n16164), .ZN(n16167) );
  NOR2_X1 U19305 ( .A1(n16165), .A2(n16181), .ZN(n16175) );
  OAI221_X1 U19306 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16168), .C2(n16179), .A(
        n16175), .ZN(n16166) );
  OAI211_X1 U19307 ( .C1(n16180), .C2(n16168), .A(n16167), .B(n16166), .ZN(
        P1_U3023) );
  NOR2_X1 U19308 ( .A1(n16170), .A2(n16169), .ZN(n16171) );
  AOI22_X1 U19309 ( .A1(n16174), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n16173), 
        .B2(n9917), .ZN(n16178) );
  AOI22_X1 U19310 ( .A1(n16176), .A2(n20260), .B1(n16175), .B2(n16179), .ZN(
        n16177) );
  OAI211_X1 U19311 ( .C1(n16180), .C2(n16179), .A(n16178), .B(n16177), .ZN(
        P1_U3024) );
  OAI22_X1 U19312 ( .A1(n16183), .A2(n16182), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16181), .ZN(n16184) );
  AOI21_X1 U19313 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16185), .A(
        n16184), .ZN(n16188) );
  INV_X1 U19314 ( .A(n16186), .ZN(n16187) );
  OAI211_X1 U19315 ( .C1(n20258), .C2(n20119), .A(n16188), .B(n16187), .ZN(
        P1_U3025) );
  INV_X1 U19316 ( .A(n16189), .ZN(n16193) );
  OAI221_X1 U19317 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20936), .C2(n20940), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20835) );
  NAND2_X1 U19318 ( .A1(n20835), .A2(n16190), .ZN(n16191) );
  AOI22_X1 U19319 ( .A1(n20834), .A2(n16193), .B1(n16192), .B2(n16191), .ZN(
        P1_U3162) );
  INV_X1 U19320 ( .A(n16194), .ZN(n16196) );
  OAI211_X1 U19321 ( .C1(n20661), .C2(n16197), .A(n16196), .B(n16195), .ZN(
        P1_U3466) );
  NAND2_X1 U19322 ( .A1(n9807), .A2(n16198), .ZN(n16213) );
  NAND2_X1 U19323 ( .A1(n16214), .A2(n16213), .ZN(n16212) );
  AND2_X1 U19324 ( .A1(n16199), .A2(n19102), .ZN(n16203) );
  INV_X1 U19325 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19974) );
  OAI22_X1 U19326 ( .A1(n16201), .A2(n16200), .B1(n19974), .B2(n19181), .ZN(
        n16202) );
  AOI211_X1 U19327 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n19193), .A(
        n16203), .B(n16202), .ZN(n16207) );
  INV_X1 U19328 ( .A(n16204), .ZN(n19199) );
  AOI22_X1 U19329 ( .A1(n16205), .A2(n19188), .B1(n19168), .B2(n19199), .ZN(
        n16206) );
  OAI211_X1 U19330 ( .C1(n16208), .C2(n16212), .A(n16207), .B(n16206), .ZN(
        P2_U2824) );
  AOI22_X1 U19331 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19193), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19166), .ZN(n16218) );
  AOI22_X1 U19332 ( .A1(n16209), .A2(n19102), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n19183), .ZN(n16217) );
  AOI22_X1 U19333 ( .A1(n16211), .A2(n19188), .B1(n19168), .B2(n16210), .ZN(
        n16216) );
  OAI211_X1 U19334 ( .C1(n16214), .C2(n16213), .A(n19190), .B(n16212), .ZN(
        n16215) );
  NAND4_X1 U19335 ( .A1(n16218), .A2(n16217), .A3(n16216), .A4(n16215), .ZN(
        P2_U2825) );
  AOI22_X1 U19336 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19193), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19166), .ZN(n16230) );
  INV_X1 U19337 ( .A(n16219), .ZN(n16220) );
  AOI22_X1 U19338 ( .A1(n16220), .A2(n19102), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n19183), .ZN(n16229) );
  OAI22_X1 U19339 ( .A1(n16222), .A2(n19157), .B1(n16221), .B2(n19179), .ZN(
        n16223) );
  INV_X1 U19340 ( .A(n16223), .ZN(n16228) );
  OAI211_X1 U19341 ( .C1(n16226), .C2(n16225), .A(n19190), .B(n16224), .ZN(
        n16227) );
  NAND4_X1 U19342 ( .A1(n16230), .A2(n16229), .A3(n16228), .A4(n16227), .ZN(
        P2_U2827) );
  INV_X1 U19343 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16231) );
  INV_X1 U19344 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19962) );
  OAI22_X1 U19345 ( .A1(n16231), .A2(n19163), .B1(n19962), .B2(n19181), .ZN(
        n16232) );
  AOI21_X1 U19346 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n19183), .A(n16232), .ZN(
        n16233) );
  OAI21_X1 U19347 ( .B1(n16234), .B2(n19157), .A(n16233), .ZN(n16235) );
  AOI21_X1 U19348 ( .B1(n16236), .B2(n19102), .A(n16235), .ZN(n16241) );
  OAI211_X1 U19349 ( .C1(n16239), .C2(n16238), .A(n19190), .B(n16237), .ZN(
        n16240) );
  OAI211_X1 U19350 ( .C1(n19179), .C2(n16242), .A(n16241), .B(n16240), .ZN(
        P2_U2829) );
  INV_X1 U19351 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16243) );
  INV_X1 U19352 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19958) );
  OAI22_X1 U19353 ( .A1(n16243), .A2(n19163), .B1(n19958), .B2(n19181), .ZN(
        n16244) );
  AOI21_X1 U19354 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n19183), .A(n16244), .ZN(
        n16245) );
  OAI21_X1 U19355 ( .B1(n16246), .B2(n19157), .A(n16245), .ZN(n16247) );
  AOI21_X1 U19356 ( .B1(n16248), .B2(n19102), .A(n16247), .ZN(n16253) );
  OAI211_X1 U19357 ( .C1(n16251), .C2(n16250), .A(n19190), .B(n16249), .ZN(
        n16252) );
  OAI211_X1 U19358 ( .C1(n19179), .C2(n16254), .A(n16253), .B(n16252), .ZN(
        P2_U2831) );
  AOI22_X1 U19359 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19193), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19166), .ZN(n16264) );
  AOI22_X1 U19360 ( .A1(n16255), .A2(n19102), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n19183), .ZN(n16263) );
  INV_X1 U19361 ( .A(n16256), .ZN(n16267) );
  AOI22_X1 U19362 ( .A1(n16257), .A2(n19188), .B1(n16267), .B2(n19168), .ZN(
        n16262) );
  OAI211_X1 U19363 ( .C1(n16260), .C2(n16259), .A(n19190), .B(n16258), .ZN(
        n16261) );
  NAND4_X1 U19364 ( .A1(n16264), .A2(n16263), .A3(n16262), .A4(n16261), .ZN(
        P2_U2832) );
  AOI22_X1 U19365 ( .A1(n16266), .A2(n16265), .B1(n19203), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16272) );
  AOI22_X1 U19366 ( .A1(n19200), .A2(BUF1_REG_23__SCAN_IN), .B1(n19197), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n16271) );
  AOI22_X1 U19367 ( .A1(n16269), .A2(n16268), .B1(n19198), .B2(n16267), .ZN(
        n16270) );
  NAND3_X1 U19368 ( .A1(n16272), .A2(n16271), .A3(n16270), .ZN(P2_U2896) );
  AOI22_X1 U19369 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19271), .B1(n19270), 
        .B2(n16273), .ZN(n16280) );
  NOR3_X1 U19370 ( .A1(n16275), .A2(n16274), .A3(n19277), .ZN(n16278) );
  NOR2_X1 U19371 ( .A1(n16276), .A2(n19278), .ZN(n16277) );
  OAI211_X1 U19372 ( .C1(n16281), .C2(n19285), .A(n16280), .B(n16279), .ZN(
        P2_U2999) );
  AOI22_X1 U19373 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16355), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19271), .ZN(n16286) );
  OAI22_X1 U19374 ( .A1(n16283), .A2(n19278), .B1(n19277), .B2(n16282), .ZN(
        n16284) );
  AOI21_X1 U19375 ( .B1(n19282), .B2(n19117), .A(n16284), .ZN(n16285) );
  OAI211_X1 U19376 ( .C1(n16366), .C2(n16287), .A(n16286), .B(n16285), .ZN(
        P2_U3000) );
  AOI22_X1 U19377 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19271), .B1(n19270), 
        .B2(n16288), .ZN(n16299) );
  AND2_X1 U19378 ( .A1(n16290), .A2(n16289), .ZN(n16291) );
  XNOR2_X1 U19379 ( .A(n16292), .B(n16291), .ZN(n16372) );
  NAND2_X1 U19380 ( .A1(n16372), .A2(n16361), .ZN(n16296) );
  OAI21_X1 U19381 ( .B1(n16316), .B2(n16368), .A(n16367), .ZN(n16294) );
  AND2_X1 U19382 ( .A1(n16294), .A2(n16293), .ZN(n16373) );
  NAND2_X1 U19383 ( .A1(n16373), .A2(n16350), .ZN(n16295) );
  OAI211_X1 U19384 ( .C1(n19317), .C2(n16376), .A(n16296), .B(n16295), .ZN(
        n16297) );
  INV_X1 U19385 ( .A(n16297), .ZN(n16298) );
  OAI211_X1 U19386 ( .C1(n16300), .C2(n19285), .A(n16299), .B(n16298), .ZN(
        P2_U3001) );
  AOI22_X1 U19387 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16355), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19287), .ZN(n16306) );
  INV_X1 U19388 ( .A(n16301), .ZN(n19128) );
  OAI22_X1 U19389 ( .A1(n16303), .A2(n19277), .B1(n16302), .B2(n19278), .ZN(
        n16304) );
  AOI21_X1 U19390 ( .B1(n19282), .B2(n19128), .A(n16304), .ZN(n16305) );
  OAI211_X1 U19391 ( .C1(n16366), .C2(n16307), .A(n16306), .B(n16305), .ZN(
        P2_U3002) );
  AOI22_X1 U19392 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19271), .B1(n19270), 
        .B2(n16308), .ZN(n16321) );
  NAND3_X1 U19393 ( .A1(n16310), .A2(n16309), .A3(n16326), .ZN(n16315) );
  INV_X1 U19394 ( .A(n16311), .ZN(n16312) );
  NOR2_X1 U19395 ( .A1(n16313), .A2(n16312), .ZN(n16314) );
  XNOR2_X1 U19396 ( .A(n16315), .B(n16314), .ZN(n16392) );
  INV_X1 U19397 ( .A(n16392), .ZN(n16319) );
  AOI21_X1 U19398 ( .B1(n16336), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16318) );
  INV_X1 U19399 ( .A(n16316), .ZN(n16317) );
  NOR2_X1 U19400 ( .A1(n16318), .A2(n16317), .ZN(n16389) );
  AOI222_X1 U19401 ( .A1(n16319), .A2(n16361), .B1(n19282), .B2(n16388), .C1(
        n16350), .C2(n16389), .ZN(n16320) );
  OAI211_X1 U19402 ( .C1(n16322), .C2(n19285), .A(n16321), .B(n16320), .ZN(
        P2_U3003) );
  AOI22_X1 U19403 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16355), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19271), .ZN(n16333) );
  XNOR2_X1 U19404 ( .A(n16323), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16403) );
  INV_X1 U19405 ( .A(n16403), .ZN(n16330) );
  NOR2_X1 U19406 ( .A1(n16325), .A2(n16324), .ZN(n16329) );
  NAND2_X1 U19407 ( .A1(n16327), .A2(n16326), .ZN(n16328) );
  XNOR2_X1 U19408 ( .A(n16329), .B(n16328), .ZN(n16405) );
  OAI22_X1 U19409 ( .A1(n16330), .A2(n19277), .B1(n16405), .B2(n19278), .ZN(
        n16331) );
  AOI21_X1 U19410 ( .B1(n19282), .B2(n16398), .A(n16331), .ZN(n16332) );
  OAI211_X1 U19411 ( .C1(n16366), .C2(n16334), .A(n16333), .B(n16332), .ZN(
        P2_U3004) );
  AOI22_X1 U19412 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19287), .B1(n19270), 
        .B2(n16335), .ZN(n16343) );
  NOR3_X1 U19413 ( .A1(n16337), .A2(n16336), .A3(n19277), .ZN(n16341) );
  OAI22_X1 U19414 ( .A1(n16339), .A2(n19278), .B1(n19317), .B2(n16338), .ZN(
        n16340) );
  NOR2_X1 U19415 ( .A1(n16341), .A2(n16340), .ZN(n16342) );
  OAI211_X1 U19416 ( .C1(n16344), .C2(n19285), .A(n16343), .B(n16342), .ZN(
        P2_U3005) );
  OAI22_X1 U19417 ( .A1(n16346), .A2(n19285), .B1(n16366), .B2(n16345), .ZN(
        n16347) );
  AOI21_X1 U19418 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n19287), .A(n16347), .ZN(
        n16353) );
  INV_X1 U19419 ( .A(n16348), .ZN(n16351) );
  AOI22_X1 U19420 ( .A1(n16351), .A2(n16350), .B1(n16361), .B2(n16349), .ZN(
        n16352) );
  OAI211_X1 U19421 ( .C1(n19317), .C2(n16354), .A(n16353), .B(n16352), .ZN(
        P2_U3007) );
  AOI22_X1 U19422 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16355), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n19287), .ZN(n16364) );
  NOR2_X1 U19423 ( .A1(n19317), .A2(n16356), .ZN(n16360) );
  NOR3_X1 U19424 ( .A1(n16358), .A2(n16357), .A3(n19277), .ZN(n16359) );
  AOI211_X1 U19425 ( .C1(n16362), .C2(n16361), .A(n16360), .B(n16359), .ZN(
        n16363) );
  OAI211_X1 U19426 ( .C1(n16366), .C2(n16365), .A(n16364), .B(n16363), .ZN(
        P2_U3009) );
  INV_X1 U19427 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19936) );
  OAI21_X1 U19428 ( .B1(n16369), .B2(n16368), .A(n16367), .ZN(n16370) );
  AOI22_X1 U19429 ( .A1(n16371), .A2(n16370), .B1(n16387), .B2(n19207), .ZN(
        n16379) );
  NAND2_X1 U19430 ( .A1(n16372), .A2(n19296), .ZN(n16375) );
  NAND2_X1 U19431 ( .A1(n16373), .A2(n16413), .ZN(n16374) );
  OAI211_X1 U19432 ( .C1(n16376), .C2(n19308), .A(n16375), .B(n16374), .ZN(
        n16377) );
  INV_X1 U19433 ( .A(n16377), .ZN(n16378) );
  OAI211_X1 U19434 ( .C1(n19936), .C2(n19150), .A(n16379), .B(n16378), .ZN(
        P2_U3033) );
  OAI211_X1 U19435 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n16393), .ZN(n16381) );
  OAI22_X1 U19436 ( .A1(n10048), .A2(n16381), .B1(n19932), .B2(n19150), .ZN(
        n16386) );
  NAND2_X1 U19437 ( .A1(n16383), .A2(n16382), .ZN(n16395) );
  NOR2_X1 U19438 ( .A1(n16395), .A2(n16384), .ZN(n16385) );
  AOI211_X1 U19439 ( .C1(n19210), .C2(n16387), .A(n16386), .B(n16385), .ZN(
        n16391) );
  AOI22_X1 U19440 ( .A1(n16389), .A2(n16413), .B1(n16412), .B2(n16388), .ZN(
        n16390) );
  OAI211_X1 U19441 ( .C1(n16392), .C2(n19314), .A(n16391), .B(n16390), .ZN(
        P2_U3035) );
  NAND2_X1 U19442 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16393), .ZN(
        n16397) );
  NAND2_X1 U19443 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19287), .ZN(n16394) );
  OAI221_X1 U19444 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16397), 
        .C1(n16396), .C2(n16395), .A(n16394), .ZN(n16402) );
  INV_X1 U19445 ( .A(n16398), .ZN(n16400) );
  OAI22_X1 U19446 ( .A1(n19308), .A2(n16400), .B1(n16399), .B2(n19301), .ZN(
        n16401) );
  AOI211_X1 U19447 ( .C1(n16403), .C2(n16413), .A(n16402), .B(n16401), .ZN(
        n16404) );
  OAI21_X1 U19448 ( .B1(n16405), .B2(n19314), .A(n16404), .ZN(P2_U3036) );
  NOR2_X1 U19449 ( .A1(n19927), .A2(n19150), .ZN(n16410) );
  OAI21_X1 U19450 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16406), .ZN(n16407) );
  OAI22_X1 U19451 ( .A1(n16408), .A2(n16407), .B1(n19301), .B2(n19146), .ZN(
        n16409) );
  AOI211_X1 U19452 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n16411), .A(
        n16410), .B(n16409), .ZN(n16416) );
  AOI22_X1 U19453 ( .A1(n16414), .A2(n16413), .B1(n16412), .B2(n19142), .ZN(
        n16415) );
  OAI211_X1 U19454 ( .C1(n16417), .C2(n19314), .A(n16416), .B(n16415), .ZN(
        P2_U3038) );
  OAI22_X1 U19455 ( .A1(n19308), .A2(n16418), .B1(n19301), .B2(n19178), .ZN(
        n16420) );
  MUX2_X1 U19456 ( .A(n19305), .B(n19311), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n16419) );
  AOI211_X1 U19457 ( .C1(n19296), .C2(n16421), .A(n16420), .B(n16419), .ZN(
        n16423) );
  OAI211_X1 U19458 ( .C1(n19303), .C2(n16424), .A(n16423), .B(n16422), .ZN(
        P2_U3046) );
  NAND2_X1 U19459 ( .A1(n16425), .A2(n16451), .ZN(n16435) );
  AND3_X1 U19460 ( .A1(n16427), .A2(n16430), .A3(n16426), .ZN(n16433) );
  NAND2_X1 U19461 ( .A1(n11897), .A2(n15766), .ZN(n16428) );
  NAND2_X1 U19462 ( .A1(n16428), .A2(n9811), .ZN(n16429) );
  AOI21_X1 U19463 ( .B1(n16431), .B2(n16430), .A(n16429), .ZN(n16432) );
  MUX2_X1 U19464 ( .A(n16433), .B(n16432), .S(n11619), .Z(n16434) );
  NAND2_X1 U19465 ( .A1(n16435), .A2(n16434), .ZN(n16445) );
  MUX2_X1 U19466 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16445), .S(
        n16474), .Z(n16477) );
  MUX2_X1 U19467 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16436), .S(
        n16474), .Z(n16476) );
  INV_X1 U19468 ( .A(n12169), .ZN(n16439) );
  NAND2_X1 U19469 ( .A1(n16439), .A2(n16438), .ZN(n16442) );
  NAND2_X1 U19470 ( .A1(n16444), .A2(n16440), .ZN(n16441) );
  OAI211_X1 U19471 ( .C1(n16444), .C2(n16443), .A(n16442), .B(n16441), .ZN(
        n20046) );
  NOR2_X1 U19472 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n16469) );
  INV_X1 U19473 ( .A(n16445), .ZN(n19986) );
  INV_X1 U19474 ( .A(n11897), .ZN(n16448) );
  OAI22_X1 U19475 ( .A1(n19998), .A2(n16448), .B1(n16447), .B2(n16446), .ZN(
        n16449) );
  AOI22_X1 U19476 ( .A1(n16452), .A2(n16451), .B1(n16450), .B2(n16449), .ZN(
        n19993) );
  INV_X1 U19477 ( .A(n19993), .ZN(n16456) );
  AOI21_X1 U19478 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11897), .A(
        n20036), .ZN(n16453) );
  OAI211_X1 U19479 ( .C1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19993), .A(
        n16454), .B(n16453), .ZN(n16455) );
  OAI211_X1 U19480 ( .C1(n20028), .C2(n16456), .A(n16474), .B(n16455), .ZN(
        n16457) );
  AOI21_X1 U19481 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n19986), .A(
        n16457), .ZN(n16461) );
  INV_X1 U19482 ( .A(n16477), .ZN(n16459) );
  OAI21_X1 U19483 ( .B1(n16461), .B2(n20019), .A(n16476), .ZN(n16458) );
  NAND2_X1 U19484 ( .A1(n16459), .A2(n16458), .ZN(n16460) );
  AOI22_X1 U19485 ( .A1(n16461), .A2(n20019), .B1(n20012), .B2(n16460), .ZN(
        n16463) );
  OAI21_X1 U19486 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n16463), .A(
        n16462), .ZN(n16464) );
  INV_X1 U19487 ( .A(n16464), .ZN(n16468) );
  INV_X1 U19488 ( .A(n16465), .ZN(n16466) );
  NAND2_X1 U19489 ( .A1(n16466), .A2(n20055), .ZN(n16467) );
  OAI211_X1 U19490 ( .C1(n16470), .C2(n16469), .A(n16468), .B(n16467), .ZN(
        n16471) );
  NOR2_X1 U19491 ( .A1(n20046), .A2(n16471), .ZN(n16472) );
  OAI21_X1 U19492 ( .B1(n16474), .B2(n16473), .A(n16472), .ZN(n16475) );
  AOI21_X1 U19493 ( .B1(n16477), .B2(n16476), .A(n16475), .ZN(n16496) );
  NAND3_X1 U19494 ( .A1(n16496), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n16478), 
        .ZN(n16480) );
  NAND2_X1 U19495 ( .A1(n16480), .A2(n16479), .ZN(n16484) );
  NOR2_X1 U19496 ( .A1(n16482), .A2(n16481), .ZN(n16483) );
  NAND2_X1 U19497 ( .A1(n16486), .A2(n16485), .ZN(n20029) );
  AOI21_X1 U19498 ( .B1(n19888), .B2(n20029), .A(n20054), .ZN(n16488) );
  NOR3_X1 U19499 ( .A1(n16489), .A2(n16488), .A3(n16487), .ZN(n16494) );
  OAI21_X1 U19500 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16491), .A(n16490), 
        .ZN(n16492) );
  OAI21_X1 U19501 ( .B1(n19888), .B2(n20057), .A(n16492), .ZN(n16493) );
  OAI211_X1 U19502 ( .C1(n16496), .C2(n16495), .A(n16494), .B(n16493), .ZN(
        P2_U3176) );
  OAI221_X1 U19503 ( .B1(n12958), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n12958), 
        .C2(n19888), .A(n16497), .ZN(P2_U3593) );
  XOR2_X1 U19504 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16498), .Z(
        n16672) );
  AOI21_X1 U19505 ( .B1(n16500), .B2(n16499), .A(n16507), .ZN(n16505) );
  INV_X1 U19506 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16673) );
  NAND2_X1 U19507 ( .A1(n18296), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16501) );
  OAI221_X1 U19508 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16503), .C1(
        n16673), .C2(n16502), .A(n16501), .ZN(n16504) );
  AOI211_X1 U19509 ( .C1(n17828), .C2(n16672), .A(n16505), .B(n16504), .ZN(
        n16510) );
  NAND2_X1 U19510 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17672), .ZN(
        n18010) );
  NOR2_X1 U19511 ( .A1(n18008), .A2(n18010), .ZN(n18000) );
  INV_X1 U19512 ( .A(n18177), .ZN(n17871) );
  INV_X1 U19513 ( .A(n18175), .ZN(n17816) );
  NOR2_X1 U19514 ( .A1(n17649), .A2(n17650), .ZN(n17635) );
  NAND3_X1 U19515 ( .A1(n16508), .A2(n17635), .A3(n16507), .ZN(n16509) );
  OAI211_X1 U19516 ( .C1(n16511), .C2(n17880), .A(n16510), .B(n16509), .ZN(
        P3_U2800) );
  AOI21_X1 U19517 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17877), .A(
        n16512), .ZN(n16530) );
  NAND2_X1 U19518 ( .A1(n17628), .A2(n18194), .ZN(n16529) );
  INV_X1 U19519 ( .A(n9829), .ZN(n18773) );
  NAND2_X1 U19520 ( .A1(n17471), .A2(n18776), .ZN(n18176) );
  OAI22_X1 U19521 ( .A1(n18773), .A2(n18131), .B1(n18124), .B2(n18176), .ZN(
        n18089) );
  NOR2_X1 U19522 ( .A1(n18011), .A2(n18089), .ZN(n18045) );
  NOR2_X1 U19523 ( .A1(n18045), .A2(n18287), .ZN(n18060) );
  NOR2_X1 U19524 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16513), .ZN(
        n17618) );
  OAI21_X1 U19525 ( .B1(n17627), .B2(n17779), .A(n16514), .ZN(n16517) );
  NOR4_X1 U19526 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17779), .A3(
        n18300), .A4(n16517), .ZN(n16516) );
  INV_X1 U19527 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18930) );
  NOR2_X1 U19528 ( .A1(n16515), .A2(n18930), .ZN(n17611) );
  AOI211_X1 U19529 ( .C1(n18060), .C2(n17618), .A(n16516), .B(n17611), .ZN(
        n16528) );
  INV_X1 U19530 ( .A(n16517), .ZN(n17616) );
  INV_X1 U19531 ( .A(n16530), .ZN(n17615) );
  NOR2_X1 U19532 ( .A1(n17616), .A2(n17615), .ZN(n17614) );
  AOI211_X1 U19533 ( .C1(n17627), .C2(n16519), .A(n17614), .B(n16518), .ZN(
        n16526) );
  AOI211_X1 U19534 ( .C1(n9829), .C2(n16522), .A(n16521), .B(n16520), .ZN(
        n16523) );
  OAI21_X1 U19535 ( .B1(n16524), .B2(n18176), .A(n16523), .ZN(n16525) );
  OAI211_X1 U19536 ( .C1(n16526), .C2(n16525), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n16515), .ZN(n16527) );
  OAI211_X1 U19537 ( .C1(n16530), .C2(n16529), .A(n16528), .B(n16527), .ZN(
        P3_U2834) );
  NOR3_X1 U19538 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16532) );
  NOR4_X1 U19539 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16531) );
  INV_X2 U19540 ( .A(n16616), .ZN(U215) );
  NAND4_X1 U19541 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16532), .A3(n16531), .A4(
        U215), .ZN(U213) );
  INV_X2 U19542 ( .A(U214), .ZN(n16581) );
  INV_X1 U19543 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16618) );
  OAI222_X1 U19544 ( .A1(U212), .A2(n19218), .B1(n16583), .B2(n19367), .C1(
        U214), .C2(n16618), .ZN(U216) );
  INV_X1 U19545 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19221) );
  INV_X1 U19546 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16534) );
  OAI222_X1 U19547 ( .A1(U212), .A2(n19221), .B1(n16583), .B2(n14535), .C1(
        U214), .C2(n16534), .ZN(U217) );
  INV_X1 U19548 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n19224) );
  INV_X1 U19549 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n16535) );
  OAI222_X1 U19550 ( .A1(U212), .A2(n19224), .B1(n16583), .B2(n14540), .C1(
        U214), .C2(n16535), .ZN(U218) );
  INV_X2 U19551 ( .A(U212), .ZN(n16580) );
  AOI22_X1 U19552 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16580), .ZN(n16536) );
  OAI21_X1 U19553 ( .B1(n16537), .B2(n16583), .A(n16536), .ZN(U219) );
  AOI22_X1 U19554 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16580), .ZN(n16538) );
  OAI21_X1 U19555 ( .B1(n14551), .B2(n16583), .A(n16538), .ZN(U220) );
  AOI22_X1 U19556 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16580), .ZN(n16539) );
  OAI21_X1 U19557 ( .B1(n15260), .B2(n16583), .A(n16539), .ZN(U221) );
  AOI22_X1 U19558 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16580), .ZN(n16540) );
  OAI21_X1 U19559 ( .B1(n14560), .B2(n16583), .A(n16540), .ZN(U222) );
  AOI22_X1 U19560 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16580), .ZN(n16541) );
  OAI21_X1 U19561 ( .B1(n14567), .B2(n16583), .A(n16541), .ZN(U223) );
  AOI22_X1 U19562 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16580), .ZN(n16542) );
  OAI21_X1 U19563 ( .B1(n19363), .B2(n16583), .A(n16542), .ZN(U224) );
  AOI22_X1 U19564 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16580), .ZN(n16543) );
  OAI21_X1 U19565 ( .B1(n14579), .B2(n16583), .A(n16543), .ZN(U225) );
  AOI22_X1 U19566 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16580), .ZN(n16544) );
  OAI21_X1 U19567 ( .B1(n20296), .B2(n16583), .A(n16544), .ZN(U226) );
  AOI22_X1 U19568 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16580), .ZN(n16545) );
  OAI21_X1 U19569 ( .B1(n19346), .B2(n16583), .A(n16545), .ZN(U227) );
  AOI22_X1 U19570 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16580), .ZN(n16546) );
  OAI21_X1 U19571 ( .B1(n14593), .B2(n16583), .A(n16546), .ZN(U228) );
  AOI22_X1 U19572 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16580), .ZN(n16547) );
  OAI21_X1 U19573 ( .B1(n15322), .B2(n16583), .A(n16547), .ZN(U229) );
  INV_X1 U19574 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20277) );
  AOI22_X1 U19575 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16580), .ZN(n16548) );
  OAI21_X1 U19576 ( .B1(n20277), .B2(n16583), .A(n16548), .ZN(U230) );
  AOI22_X1 U19577 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16580), .ZN(n16549) );
  OAI21_X1 U19578 ( .B1(n20268), .B2(n16583), .A(n16549), .ZN(U231) );
  INV_X1 U19579 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16551) );
  AOI22_X1 U19580 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16580), .ZN(n16550) );
  OAI21_X1 U19581 ( .B1(n16551), .B2(n16583), .A(n16550), .ZN(U232) );
  INV_X1 U19582 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16553) );
  AOI22_X1 U19583 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16580), .ZN(n16552) );
  OAI21_X1 U19584 ( .B1(n16553), .B2(n16583), .A(n16552), .ZN(U233) );
  INV_X1 U19585 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16555) );
  AOI22_X1 U19586 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16580), .ZN(n16554) );
  OAI21_X1 U19587 ( .B1(n16555), .B2(n16583), .A(n16554), .ZN(U234) );
  INV_X1 U19588 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16557) );
  AOI22_X1 U19589 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16580), .ZN(n16556) );
  OAI21_X1 U19590 ( .B1(n16557), .B2(n16583), .A(n16556), .ZN(U235) );
  AOI22_X1 U19591 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16580), .ZN(n16558) );
  OAI21_X1 U19592 ( .B1(n16559), .B2(n16583), .A(n16558), .ZN(U236) );
  AOI22_X1 U19593 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16580), .ZN(n16560) );
  OAI21_X1 U19594 ( .B1(n16561), .B2(n16583), .A(n16560), .ZN(U237) );
  AOI22_X1 U19595 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16580), .ZN(n16562) );
  OAI21_X1 U19596 ( .B1(n16563), .B2(n16583), .A(n16562), .ZN(U238) );
  AOI22_X1 U19597 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16580), .ZN(n16564) );
  OAI21_X1 U19598 ( .B1(n16565), .B2(n16583), .A(n16564), .ZN(U239) );
  INV_X1 U19599 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16567) );
  AOI22_X1 U19600 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16580), .ZN(n16566) );
  OAI21_X1 U19601 ( .B1(n16567), .B2(n16583), .A(n16566), .ZN(U240) );
  INV_X1 U19602 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16569) );
  AOI22_X1 U19603 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16580), .ZN(n16568) );
  OAI21_X1 U19604 ( .B1(n16569), .B2(n16583), .A(n16568), .ZN(U241) );
  INV_X1 U19605 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16571) );
  AOI22_X1 U19606 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16580), .ZN(n16570) );
  OAI21_X1 U19607 ( .B1(n16571), .B2(n16583), .A(n16570), .ZN(U242) );
  INV_X1 U19608 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16573) );
  AOI22_X1 U19609 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16580), .ZN(n16572) );
  OAI21_X1 U19610 ( .B1(n16573), .B2(n16583), .A(n16572), .ZN(U243) );
  INV_X1 U19611 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16575) );
  AOI22_X1 U19612 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16580), .ZN(n16574) );
  OAI21_X1 U19613 ( .B1(n16575), .B2(n16583), .A(n16574), .ZN(U244) );
  AOI22_X1 U19614 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16580), .ZN(n16576) );
  OAI21_X1 U19615 ( .B1(n16577), .B2(n16583), .A(n16576), .ZN(U245) );
  AOI22_X1 U19616 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16580), .ZN(n16578) );
  OAI21_X1 U19617 ( .B1(n16579), .B2(n16583), .A(n16578), .ZN(U246) );
  AOI22_X1 U19618 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16581), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16580), .ZN(n16582) );
  OAI21_X1 U19619 ( .B1(n16584), .B2(n16583), .A(n16582), .ZN(U247) );
  OAI22_X1 U19620 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16616), .ZN(n16585) );
  INV_X1 U19621 ( .A(n16585), .ZN(U251) );
  OAI22_X1 U19622 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16616), .ZN(n16586) );
  INV_X1 U19623 ( .A(n16586), .ZN(U252) );
  INV_X1 U19624 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16587) );
  INV_X1 U19625 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18321) );
  AOI22_X1 U19626 ( .A1(n16616), .A2(n16587), .B1(n18321), .B2(U215), .ZN(U253) );
  INV_X1 U19627 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16588) );
  INV_X1 U19628 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18326) );
  AOI22_X1 U19629 ( .A1(n16616), .A2(n16588), .B1(n18326), .B2(U215), .ZN(U254) );
  INV_X1 U19630 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16589) );
  INV_X1 U19631 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18331) );
  AOI22_X1 U19632 ( .A1(n16616), .A2(n16589), .B1(n18331), .B2(U215), .ZN(U255) );
  INV_X1 U19633 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16590) );
  INV_X1 U19634 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18336) );
  AOI22_X1 U19635 ( .A1(n16616), .A2(n16590), .B1(n18336), .B2(U215), .ZN(U256) );
  INV_X1 U19636 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16591) );
  INV_X1 U19637 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18341) );
  AOI22_X1 U19638 ( .A1(n16612), .A2(n16591), .B1(n18341), .B2(U215), .ZN(U257) );
  INV_X1 U19639 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16592) );
  INV_X1 U19640 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18346) );
  AOI22_X1 U19641 ( .A1(n16616), .A2(n16592), .B1(n18346), .B2(U215), .ZN(U258) );
  OAI22_X1 U19642 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16616), .ZN(n16593) );
  INV_X1 U19643 ( .A(n16593), .ZN(U259) );
  INV_X1 U19644 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16594) );
  INV_X1 U19645 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17464) );
  AOI22_X1 U19646 ( .A1(n16612), .A2(n16594), .B1(n17464), .B2(U215), .ZN(U260) );
  INV_X1 U19647 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16595) );
  INV_X1 U19648 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U19649 ( .A1(n16612), .A2(n16595), .B1(n17458), .B2(U215), .ZN(U261) );
  OAI22_X1 U19650 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16616), .ZN(n16596) );
  INV_X1 U19651 ( .A(n16596), .ZN(U262) );
  INV_X1 U19652 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16597) );
  INV_X1 U19653 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U19654 ( .A1(n16612), .A2(n16597), .B1(n17451), .B2(U215), .ZN(U263) );
  INV_X1 U19655 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16598) );
  INV_X1 U19656 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U19657 ( .A1(n16616), .A2(n16598), .B1(n17446), .B2(U215), .ZN(U264) );
  OAI22_X1 U19658 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16616), .ZN(n16599) );
  INV_X1 U19659 ( .A(n16599), .ZN(U265) );
  OAI22_X1 U19660 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16612), .ZN(n16600) );
  INV_X1 U19661 ( .A(n16600), .ZN(U266) );
  OAI22_X1 U19662 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16616), .ZN(n16601) );
  INV_X1 U19663 ( .A(n16601), .ZN(U267) );
  OAI22_X1 U19664 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16616), .ZN(n16602) );
  INV_X1 U19665 ( .A(n16602), .ZN(U268) );
  OAI22_X1 U19666 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16616), .ZN(n16603) );
  INV_X1 U19667 ( .A(n16603), .ZN(U269) );
  OAI22_X1 U19668 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16616), .ZN(n16604) );
  INV_X1 U19669 ( .A(n16604), .ZN(U270) );
  INV_X1 U19670 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16605) );
  INV_X1 U19671 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19345) );
  AOI22_X1 U19672 ( .A1(n16612), .A2(n16605), .B1(n19345), .B2(U215), .ZN(U271) );
  OAI22_X1 U19673 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16612), .ZN(n16606) );
  INV_X1 U19674 ( .A(n16606), .ZN(U272) );
  OAI22_X1 U19675 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16612), .ZN(n16608) );
  INV_X1 U19676 ( .A(n16608), .ZN(U273) );
  INV_X1 U19677 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16609) );
  INV_X1 U19678 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19362) );
  AOI22_X1 U19679 ( .A1(n16616), .A2(n16609), .B1(n19362), .B2(U215), .ZN(U274) );
  INV_X1 U19680 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16610) );
  INV_X1 U19681 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n19319) );
  AOI22_X1 U19682 ( .A1(n16612), .A2(n16610), .B1(n19319), .B2(U215), .ZN(U275) );
  INV_X1 U19683 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16611) );
  INV_X1 U19684 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n19331) );
  AOI22_X1 U19685 ( .A1(n16612), .A2(n16611), .B1(n19331), .B2(U215), .ZN(U276) );
  INV_X1 U19686 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16613) );
  AOI22_X1 U19687 ( .A1(n16616), .A2(n16613), .B1(n15259), .B2(U215), .ZN(U277) );
  INV_X1 U19688 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16614) );
  INV_X1 U19689 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19340) );
  AOI22_X1 U19690 ( .A1(n16616), .A2(n16614), .B1(n19340), .B2(U215), .ZN(U278) );
  INV_X1 U19691 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16615) );
  INV_X1 U19692 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17364) );
  AOI22_X1 U19693 ( .A1(n16616), .A2(n16615), .B1(n17364), .B2(U215), .ZN(U279) );
  INV_X1 U19694 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19352) );
  AOI22_X1 U19695 ( .A1(n16616), .A2(n19224), .B1(n19352), .B2(U215), .ZN(U280) );
  INV_X1 U19696 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19358) );
  AOI22_X1 U19697 ( .A1(n16616), .A2(n19221), .B1(n19358), .B2(U215), .ZN(U281) );
  INV_X1 U19698 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19365) );
  AOI22_X1 U19699 ( .A1(n16616), .A2(n19218), .B1(n19365), .B2(U215), .ZN(U282) );
  INV_X1 U19700 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16617) );
  AOI222_X1 U19701 ( .A1(n16618), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19218), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16617), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16619) );
  INV_X2 U19702 ( .A(n16621), .ZN(n16620) );
  INV_X1 U19703 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18894) );
  INV_X1 U19704 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19931) );
  AOI22_X1 U19705 ( .A1(n16620), .A2(n18894), .B1(n19931), .B2(n16621), .ZN(
        U347) );
  INV_X1 U19706 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18892) );
  INV_X1 U19707 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19930) );
  AOI22_X1 U19708 ( .A1(n16620), .A2(n18892), .B1(n19930), .B2(n16621), .ZN(
        U348) );
  INV_X1 U19709 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18890) );
  INV_X1 U19710 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19928) );
  AOI22_X1 U19711 ( .A1(n16620), .A2(n18890), .B1(n19928), .B2(n16621), .ZN(
        U349) );
  INV_X1 U19712 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18888) );
  INV_X1 U19713 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19926) );
  AOI22_X1 U19714 ( .A1(n16620), .A2(n18888), .B1(n19926), .B2(n16621), .ZN(
        U350) );
  INV_X1 U19715 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18886) );
  INV_X1 U19716 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19925) );
  AOI22_X1 U19717 ( .A1(n16620), .A2(n18886), .B1(n19925), .B2(n16621), .ZN(
        U351) );
  INV_X1 U19718 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18884) );
  INV_X1 U19719 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19923) );
  AOI22_X1 U19720 ( .A1(n16620), .A2(n18884), .B1(n19923), .B2(n16621), .ZN(
        U352) );
  INV_X1 U19721 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18882) );
  INV_X1 U19722 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19921) );
  AOI22_X1 U19723 ( .A1(n16620), .A2(n18882), .B1(n19921), .B2(n16621), .ZN(
        U353) );
  INV_X1 U19724 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18880) );
  AOI22_X1 U19725 ( .A1(n16620), .A2(n18880), .B1(n19918), .B2(n16621), .ZN(
        U354) );
  INV_X1 U19726 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18932) );
  INV_X1 U19727 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19969) );
  AOI22_X1 U19728 ( .A1(n16620), .A2(n18932), .B1(n19969), .B2(n16621), .ZN(
        U356) );
  INV_X1 U19729 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18929) );
  INV_X1 U19730 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19967) );
  AOI22_X1 U19731 ( .A1(n16620), .A2(n18929), .B1(n19967), .B2(n16621), .ZN(
        U357) );
  INV_X1 U19732 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18928) );
  INV_X1 U19733 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19964) );
  AOI22_X1 U19734 ( .A1(n16620), .A2(n18928), .B1(n19964), .B2(n16621), .ZN(
        U358) );
  INV_X1 U19735 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18926) );
  INV_X1 U19736 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19963) );
  AOI22_X1 U19737 ( .A1(n16620), .A2(n18926), .B1(n19963), .B2(n16621), .ZN(
        U359) );
  INV_X1 U19738 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18924) );
  INV_X1 U19739 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19961) );
  AOI22_X1 U19740 ( .A1(n16620), .A2(n18924), .B1(n19961), .B2(n16621), .ZN(
        U360) );
  INV_X1 U19741 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18922) );
  INV_X1 U19742 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19959) );
  AOI22_X1 U19743 ( .A1(n16620), .A2(n18922), .B1(n19959), .B2(n16621), .ZN(
        U361) );
  INV_X1 U19744 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18919) );
  INV_X1 U19745 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19957) );
  AOI22_X1 U19746 ( .A1(n16620), .A2(n18919), .B1(n19957), .B2(n16621), .ZN(
        U362) );
  INV_X1 U19747 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18918) );
  INV_X1 U19748 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19955) );
  AOI22_X1 U19749 ( .A1(n16620), .A2(n18918), .B1(n19955), .B2(n16621), .ZN(
        U363) );
  INV_X1 U19750 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18915) );
  INV_X1 U19751 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19953) );
  AOI22_X1 U19752 ( .A1(n16620), .A2(n18915), .B1(n19953), .B2(n16621), .ZN(
        U364) );
  INV_X1 U19753 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18878) );
  INV_X1 U19754 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19916) );
  AOI22_X1 U19755 ( .A1(n16620), .A2(n18878), .B1(n19916), .B2(n16621), .ZN(
        U365) );
  INV_X1 U19756 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18914) );
  INV_X1 U19757 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19951) );
  AOI22_X1 U19758 ( .A1(n16620), .A2(n18914), .B1(n19951), .B2(n16621), .ZN(
        U366) );
  INV_X1 U19759 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18911) );
  INV_X1 U19760 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19949) );
  AOI22_X1 U19761 ( .A1(n16620), .A2(n18911), .B1(n19949), .B2(n16621), .ZN(
        U367) );
  INV_X1 U19762 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18910) );
  INV_X1 U19763 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19947) );
  AOI22_X1 U19764 ( .A1(n16620), .A2(n18910), .B1(n19947), .B2(n16621), .ZN(
        U368) );
  INV_X1 U19765 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18908) );
  INV_X1 U19766 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19945) );
  AOI22_X1 U19767 ( .A1(n16620), .A2(n18908), .B1(n19945), .B2(n16621), .ZN(
        U369) );
  INV_X1 U19768 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18906) );
  INV_X1 U19769 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19943) );
  AOI22_X1 U19770 ( .A1(n16620), .A2(n18906), .B1(n19943), .B2(n16621), .ZN(
        U370) );
  INV_X1 U19771 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18904) );
  INV_X1 U19772 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19941) );
  AOI22_X1 U19773 ( .A1(n16620), .A2(n18904), .B1(n19941), .B2(n16621), .ZN(
        U371) );
  INV_X1 U19774 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18902) );
  INV_X1 U19775 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19939) );
  AOI22_X1 U19776 ( .A1(n16620), .A2(n18902), .B1(n19939), .B2(n16621), .ZN(
        U372) );
  INV_X1 U19777 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18900) );
  INV_X1 U19778 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19937) );
  AOI22_X1 U19779 ( .A1(n16620), .A2(n18900), .B1(n19937), .B2(n16621), .ZN(
        U373) );
  INV_X1 U19780 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18898) );
  INV_X1 U19781 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19935) );
  AOI22_X1 U19782 ( .A1(n16620), .A2(n18898), .B1(n19935), .B2(n16621), .ZN(
        U374) );
  INV_X1 U19783 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18896) );
  INV_X1 U19784 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19933) );
  AOI22_X1 U19785 ( .A1(n16620), .A2(n18896), .B1(n19933), .B2(n16621), .ZN(
        U375) );
  INV_X1 U19786 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18876) );
  INV_X1 U19787 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19915) );
  AOI22_X1 U19788 ( .A1(n16620), .A2(n18876), .B1(n19915), .B2(n16621), .ZN(
        U376) );
  INV_X1 U19789 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16622) );
  INV_X1 U19790 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18875) );
  NAND2_X1 U19791 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18875), .ZN(n18867) );
  AOI22_X1 U19792 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18867), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18873), .ZN(n18951) );
  OAI21_X1 U19793 ( .B1(n18873), .B2(n16622), .A(n18948), .ZN(P3_U2633) );
  NAND2_X1 U19794 ( .A1(n18840), .A2(n18954), .ZN(n16626) );
  INV_X1 U19795 ( .A(n18851), .ZN(n16625) );
  INV_X1 U19796 ( .A(n16629), .ZN(n16623) );
  OAI21_X1 U19797 ( .B1(n16623), .B2(n17540), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16624) );
  OAI21_X1 U19798 ( .B1(n16626), .B2(n16625), .A(n16624), .ZN(P3_U2634) );
  AOI21_X1 U19799 ( .B1(n18873), .B2(n18875), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16627) );
  AOI22_X1 U19800 ( .A1(n18936), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16627), 
        .B2(n18997), .ZN(P3_U2635) );
  NOR2_X1 U19801 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18861) );
  OAI21_X1 U19802 ( .B1(n18861), .B2(BS16), .A(n18951), .ZN(n18949) );
  OAI21_X1 U19803 ( .B1(n18951), .B2(n19007), .A(n18949), .ZN(P3_U2636) );
  AND3_X1 U19804 ( .A1(n18779), .A2(n16629), .A3(n16628), .ZN(n18780) );
  NOR2_X1 U19805 ( .A1(n18780), .A2(n18846), .ZN(n18999) );
  OAI21_X1 U19806 ( .B1(n18999), .B2(n18305), .A(n16630), .ZN(P3_U2637) );
  NOR4_X1 U19807 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16634) );
  NOR4_X1 U19808 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16633) );
  NOR4_X1 U19809 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16632) );
  NOR4_X1 U19810 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16631) );
  NAND4_X1 U19811 ( .A1(n16634), .A2(n16633), .A3(n16632), .A4(n16631), .ZN(
        n16640) );
  NOR4_X1 U19812 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16638) );
  AOI211_X1 U19813 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16637) );
  NOR4_X1 U19814 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16636) );
  NOR4_X1 U19815 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16635) );
  NAND4_X1 U19816 ( .A1(n16638), .A2(n16637), .A3(n16636), .A4(n16635), .ZN(
        n16639) );
  NOR2_X1 U19817 ( .A1(n16640), .A2(n16639), .ZN(n18996) );
  INV_X1 U19818 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18944) );
  NOR3_X1 U19819 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16642) );
  OAI21_X1 U19820 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16642), .A(n18996), .ZN(
        n16641) );
  OAI21_X1 U19821 ( .B1(n18996), .B2(n18944), .A(n16641), .ZN(P3_U2638) );
  INV_X1 U19822 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18989) );
  INV_X1 U19823 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18950) );
  AOI21_X1 U19824 ( .B1(n18989), .B2(n18950), .A(n16642), .ZN(n16643) );
  INV_X1 U19825 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18941) );
  INV_X1 U19826 ( .A(n18996), .ZN(n18991) );
  AOI22_X1 U19827 ( .A1(n18996), .A2(n16643), .B1(n18941), .B2(n18991), .ZN(
        P3_U2639) );
  NOR4_X4 U19828 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n18966), .ZN(n17006) );
  NOR2_X1 U19829 ( .A1(n18199), .A2(n17006), .ZN(n16976) );
  NOR2_X2 U19830 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18954), .ZN(n18849) );
  NAND2_X1 U19831 ( .A1(n18851), .A2(n18849), .ZN(n18844) );
  INV_X1 U19832 ( .A(n19009), .ZN(n18860) );
  AOI211_X1 U19833 ( .C1(n19008), .C2(n19006), .A(n18860), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16644) );
  AOI211_X4 U19834 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16646), .A(n16644), .B(
        n19021), .ZN(n17024) );
  INV_X1 U19835 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18938) );
  INV_X1 U19836 ( .A(n16644), .ZN(n18838) );
  INV_X1 U19837 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18923) );
  INV_X1 U19838 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18920) );
  INV_X1 U19839 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18916) );
  INV_X1 U19840 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18912) );
  INV_X1 U19841 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18909) );
  INV_X1 U19842 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18901) );
  INV_X1 U19843 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18897) );
  INV_X1 U19844 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18893) );
  INV_X1 U19845 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18889) );
  INV_X1 U19846 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18885) );
  NAND3_X1 U19847 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16981) );
  NOR2_X1 U19848 ( .A1(n18881), .A2(n16981), .ZN(n16953) );
  NAND2_X1 U19849 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16953), .ZN(n16933) );
  NOR2_X1 U19850 ( .A1(n18885), .A2(n16933), .ZN(n16934) );
  NAND2_X1 U19851 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16934), .ZN(n16921) );
  NOR2_X1 U19852 ( .A1(n18889), .A2(n16921), .ZN(n16901) );
  NAND2_X1 U19853 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16901), .ZN(n16896) );
  NOR2_X1 U19854 ( .A1(n18893), .A2(n16896), .ZN(n16881) );
  NAND2_X1 U19855 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16881), .ZN(n16871) );
  NOR2_X1 U19856 ( .A1(n18897), .A2(n16871), .ZN(n16856) );
  NAND2_X1 U19857 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16856), .ZN(n16844) );
  NOR2_X1 U19858 ( .A1(n18901), .A2(n16844), .ZN(n16845) );
  NAND4_X1 U19859 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .A4(n16845), .ZN(n16790) );
  NOR3_X1 U19860 ( .A1(n18912), .A2(n18909), .A3(n16790), .ZN(n16784) );
  NAND2_X1 U19861 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16784), .ZN(n16758) );
  NOR2_X1 U19862 ( .A1(n18916), .A2(n16758), .ZN(n16757) );
  NAND2_X1 U19863 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16757), .ZN(n16744) );
  NOR2_X1 U19864 ( .A1(n18920), .A2(n16744), .ZN(n16736) );
  NAND2_X1 U19865 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16736), .ZN(n16727) );
  NOR2_X1 U19866 ( .A1(n18923), .A2(n16727), .ZN(n16712) );
  NAND2_X1 U19867 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16712), .ZN(n16661) );
  NAND4_X1 U19868 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16696), .ZN(n16663) );
  NOR3_X1 U19869 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18938), .A3(n16663), 
        .ZN(n16645) );
  AOI21_X1 U19870 ( .B1(n17024), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16645), .ZN(
        n16668) );
  NAND2_X1 U19871 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16646), .ZN(n16647) );
  AOI211_X4 U19872 ( .C1(n19007), .C2(n19009), .A(n19021), .B(n16647), .ZN(
        n17023) );
  NOR3_X1 U19873 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16996) );
  INV_X1 U19874 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17326) );
  NAND2_X1 U19875 ( .A1(n16996), .A2(n17326), .ZN(n16992) );
  NOR2_X1 U19876 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16992), .ZN(n16970) );
  INV_X1 U19877 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16961) );
  NAND2_X1 U19878 ( .A1(n16970), .A2(n16961), .ZN(n16960) );
  NAND2_X1 U19879 ( .A1(n16943), .A2(n17314), .ZN(n16939) );
  INV_X1 U19880 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16911) );
  NAND2_X1 U19881 ( .A1(n16920), .A2(n16911), .ZN(n16910) );
  NAND2_X1 U19882 ( .A1(n16897), .A2(n16648), .ZN(n16883) );
  INV_X1 U19883 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16862) );
  NAND2_X1 U19884 ( .A1(n16876), .A2(n16862), .ZN(n16861) );
  INV_X1 U19885 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16840) );
  NAND2_X1 U19886 ( .A1(n16846), .A2(n16840), .ZN(n16839) );
  INV_X1 U19887 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16821) );
  NAND2_X1 U19888 ( .A1(n16825), .A2(n16821), .ZN(n16818) );
  INV_X1 U19889 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17157) );
  NAND2_X1 U19890 ( .A1(n16803), .A2(n17157), .ZN(n16792) );
  NAND2_X1 U19891 ( .A1(n16781), .A2(n16778), .ZN(n16770) );
  NAND2_X1 U19892 ( .A1(n16759), .A2(n16753), .ZN(n16752) );
  NAND2_X1 U19893 ( .A1(n16723), .A2(n17035), .ZN(n16714) );
  NOR2_X1 U19894 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16714), .ZN(n16713) );
  INV_X1 U19895 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17078) );
  NAND2_X1 U19896 ( .A1(n16713), .A2(n17078), .ZN(n16707) );
  NOR2_X1 U19897 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16707), .ZN(n16691) );
  INV_X1 U19898 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16687) );
  NAND2_X1 U19899 ( .A1(n16691), .A2(n16687), .ZN(n16670) );
  NOR2_X1 U19900 ( .A1(n17016), .A2(n16670), .ZN(n16676) );
  INV_X1 U19901 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17041) );
  INV_X1 U19902 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16722) );
  NOR2_X1 U19903 ( .A1(n17975), .A2(n17653), .ZN(n16655) );
  INV_X1 U19904 ( .A(n16655), .ZN(n16656) );
  NOR2_X1 U19905 ( .A1(n17654), .A2(n16656), .ZN(n17620) );
  INV_X1 U19906 ( .A(n17620), .ZN(n16653) );
  NOR2_X1 U19907 ( .A1(n16722), .A2(n16653), .ZN(n16652) );
  NAND2_X1 U19908 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16652), .ZN(
        n16651) );
  AOI21_X1 U19909 ( .B1(n16650), .B2(n16651), .A(n16649), .ZN(n17613) );
  OAI21_X1 U19910 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16652), .A(
        n16651), .ZN(n17630) );
  INV_X1 U19911 ( .A(n17630), .ZN(n16703) );
  AOI21_X1 U19912 ( .B1(n16722), .B2(n16653), .A(n16652), .ZN(n17641) );
  INV_X1 U19913 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17668) );
  NOR2_X1 U19914 ( .A1(n17668), .A2(n16656), .ZN(n16654) );
  OAI21_X1 U19915 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16654), .A(
        n16653), .ZN(n17656) );
  INV_X1 U19916 ( .A(n17656), .ZN(n16726) );
  OAI22_X1 U19917 ( .A1(n17668), .A2(n16655), .B1(n16656), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17664) );
  NOR2_X1 U19918 ( .A1(n17975), .A2(n17698), .ZN(n16659) );
  NAND2_X1 U19919 ( .A1(n9918), .A2(n16659), .ZN(n17685) );
  INV_X1 U19920 ( .A(n17685), .ZN(n16657) );
  OAI21_X1 U19921 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n16657), .A(
        n16656), .ZN(n17681) );
  INV_X1 U19922 ( .A(n17681), .ZN(n16747) );
  INV_X1 U19923 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17699) );
  NAND2_X1 U19924 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16659), .ZN(
        n16658) );
  AOI21_X1 U19925 ( .B1(n17699), .B2(n16658), .A(n16657), .ZN(n17697) );
  OAI21_X1 U19926 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n16659), .A(
        n16658), .ZN(n17713) );
  INV_X1 U19927 ( .A(n17713), .ZN(n16769) );
  INV_X1 U19928 ( .A(n17737), .ZN(n16660) );
  INV_X1 U19929 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16826) );
  INV_X1 U19930 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17796) );
  INV_X1 U19931 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17911) );
  NAND2_X1 U19932 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17906), .ZN(
        n16954) );
  NOR2_X1 U19933 ( .A1(n17911), .A2(n16954), .ZN(n16942) );
  AND2_X1 U19934 ( .A1(n17794), .A2(n16942), .ZN(n16893) );
  NAND2_X1 U19935 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16893), .ZN(
        n16885) );
  INV_X1 U19936 ( .A(n16885), .ZN(n17808) );
  NAND2_X1 U19937 ( .A1(n17807), .A2(n17808), .ZN(n16860) );
  NOR2_X1 U19938 ( .A1(n17796), .A2(n16860), .ZN(n17769) );
  NAND2_X1 U19939 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17769), .ZN(
        n16833) );
  NOR2_X1 U19940 ( .A1(n16826), .A2(n16833), .ZN(n16822) );
  NAND2_X1 U19941 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16822), .ZN(
        n16809) );
  INV_X1 U19942 ( .A(n16809), .ZN(n17734) );
  NAND2_X1 U19943 ( .A1(n16660), .A2(n17734), .ZN(n17694) );
  AOI21_X1 U19944 ( .B1(n10031), .B2(n17694), .A(n16659), .ZN(n17725) );
  NOR2_X1 U19945 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16809), .ZN(
        n16800) );
  AOI21_X1 U19946 ( .B1(n16660), .B2(n16800), .A(n16985), .ZN(n16780) );
  NOR2_X1 U19947 ( .A1(n17725), .A2(n16780), .ZN(n16779) );
  NOR2_X1 U19948 ( .A1(n16779), .A2(n16894), .ZN(n16768) );
  NOR2_X1 U19949 ( .A1(n16769), .A2(n16768), .ZN(n16767) );
  NOR2_X1 U19950 ( .A1(n16767), .A2(n16894), .ZN(n16761) );
  NOR2_X1 U19951 ( .A1(n17697), .A2(n16761), .ZN(n16760) );
  NOR2_X1 U19952 ( .A1(n16738), .A2(n16894), .ZN(n16725) );
  NOR2_X1 U19953 ( .A1(n16726), .A2(n16725), .ZN(n16724) );
  NOR2_X1 U19954 ( .A1(n16724), .A2(n16985), .ZN(n16716) );
  NOR2_X1 U19955 ( .A1(n17641), .A2(n16716), .ZN(n16715) );
  NOR2_X1 U19956 ( .A1(n16692), .A2(n16894), .ZN(n16680) );
  NOR2_X1 U19957 ( .A1(n16894), .A2(n18852), .ZN(n17012) );
  INV_X1 U19958 ( .A(n17012), .ZN(n16944) );
  NOR3_X1 U19959 ( .A1(n16672), .A2(n16671), .A3(n16944), .ZN(n16666) );
  NAND3_X1 U19960 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16662) );
  AND2_X1 U19961 ( .A1(n16999), .A2(n16661), .ZN(n16711) );
  NOR2_X1 U19962 ( .A1(n17019), .A2(n16711), .ZN(n16710) );
  INV_X1 U19963 ( .A(n16710), .ZN(n16719) );
  AOI21_X1 U19964 ( .B1(n16999), .B2(n16662), .A(n16719), .ZN(n16690) );
  NOR2_X1 U19965 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16663), .ZN(n16675) );
  INV_X1 U19966 ( .A(n16675), .ZN(n16664) );
  AOI21_X1 U19967 ( .B1(n16690), .B2(n16664), .A(n18935), .ZN(n16665) );
  AOI211_X1 U19968 ( .C1(n16676), .C2(n17041), .A(n16666), .B(n16665), .ZN(
        n16667) );
  OAI211_X1 U19969 ( .C1(n16669), .C2(n16965), .A(n16668), .B(n16667), .ZN(
        P3_U2640) );
  NAND2_X1 U19970 ( .A1(n17023), .A2(n16670), .ZN(n16685) );
  OAI22_X1 U19971 ( .A1(n16690), .A2(n18938), .B1(n16673), .B2(n16965), .ZN(
        n16674) );
  OAI21_X1 U19972 ( .B1(n17024), .B2(n16676), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16677) );
  OAI211_X1 U19973 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16685), .A(n16678), .B(
        n16677), .ZN(P3_U2641) );
  INV_X1 U19974 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18931) );
  AOI211_X1 U19975 ( .C1(n16681), .C2(n16680), .A(n16679), .B(n18852), .ZN(
        n16684) );
  NAND3_X1 U19976 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16696), .ZN(n16682) );
  OAI22_X1 U19977 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16682), .B1(n10032), 
        .B2(n16965), .ZN(n16683) );
  AOI211_X1 U19978 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17024), .A(n16684), .B(
        n16683), .ZN(n16689) );
  INV_X1 U19979 ( .A(n16685), .ZN(n16686) );
  OAI21_X1 U19980 ( .B1(n16691), .B2(n16687), .A(n16686), .ZN(n16688) );
  OAI211_X1 U19981 ( .C1(n16690), .C2(n18931), .A(n16689), .B(n16688), .ZN(
        P3_U2642) );
  AOI22_X1 U19982 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17011), .B1(
        n17024), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16700) );
  AOI211_X1 U19983 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16707), .A(n16691), .B(
        n17016), .ZN(n16695) );
  AOI211_X1 U19984 ( .C1(n17613), .C2(n16693), .A(n16692), .B(n18852), .ZN(
        n16694) );
  NOR2_X1 U19985 ( .A1(n16695), .A2(n16694), .ZN(n16699) );
  INV_X1 U19986 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18927) );
  AND2_X1 U19987 ( .A1(n18927), .A2(n16696), .ZN(n16706) );
  OAI21_X1 U19988 ( .B1(n16706), .B2(n16719), .A(P3_REIP_REG_28__SCAN_IN), 
        .ZN(n16698) );
  NAND3_X1 U19989 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16696), .A3(n18930), 
        .ZN(n16697) );
  NAND4_X1 U19990 ( .A1(n16700), .A2(n16699), .A3(n16698), .A4(n16697), .ZN(
        P3_U2643) );
  AOI211_X1 U19991 ( .C1(n16703), .C2(n16702), .A(n16701), .B(n18852), .ZN(
        n16705) );
  OAI22_X1 U19992 ( .A1(n17610), .A2(n16965), .B1(n17013), .B2(n17078), .ZN(
        n16704) );
  NOR3_X1 U19993 ( .A1(n16706), .A2(n16705), .A3(n16704), .ZN(n16709) );
  OAI211_X1 U19994 ( .C1(n16713), .C2(n17078), .A(n17023), .B(n16707), .ZN(
        n16708) );
  OAI211_X1 U19995 ( .C1(n16710), .C2(n18927), .A(n16709), .B(n16708), .ZN(
        P3_U2644) );
  AOI22_X1 U19996 ( .A1(n17024), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16712), 
        .B2(n16711), .ZN(n16721) );
  AOI211_X1 U19997 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16714), .A(n16713), .B(
        n17016), .ZN(n16718) );
  AOI211_X1 U19998 ( .C1(n17641), .C2(n16716), .A(n16715), .B(n18852), .ZN(
        n16717) );
  AOI211_X1 U19999 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16719), .A(n16718), 
        .B(n16717), .ZN(n16720) );
  OAI211_X1 U20000 ( .C1(n16722), .C2(n16965), .A(n16721), .B(n16720), .ZN(
        P3_U2645) );
  OR2_X1 U20001 ( .A1(n17016), .A2(n16723), .ZN(n16737) );
  AOI21_X1 U20002 ( .B1(n17023), .B2(n16723), .A(n17024), .ZN(n16734) );
  AOI211_X1 U20003 ( .C1(n16726), .C2(n16725), .A(n16724), .B(n18852), .ZN(
        n16732) );
  NOR2_X1 U20004 ( .A1(n17025), .A2(n16727), .ZN(n16730) );
  INV_X1 U20005 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18921) );
  OAI21_X1 U20006 ( .B1(n16736), .B2(n17025), .A(n17028), .ZN(n16751) );
  AOI21_X1 U20007 ( .B1(n16999), .B2(n18921), .A(n16751), .ZN(n16728) );
  INV_X1 U20008 ( .A(n16728), .ZN(n16729) );
  MUX2_X1 U20009 ( .A(n16730), .B(n16729), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n16731) );
  AOI211_X1 U20010 ( .C1(n17011), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16732), .B(n16731), .ZN(n16733) );
  OAI221_X1 U20011 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16737), .C1(n17035), 
        .C2(n16734), .A(n16733), .ZN(P3_U2646) );
  NOR2_X1 U20012 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17025), .ZN(n16735) );
  AOI22_X1 U20013 ( .A1(n17024), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16736), 
        .B2(n16735), .ZN(n16743) );
  AOI21_X1 U20014 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16752), .A(n16737), .ZN(
        n16741) );
  AOI211_X1 U20015 ( .C1(n17664), .C2(n16739), .A(n16738), .B(n18852), .ZN(
        n16740) );
  AOI211_X1 U20016 ( .C1(n16751), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16741), 
        .B(n16740), .ZN(n16742) );
  OAI211_X1 U20017 ( .C1(n17668), .C2(n16965), .A(n16743), .B(n16742), .ZN(
        P3_U2647) );
  OAI21_X1 U20018 ( .B1(n17025), .B2(n16744), .A(n18920), .ZN(n16750) );
  AOI211_X1 U20019 ( .C1(n16747), .C2(n16746), .A(n16745), .B(n18852), .ZN(
        n16749) );
  INV_X1 U20020 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17684) );
  OAI22_X1 U20021 ( .A1(n17684), .A2(n16965), .B1(n17013), .B2(n16753), .ZN(
        n16748) );
  AOI211_X1 U20022 ( .C1(n16751), .C2(n16750), .A(n16749), .B(n16748), .ZN(
        n16755) );
  OAI211_X1 U20023 ( .C1(n16759), .C2(n16753), .A(n17023), .B(n16752), .ZN(
        n16754) );
  NAND2_X1 U20024 ( .A1(n16755), .A2(n16754), .ZN(P3_U2648) );
  NOR2_X1 U20025 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17025), .ZN(n16756) );
  AOI22_X1 U20026 ( .A1(n17024), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n16757), 
        .B2(n16756), .ZN(n16766) );
  INV_X1 U20027 ( .A(n16758), .ZN(n16775) );
  OAI221_X1 U20028 ( .B1(n17025), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n17025), 
        .C2(n16775), .A(n17028), .ZN(n16764) );
  AOI211_X1 U20029 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16770), .A(n16759), .B(
        n17016), .ZN(n16763) );
  AOI211_X1 U20030 ( .C1(n17697), .C2(n16761), .A(n16760), .B(n18852), .ZN(
        n16762) );
  AOI211_X1 U20031 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16764), .A(n16763), 
        .B(n16762), .ZN(n16765) );
  OAI211_X1 U20032 ( .C1(n17699), .C2(n16965), .A(n16766), .B(n16765), .ZN(
        P3_U2649) );
  NOR2_X1 U20033 ( .A1(n17025), .A2(n16775), .ZN(n16785) );
  NOR2_X1 U20034 ( .A1(n17019), .A2(n16785), .ZN(n16788) );
  INV_X1 U20035 ( .A(n16788), .ZN(n16774) );
  AOI211_X1 U20036 ( .C1(n16769), .C2(n16768), .A(n16767), .B(n18852), .ZN(
        n16773) );
  INV_X1 U20037 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17716) );
  OAI211_X1 U20038 ( .C1(n16781), .C2(n16778), .A(n17023), .B(n16770), .ZN(
        n16771) );
  OAI21_X1 U20039 ( .B1(n16965), .B2(n17716), .A(n16771), .ZN(n16772) );
  AOI211_X1 U20040 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16774), .A(n16773), 
        .B(n16772), .ZN(n16777) );
  NAND3_X1 U20041 ( .A1(n16999), .A2(n16775), .A3(n18916), .ZN(n16776) );
  OAI211_X1 U20042 ( .C1(n16778), .C2(n17013), .A(n16777), .B(n16776), .ZN(
        P3_U2650) );
  INV_X1 U20043 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18913) );
  AOI22_X1 U20044 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17011), .B1(
        n17024), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16787) );
  AOI211_X1 U20045 ( .C1(n17725), .C2(n16780), .A(n16779), .B(n18852), .ZN(
        n16783) );
  AOI211_X1 U20046 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16792), .A(n16781), .B(
        n17016), .ZN(n16782) );
  AOI211_X1 U20047 ( .C1(n16785), .C2(n16784), .A(n16783), .B(n16782), .ZN(
        n16786) );
  OAI211_X1 U20048 ( .C1(n16788), .C2(n18913), .A(n16787), .B(n16786), .ZN(
        P3_U2651) );
  INV_X1 U20049 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17748) );
  NOR2_X1 U20050 ( .A1(n17748), .A2(n16809), .ZN(n16799) );
  OAI21_X1 U20051 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16799), .A(
        n17694), .ZN(n17740) );
  INV_X1 U20052 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16987) );
  AOI21_X1 U20053 ( .B1(n16799), .B2(n16987), .A(n16894), .ZN(n16789) );
  XOR2_X1 U20054 ( .A(n17740), .B(n16789), .Z(n16797) );
  AOI21_X1 U20055 ( .B1(n16790), .B2(n16999), .A(n17019), .ZN(n16808) );
  INV_X1 U20056 ( .A(n16808), .ZN(n16817) );
  NOR3_X1 U20057 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17025), .A3(n16790), 
        .ZN(n16798) );
  NOR4_X1 U20058 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n17025), .A3(n18909), 
        .A4(n16790), .ZN(n16791) );
  AOI211_X1 U20059 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17011), .A(
        n18199), .B(n16791), .ZN(n16794) );
  OAI211_X1 U20060 ( .C1(n16803), .C2(n17157), .A(n17023), .B(n16792), .ZN(
        n16793) );
  OAI211_X1 U20061 ( .C1(n17157), .C2(n17013), .A(n16794), .B(n16793), .ZN(
        n16795) );
  AOI221_X1 U20062 ( .B1(n16817), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n16798), 
        .C2(P3_REIP_REG_19__SCAN_IN), .A(n16795), .ZN(n16796) );
  OAI21_X1 U20063 ( .B1(n18852), .B2(n16797), .A(n16796), .ZN(P3_U2652) );
  AOI211_X1 U20064 ( .C1(n17024), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18199), .B(
        n16798), .ZN(n16807) );
  AOI21_X1 U20065 ( .B1(n17748), .B2(n16809), .A(n16799), .ZN(n16802) );
  NOR2_X1 U20066 ( .A1(n16800), .A2(n16985), .ZN(n16812) );
  INV_X1 U20067 ( .A(n16802), .ZN(n17745) );
  INV_X1 U20068 ( .A(n16812), .ZN(n16801) );
  AOI221_X1 U20069 ( .B1(n16802), .B2(n16812), .C1(n17745), .C2(n16801), .A(
        n18852), .ZN(n16805) );
  AOI211_X1 U20070 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16818), .A(n16803), .B(
        n17016), .ZN(n16804) );
  AOI211_X1 U20071 ( .C1(n17011), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16805), .B(n16804), .ZN(n16806) );
  OAI211_X1 U20072 ( .C1(n18909), .C2(n16808), .A(n16807), .B(n16806), .ZN(
        P3_U2653) );
  INV_X1 U20073 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18905) );
  NOR3_X1 U20074 ( .A1(n17025), .A2(n18901), .A3(n16844), .ZN(n16838) );
  NAND2_X1 U20075 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16838), .ZN(n16832) );
  NOR3_X1 U20076 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n18905), .A3(n16832), 
        .ZN(n16816) );
  OAI21_X1 U20077 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16822), .A(
        n16809), .ZN(n17761) );
  INV_X1 U20078 ( .A(n17761), .ZN(n16813) );
  AOI21_X1 U20079 ( .B1(n16822), .B2(n16987), .A(n17761), .ZN(n16810) );
  AOI21_X1 U20080 ( .B1(n16931), .B2(n16810), .A(n18852), .ZN(n16811) );
  OAI21_X1 U20081 ( .B1(n16813), .B2(n16812), .A(n16811), .ZN(n16814) );
  OAI211_X1 U20082 ( .C1(n10030), .C2(n16965), .A(n16515), .B(n16814), .ZN(
        n16815) );
  AOI211_X1 U20083 ( .C1(n16817), .C2(P3_REIP_REG_17__SCAN_IN), .A(n16816), 
        .B(n16815), .ZN(n16820) );
  OAI211_X1 U20084 ( .C1(n16825), .C2(n16821), .A(n17023), .B(n16818), .ZN(
        n16819) );
  OAI211_X1 U20085 ( .C1(n16821), .C2(n17013), .A(n16820), .B(n16819), .ZN(
        P3_U2654) );
  INV_X1 U20086 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18903) );
  OAI21_X1 U20087 ( .B1(n16845), .B2(n17025), .A(n17028), .ZN(n16851) );
  AOI21_X1 U20088 ( .B1(n16838), .B2(n18903), .A(n16851), .ZN(n16831) );
  AOI21_X1 U20089 ( .B1(n16826), .B2(n16833), .A(n16822), .ZN(n17770) );
  INV_X1 U20090 ( .A(n16833), .ZN(n16823) );
  AOI21_X1 U20091 ( .B1(n16823), .B2(n16987), .A(n16894), .ZN(n16835) );
  OAI21_X1 U20092 ( .B1(n17770), .B2(n16835), .A(n17006), .ZN(n16824) );
  AOI21_X1 U20093 ( .B1(n17770), .B2(n16835), .A(n16824), .ZN(n16829) );
  AOI211_X1 U20094 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16839), .A(n16825), .B(
        n17016), .ZN(n16828) );
  OAI22_X1 U20095 ( .A1(n16826), .A2(n16965), .B1(n17013), .B2(n17206), .ZN(
        n16827) );
  NOR4_X1 U20096 ( .A1(n18296), .A2(n16829), .A3(n16828), .A4(n16827), .ZN(
        n16830) );
  OAI221_X1 U20097 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16832), .C1(n18905), 
        .C2(n16831), .A(n16830), .ZN(P3_U2655) );
  NAND2_X1 U20098 ( .A1(n17006), .A2(n16894), .ZN(n17010) );
  OAI21_X1 U20099 ( .B1(n16894), .B2(n16987), .A(n17006), .ZN(n17022) );
  OAI21_X1 U20100 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17769), .A(
        n16833), .ZN(n17782) );
  AOI211_X1 U20101 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17010), .A(
        n17022), .B(n17782), .ZN(n16834) );
  AOI21_X1 U20102 ( .B1(n17011), .B2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16834), .ZN(n16843) );
  NAND3_X1 U20103 ( .A1(n17006), .A2(n16835), .A3(n17782), .ZN(n16836) );
  OAI211_X1 U20104 ( .C1(n17013), .C2(n16840), .A(n16515), .B(n16836), .ZN(
        n16837) );
  AOI221_X1 U20105 ( .B1(n16851), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n16838), 
        .C2(n18903), .A(n16837), .ZN(n16842) );
  OAI211_X1 U20106 ( .C1(n16846), .C2(n16840), .A(n17023), .B(n16839), .ZN(
        n16841) );
  NAND3_X1 U20107 ( .A1(n16843), .A2(n16842), .A3(n16841), .ZN(P3_U2656) );
  AOI22_X1 U20108 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17011), .B1(
        n17024), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16855) );
  NOR2_X1 U20109 ( .A1(n17025), .A2(n16844), .ZN(n16849) );
  INV_X1 U20110 ( .A(n16845), .ZN(n16848) );
  AOI211_X1 U20111 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16861), .A(n16846), .B(
        n17016), .ZN(n16847) );
  AOI211_X1 U20112 ( .C1(n16849), .C2(n16848), .A(n18199), .B(n16847), .ZN(
        n16854) );
  AOI21_X1 U20113 ( .B1(n17796), .B2(n16860), .A(n17769), .ZN(n17799) );
  NOR2_X1 U20114 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17975), .ZN(
        n17007) );
  INV_X1 U20115 ( .A(n17007), .ZN(n16972) );
  NOR2_X1 U20116 ( .A1(n17872), .A2(n16972), .ZN(n16945) );
  INV_X1 U20117 ( .A(n16945), .ZN(n16930) );
  OAI21_X1 U20118 ( .B1(n16850), .B2(n16930), .A(n16931), .ZN(n16887) );
  OAI21_X1 U20119 ( .B1(n17807), .B2(n16985), .A(n16887), .ZN(n16868) );
  XOR2_X1 U20120 ( .A(n17799), .B(n16868), .Z(n16852) );
  AOI22_X1 U20121 ( .A1(n17006), .A2(n16852), .B1(P3_REIP_REG_14__SCAN_IN), 
        .B2(n16851), .ZN(n16853) );
  NAND3_X1 U20122 ( .A1(n16855), .A2(n16854), .A3(n16853), .ZN(P3_U2657) );
  AOI21_X1 U20123 ( .B1(n16999), .B2(n16871), .A(n17019), .ZN(n16891) );
  OAI21_X1 U20124 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17025), .A(n16891), 
        .ZN(n16867) );
  NAND2_X1 U20125 ( .A1(n16999), .A2(n16856), .ZN(n16857) );
  OAI22_X1 U20126 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16857), .B1(n17013), 
        .B2(n16862), .ZN(n16866) );
  NOR2_X1 U20127 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18852), .ZN(
        n16859) );
  INV_X1 U20128 ( .A(n17010), .ZN(n16858) );
  AOI21_X1 U20129 ( .B1(n16859), .B2(n17813), .A(n16858), .ZN(n16864) );
  NOR2_X1 U20130 ( .A1(n17824), .A2(n16885), .ZN(n16873) );
  OAI21_X1 U20131 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16873), .A(
        n16860), .ZN(n17811) );
  OAI211_X1 U20132 ( .C1(n16876), .C2(n16862), .A(n17023), .B(n16861), .ZN(
        n16863) );
  OAI211_X1 U20133 ( .C1(n16864), .C2(n17811), .A(n16515), .B(n16863), .ZN(
        n16865) );
  AOI211_X1 U20134 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16867), .A(n16866), 
        .B(n16865), .ZN(n16870) );
  NAND3_X1 U20135 ( .A1(n17006), .A2(n17811), .A3(n16868), .ZN(n16869) );
  OAI211_X1 U20136 ( .C1(n16965), .C2(n17813), .A(n16870), .B(n16869), .ZN(
        P3_U2658) );
  NOR3_X1 U20137 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17025), .A3(n16871), 
        .ZN(n16872) );
  AOI211_X1 U20138 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17011), .A(
        n18199), .B(n16872), .ZN(n16880) );
  AOI21_X1 U20139 ( .B1(n17824), .B2(n16885), .A(n16873), .ZN(n17827) );
  INV_X1 U20140 ( .A(n16887), .ZN(n16875) );
  INV_X1 U20141 ( .A(n17827), .ZN(n16874) );
  AOI221_X1 U20142 ( .B1(n17827), .B2(n16875), .C1(n16874), .C2(n16887), .A(
        n18852), .ZN(n16878) );
  AOI211_X1 U20143 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16883), .A(n16876), .B(
        n17016), .ZN(n16877) );
  AOI211_X1 U20144 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17024), .A(n16878), .B(
        n16877), .ZN(n16879) );
  OAI211_X1 U20145 ( .C1(n18897), .C2(n16891), .A(n16880), .B(n16879), .ZN(
        P3_U2659) );
  AOI21_X1 U20146 ( .B1(n16999), .B2(n16881), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16892) );
  INV_X1 U20147 ( .A(n16897), .ZN(n16882) );
  AOI21_X1 U20148 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n16882), .A(n17016), .ZN(
        n16884) );
  AOI22_X1 U20149 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17011), .B1(
        n16884), .B2(n16883), .ZN(n16890) );
  OAI21_X1 U20150 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16893), .A(
        n16885), .ZN(n17846) );
  NOR3_X1 U20151 ( .A1(n17873), .A2(n16908), .A3(n16930), .ZN(n16895) );
  OAI221_X1 U20152 ( .B1(n17846), .B2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C1(
        n17846), .C2(n16895), .A(n17006), .ZN(n16886) );
  AOI22_X1 U20153 ( .A1(n17846), .A2(n16887), .B1(n17010), .B2(n16886), .ZN(
        n16888) );
  AOI211_X1 U20154 ( .C1(n17024), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18199), .B(
        n16888), .ZN(n16889) );
  OAI211_X1 U20155 ( .C1(n16892), .C2(n16891), .A(n16890), .B(n16889), .ZN(
        P3_U2660) );
  INV_X1 U20156 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17876) );
  INV_X1 U20157 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17886) );
  OR3_X1 U20158 ( .A1(n17975), .A2(n17872), .A3(n17886), .ZN(n16929) );
  NOR2_X1 U20159 ( .A1(n17876), .A2(n16929), .ZN(n16918) );
  NAND2_X1 U20160 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16918), .ZN(
        n16905) );
  AOI21_X1 U20161 ( .B1(n17849), .B2(n16905), .A(n16893), .ZN(n17847) );
  NOR2_X1 U20162 ( .A1(n16895), .A2(n16894), .ZN(n16907) );
  XNOR2_X1 U20163 ( .A(n17847), .B(n16907), .ZN(n16904) );
  NOR3_X1 U20164 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n17025), .A3(n16896), 
        .ZN(n16900) );
  AOI211_X1 U20165 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16910), .A(n16897), .B(
        n17016), .ZN(n16899) );
  INV_X1 U20166 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17270) );
  OAI22_X1 U20167 ( .A1(n17849), .A2(n16965), .B1(n17013), .B2(n17270), .ZN(
        n16898) );
  NOR4_X1 U20168 ( .A1(n18296), .A2(n16900), .A3(n16899), .A4(n16898), .ZN(
        n16903) );
  NOR4_X1 U20169 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17025), .A3(n18889), .A4(
        n16921), .ZN(n16909) );
  OAI21_X1 U20170 ( .B1(n16901), .B2(n17025), .A(n17028), .ZN(n16922) );
  OAI21_X1 U20171 ( .B1(n16909), .B2(n16922), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16902) );
  OAI211_X1 U20172 ( .C1(n18852), .C2(n16904), .A(n16903), .B(n16902), .ZN(
        P3_U2661) );
  OAI21_X1 U20173 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16918), .A(
        n16905), .ZN(n17865) );
  NOR2_X1 U20174 ( .A1(n17873), .A2(n16930), .ZN(n16906) );
  AOI22_X1 U20175 ( .A1(n16907), .A2(n17865), .B1(n16906), .B2(n16908), .ZN(
        n16917) );
  OAI22_X1 U20176 ( .A1(n16908), .A2(n16965), .B1(n17013), .B2(n16911), .ZN(
        n16915) );
  INV_X1 U20177 ( .A(n16909), .ZN(n16913) );
  OAI211_X1 U20178 ( .C1(n16920), .C2(n16911), .A(n17023), .B(n16910), .ZN(
        n16912) );
  OAI211_X1 U20179 ( .C1(n17010), .C2(n17865), .A(n16913), .B(n16912), .ZN(
        n16914) );
  AOI211_X1 U20180 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n16922), .A(n16915), .B(
        n16914), .ZN(n16916) );
  OAI211_X1 U20181 ( .C1(n16917), .C2(n18852), .A(n16916), .B(n16515), .ZN(
        P3_U2662) );
  OAI21_X1 U20182 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16929), .A(
        n16931), .ZN(n16919) );
  AOI21_X1 U20183 ( .B1(n17876), .B2(n16929), .A(n16918), .ZN(n17883) );
  XOR2_X1 U20184 ( .A(n16919), .B(n17883), .Z(n16928) );
  AOI211_X1 U20185 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16939), .A(n16920), .B(
        n17016), .ZN(n16926) );
  NOR2_X1 U20186 ( .A1(n17025), .A2(n16921), .ZN(n16923) );
  OAI21_X1 U20187 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n16923), .A(n16922), .ZN(
        n16924) );
  OAI211_X1 U20188 ( .C1(n17013), .C2(n13776), .A(n16515), .B(n16924), .ZN(
        n16925) );
  AOI211_X1 U20189 ( .C1(n17011), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16926), .B(n16925), .ZN(n16927) );
  OAI21_X1 U20190 ( .B1(n16928), .B2(n18852), .A(n16927), .ZN(P3_U2663) );
  OAI21_X1 U20191 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16942), .A(
        n16929), .ZN(n17897) );
  NAND2_X1 U20192 ( .A1(n16931), .A2(n16930), .ZN(n16932) );
  XOR2_X1 U20193 ( .A(n17897), .B(n16932), .Z(n16938) );
  AOI21_X1 U20194 ( .B1(n16999), .B2(n16933), .A(n17019), .ZN(n16958) );
  OR3_X1 U20195 ( .A1(n17025), .A2(n16933), .A3(P3_REIP_REG_6__SCAN_IN), .ZN(
        n16951) );
  INV_X1 U20196 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18887) );
  AOI21_X1 U20197 ( .B1(n16958), .B2(n16951), .A(n18887), .ZN(n16937) );
  NAND3_X1 U20198 ( .A1(n16999), .A2(n16934), .A3(n18887), .ZN(n16935) );
  OAI211_X1 U20199 ( .C1(n17886), .C2(n16965), .A(n16515), .B(n16935), .ZN(
        n16936) );
  AOI211_X1 U20200 ( .C1(n17006), .C2(n16938), .A(n16937), .B(n16936), .ZN(
        n16941) );
  OAI211_X1 U20201 ( .C1(n16943), .C2(n17314), .A(n17023), .B(n16939), .ZN(
        n16940) );
  OAI211_X1 U20202 ( .C1(n17314), .C2(n17013), .A(n16941), .B(n16940), .ZN(
        P3_U2664) );
  AOI21_X1 U20203 ( .B1(n17911), .B2(n16954), .A(n16942), .ZN(n17914) );
  AOI21_X1 U20204 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17010), .A(
        n17022), .ZN(n16950) );
  AOI211_X1 U20205 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16960), .A(n16943), .B(
        n17016), .ZN(n16947) );
  NOR3_X1 U20206 ( .A1(n17914), .A2(n16945), .A3(n16944), .ZN(n16946) );
  AOI211_X1 U20207 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17024), .A(n16947), .B(
        n16946), .ZN(n16948) );
  OAI211_X1 U20208 ( .C1(n16958), .C2(n18885), .A(n16948), .B(n16515), .ZN(
        n16949) );
  AOI21_X1 U20209 ( .B1(n17914), .B2(n16950), .A(n16949), .ZN(n16952) );
  OAI211_X1 U20210 ( .C1(n16965), .C2(n17911), .A(n16952), .B(n16951), .ZN(
        P3_U2665) );
  INV_X1 U20211 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16964) );
  AOI21_X1 U20212 ( .B1(n16999), .B2(n16953), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16957) );
  NAND2_X1 U20213 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17916), .ZN(
        n16967) );
  INV_X1 U20214 ( .A(n16954), .ZN(n16955) );
  AOI21_X1 U20215 ( .B1(n16964), .B2(n16967), .A(n16955), .ZN(n17922) );
  AOI21_X1 U20216 ( .B1(n17916), .B2(n17007), .A(n16985), .ZN(n16974) );
  XNOR2_X1 U20217 ( .A(n17922), .B(n16974), .ZN(n16956) );
  OAI22_X1 U20218 ( .A1(n16958), .A2(n16957), .B1(n18852), .B2(n16956), .ZN(
        n16959) );
  AOI211_X1 U20219 ( .C1(n17024), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18199), .B(
        n16959), .ZN(n16963) );
  OAI211_X1 U20220 ( .C1(n16970), .C2(n16961), .A(n17023), .B(n16960), .ZN(
        n16962) );
  OAI211_X1 U20221 ( .C1(n16965), .C2(n16964), .A(n16963), .B(n16962), .ZN(
        P3_U2666) );
  NOR2_X1 U20222 ( .A1(n17975), .A2(n16966), .ZN(n16983) );
  OAI21_X1 U20223 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16983), .A(
        n16967), .ZN(n17937) );
  NAND2_X1 U20224 ( .A1(n18314), .A2(n19023), .ZN(n17015) );
  AOI21_X1 U20225 ( .B1(n11489), .B2(n18783), .A(n17015), .ZN(n16969) );
  NOR3_X1 U20226 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17025), .A3(n16981), .ZN(
        n16968) );
  AOI211_X1 U20227 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17024), .A(n16969), .B(
        n16968), .ZN(n16980) );
  AOI211_X1 U20228 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16992), .A(n16970), .B(
        n17016), .ZN(n16978) );
  NAND2_X1 U20229 ( .A1(n17945), .A2(n16971), .ZN(n17930) );
  OAI21_X1 U20230 ( .B1(n17930), .B2(n16972), .A(n16515), .ZN(n16973) );
  AOI21_X1 U20231 ( .B1(n16974), .B2(n17937), .A(n16973), .ZN(n16975) );
  AOI21_X1 U20232 ( .B1(n16999), .B2(n16981), .A(n17019), .ZN(n16989) );
  OAI22_X1 U20233 ( .A1(n16976), .A2(n16975), .B1(n16989), .B2(n18881), .ZN(
        n16977) );
  AOI211_X1 U20234 ( .C1(n17011), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16978), .B(n16977), .ZN(n16979) );
  OAI211_X1 U20235 ( .C1(n17937), .C2(n17010), .A(n16980), .B(n16979), .ZN(
        P3_U2667) );
  NAND2_X1 U20236 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16998) );
  NAND2_X1 U20237 ( .A1(n16999), .A2(n16981), .ZN(n16982) );
  OAI21_X1 U20238 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18794), .A(
        n11489), .ZN(n18955) );
  OAI22_X1 U20239 ( .A1(n16998), .A2(n16982), .B1(n17015), .B2(n18955), .ZN(
        n16991) );
  INV_X1 U20240 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18879) );
  NAND2_X1 U20241 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16995) );
  AOI21_X1 U20242 ( .B1(n16984), .B2(n16995), .A(n16983), .ZN(n17948) );
  INV_X1 U20243 ( .A(n16995), .ZN(n16986) );
  AOI21_X1 U20244 ( .B1(n16987), .B2(n16986), .A(n16985), .ZN(n17005) );
  XNOR2_X1 U20245 ( .A(n17948), .B(n17005), .ZN(n16988) );
  OAI22_X1 U20246 ( .A1(n16989), .A2(n18879), .B1(n18852), .B2(n16988), .ZN(
        n16990) );
  AOI211_X1 U20247 ( .C1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n17011), .A(
        n16991), .B(n16990), .ZN(n16994) );
  OAI211_X1 U20248 ( .C1(n16996), .C2(n17326), .A(n17023), .B(n16992), .ZN(
        n16993) );
  OAI211_X1 U20249 ( .C1(n17326), .C2(n17013), .A(n16994), .B(n16993), .ZN(
        P3_U2668) );
  OAI21_X1 U20250 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16995), .ZN(n17965) );
  INV_X1 U20251 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17343) );
  INV_X1 U20252 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17337) );
  NAND2_X1 U20253 ( .A1(n17343), .A2(n17337), .ZN(n16997) );
  AOI211_X1 U20254 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16997), .A(n16996), .B(
        n17016), .ZN(n17004) );
  NAND2_X1 U20255 ( .A1(n18972), .A2(n11307), .ZN(n18793) );
  INV_X1 U20256 ( .A(n18793), .ZN(n18784) );
  NOR2_X1 U20257 ( .A1(n18794), .A2(n18784), .ZN(n18969) );
  INV_X1 U20258 ( .A(n17015), .ZN(n17026) );
  AOI22_X1 U20259 ( .A1(n17019), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18969), 
        .B2(n17026), .ZN(n17001) );
  OAI211_X1 U20260 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16999), .B(n16998), .ZN(n17000) );
  OAI211_X1 U20261 ( .C1(n17002), .C2(n17013), .A(n17001), .B(n17000), .ZN(
        n17003) );
  AOI211_X1 U20262 ( .C1(n17011), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17004), .B(n17003), .ZN(n17009) );
  OAI211_X1 U20263 ( .C1(n17007), .C2(n17965), .A(n17006), .B(n17005), .ZN(
        n17008) );
  OAI211_X1 U20264 ( .C1(n17010), .C2(n17965), .A(n17009), .B(n17008), .ZN(
        P3_U2669) );
  AOI21_X1 U20265 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17012), .A(
        n17011), .ZN(n17021) );
  OAI22_X1 U20266 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17025), .B1(n17013), 
        .B2(n17337), .ZN(n17018) );
  OAI21_X1 U20267 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17332), .ZN(n17339) );
  NAND2_X1 U20268 ( .A1(n17014), .A2(n11307), .ZN(n18973) );
  OAI22_X1 U20269 ( .A1(n17016), .A2(n17339), .B1(n18973), .B2(n17015), .ZN(
        n17017) );
  AOI211_X1 U20270 ( .C1(n17019), .C2(P3_REIP_REG_1__SCAN_IN), .A(n17018), .B(
        n17017), .ZN(n17020) );
  OAI221_X1 U20271 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17022), .C1(
        n17975), .C2(n17021), .A(n17020), .ZN(P3_U2670) );
  NOR2_X1 U20272 ( .A1(n17024), .A2(n17023), .ZN(n17031) );
  NAND2_X1 U20273 ( .A1(n17028), .A2(n17025), .ZN(n17027) );
  AOI22_X1 U20274 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17027), .B1(n17026), 
        .B2(n18987), .ZN(n17030) );
  NAND3_X1 U20275 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18956), .A3(
        n17028), .ZN(n17029) );
  OAI211_X1 U20276 ( .C1(n17031), .C2(n17343), .A(n17030), .B(n17029), .ZN(
        P3_U2671) );
  INV_X1 U20277 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17033) );
  NOR2_X1 U20278 ( .A1(n17033), .A2(n17032), .ZN(n17112) );
  INV_X1 U20279 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17036) );
  NAND4_X1 U20280 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17034)
         );
  NOR3_X1 U20281 ( .A1(n17036), .A2(n17035), .A3(n17034), .ZN(n17037) );
  NAND4_X1 U20282 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17073), .A3(n17112), 
        .A4(n17037), .ZN(n17040) );
  NOR2_X1 U20283 ( .A1(n17041), .A2(n17040), .ZN(n17068) );
  NAND2_X1 U20284 ( .A1(n17336), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17039) );
  NAND2_X1 U20285 ( .A1(n17068), .A2(n18350), .ZN(n17038) );
  OAI22_X1 U20286 ( .A1(n17068), .A2(n17039), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17038), .ZN(P3_U2672) );
  NAND2_X1 U20287 ( .A1(n17041), .A2(n17040), .ZN(n17042) );
  NAND2_X1 U20288 ( .A1(n17042), .A2(n17336), .ZN(n17067) );
  AOI22_X1 U20289 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11378), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20290 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20291 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17043) );
  OAI211_X1 U20292 ( .C1(n17296), .C2(n17045), .A(n17044), .B(n17043), .ZN(
        n17051) );
  AOI22_X1 U20293 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20294 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20295 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9809), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17047) );
  NAND2_X1 U20296 ( .A1(n9804), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n17046) );
  NAND4_X1 U20297 ( .A1(n17049), .A2(n17048), .A3(n17047), .A4(n17046), .ZN(
        n17050) );
  AOI211_X1 U20298 ( .C1(n9810), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17051), .B(n17050), .ZN(n17052) );
  OAI211_X1 U20299 ( .C1(n10327), .C2(n18759), .A(n17053), .B(n17052), .ZN(
        n17070) );
  NAND2_X1 U20300 ( .A1(n17071), .A2(n17070), .ZN(n17069) );
  AOI22_X1 U20301 ( .A1(n11309), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17297), .ZN(n17065) );
  OAI22_X1 U20302 ( .A1(n17172), .A2(n17054), .B1(n13764), .B2(n18397), .ZN(
        n17062) );
  AOI22_X1 U20303 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11331), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n11378), .ZN(n17060) );
  AOI22_X1 U20304 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17292), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n15791), .ZN(n17056) );
  AOI22_X1 U20305 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17298), .ZN(n17055) );
  OAI211_X1 U20306 ( .C1(n17057), .C2(n17296), .A(n17056), .B(n17055), .ZN(
        n17058) );
  AOI21_X1 U20307 ( .B1(n9809), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(n17058), .ZN(n17059) );
  OAI211_X1 U20308 ( .C1(n17220), .C2(n11450), .A(n17060), .B(n17059), .ZN(
        n17061) );
  AOI211_X1 U20309 ( .C1(n9810), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n17062), .B(n17061), .ZN(n17064) );
  AOI22_X1 U20310 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17117), .ZN(n17063) );
  NAND3_X1 U20311 ( .A1(n17065), .A2(n17064), .A3(n17063), .ZN(n17066) );
  XOR2_X1 U20312 ( .A(n17069), .B(n17066), .Z(n17352) );
  OAI22_X1 U20313 ( .A1(n17068), .A2(n17067), .B1(n17352), .B2(n17336), .ZN(
        P3_U2673) );
  OAI21_X1 U20314 ( .B1(n17071), .B2(n17070), .A(n17069), .ZN(n17359) );
  NOR2_X1 U20315 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17079), .ZN(n17072) );
  AOI22_X1 U20316 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17074), .B1(n17073), 
        .B2(n17072), .ZN(n17075) );
  OAI21_X1 U20317 ( .B1(n17324), .B2(n17359), .A(n17075), .ZN(P3_U2674) );
  OAI211_X1 U20318 ( .C1(n17367), .C2(n17366), .A(n17341), .B(n17365), .ZN(
        n17076) );
  OAI221_X1 U20319 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17079), .C1(n17078), 
        .C2(n17077), .A(n17076), .ZN(P3_U2676) );
  AOI21_X1 U20320 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17336), .A(n17088), .ZN(
        n17081) );
  XNOR2_X1 U20321 ( .A(n17080), .B(n17084), .ZN(n17376) );
  OAI22_X1 U20322 ( .A1(n17082), .A2(n17081), .B1(n17336), .B2(n17376), .ZN(
        P3_U2677) );
  INV_X1 U20323 ( .A(n17083), .ZN(n17091) );
  AOI21_X1 U20324 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17336), .A(n17091), .ZN(
        n17087) );
  OAI21_X1 U20325 ( .B1(n17086), .B2(n17085), .A(n17084), .ZN(n17381) );
  OAI22_X1 U20326 ( .A1(n17088), .A2(n17087), .B1(n17336), .B2(n17381), .ZN(
        P3_U2678) );
  AOI21_X1 U20327 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17336), .A(n17097), .ZN(
        n17090) );
  XNOR2_X1 U20328 ( .A(n17089), .B(n17093), .ZN(n17386) );
  OAI22_X1 U20329 ( .A1(n17091), .A2(n17090), .B1(n17336), .B2(n17386), .ZN(
        P3_U2679) );
  INV_X1 U20330 ( .A(n17092), .ZN(n17111) );
  AOI21_X1 U20331 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17336), .A(n17111), .ZN(
        n17096) );
  OAI21_X1 U20332 ( .B1(n17095), .B2(n17094), .A(n17093), .ZN(n17391) );
  OAI22_X1 U20333 ( .A1(n17097), .A2(n17096), .B1(n17324), .B2(n17391), .ZN(
        P3_U2680) );
  AOI21_X1 U20334 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17336), .A(n17098), .ZN(
        n17110) );
  AOI22_X1 U20335 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17108) );
  AOI22_X1 U20336 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U20337 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9810), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17106) );
  OAI22_X1 U20338 ( .A1(n9858), .A2(n18582), .B1(n17307), .B2(n18345), .ZN(
        n17104) );
  AOI22_X1 U20339 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11392), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20340 ( .A1(n11309), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20341 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17100) );
  NAND2_X1 U20342 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n17099) );
  NAND4_X1 U20343 ( .A1(n17102), .A2(n17101), .A3(n17100), .A4(n17099), .ZN(
        n17103) );
  AOI211_X1 U20344 ( .C1(n17298), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17104), .B(n17103), .ZN(n17105) );
  NAND4_X1 U20345 ( .A1(n17108), .A2(n17107), .A3(n17106), .A4(n17105), .ZN(
        n17392) );
  INV_X1 U20346 ( .A(n17392), .ZN(n17109) );
  OAI22_X1 U20347 ( .A1(n17111), .A2(n17110), .B1(n17109), .B2(n17336), .ZN(
        P3_U2681) );
  NOR2_X1 U20348 ( .A1(n17341), .A2(n17112), .ZN(n17140) );
  AOI22_X1 U20349 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17113) );
  OAI21_X1 U20350 ( .B1(n11376), .B2(n17114), .A(n17113), .ZN(n17126) );
  AOI22_X1 U20351 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11392), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U20352 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9810), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17115) );
  OAI21_X1 U20353 ( .B1(n17172), .B2(n17116), .A(n17115), .ZN(n17122) );
  AOI22_X1 U20354 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20355 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17118) );
  OAI211_X1 U20356 ( .C1(n13764), .C2(n17120), .A(n17119), .B(n17118), .ZN(
        n17121) );
  AOI211_X1 U20357 ( .C1(n17276), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17122), .B(n17121), .ZN(n17123) );
  OAI211_X1 U20358 ( .C1(n17307), .C2(n18340), .A(n17124), .B(n17123), .ZN(
        n17125) );
  AOI211_X1 U20359 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n17126), .B(n17125), .ZN(n17399) );
  INV_X1 U20360 ( .A(n17399), .ZN(n17127) );
  AOI22_X1 U20361 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17140), .B1(n17341), 
        .B2(n17127), .ZN(n17128) );
  OAI21_X1 U20362 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17129), .A(n17128), .ZN(
        P3_U2682) );
  AOI22_X1 U20363 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17139) );
  INV_X1 U20364 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18388) );
  AOI22_X1 U20365 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20366 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17130) );
  OAI211_X1 U20367 ( .C1(n11489), .C2(n18388), .A(n17131), .B(n17130), .ZN(
        n17137) );
  AOI22_X1 U20368 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20369 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20370 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17133) );
  NAND2_X1 U20371 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n17132) );
  NAND4_X1 U20372 ( .A1(n17135), .A2(n17134), .A3(n17133), .A4(n17132), .ZN(
        n17136) );
  AOI211_X1 U20373 ( .C1(n17276), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17137), .B(n17136), .ZN(n17138) );
  OAI211_X1 U20374 ( .C1(n17307), .C2(n18335), .A(n17139), .B(n17138), .ZN(
        n17403) );
  INV_X1 U20375 ( .A(n17403), .ZN(n17143) );
  OAI21_X1 U20376 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17141), .A(n17140), .ZN(
        n17142) );
  OAI21_X1 U20377 ( .B1(n17143), .B2(n17324), .A(n17142), .ZN(P3_U2683) );
  AOI22_X1 U20378 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17144) );
  OAI21_X1 U20379 ( .B1(n17145), .B2(n17257), .A(n17144), .ZN(n17155) );
  AOI22_X1 U20380 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9804), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17153) );
  OAI22_X1 U20381 ( .A1(n11376), .A2(n17146), .B1(n17307), .B2(n18330), .ZN(
        n17151) );
  AOI22_X1 U20382 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20383 ( .A1(n11309), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20384 ( .A1(n17276), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17147) );
  NAND3_X1 U20385 ( .A1(n17149), .A2(n17148), .A3(n17147), .ZN(n17150) );
  AOI211_X1 U20386 ( .C1(n17117), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n17151), .B(n17150), .ZN(n17152) );
  OAI211_X1 U20387 ( .C1(n11489), .C2(n18385), .A(n17153), .B(n17152), .ZN(
        n17154) );
  AOI211_X1 U20388 ( .C1(n11331), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17155), .B(n17154), .ZN(n17413) );
  INV_X1 U20389 ( .A(n17156), .ZN(n17158) );
  OAI33_X1 U20390 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17393), .A3(n17158), 
        .B1(n17157), .B2(n17341), .B3(n17156), .ZN(n17159) );
  INV_X1 U20391 ( .A(n17159), .ZN(n17160) );
  OAI21_X1 U20392 ( .B1(n17413), .B2(n17324), .A(n17160), .ZN(P3_U2684) );
  AOI22_X1 U20393 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17161) );
  OAI21_X1 U20394 ( .B1(n10327), .B2(n17162), .A(n17161), .ZN(n17174) );
  INV_X1 U20395 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17171) );
  AOI22_X1 U20396 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17170) );
  AOI22_X1 U20397 ( .A1(n17276), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9809), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17163) );
  OAI21_X1 U20398 ( .B1(n17307), .B2(n18325), .A(n17163), .ZN(n17168) );
  INV_X1 U20399 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20400 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11518), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20401 ( .A1(n11309), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11331), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17164) );
  OAI211_X1 U20402 ( .C1(n10328), .C2(n17166), .A(n17165), .B(n17164), .ZN(
        n17167) );
  AOI211_X1 U20403 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17168), .B(n17167), .ZN(n17169) );
  OAI211_X1 U20404 ( .C1(n17172), .C2(n17171), .A(n17170), .B(n17169), .ZN(
        n17173) );
  AOI211_X1 U20405 ( .C1(n9808), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n17174), .B(n17173), .ZN(n17417) );
  INV_X1 U20406 ( .A(n17192), .ZN(n17175) );
  OAI33_X1 U20407 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17393), .A3(n17192), 
        .B1(n17176), .B2(n17341), .B3(n17175), .ZN(n17177) );
  INV_X1 U20408 ( .A(n17177), .ZN(n17178) );
  OAI21_X1 U20409 ( .B1(n17417), .B2(n17324), .A(n17178), .ZN(P3_U2685) );
  AOI22_X1 U20410 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17179) );
  OAI21_X1 U20411 ( .B1(n11376), .B2(n17301), .A(n17179), .ZN(n17190) );
  AOI22_X1 U20412 ( .A1(n11378), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20413 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17180) );
  OAI21_X1 U20414 ( .B1(n17296), .B2(n17181), .A(n17180), .ZN(n17186) );
  AOI22_X1 U20415 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U20416 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17182) );
  OAI211_X1 U20417 ( .C1(n10328), .C2(n17184), .A(n17183), .B(n17182), .ZN(
        n17185) );
  AOI211_X1 U20418 ( .C1(n9809), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n17186), .B(n17185), .ZN(n17187) );
  OAI211_X1 U20419 ( .C1(n11340), .C2(n18723), .A(n17188), .B(n17187), .ZN(
        n17189) );
  AOI211_X1 U20420 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n17190), .B(n17189), .ZN(n17423) );
  OAI211_X1 U20421 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n17193), .A(n17192), .B(
        n17336), .ZN(n17194) );
  OAI21_X1 U20422 ( .B1(n17423), .B2(n17324), .A(n17194), .ZN(P3_U2686) );
  AOI22_X1 U20423 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17195) );
  OAI21_X1 U20424 ( .B1(n11340), .B2(n18716), .A(n17195), .ZN(n17205) );
  AOI22_X1 U20425 ( .A1(n11309), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20426 ( .A1(n17276), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17196) );
  OAI21_X1 U20427 ( .B1(n17307), .B2(n18317), .A(n17196), .ZN(n17200) );
  INV_X1 U20428 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18378) );
  AOI22_X1 U20429 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U20430 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17197) );
  OAI211_X1 U20431 ( .C1(n11489), .C2(n18378), .A(n17198), .B(n17197), .ZN(
        n17199) );
  AOI211_X1 U20432 ( .C1(n9804), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17200), .B(n17199), .ZN(n17201) );
  OAI211_X1 U20433 ( .C1(n17172), .C2(n17203), .A(n17202), .B(n17201), .ZN(
        n17204) );
  AOI211_X1 U20434 ( .C1(n11331), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n17205), .B(n17204), .ZN(n17430) );
  NAND3_X1 U20435 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17324), .A3(n17221), 
        .ZN(n17208) );
  NAND4_X1 U20436 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17227), .A4(n17206), .ZN(n17207) );
  OAI211_X1 U20437 ( .C1(n17430), .C2(n17336), .A(n17208), .B(n17207), .ZN(
        P3_U2687) );
  AOI22_X1 U20438 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17243), .B1(
        n11331), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20439 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n15791), .ZN(n17209) );
  OAI21_X1 U20440 ( .B1(n11376), .B2(n18397), .A(n17209), .ZN(n17216) );
  OAI22_X1 U20441 ( .A1(n13764), .A2(n18354), .B1(n18771), .B2(n17307), .ZN(
        n17210) );
  AOI21_X1 U20442 ( .B1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17276), .A(
        n17210), .ZN(n17214) );
  AOI22_X1 U20443 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17293), .ZN(n17213) );
  AOI22_X1 U20444 ( .A1(n11309), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20445 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n9809), .B1(n9810), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17211) );
  NAND4_X1 U20446 ( .A1(n17214), .A2(n17213), .A3(n17212), .A4(n17211), .ZN(
        n17215) );
  AOI211_X1 U20447 ( .C1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .C2(n17297), .A(
        n17216), .B(n17215), .ZN(n17217) );
  OAI211_X1 U20448 ( .C1(n17220), .C2(n17219), .A(n17218), .B(n17217), .ZN(
        n17434) );
  INV_X1 U20449 ( .A(n17434), .ZN(n17224) );
  OAI211_X1 U20450 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17222), .A(n17221), .B(
        n17324), .ZN(n17223) );
  OAI21_X1 U20451 ( .B1(n17224), .B2(n17324), .A(n17223), .ZN(P3_U2688) );
  AOI22_X1 U20452 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17227), .B1(n17226), 
        .B2(n17225), .ZN(n17239) );
  AOI22_X1 U20453 ( .A1(n17276), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20454 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20455 ( .A1(n17297), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17229) );
  OAI211_X1 U20456 ( .C1(n13764), .C2(n18345), .A(n17230), .B(n17229), .ZN(
        n17236) );
  AOI22_X1 U20457 ( .A1(n11309), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20458 ( .A1(n9808), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20459 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17232) );
  NAND2_X1 U20460 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n17231) );
  NAND4_X1 U20461 ( .A1(n17234), .A2(n17233), .A3(n17232), .A4(n17231), .ZN(
        n17235) );
  AOI211_X1 U20462 ( .C1(n9809), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17236), .B(n17235), .ZN(n17237) );
  OAI211_X1 U20463 ( .C1(n17307), .C2(n18759), .A(n17238), .B(n17237), .ZN(
        n17439) );
  MUX2_X1 U20464 ( .A(n17239), .B(n17439), .S(n17341), .Z(P3_U2689) );
  AOI22_X1 U20465 ( .A1(n11309), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11518), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17240) );
  OAI21_X1 U20466 ( .B1(n17242), .B2(n17241), .A(n17240), .ZN(n17254) );
  AOI22_X1 U20467 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11378), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17252) );
  INV_X1 U20468 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17245) );
  AOI22_X1 U20469 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9809), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17244) );
  OAI21_X1 U20470 ( .B1(n17296), .B2(n17245), .A(n17244), .ZN(n17250) );
  AOI22_X1 U20471 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20472 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17246) );
  OAI211_X1 U20473 ( .C1(n10328), .C2(n17248), .A(n17247), .B(n17246), .ZN(
        n17249) );
  AOI211_X1 U20474 ( .C1(n9804), .C2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n17250), .B(n17249), .ZN(n17251) );
  OAI211_X1 U20475 ( .C1(n17291), .C2(n18575), .A(n17252), .B(n17251), .ZN(
        n17253) );
  AOI211_X1 U20476 ( .C1(n9808), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n17254), .B(n17253), .ZN(n17448) );
  NAND3_X1 U20477 ( .A1(n17256), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17324), 
        .ZN(n17255) );
  OAI221_X1 U20478 ( .B1(n17256), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17336), 
        .C2(n17448), .A(n17255), .ZN(P3_U2691) );
  AOI22_X1 U20479 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11392), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U20480 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17267) );
  OAI22_X1 U20481 ( .A1(n11340), .A2(n17258), .B1(n10327), .B2(n17257), .ZN(
        n17265) );
  AOI22_X1 U20482 ( .A1(n17276), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U20483 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U20484 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17259) );
  OAI211_X1 U20485 ( .C1(n13764), .C2(n18330), .A(n17260), .B(n17259), .ZN(
        n17261) );
  AOI21_X1 U20486 ( .B1(n9809), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(n17261), .ZN(n17262) );
  OAI211_X1 U20487 ( .C1(n17307), .C2(n18737), .A(n17263), .B(n17262), .ZN(
        n17264) );
  AOI211_X1 U20488 ( .C1(n17243), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n17265), .B(n17264), .ZN(n17266) );
  NAND3_X1 U20489 ( .A1(n17268), .A2(n17267), .A3(n17266), .ZN(n17452) );
  INV_X1 U20490 ( .A(n17452), .ZN(n17273) );
  NOR2_X1 U20491 ( .A1(n13776), .A2(n17269), .ZN(n17311) );
  NAND2_X1 U20492 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17311), .ZN(n17310) );
  NOR2_X1 U20493 ( .A1(n17270), .A2(n17310), .ZN(n17289) );
  OAI21_X1 U20494 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17289), .A(n17324), .ZN(
        n17271) );
  OAI22_X1 U20495 ( .A1(n17273), .A2(n17324), .B1(n17272), .B2(n17271), .ZN(
        P3_U2692) );
  AOI22_X1 U20496 ( .A1(n11331), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17117), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17274) );
  OAI21_X1 U20497 ( .B1(n10327), .B2(n17275), .A(n17274), .ZN(n17286) );
  AOI22_X1 U20498 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15791), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17284) );
  INV_X1 U20499 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17278) );
  AOI22_X1 U20500 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17276), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17277) );
  OAI21_X1 U20501 ( .B1(n11489), .B2(n17278), .A(n17277), .ZN(n17282) );
  AOI22_X1 U20502 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14282), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20503 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17279) );
  OAI211_X1 U20504 ( .C1(n13764), .C2(n18325), .A(n17280), .B(n17279), .ZN(
        n17281) );
  AOI211_X1 U20505 ( .C1(n9810), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17282), .B(n17281), .ZN(n17283) );
  OAI211_X1 U20506 ( .C1(n17307), .C2(n18730), .A(n17284), .B(n17283), .ZN(
        n17285) );
  AOI211_X1 U20507 ( .C1(n9808), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n17286), .B(n17285), .ZN(n17455) );
  INV_X1 U20508 ( .A(n17310), .ZN(n17287) );
  OAI21_X1 U20509 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17287), .A(n17324), .ZN(
        n17288) );
  OAI22_X1 U20510 ( .A1(n17455), .A2(n17336), .B1(n17289), .B2(n17288), .ZN(
        P3_U2693) );
  AOI22_X1 U20511 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11331), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17290) );
  OAI21_X1 U20512 ( .B1(n17291), .B2(n18568), .A(n17290), .ZN(n17309) );
  AOI22_X1 U20513 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17306) );
  INV_X1 U20514 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20515 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9809), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17294) );
  OAI21_X1 U20516 ( .B1(n17296), .B2(n17295), .A(n17294), .ZN(n17303) );
  AOI22_X1 U20517 ( .A1(n17117), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17297), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20518 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17299) );
  OAI211_X1 U20519 ( .C1(n10328), .C2(n17301), .A(n17300), .B(n17299), .ZN(
        n17302) );
  AOI211_X1 U20520 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n17303), .B(n17302), .ZN(n17305) );
  OAI211_X1 U20521 ( .C1(n17307), .C2(n18723), .A(n17306), .B(n17305), .ZN(
        n17308) );
  AOI211_X1 U20522 ( .C1(n9808), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n17309), .B(n17308), .ZN(n17461) );
  OAI21_X1 U20523 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17311), .A(n17310), .ZN(
        n17312) );
  AOI22_X1 U20524 ( .A1(n17341), .A2(n17461), .B1(n17312), .B2(n17324), .ZN(
        P3_U2694) );
  OAI33_X1 U20525 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17393), .A3(n17315), .B1(
        n17314), .B2(n17341), .B3(n17313), .ZN(n17316) );
  AOI21_X1 U20526 ( .B1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17341), .A(
        n17316), .ZN(n17317) );
  INV_X1 U20527 ( .A(n17317), .ZN(P3_U2696) );
  AOI21_X1 U20528 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17322), .A(n17341), .ZN(
        n17321) );
  AOI22_X1 U20529 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17341), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17321), .ZN(n17320) );
  INV_X1 U20530 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17318) );
  NAND4_X1 U20531 ( .A1(n18350), .A2(P3_EBX_REG_5__SCAN_IN), .A3(n17322), .A4(
        n17318), .ZN(n17319) );
  NAND2_X1 U20532 ( .A1(n17320), .A2(n17319), .ZN(P3_U2697) );
  OAI21_X1 U20533 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17322), .A(n17321), .ZN(
        n17323) );
  OAI21_X1 U20534 ( .B1(n17324), .B2(n18340), .A(n17323), .ZN(P3_U2698) );
  INV_X1 U20535 ( .A(n17338), .ZN(n17340) );
  NAND2_X1 U20536 ( .A1(n17325), .A2(n17340), .ZN(n17329) );
  NOR2_X1 U20537 ( .A1(n17326), .A2(n17329), .ZN(n17331) );
  AOI21_X1 U20538 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17336), .A(n17331), .ZN(
        n17327) );
  OAI22_X1 U20539 ( .A1(n17328), .A2(n17327), .B1(n18335), .B2(n17336), .ZN(
        P3_U2699) );
  INV_X1 U20540 ( .A(n17329), .ZN(n17334) );
  AOI21_X1 U20541 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17336), .A(n17334), .ZN(
        n17330) );
  OAI22_X1 U20542 ( .A1(n17331), .A2(n17330), .B1(n18330), .B2(n17336), .ZN(
        P3_U2700) );
  INV_X1 U20543 ( .A(n17332), .ZN(n17333) );
  AOI221_X1 U20544 ( .B1(n17333), .B2(n17344), .C1(n17393), .C2(n17344), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17335) );
  AOI211_X1 U20545 ( .C1(n17341), .C2(n18325), .A(n17335), .B(n17334), .ZN(
        P3_U2701) );
  OAI222_X1 U20546 ( .A1(n17339), .A2(n17338), .B1(n17337), .B2(n17344), .C1(
        n18320), .C2(n17336), .ZN(P3_U2702) );
  AOI22_X1 U20547 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17341), .B1(
        n17340), .B2(n17343), .ZN(n17342) );
  OAI21_X1 U20548 ( .B1(n17344), .B2(n17343), .A(n17342), .ZN(P3_U2703) );
  INV_X1 U20549 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17566) );
  INV_X1 U20550 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17562) );
  INV_X1 U20551 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17556) );
  INV_X1 U20552 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17609) );
  NAND2_X1 U20553 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17487) );
  NAND4_X1 U20554 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n17345) );
  NOR2_X1 U20555 ( .A1(n17487), .A2(n17345), .ZN(n17469) );
  NAND3_X1 U20556 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(n17469), .ZN(n17431) );
  INV_X1 U20557 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17590) );
  NAND2_X1 U20558 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .ZN(n17437) );
  NAND4_X1 U20559 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n17346)
         );
  NOR3_X1 U20560 ( .A1(n17590), .A2(n17437), .A3(n17346), .ZN(n17432) );
  INV_X1 U20561 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17554) );
  INV_X1 U20562 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17552) );
  NOR2_X1 U20563 ( .A1(n17554), .A2(n17552), .ZN(n17347) );
  NAND4_X1 U20564 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n17347), .ZN(n17398) );
  NOR3_X2 U20565 ( .A1(n17556), .A2(n17426), .A3(n17398), .ZN(n17388) );
  NAND2_X1 U20566 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17388), .ZN(n17387) );
  NOR2_X2 U20567 ( .A1(n17562), .A2(n17382), .ZN(n17377) );
  NAND2_X1 U20568 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17377), .ZN(n17373) );
  INV_X1 U20569 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17572) );
  OR2_X1 U20570 ( .A1(n9861), .A2(n17572), .ZN(n17350) );
  NAND2_X1 U20571 ( .A1(n17488), .A2(n9861), .ZN(n17355) );
  OAI21_X1 U20572 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17486), .A(n17355), .ZN(
        n17348) );
  AOI22_X1 U20573 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17424), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17348), .ZN(n17349) );
  OAI21_X1 U20574 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17350), .A(n17349), .ZN(
        P3_U2704) );
  OAI22_X1 U20575 ( .A1(n17352), .A2(n17490), .B1(n19358), .B2(n17407), .ZN(
        n17353) );
  AOI21_X1 U20576 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17425), .A(n17353), .ZN(
        n17354) );
  OAI221_X1 U20577 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n9861), .C1(n17572), 
        .C2(n17355), .A(n17354), .ZN(P3_U2705) );
  AOI22_X1 U20578 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17424), .ZN(n17358) );
  OAI211_X1 U20579 ( .C1(n17356), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17488), .B(
        n9861), .ZN(n17357) );
  OAI211_X1 U20580 ( .C1(n17359), .C2(n17490), .A(n17358), .B(n17357), .ZN(
        P3_U2706) );
  AOI22_X1 U20581 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17425), .B1(n17497), .B2(
        n17360), .ZN(n17363) );
  OAI211_X1 U20582 ( .C1(n17368), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17488), .B(
        n17361), .ZN(n17362) );
  OAI211_X1 U20583 ( .C1(n17407), .C2(n17364), .A(n17363), .B(n17362), .ZN(
        P3_U2707) );
  OAI21_X1 U20584 ( .B1(n17367), .B2(n17366), .A(n17365), .ZN(n17372) );
  AOI22_X1 U20585 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17424), .ZN(n17371) );
  AOI211_X1 U20586 ( .C1(n17566), .C2(n17373), .A(n17368), .B(n17408), .ZN(
        n17369) );
  INV_X1 U20587 ( .A(n17369), .ZN(n17370) );
  OAI211_X1 U20588 ( .C1(n17372), .C2(n17490), .A(n17371), .B(n17370), .ZN(
        P3_U2708) );
  AOI22_X1 U20589 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17424), .ZN(n17375) );
  OAI211_X1 U20590 ( .C1(n17377), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17488), .B(
        n17373), .ZN(n17374) );
  OAI211_X1 U20591 ( .C1(n17376), .C2(n17490), .A(n17375), .B(n17374), .ZN(
        P3_U2709) );
  AOI22_X1 U20592 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17424), .ZN(n17380) );
  AOI211_X1 U20593 ( .C1(n17562), .C2(n17382), .A(n17377), .B(n17408), .ZN(
        n17378) );
  INV_X1 U20594 ( .A(n17378), .ZN(n17379) );
  OAI211_X1 U20595 ( .C1(n17381), .C2(n17490), .A(n17380), .B(n17379), .ZN(
        P3_U2710) );
  AOI22_X1 U20596 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17424), .ZN(n17385) );
  OAI211_X1 U20597 ( .C1(n17383), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17488), .B(
        n17382), .ZN(n17384) );
  OAI211_X1 U20598 ( .C1(n17386), .C2(n17490), .A(n17385), .B(n17384), .ZN(
        P3_U2711) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17424), .ZN(n17390) );
  OAI211_X1 U20600 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17388), .A(n17488), .B(
        n17387), .ZN(n17389) );
  OAI211_X1 U20601 ( .C1(n17391), .C2(n17490), .A(n17390), .B(n17389), .ZN(
        P3_U2712) );
  NOR2_X1 U20602 ( .A1(n17393), .A2(n17426), .ZN(n17420) );
  NAND2_X1 U20603 ( .A1(n17420), .A2(n17556), .ZN(n17397) );
  AOI22_X1 U20604 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17424), .B1(n17497), .B2(
        n17392), .ZN(n17396) );
  INV_X1 U20605 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17550) );
  INV_X1 U20606 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17546) );
  NAND2_X1 U20607 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17418), .ZN(n17414) );
  NAND2_X1 U20608 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17409), .ZN(n17404) );
  NAND2_X1 U20609 ( .A1(n17488), .A2(n17404), .ZN(n17402) );
  OAI21_X1 U20610 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17486), .A(n17402), .ZN(
        n17394) );
  AOI22_X1 U20611 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17425), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17394), .ZN(n17395) );
  OAI211_X1 U20612 ( .C1(n17398), .C2(n17397), .A(n17396), .B(n17395), .ZN(
        P3_U2713) );
  INV_X1 U20613 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19351) );
  OAI22_X1 U20614 ( .A1(n17399), .A2(n17490), .B1(n19351), .B2(n17407), .ZN(
        n17400) );
  AOI21_X1 U20615 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17425), .A(n17400), .ZN(
        n17401) );
  OAI221_X1 U20616 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17404), .C1(n17554), 
        .C2(n17402), .A(n17401), .ZN(P3_U2714) );
  AOI22_X1 U20617 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17425), .B1(n17497), .B2(
        n17403), .ZN(n17406) );
  OAI211_X1 U20618 ( .C1(n17409), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17488), .B(
        n17404), .ZN(n17405) );
  OAI211_X1 U20619 ( .C1(n17407), .C2(n19345), .A(n17406), .B(n17405), .ZN(
        P3_U2715) );
  AOI22_X1 U20620 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17424), .ZN(n17412) );
  AOI211_X1 U20621 ( .C1(n17550), .C2(n17414), .A(n17409), .B(n17408), .ZN(
        n17410) );
  INV_X1 U20622 ( .A(n17410), .ZN(n17411) );
  OAI211_X1 U20623 ( .C1(n17413), .C2(n17490), .A(n17412), .B(n17411), .ZN(
        P3_U2716) );
  AOI22_X1 U20624 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17424), .ZN(n17416) );
  OAI211_X1 U20625 ( .C1(n17418), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17488), .B(
        n17414), .ZN(n17415) );
  OAI211_X1 U20626 ( .C1(n17417), .C2(n17490), .A(n17416), .B(n17415), .ZN(
        P3_U2717) );
  AOI22_X1 U20627 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17424), .ZN(n17422) );
  INV_X1 U20628 ( .A(n17418), .ZN(n17419) );
  OAI211_X1 U20629 ( .C1(n17420), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17488), .B(
        n17419), .ZN(n17421) );
  OAI211_X1 U20630 ( .C1(n17423), .C2(n17490), .A(n17422), .B(n17421), .ZN(
        P3_U2718) );
  AOI22_X1 U20631 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17425), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17424), .ZN(n17429) );
  OAI211_X1 U20632 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17427), .A(n17488), .B(
        n17426), .ZN(n17428) );
  OAI211_X1 U20633 ( .C1(n17430), .C2(n17490), .A(n17429), .B(n17428), .ZN(
        P3_U2719) );
  NAND2_X1 U20634 ( .A1(n17432), .A2(n17473), .ZN(n17436) );
  NAND2_X1 U20635 ( .A1(n17488), .A2(n17433), .ZN(n17441) );
  AOI22_X1 U20636 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17498), .B1(n17497), .B2(
        n17434), .ZN(n17435) );
  OAI221_X1 U20637 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17436), .C1(n17609), 
        .C2(n17441), .A(n17435), .ZN(P3_U2720) );
  NAND2_X1 U20638 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n17438) );
  NAND2_X1 U20639 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17473), .ZN(n17459) );
  NOR2_X1 U20640 ( .A1(n17437), .A2(n17459), .ZN(n17447) );
  INV_X1 U20641 ( .A(n17447), .ZN(n17454) );
  NOR2_X1 U20642 ( .A1(n17438), .A2(n17454), .ZN(n17450) );
  NAND2_X1 U20643 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17450), .ZN(n17442) );
  INV_X1 U20644 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17604) );
  AOI22_X1 U20645 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17498), .B1(n17497), .B2(
        n17439), .ZN(n17440) );
  OAI221_X1 U20646 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17442), .C1(n17604), 
        .C2(n17441), .A(n17440), .ZN(P3_U2721) );
  INV_X1 U20647 ( .A(n17442), .ZN(n17445) );
  AOI21_X1 U20648 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17488), .A(n17450), .ZN(
        n17444) );
  OAI222_X1 U20649 ( .A1(n17493), .A2(n17446), .B1(n17445), .B2(n17444), .C1(
        n17490), .C2(n17443), .ZN(P3_U2722) );
  AOI22_X1 U20650 ( .A1(n17447), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17488), .ZN(n17449) );
  OAI222_X1 U20651 ( .A1(n17493), .A2(n17451), .B1(n17450), .B2(n17449), .C1(
        n17490), .C2(n17448), .ZN(P3_U2723) );
  INV_X1 U20652 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17596) );
  NAND2_X1 U20653 ( .A1(n17488), .A2(n17454), .ZN(n17457) );
  AOI22_X1 U20654 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17498), .B1(n17497), .B2(
        n17452), .ZN(n17453) );
  OAI221_X1 U20655 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17454), .C1(n17596), 
        .C2(n17457), .A(n17453), .ZN(P3_U2724) );
  INV_X1 U20656 ( .A(n17459), .ZN(n17460) );
  AOI21_X1 U20657 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17460), .A(
        P3_EAX_REG_10__SCAN_IN), .ZN(n17456) );
  OAI222_X1 U20658 ( .A1(n17493), .A2(n17458), .B1(n17457), .B2(n17456), .C1(
        n17490), .C2(n17455), .ZN(P3_U2725) );
  INV_X1 U20659 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17592) );
  NOR2_X1 U20660 ( .A1(n17592), .A2(n17459), .ZN(n17463) );
  AOI21_X1 U20661 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17488), .A(n17460), .ZN(
        n17462) );
  OAI222_X1 U20662 ( .A1(n17493), .A2(n17464), .B1(n17463), .B2(n17462), .C1(
        n17490), .C2(n17461), .ZN(P3_U2726) );
  AOI22_X1 U20663 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17498), .B1(n17497), .B2(
        n17465), .ZN(n17468) );
  OAI221_X1 U20664 ( .B1(n17466), .B2(P3_EAX_REG_8__SCAN_IN), .C1(n9981), .C2(
        n17590), .A(n17488), .ZN(n17467) );
  NAND2_X1 U20665 ( .A1(n17468), .A2(n17467), .ZN(P3_U2727) );
  INV_X1 U20666 ( .A(n17469), .ZN(n17470) );
  NOR2_X1 U20667 ( .A1(n17470), .A2(n17486), .ZN(n17478) );
  AOI22_X1 U20668 ( .A1(n17478), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17488), .ZN(n17472) );
  OAI222_X1 U20669 ( .A1(n17493), .A2(n18346), .B1(n17473), .B2(n17472), .C1(
        n17490), .C2(n17471), .ZN(P3_U2728) );
  AND2_X1 U20670 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17478), .ZN(n17475) );
  AOI21_X1 U20671 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17488), .A(n17478), .ZN(
        n17474) );
  OAI222_X1 U20672 ( .A1(n18341), .A2(n17493), .B1(n17475), .B2(n17474), .C1(
        n17490), .C2(n17902), .ZN(P3_U2729) );
  INV_X1 U20673 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17582) );
  INV_X1 U20674 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17578) );
  NOR3_X1 U20675 ( .A1(n17578), .A2(n17487), .A3(n17486), .ZN(n17492) );
  NAND2_X1 U20676 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17492), .ZN(n17479) );
  NOR2_X1 U20677 ( .A1(n17582), .A2(n17479), .ZN(n17482) );
  AOI21_X1 U20678 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17488), .A(n17482), .ZN(
        n17477) );
  OAI222_X1 U20679 ( .A1(n18336), .A2(n17493), .B1(n17478), .B2(n17477), .C1(
        n17490), .C2(n17476), .ZN(P3_U2730) );
  INV_X1 U20680 ( .A(n17479), .ZN(n17485) );
  AOI21_X1 U20681 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17488), .A(n17485), .ZN(
        n17481) );
  OAI222_X1 U20682 ( .A1(n18331), .A2(n17493), .B1(n17482), .B2(n17481), .C1(
        n17490), .C2(n17480), .ZN(P3_U2731) );
  AOI21_X1 U20683 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17488), .A(n17492), .ZN(
        n17484) );
  OAI222_X1 U20684 ( .A1(n18326), .A2(n17493), .B1(n17485), .B2(n17484), .C1(
        n17490), .C2(n17483), .ZN(P3_U2732) );
  NOR2_X1 U20685 ( .A1(n17487), .A2(n17486), .ZN(n17501) );
  AOI21_X1 U20686 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17488), .A(n17501), .ZN(
        n17491) );
  OAI222_X1 U20687 ( .A1(n18321), .A2(n17493), .B1(n17492), .B2(n17491), .C1(
        n17490), .C2(n17489), .ZN(P3_U2733) );
  NOR2_X1 U20688 ( .A1(n17494), .A2(n17574), .ZN(n17495) );
  OAI21_X1 U20689 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17495), .A(n17488), .ZN(
        n17500) );
  AOI22_X1 U20690 ( .A1(n17498), .A2(BUF2_REG_1__SCAN_IN), .B1(n17497), .B2(
        n17496), .ZN(n17499) );
  OAI21_X1 U20691 ( .B1(n17501), .B2(n17500), .A(n17499), .ZN(P3_U2734) );
  NOR2_X2 U20692 ( .A1(n18966), .A2(n17980), .ZN(n19001) );
  NOR2_X4 U20693 ( .A1(n19001), .A2(n17521), .ZN(n17518) );
  AND2_X1 U20694 ( .A1(n17518), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AOI22_X1 U20695 ( .A1(n19001), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17518), .ZN(n17504) );
  OAI21_X1 U20696 ( .B1(n17572), .B2(n17520), .A(n17504), .ZN(P3_U2737) );
  INV_X1 U20697 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17570) );
  AOI22_X1 U20698 ( .A1(n19001), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17505) );
  OAI21_X1 U20699 ( .B1(n17570), .B2(n17520), .A(n17505), .ZN(P3_U2738) );
  INV_X1 U20700 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17568) );
  AOI22_X1 U20701 ( .A1(n19001), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17506) );
  OAI21_X1 U20702 ( .B1(n17568), .B2(n17520), .A(n17506), .ZN(P3_U2739) );
  AOI22_X1 U20703 ( .A1(n19001), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17507) );
  OAI21_X1 U20704 ( .B1(n17566), .B2(n17520), .A(n17507), .ZN(P3_U2740) );
  INV_X1 U20705 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17564) );
  AOI22_X1 U20706 ( .A1(n19001), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17508) );
  OAI21_X1 U20707 ( .B1(n17564), .B2(n17520), .A(n17508), .ZN(P3_U2741) );
  AOI22_X1 U20708 ( .A1(n19001), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17509) );
  OAI21_X1 U20709 ( .B1(n17562), .B2(n17520), .A(n17509), .ZN(P3_U2742) );
  INV_X1 U20710 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17560) );
  AOI22_X1 U20711 ( .A1(n19001), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17510) );
  OAI21_X1 U20712 ( .B1(n17560), .B2(n17520), .A(n17510), .ZN(P3_U2743) );
  INV_X1 U20713 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17558) );
  CLKBUF_X1 U20714 ( .A(n19001), .Z(n17537) );
  AOI22_X1 U20715 ( .A1(n17537), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17511) );
  OAI21_X1 U20716 ( .B1(n17558), .B2(n17520), .A(n17511), .ZN(P3_U2744) );
  AOI22_X1 U20717 ( .A1(n17537), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17512) );
  OAI21_X1 U20718 ( .B1(n17556), .B2(n17520), .A(n17512), .ZN(P3_U2745) );
  AOI22_X1 U20719 ( .A1(n17537), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17513) );
  OAI21_X1 U20720 ( .B1(n17554), .B2(n17520), .A(n17513), .ZN(P3_U2746) );
  AOI22_X1 U20721 ( .A1(n17537), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17514) );
  OAI21_X1 U20722 ( .B1(n17552), .B2(n17520), .A(n17514), .ZN(P3_U2747) );
  AOI22_X1 U20723 ( .A1(n17537), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17515) );
  OAI21_X1 U20724 ( .B1(n17550), .B2(n17520), .A(n17515), .ZN(P3_U2748) );
  INV_X1 U20725 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17548) );
  AOI22_X1 U20726 ( .A1(n17537), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17516) );
  OAI21_X1 U20727 ( .B1(n17548), .B2(n17520), .A(n17516), .ZN(P3_U2749) );
  AOI22_X1 U20728 ( .A1(n17537), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17517) );
  OAI21_X1 U20729 ( .B1(n17546), .B2(n17520), .A(n17517), .ZN(P3_U2750) );
  INV_X1 U20730 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17544) );
  AOI22_X1 U20731 ( .A1(n17537), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17519) );
  OAI21_X1 U20732 ( .B1(n17544), .B2(n17520), .A(n17519), .ZN(P3_U2751) );
  AOI22_X1 U20733 ( .A1(n17537), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17522) );
  OAI21_X1 U20734 ( .B1(n17609), .B2(n17539), .A(n17522), .ZN(P3_U2752) );
  AOI22_X1 U20735 ( .A1(n17537), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17523) );
  OAI21_X1 U20736 ( .B1(n17604), .B2(n17539), .A(n17523), .ZN(P3_U2753) );
  INV_X1 U20737 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17602) );
  AOI22_X1 U20738 ( .A1(n17537), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17524) );
  OAI21_X1 U20739 ( .B1(n17602), .B2(n17539), .A(n17524), .ZN(P3_U2754) );
  INV_X1 U20740 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17600) );
  AOI22_X1 U20741 ( .A1(n17537), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17525) );
  OAI21_X1 U20742 ( .B1(n17600), .B2(n17539), .A(n17525), .ZN(P3_U2755) );
  AOI22_X1 U20743 ( .A1(n17537), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17526) );
  OAI21_X1 U20744 ( .B1(n17596), .B2(n17539), .A(n17526), .ZN(P3_U2756) );
  INV_X1 U20745 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17594) );
  AOI22_X1 U20746 ( .A1(n17537), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17527) );
  OAI21_X1 U20747 ( .B1(n17594), .B2(n17539), .A(n17527), .ZN(P3_U2757) );
  AOI22_X1 U20748 ( .A1(n17537), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17528) );
  OAI21_X1 U20749 ( .B1(n17592), .B2(n17539), .A(n17528), .ZN(P3_U2758) );
  AOI22_X1 U20750 ( .A1(n17537), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17529) );
  OAI21_X1 U20751 ( .B1(n17590), .B2(n17539), .A(n17529), .ZN(P3_U2759) );
  INV_X1 U20752 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17588) );
  AOI22_X1 U20753 ( .A1(n17537), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17530) );
  OAI21_X1 U20754 ( .B1(n17588), .B2(n17539), .A(n17530), .ZN(P3_U2760) );
  INV_X1 U20755 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17586) );
  AOI22_X1 U20756 ( .A1(n17537), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17531) );
  OAI21_X1 U20757 ( .B1(n17586), .B2(n17539), .A(n17531), .ZN(P3_U2761) );
  INV_X1 U20758 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17584) );
  AOI22_X1 U20759 ( .A1(n17537), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17532) );
  OAI21_X1 U20760 ( .B1(n17584), .B2(n17539), .A(n17532), .ZN(P3_U2762) );
  AOI22_X1 U20761 ( .A1(n17537), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U20762 ( .B1(n17582), .B2(n17539), .A(n17533), .ZN(P3_U2763) );
  INV_X1 U20763 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17580) );
  AOI22_X1 U20764 ( .A1(n17537), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17534) );
  OAI21_X1 U20765 ( .B1(n17580), .B2(n17539), .A(n17534), .ZN(P3_U2764) );
  AOI22_X1 U20766 ( .A1(n17537), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U20767 ( .B1(n17578), .B2(n17539), .A(n17535), .ZN(P3_U2765) );
  INV_X1 U20768 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17576) );
  AOI22_X1 U20769 ( .A1(n17537), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17536) );
  OAI21_X1 U20770 ( .B1(n17576), .B2(n17539), .A(n17536), .ZN(P3_U2766) );
  AOI22_X1 U20771 ( .A1(n17537), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17518), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17538) );
  OAI21_X1 U20772 ( .B1(n17574), .B2(n17539), .A(n17538), .ZN(P3_U2767) );
  AOI22_X1 U20773 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17606), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17597), .ZN(n17543) );
  OAI21_X1 U20774 ( .B1(n17544), .B2(n17608), .A(n17543), .ZN(P3_U2768) );
  AOI22_X1 U20775 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17606), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17597), .ZN(n17545) );
  OAI21_X1 U20776 ( .B1(n17546), .B2(n17608), .A(n17545), .ZN(P3_U2769) );
  AOI22_X1 U20777 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17606), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17597), .ZN(n17547) );
  OAI21_X1 U20778 ( .B1(n17548), .B2(n17608), .A(n17547), .ZN(P3_U2770) );
  AOI22_X1 U20779 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17598), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17597), .ZN(n17549) );
  OAI21_X1 U20780 ( .B1(n17550), .B2(n17608), .A(n17549), .ZN(P3_U2771) );
  AOI22_X1 U20781 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17598), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17597), .ZN(n17551) );
  OAI21_X1 U20782 ( .B1(n17552), .B2(n17608), .A(n17551), .ZN(P3_U2772) );
  AOI22_X1 U20783 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17598), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17597), .ZN(n17553) );
  OAI21_X1 U20784 ( .B1(n17554), .B2(n17608), .A(n17553), .ZN(P3_U2773) );
  AOI22_X1 U20785 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17598), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17597), .ZN(n17555) );
  OAI21_X1 U20786 ( .B1(n17556), .B2(n17608), .A(n17555), .ZN(P3_U2774) );
  AOI22_X1 U20787 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17598), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17597), .ZN(n17557) );
  OAI21_X1 U20788 ( .B1(n17558), .B2(n17608), .A(n17557), .ZN(P3_U2775) );
  AOI22_X1 U20789 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17598), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17597), .ZN(n17559) );
  OAI21_X1 U20790 ( .B1(n17560), .B2(n17608), .A(n17559), .ZN(P3_U2776) );
  AOI22_X1 U20791 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17598), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17597), .ZN(n17561) );
  OAI21_X1 U20792 ( .B1(n17562), .B2(n17608), .A(n17561), .ZN(P3_U2777) );
  AOI22_X1 U20793 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17598), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17597), .ZN(n17563) );
  OAI21_X1 U20794 ( .B1(n17564), .B2(n17608), .A(n17563), .ZN(P3_U2778) );
  AOI22_X1 U20795 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17598), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17597), .ZN(n17565) );
  OAI21_X1 U20796 ( .B1(n17566), .B2(n17608), .A(n17565), .ZN(P3_U2779) );
  AOI22_X1 U20797 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17606), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17597), .ZN(n17567) );
  OAI21_X1 U20798 ( .B1(n17568), .B2(n17608), .A(n17567), .ZN(P3_U2780) );
  AOI22_X1 U20799 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17606), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17597), .ZN(n17569) );
  OAI21_X1 U20800 ( .B1(n17570), .B2(n17608), .A(n17569), .ZN(P3_U2781) );
  AOI22_X1 U20801 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17606), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17597), .ZN(n17571) );
  OAI21_X1 U20802 ( .B1(n17572), .B2(n17608), .A(n17571), .ZN(P3_U2782) );
  AOI22_X1 U20803 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17597), .ZN(n17573) );
  OAI21_X1 U20804 ( .B1(n17574), .B2(n17608), .A(n17573), .ZN(P3_U2783) );
  AOI22_X1 U20805 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17597), .ZN(n17575) );
  OAI21_X1 U20806 ( .B1(n17576), .B2(n17608), .A(n17575), .ZN(P3_U2784) );
  AOI22_X1 U20807 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17597), .ZN(n17577) );
  OAI21_X1 U20808 ( .B1(n17578), .B2(n17608), .A(n17577), .ZN(P3_U2785) );
  AOI22_X1 U20809 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17597), .ZN(n17579) );
  OAI21_X1 U20810 ( .B1(n17580), .B2(n17608), .A(n17579), .ZN(P3_U2786) );
  AOI22_X1 U20811 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17605), .ZN(n17581) );
  OAI21_X1 U20812 ( .B1(n17582), .B2(n17608), .A(n17581), .ZN(P3_U2787) );
  AOI22_X1 U20813 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17605), .ZN(n17583) );
  OAI21_X1 U20814 ( .B1(n17584), .B2(n17608), .A(n17583), .ZN(P3_U2788) );
  AOI22_X1 U20815 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17605), .ZN(n17585) );
  OAI21_X1 U20816 ( .B1(n17586), .B2(n17608), .A(n17585), .ZN(P3_U2789) );
  AOI22_X1 U20817 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17605), .ZN(n17587) );
  OAI21_X1 U20818 ( .B1(n17588), .B2(n17608), .A(n17587), .ZN(P3_U2790) );
  AOI22_X1 U20819 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17605), .ZN(n17589) );
  OAI21_X1 U20820 ( .B1(n17590), .B2(n17608), .A(n17589), .ZN(P3_U2791) );
  AOI22_X1 U20821 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17605), .ZN(n17591) );
  OAI21_X1 U20822 ( .B1(n17592), .B2(n17608), .A(n17591), .ZN(P3_U2792) );
  AOI22_X1 U20823 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17598), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17597), .ZN(n17593) );
  OAI21_X1 U20824 ( .B1(n17594), .B2(n17608), .A(n17593), .ZN(P3_U2793) );
  AOI22_X1 U20825 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17605), .ZN(n17595) );
  OAI21_X1 U20826 ( .B1(n17596), .B2(n17608), .A(n17595), .ZN(P3_U2794) );
  AOI22_X1 U20827 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17598), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17597), .ZN(n17599) );
  OAI21_X1 U20828 ( .B1(n17600), .B2(n17608), .A(n17599), .ZN(P3_U2795) );
  AOI22_X1 U20829 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17605), .ZN(n17601) );
  OAI21_X1 U20830 ( .B1(n17602), .B2(n17608), .A(n17601), .ZN(P3_U2796) );
  AOI22_X1 U20831 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17605), .ZN(n17603) );
  OAI21_X1 U20832 ( .B1(n17604), .B2(n17608), .A(n17603), .ZN(P3_U2797) );
  AOI22_X1 U20833 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17606), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17605), .ZN(n17607) );
  OAI21_X1 U20834 ( .B1(n17609), .B2(n17608), .A(n17607), .ZN(P3_U2798) );
  NOR4_X1 U20835 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17736), .A3(
        n17610), .A4(n17622), .ZN(n17612) );
  AOI211_X1 U20836 ( .C1(n17828), .C2(n17613), .A(n17612), .B(n17611), .ZN(
        n17626) );
  AOI211_X1 U20837 ( .C1(n17616), .C2(n17615), .A(n17614), .B(n17880), .ZN(
        n17617) );
  AOI21_X1 U20838 ( .B1(n10079), .B2(n17618), .A(n17617), .ZN(n17625) );
  INV_X1 U20839 ( .A(n17985), .ZN(n17619) );
  AOI22_X1 U20840 ( .A1(n17703), .A2(n17991), .B1(n17962), .B2(n17619), .ZN(
        n17648) );
  NAND2_X1 U20841 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17648), .ZN(
        n17634) );
  OAI211_X1 U20842 ( .C1(n17703), .C2(n17962), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17634), .ZN(n17624) );
  NOR3_X1 U20843 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17736), .A3(
        n17622), .ZN(n17632) );
  OAI21_X1 U20844 ( .B1(n17620), .B2(n17980), .A(n17979), .ZN(n17621) );
  AOI21_X1 U20845 ( .B1(n18855), .B2(n17622), .A(n17621), .ZN(n17645) );
  OAI21_X1 U20846 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17721), .A(
        n17645), .ZN(n17633) );
  OAI21_X1 U20847 ( .B1(n17632), .B2(n17633), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17623) );
  NAND4_X1 U20848 ( .A1(n17626), .A2(n17625), .A3(n17624), .A4(n17623), .ZN(
        P3_U2802) );
  NOR2_X1 U20849 ( .A1(n17628), .A2(n17627), .ZN(n17629) );
  XNOR2_X1 U20850 ( .A(n17629), .B(n17779), .ZN(n17998) );
  INV_X1 U20851 ( .A(n17828), .ZN(n17812) );
  OAI22_X1 U20852 ( .A1(n16515), .A2(n18927), .B1(n17812), .B2(n17630), .ZN(
        n17631) );
  AOI211_X1 U20853 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17633), .A(
        n17632), .B(n17631), .ZN(n17637) );
  OAI21_X1 U20854 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17635), .A(
        n17634), .ZN(n17636) );
  OAI211_X1 U20855 ( .C1(n17998), .C2(n17880), .A(n17637), .B(n17636), .ZN(
        P3_U2803) );
  OAI21_X1 U20856 ( .B1(n17639), .B2(n17649), .A(n17638), .ZN(n18001) );
  AOI21_X1 U20857 ( .B1(n17640), .B2(n18708), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17644) );
  INV_X1 U20858 ( .A(n17721), .ZN(n17642) );
  OAI21_X1 U20859 ( .B1(n17828), .B2(n17642), .A(n17641), .ZN(n17643) );
  NAND2_X1 U20860 ( .A1(n18296), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18002) );
  OAI211_X1 U20861 ( .C1(n17645), .C2(n17644), .A(n17643), .B(n18002), .ZN(
        n17646) );
  AOI21_X1 U20862 ( .B1(n17852), .B2(n18001), .A(n17646), .ZN(n17647) );
  OAI221_X1 U20863 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17650), 
        .C1(n17649), .C2(n17648), .A(n17647), .ZN(P3_U2804) );
  INV_X1 U20864 ( .A(n18131), .ZN(n17787) );
  NAND2_X1 U20865 ( .A1(n17787), .A2(n17672), .ZN(n18024) );
  NOR2_X1 U20866 ( .A1(n18024), .A2(n17676), .ZN(n17651) );
  XNOR2_X1 U20867 ( .A(n17651), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18022) );
  AND2_X1 U20868 ( .A1(n17653), .A2(n18708), .ZN(n17652) );
  AOI211_X1 U20869 ( .C1(n17693), .C2(n17685), .A(n17946), .B(n17652), .ZN(
        n17683) );
  OAI21_X1 U20870 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17721), .A(
        n17683), .ZN(n17667) );
  NOR2_X1 U20871 ( .A1(n17736), .A2(n17653), .ZN(n17669) );
  OAI211_X1 U20872 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17669), .B(n17654), .ZN(n17655) );
  NAND2_X1 U20873 ( .A1(n18296), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18006) );
  OAI211_X1 U20874 ( .C1(n17812), .C2(n17656), .A(n17655), .B(n18006), .ZN(
        n17657) );
  AOI21_X1 U20875 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17667), .A(
        n17657), .ZN(n17663) );
  NOR2_X1 U20876 ( .A1(n18010), .A2(n18124), .ZN(n17658) );
  XNOR2_X1 U20877 ( .A(n17658), .B(n18008), .ZN(n18019) );
  OAI21_X1 U20878 ( .B1(n17877), .B2(n17660), .A(n17659), .ZN(n17661) );
  XNOR2_X1 U20879 ( .A(n17661), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18018) );
  AOI22_X1 U20880 ( .A1(n17703), .A2(n18019), .B1(n17852), .B2(n18018), .ZN(
        n17662) );
  OAI211_X1 U20881 ( .C1(n17984), .C2(n18022), .A(n17663), .B(n17662), .ZN(
        P3_U2805) );
  AOI22_X1 U20882 ( .A1(n17703), .A2(n18026), .B1(n17962), .B2(n18024), .ZN(
        n17690) );
  AOI22_X1 U20883 ( .A1(n18296), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17828), 
        .B2(n17664), .ZN(n17665) );
  INV_X1 U20884 ( .A(n17665), .ZN(n17666) );
  AOI221_X1 U20885 ( .B1(n17669), .B2(n17668), .C1(n17667), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17666), .ZN(n17675) );
  OAI21_X1 U20886 ( .B1(n17671), .B2(n17676), .A(n17670), .ZN(n18034) );
  INV_X1 U20887 ( .A(n17672), .ZN(n17673) );
  NOR2_X1 U20888 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17673), .ZN(
        n18033) );
  AOI22_X1 U20889 ( .A1(n17852), .A2(n18034), .B1(n10079), .B2(n18033), .ZN(
        n17674) );
  OAI211_X1 U20890 ( .C1(n17690), .C2(n17676), .A(n17675), .B(n17674), .ZN(
        P3_U2806) );
  NAND2_X1 U20891 ( .A1(n18007), .A2(n10079), .ZN(n17692) );
  OAI22_X1 U20892 ( .A1(n17677), .A2(n17704), .B1(n17877), .B2(n18059), .ZN(
        n17678) );
  NOR2_X1 U20893 ( .A1(n17678), .A2(n17727), .ZN(n17679) );
  XNOR2_X1 U20894 ( .A(n17679), .B(n17691), .ZN(n18039) );
  AOI21_X1 U20895 ( .B1(n17680), .B2(n18708), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17682) );
  OAI22_X1 U20896 ( .A1(n17683), .A2(n17682), .B1(n17812), .B2(n17681), .ZN(
        n17688) );
  NAND2_X1 U20897 ( .A1(n17642), .A2(n17684), .ZN(n17686) );
  OAI22_X1 U20898 ( .A1(n16515), .A2(n18920), .B1(n17686), .B2(n17685), .ZN(
        n17687) );
  AOI211_X1 U20899 ( .C1(n17852), .C2(n18039), .A(n17688), .B(n17687), .ZN(
        n17689) );
  OAI221_X1 U20900 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17692), 
        .C1(n17691), .C2(n17690), .A(n17689), .ZN(P3_U2807) );
  AOI21_X1 U20901 ( .B1(n17694), .B2(n17693), .A(n17946), .ZN(n17695) );
  INV_X1 U20902 ( .A(n17695), .ZN(n17696) );
  AOI21_X1 U20903 ( .B1(n18855), .B2(n17698), .A(n17696), .ZN(n17723) );
  OAI21_X1 U20904 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17721), .A(
        n17723), .ZN(n17715) );
  AOI22_X1 U20905 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17715), .B1(
        n17828), .B2(n17697), .ZN(n17709) );
  NOR2_X1 U20906 ( .A1(n17736), .A2(n17698), .ZN(n17717) );
  AOI21_X1 U20907 ( .B1(n17716), .B2(n17699), .A(n9918), .ZN(n17700) );
  AOI22_X1 U20908 ( .A1(n18296), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17717), 
        .B2(n17700), .ZN(n17708) );
  NOR2_X1 U20909 ( .A1(n17703), .A2(n17962), .ZN(n17726) );
  NAND2_X1 U20910 ( .A1(n10007), .A2(n17702), .ZN(n18044) );
  INV_X1 U20911 ( .A(n18044), .ZN(n18048) );
  AOI22_X1 U20912 ( .A1(n17703), .A2(n18124), .B1(n17962), .B2(n18131), .ZN(
        n17777) );
  OAI21_X1 U20913 ( .B1(n17726), .B2(n18048), .A(n17777), .ZN(n17718) );
  OAI221_X1 U20914 ( .B1(n17704), .B2(n11422), .C1(n17704), .C2(n18048), .A(
        n11427), .ZN(n17705) );
  XNOR2_X1 U20915 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17705), .ZN(
        n18043) );
  AOI22_X1 U20916 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17718), .B1(
        n17852), .B2(n18043), .ZN(n17707) );
  NAND3_X1 U20917 ( .A1(n10079), .A2(n18048), .A3(n18059), .ZN(n17706) );
  NAND4_X1 U20918 ( .A1(n17709), .A2(n17708), .A3(n17707), .A4(n17706), .ZN(
        P3_U2808) );
  NAND3_X1 U20919 ( .A1(n17877), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17710), .ZN(n17731) );
  INV_X1 U20920 ( .A(n17752), .ZN(n17732) );
  OAI22_X1 U20921 ( .A1(n18062), .A2(n17731), .B1(n17732), .B2(n17711), .ZN(
        n17712) );
  XNOR2_X1 U20922 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17712), .ZN(
        n18069) );
  OAI22_X1 U20923 ( .A1(n16515), .A2(n18916), .B1(n17812), .B2(n17713), .ZN(
        n17714) );
  AOI221_X1 U20924 ( .B1(n17717), .B2(n17716), .C1(n17715), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17714), .ZN(n17720) );
  NOR2_X1 U20925 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18062), .ZN(
        n18061) );
  NAND2_X1 U20926 ( .A1(n10007), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18063) );
  NOR2_X1 U20927 ( .A1(n17778), .A2(n18063), .ZN(n17743) );
  AOI22_X1 U20928 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17718), .B1(
        n18061), .B2(n17743), .ZN(n17719) );
  OAI211_X1 U20929 ( .C1(n18069), .C2(n17880), .A(n17720), .B(n17719), .ZN(
        P3_U2809) );
  INV_X1 U20930 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18080) );
  NOR2_X1 U20931 ( .A1(n18080), .A2(n18063), .ZN(n18073) );
  NAND2_X1 U20932 ( .A1(n18073), .A2(n18050), .ZN(n18079) );
  AOI21_X1 U20933 ( .B1(n9926), .B2(n18708), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17722) );
  OAI22_X1 U20934 ( .A1(n17723), .A2(n17722), .B1(n16515), .B2(n18913), .ZN(
        n17724) );
  AOI221_X1 U20935 ( .B1(n17828), .B2(n17725), .C1(n17642), .C2(n17725), .A(
        n17724), .ZN(n17730) );
  OAI21_X1 U20936 ( .B1(n17726), .B2(n18073), .A(n17777), .ZN(n17742) );
  AOI221_X1 U20937 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17731), 
        .C1(n18080), .C2(n17750), .A(n17727), .ZN(n17728) );
  XNOR2_X1 U20938 ( .A(n17728), .B(n18050), .ZN(n18070) );
  AOI22_X1 U20939 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17742), .B1(
        n17852), .B2(n18070), .ZN(n17729) );
  OAI211_X1 U20940 ( .C1(n17778), .C2(n18079), .A(n17730), .B(n17729), .ZN(
        P3_U2810) );
  OAI21_X1 U20941 ( .B1(n17750), .B2(n17732), .A(n17731), .ZN(n17733) );
  XNOR2_X1 U20942 ( .A(n17733), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18085) );
  AOI21_X1 U20943 ( .B1(n18855), .B2(n17735), .A(n17946), .ZN(n17759) );
  OAI21_X1 U20944 ( .B1(n17734), .B2(n17980), .A(n17759), .ZN(n17747) );
  AOI22_X1 U20945 ( .A1(n18296), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17747), .ZN(n17739) );
  NOR2_X1 U20946 ( .A1(n17736), .A2(n17735), .ZN(n17749) );
  OAI211_X1 U20947 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17749), .B(n17737), .ZN(n17738) );
  OAI211_X1 U20948 ( .C1(n17812), .C2(n17740), .A(n17739), .B(n17738), .ZN(
        n17741) );
  AOI221_X1 U20949 ( .B1(n17743), .B2(n18080), .C1(n17742), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17741), .ZN(n17744) );
  OAI21_X1 U20950 ( .B1(n18085), .B2(n17880), .A(n17744), .ZN(P3_U2811) );
  NAND2_X1 U20951 ( .A1(n10007), .A2(n17751), .ZN(n18100) );
  OAI22_X1 U20952 ( .A1(n16515), .A2(n18909), .B1(n17812), .B2(n17745), .ZN(
        n17746) );
  AOI221_X1 U20953 ( .B1(n17749), .B2(n17748), .C1(n17747), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17746), .ZN(n17755) );
  OAI21_X1 U20954 ( .B1(n10007), .B2(n17778), .A(n17777), .ZN(n17763) );
  OAI21_X1 U20955 ( .B1(n17779), .B2(n17751), .A(n17750), .ZN(n17753) );
  XNOR2_X1 U20956 ( .A(n17753), .B(n17752), .ZN(n18096) );
  AOI22_X1 U20957 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17763), .B1(
        n17852), .B2(n18096), .ZN(n17754) );
  OAI211_X1 U20958 ( .C1(n17778), .C2(n18100), .A(n17755), .B(n17754), .ZN(
        P3_U2812) );
  AOI21_X1 U20959 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17757), .A(
        n17756), .ZN(n18107) );
  AOI21_X1 U20960 ( .B1(n17758), .B2(n18708), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17760) );
  OAI22_X1 U20961 ( .A1(n17966), .A2(n17761), .B1(n17760), .B2(n17759), .ZN(
        n17762) );
  AOI21_X1 U20962 ( .B1(n18199), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17762), 
        .ZN(n17765) );
  NOR2_X1 U20963 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18116), .ZN(
        n18103) );
  AOI22_X1 U20964 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17763), .B1(
        n10079), .B2(n18103), .ZN(n17764) );
  OAI211_X1 U20965 ( .C1(n18107), .C2(n17880), .A(n17765), .B(n17764), .ZN(
        P3_U2813) );
  OAI21_X1 U20966 ( .B1(n17779), .B2(n11422), .A(n17766), .ZN(n17767) );
  XNOR2_X1 U20967 ( .A(n17767), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n18118) );
  AOI21_X1 U20968 ( .B1(n18855), .B2(n17768), .A(n17946), .ZN(n17795) );
  OAI21_X1 U20969 ( .B1(n17769), .B2(n17980), .A(n17795), .ZN(n17784) );
  AOI22_X1 U20970 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17784), .B1(
        n17828), .B2(n17770), .ZN(n17774) );
  INV_X1 U20971 ( .A(n17807), .ZN(n17797) );
  NAND2_X1 U20972 ( .A1(n17809), .A2(n17771), .ZN(n17825) );
  NOR3_X1 U20973 ( .A1(n17797), .A2(n17796), .A3(n17825), .ZN(n17786) );
  OAI211_X1 U20974 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17786), .B(n17772), .ZN(n17773) );
  OAI211_X1 U20975 ( .C1(n18905), .C2(n16515), .A(n17774), .B(n17773), .ZN(
        n17775) );
  AOI21_X1 U20976 ( .B1(n17852), .B2(n18118), .A(n17775), .ZN(n17776) );
  OAI221_X1 U20977 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17778), 
        .C1(n18116), .C2(n17777), .A(n17776), .ZN(P3_U2814) );
  NOR4_X1 U20978 ( .A1(n17780), .A2(n18212), .A3(n17779), .A4(n18210), .ZN(
        n17839) );
  NAND2_X1 U20979 ( .A1(n18155), .A2(n17839), .ZN(n17830) );
  NOR2_X1 U20980 ( .A1(n11418), .A2(n17830), .ZN(n17817) );
  NAND2_X1 U20981 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17819), .ZN(
        n18163) );
  OAI221_X1 U20982 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17803), 
        .C1(n18139), .C2(n17817), .A(n18163), .ZN(n17781) );
  XNOR2_X1 U20983 ( .A(n18112), .B(n17781), .ZN(n18134) );
  INV_X1 U20984 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17785) );
  OAI22_X1 U20985 ( .A1(n16515), .A2(n18903), .B1(n17812), .B2(n17782), .ZN(
        n17783) );
  AOI221_X1 U20986 ( .B1(n17786), .B2(n17785), .C1(n17784), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17783), .ZN(n17791) );
  NOR2_X1 U20987 ( .A1(n11422), .A2(n17885), .ZN(n17789) );
  NAND2_X1 U20988 ( .A1(n17792), .A2(n18112), .ZN(n18123) );
  NOR2_X1 U20989 ( .A1(n17787), .A2(n17984), .ZN(n17788) );
  NAND3_X1 U20990 ( .A1(n18144), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n18175), .ZN(n17800) );
  NAND2_X1 U20991 ( .A1(n18112), .A2(n17800), .ZN(n18130) );
  AOI22_X1 U20992 ( .A1(n17789), .A2(n18123), .B1(n17788), .B2(n18130), .ZN(
        n17790) );
  OAI211_X1 U20993 ( .C1(n17880), .C2(n18134), .A(n17791), .B(n17790), .ZN(
        P3_U2815) );
  NOR2_X1 U20994 ( .A1(n17871), .A2(n18137), .ZN(n18157) );
  OAI221_X1 U20995 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18157), .A(n17792), .ZN(
        n18149) );
  INV_X1 U20996 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17836) );
  NAND3_X1 U20997 ( .A1(n17906), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18708), .ZN(n17887) );
  INV_X1 U20998 ( .A(n17887), .ZN(n17793) );
  NAND2_X1 U20999 ( .A1(n17794), .A2(n17793), .ZN(n17851) );
  OR2_X1 U21000 ( .A1(n17836), .A2(n17851), .ZN(n17838) );
  AOI221_X1 U21001 ( .B1(n17797), .B2(n17796), .C1(n17838), .C2(n17796), .A(
        n17795), .ZN(n17798) );
  NOR2_X1 U21002 ( .A1(n16515), .A2(n18901), .ZN(n18141) );
  AOI211_X1 U21003 ( .C1(n17799), .C2(n17971), .A(n17798), .B(n18141), .ZN(
        n17806) );
  NAND2_X1 U21004 ( .A1(n18144), .A2(n18175), .ZN(n17802) );
  INV_X1 U21005 ( .A(n17800), .ZN(n17801) );
  AOI21_X1 U21006 ( .B1(n18139), .B2(n17802), .A(n17801), .ZN(n18146) );
  OAI21_X1 U21007 ( .B1(n17803), .B2(n17817), .A(n18163), .ZN(n17804) );
  XNOR2_X1 U21008 ( .A(n17804), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18145) );
  AOI22_X1 U21009 ( .A1(n17962), .A2(n18146), .B1(n17852), .B2(n18145), .ZN(
        n17805) );
  OAI211_X1 U21010 ( .C1(n17885), .C2(n18149), .A(n17806), .B(n17805), .ZN(
        P3_U2816) );
  NAND2_X1 U21011 ( .A1(n18155), .A2(n17867), .ZN(n17835) );
  AOI211_X1 U21012 ( .C1(n17824), .C2(n17813), .A(n17807), .B(n17825), .ZN(
        n17815) );
  OAI22_X1 U21013 ( .A1(n17809), .A2(n17944), .B1(n17808), .B2(n17980), .ZN(
        n17810) );
  NOR2_X1 U21014 ( .A1(n17946), .A2(n17810), .ZN(n17823) );
  OAI22_X1 U21015 ( .A1(n17823), .A2(n17813), .B1(n17812), .B2(n17811), .ZN(
        n17814) );
  AOI211_X1 U21016 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18296), .A(n17815), 
        .B(n17814), .ZN(n17822) );
  NOR2_X1 U21017 ( .A1(n17816), .A2(n18137), .ZN(n18156) );
  OAI22_X1 U21018 ( .A1(n18157), .A2(n17885), .B1(n18156), .B2(n17984), .ZN(
        n17832) );
  INV_X1 U21019 ( .A(n17817), .ZN(n17818) );
  OAI21_X1 U21020 ( .B1(n17829), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17818), .ZN(n17820) );
  XNOR2_X1 U21021 ( .A(n17820), .B(n17819), .ZN(n18153) );
  AOI22_X1 U21022 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17832), .B1(
        n17852), .B2(n18153), .ZN(n17821) );
  OAI211_X1 U21023 ( .C1(n18163), .C2(n17835), .A(n17822), .B(n17821), .ZN(
        P3_U2817) );
  NAND2_X1 U21024 ( .A1(n18296), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18171) );
  OAI221_X1 U21025 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17825), .C1(
        n17824), .C2(n17823), .A(n18171), .ZN(n17826) );
  AOI21_X1 U21026 ( .B1(n17828), .B2(n17827), .A(n17826), .ZN(n17834) );
  NAND2_X1 U21027 ( .A1(n17830), .A2(n17829), .ZN(n17831) );
  XNOR2_X1 U21028 ( .A(n17831), .B(n11418), .ZN(n18170) );
  AOI22_X1 U21029 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17832), .B1(
        n17852), .B2(n18170), .ZN(n17833) );
  OAI211_X1 U21030 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17835), .A(
        n17834), .B(n17833), .ZN(P3_U2818) );
  OAI21_X1 U21031 ( .B1(n17976), .B2(n17836), .A(n17851), .ZN(n17837) );
  AOI22_X1 U21032 ( .A1(n18296), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17838), 
        .B2(n17837), .ZN(n17845) );
  NOR2_X1 U21033 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18182), .ZN(
        n18173) );
  OAI22_X1 U21034 ( .A1(n18177), .A2(n17885), .B1(n17984), .B2(n18175), .ZN(
        n17868) );
  AOI21_X1 U21035 ( .B1(n18182), .B2(n17867), .A(n17868), .ZN(n17856) );
  INV_X1 U21036 ( .A(n17839), .ZN(n17859) );
  NOR2_X1 U21037 ( .A1(n18198), .A2(n17859), .ZN(n17858) );
  AOI21_X1 U21038 ( .B1(n17858), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17840), .ZN(n17841) );
  XNOR2_X1 U21039 ( .A(n17841), .B(n17842), .ZN(n18187) );
  OAI22_X1 U21040 ( .A1(n17856), .A2(n17842), .B1(n18187), .B2(n17880), .ZN(
        n17843) );
  AOI21_X1 U21041 ( .B1(n18173), .B2(n17867), .A(n17843), .ZN(n17844) );
  OAI211_X1 U21042 ( .C1(n17966), .C2(n17846), .A(n17845), .B(n17844), .ZN(
        P3_U2819) );
  AOI21_X1 U21043 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17867), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17855) );
  AOI22_X1 U21044 ( .A1(n18296), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17847), 
        .B2(n17971), .ZN(n17854) );
  NOR2_X1 U21045 ( .A1(n17858), .A2(n9884), .ZN(n17848) );
  XNOR2_X1 U21046 ( .A(n17848), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18193) );
  NOR2_X1 U21047 ( .A1(n17873), .A2(n17887), .ZN(n17862) );
  NAND2_X1 U21048 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17862), .ZN(
        n17861) );
  OAI21_X1 U21049 ( .B1(n17976), .B2(n17849), .A(n17861), .ZN(n17850) );
  AOI22_X1 U21050 ( .A1(n17852), .A2(n18193), .B1(n17851), .B2(n17850), .ZN(
        n17853) );
  OAI211_X1 U21051 ( .C1(n17856), .C2(n17855), .A(n17854), .B(n17853), .ZN(
        P3_U2820) );
  AOI211_X1 U21052 ( .C1(n18198), .C2(n17859), .A(n17858), .B(n17857), .ZN(
        n17860) );
  NOR2_X1 U21053 ( .A1(n9884), .A2(n17860), .ZN(n18206) );
  INV_X1 U21054 ( .A(n17976), .ZN(n17907) );
  OAI211_X1 U21055 ( .C1(n17862), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17907), .B(n17861), .ZN(n17864) );
  NAND2_X1 U21056 ( .A1(n18296), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17863) );
  OAI211_X1 U21057 ( .C1(n17966), .C2(n17865), .A(n17864), .B(n17863), .ZN(
        n17866) );
  AOI221_X1 U21058 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17868), .C1(
        n18198), .C2(n17867), .A(n17866), .ZN(n17869) );
  OAI21_X1 U21059 ( .B1(n18206), .B2(n17880), .A(n17869), .ZN(P3_U2821) );
  NAND2_X1 U21060 ( .A1(n17871), .A2(n17870), .ZN(n18217) );
  AOI21_X1 U21061 ( .B1(n18855), .B2(n17872), .A(n17946), .ZN(n17888) );
  NOR2_X1 U21062 ( .A1(n17872), .A2(n17886), .ZN(n17874) );
  OAI211_X1 U21063 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17874), .A(
        n18708), .B(n17873), .ZN(n17875) );
  NAND2_X1 U21064 ( .A1(n18296), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18214) );
  OAI211_X1 U21065 ( .C1(n17888), .C2(n17876), .A(n17875), .B(n18214), .ZN(
        n17882) );
  XNOR2_X1 U21066 ( .A(n17877), .B(n18217), .ZN(n18224) );
  OAI21_X1 U21067 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17879), .A(
        n17878), .ZN(n18216) );
  OAI22_X1 U21068 ( .A1(n18224), .A2(n17880), .B1(n17984), .B2(n18216), .ZN(
        n17881) );
  AOI211_X1 U21069 ( .C1(n17883), .C2(n17971), .A(n17882), .B(n17881), .ZN(
        n17884) );
  OAI21_X1 U21070 ( .B1(n17885), .B2(n18217), .A(n17884), .ZN(P3_U2822) );
  AOI22_X1 U21071 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17888), .B1(
        n17887), .B2(n17886), .ZN(n17889) );
  AOI21_X1 U21072 ( .B1(n18199), .B2(P3_REIP_REG_7__SCAN_IN), .A(n17889), .ZN(
        n17896) );
  AOI21_X1 U21073 ( .B1(n18210), .B2(n17891), .A(n17890), .ZN(n18227) );
  NOR2_X1 U21074 ( .A1(n17893), .A2(n17892), .ZN(n17894) );
  XNOR2_X1 U21075 ( .A(n17894), .B(n18210), .ZN(n18226) );
  AOI22_X1 U21076 ( .A1(n17972), .A2(n18227), .B1(n17962), .B2(n18226), .ZN(
        n17895) );
  OAI211_X1 U21077 ( .C1(n17966), .C2(n17897), .A(n17896), .B(n17895), .ZN(
        P3_U2823) );
  AOI22_X1 U21078 ( .A1(n17900), .A2(n17919), .B1(n17899), .B2(n17898), .ZN(
        n17905) );
  AOI22_X1 U21079 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17903), .B1(
        n17902), .B2(n17901), .ZN(n17904) );
  XNOR2_X1 U21080 ( .A(n17905), .B(n17904), .ZN(n18241) );
  NAND2_X1 U21081 ( .A1(n17906), .A2(n18708), .ZN(n17912) );
  NAND2_X1 U21082 ( .A1(n17907), .A2(n17912), .ZN(n17925) );
  AOI21_X1 U21083 ( .B1(n17909), .B2(n17908), .A(n9910), .ZN(n18238) );
  AOI22_X1 U21084 ( .A1(n17972), .A2(n18238), .B1(n18296), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n17910) );
  OAI221_X1 U21085 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17912), .C1(
        n17911), .C2(n17925), .A(n17910), .ZN(n17913) );
  AOI21_X1 U21086 ( .B1(n17914), .B2(n17971), .A(n17913), .ZN(n17915) );
  OAI21_X1 U21087 ( .B1(n18241), .B2(n17984), .A(n17915), .ZN(P3_U2824) );
  AOI21_X1 U21088 ( .B1(n17916), .B2(n17979), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17926) );
  AOI21_X1 U21089 ( .B1(n18246), .B2(n17918), .A(n17917), .ZN(n18243) );
  AOI22_X1 U21090 ( .A1(n17972), .A2(n18243), .B1(n18296), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17924) );
  AOI21_X1 U21091 ( .B1(n17921), .B2(n17920), .A(n17919), .ZN(n18242) );
  AOI22_X1 U21092 ( .A1(n17962), .A2(n18242), .B1(n17922), .B2(n17971), .ZN(
        n17923) );
  OAI211_X1 U21093 ( .C1(n17926), .C2(n17925), .A(n17924), .B(n17923), .ZN(
        P3_U2825) );
  AOI21_X1 U21094 ( .B1(n17929), .B2(n17928), .A(n17927), .ZN(n18255) );
  OAI22_X1 U21095 ( .A1(n16515), .A2(n18881), .B1(n18348), .B2(n17930), .ZN(
        n17931) );
  AOI21_X1 U21096 ( .B1(n17962), .B2(n18255), .A(n17931), .ZN(n17936) );
  AOI21_X1 U21097 ( .B1(n17934), .B2(n17933), .A(n17932), .ZN(n18253) );
  OAI21_X1 U21098 ( .B1(n17945), .B2(n17944), .A(n17979), .ZN(n17949) );
  AOI22_X1 U21099 ( .A1(n17972), .A2(n18253), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17949), .ZN(n17935) );
  OAI211_X1 U21100 ( .C1(n17966), .C2(n17937), .A(n17936), .B(n17935), .ZN(
        P3_U2826) );
  AOI21_X1 U21101 ( .B1(n17940), .B2(n17939), .A(n17938), .ZN(n18260) );
  AOI22_X1 U21102 ( .A1(n17962), .A2(n18260), .B1(n18296), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17952) );
  AOI21_X1 U21103 ( .B1(n17943), .B2(n17942), .A(n17941), .ZN(n18261) );
  NOR2_X1 U21104 ( .A1(n17945), .A2(n17944), .ZN(n17947) );
  NOR2_X1 U21105 ( .A1(n17946), .A2(n17960), .ZN(n17959) );
  AOI22_X1 U21106 ( .A1(n17972), .A2(n18261), .B1(n17947), .B2(n17959), .ZN(
        n17951) );
  AOI22_X1 U21107 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17949), .B1(
        n17948), .B2(n17971), .ZN(n17950) );
  NAND3_X1 U21108 ( .A1(n17952), .A2(n17951), .A3(n17950), .ZN(P3_U2827) );
  AOI21_X1 U21109 ( .B1(n17955), .B2(n17954), .A(n17953), .ZN(n18278) );
  AOI22_X1 U21110 ( .A1(n17972), .A2(n18278), .B1(n18296), .B2(
        P3_REIP_REG_2__SCAN_IN), .ZN(n17964) );
  AOI21_X1 U21111 ( .B1(n17958), .B2(n17957), .A(n17956), .ZN(n18276) );
  AOI21_X1 U21112 ( .B1(n17960), .B2(n18348), .A(n17959), .ZN(n17961) );
  AOI21_X1 U21113 ( .B1(n17962), .B2(n18276), .A(n17961), .ZN(n17963) );
  OAI211_X1 U21114 ( .C1(n17966), .C2(n17965), .A(n17964), .B(n17963), .ZN(
        P3_U2828) );
  NOR2_X1 U21115 ( .A1(n17978), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17967) );
  XOR2_X1 U21116 ( .A(n17967), .B(n17970), .Z(n18292) );
  OAI22_X1 U21117 ( .A1(n17984), .A2(n18292), .B1(n16515), .B2(n18989), .ZN(
        n17968) );
  INV_X1 U21118 ( .A(n17968), .ZN(n17974) );
  AOI21_X1 U21119 ( .B1(n17977), .B2(n17970), .A(n17969), .ZN(n18286) );
  AOI22_X1 U21120 ( .A1(n17972), .A2(n18286), .B1(n17975), .B2(n17971), .ZN(
        n17973) );
  OAI211_X1 U21121 ( .C1(n17976), .C2(n17975), .A(n17974), .B(n17973), .ZN(
        P3_U2829) );
  OAI21_X1 U21122 ( .B1(n17978), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17977), .ZN(n18301) );
  INV_X1 U21123 ( .A(n18301), .ZN(n18303) );
  NAND3_X1 U21124 ( .A1(n18966), .A2(n17980), .A3(n17979), .ZN(n17981) );
  AOI22_X1 U21125 ( .A1(n18296), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17981), .ZN(n17982) );
  OAI221_X1 U21126 ( .B1(n18303), .B2(n17984), .C1(n18301), .C2(n17983), .A(
        n17982), .ZN(P3_U2830) );
  NOR2_X1 U21127 ( .A1(n17985), .A2(n18773), .ZN(n17990) );
  OAI22_X1 U21128 ( .A1(n18814), .A2(n18059), .B1(n17986), .B2(n18111), .ZN(
        n18053) );
  NAND3_X1 U21129 ( .A1(n18048), .A2(n18090), .A3(n18053), .ZN(n18025) );
  INV_X1 U21130 ( .A(n18271), .ZN(n18095) );
  OAI21_X1 U21131 ( .B1(n18009), .B2(n18025), .A(n18095), .ZN(n18014) );
  OAI211_X1 U21132 ( .C1(n18271), .C2(n17988), .A(n18014), .B(n17987), .ZN(
        n17989) );
  AOI211_X1 U21133 ( .C1(n18125), .C2(n17991), .A(n17990), .B(n17989), .ZN(
        n18005) );
  NOR3_X1 U21134 ( .A1(n18045), .A2(n18059), .A3(n18044), .ZN(n18038) );
  NAND3_X1 U21135 ( .A1(n18038), .A2(n17992), .A3(n17994), .ZN(n17993) );
  OAI21_X1 U21136 ( .B1(n18005), .B2(n17994), .A(n17993), .ZN(n17995) );
  AOI22_X1 U21137 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18289), .B1(
        n18293), .B2(n17995), .ZN(n17997) );
  NAND2_X1 U21138 ( .A1(n18296), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17996) );
  OAI211_X1 U21139 ( .C1(n17998), .C2(n18223), .A(n17997), .B(n17996), .ZN(
        P3_U2835) );
  INV_X1 U21140 ( .A(n18045), .ZN(n17999) );
  OAI221_X1 U21141 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18000), 
        .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17999), .A(n18293), .ZN(
        n18004) );
  AOI22_X1 U21142 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18289), .B1(
        n18194), .B2(n18001), .ZN(n18003) );
  OAI211_X1 U21143 ( .C1(n18005), .C2(n18004), .A(n18003), .B(n18002), .ZN(
        P3_U2836) );
  INV_X1 U21144 ( .A(n18006), .ZN(n18017) );
  INV_X1 U21145 ( .A(n18047), .ZN(n18091) );
  AOI21_X1 U21146 ( .B1(n18007), .B2(n18091), .A(n18809), .ZN(n18023) );
  AOI211_X1 U21147 ( .C1(n10076), .C2(n18009), .A(n18023), .B(n18008), .ZN(
        n18015) );
  INV_X1 U21148 ( .A(n18010), .ZN(n18012) );
  AOI21_X1 U21149 ( .B1(n18012), .B2(n18011), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18013) );
  AOI211_X1 U21150 ( .C1(n18015), .C2(n18014), .A(n18013), .B(n18287), .ZN(
        n18016) );
  AOI211_X1 U21151 ( .C1(n18289), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18017), .B(n18016), .ZN(n18021) );
  AOI22_X1 U21152 ( .A1(n18150), .A2(n18019), .B1(n18194), .B2(n18018), .ZN(
        n18020) );
  OAI211_X1 U21153 ( .C1(n18302), .C2(n18022), .A(n18021), .B(n18020), .ZN(
        P3_U2837) );
  INV_X1 U21154 ( .A(n18023), .ZN(n18030) );
  INV_X1 U21155 ( .A(n18024), .ZN(n18028) );
  AOI22_X1 U21156 ( .A1(n18125), .A2(n18026), .B1(n18095), .B2(n18025), .ZN(
        n18027) );
  OAI211_X1 U21157 ( .C1(n18028), .C2(n18773), .A(n18027), .B(n18236), .ZN(
        n18032) );
  INV_X1 U21158 ( .A(n18032), .ZN(n18029) );
  NAND3_X1 U21159 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18030), .A3(
        n18029), .ZN(n18031) );
  NAND2_X1 U21160 ( .A1(n16515), .A2(n18031), .ZN(n18041) );
  OAI21_X1 U21161 ( .B1(n18235), .B2(n18032), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18037) );
  AOI22_X1 U21162 ( .A1(n18194), .A2(n18034), .B1(n18060), .B2(n18033), .ZN(
        n18036) );
  NAND2_X1 U21163 ( .A1(n18199), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18035) );
  OAI211_X1 U21164 ( .C1(n18041), .C2(n18037), .A(n18036), .B(n18035), .ZN(
        P3_U2838) );
  AOI21_X1 U21165 ( .B1(n18038), .B2(n18236), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18042) );
  AOI22_X1 U21166 ( .A1(n18199), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18194), 
        .B2(n18039), .ZN(n18040) );
  OAI21_X1 U21167 ( .B1(n18042), .B2(n18041), .A(n18040), .ZN(P3_U2839) );
  AOI22_X1 U21168 ( .A1(n18199), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n18194), 
        .B2(n18043), .ZN(n18058) );
  NOR2_X1 U21169 ( .A1(n18045), .A2(n18044), .ZN(n18056) );
  NOR2_X1 U21170 ( .A1(n9829), .A2(n18125), .ZN(n18174) );
  INV_X1 U21171 ( .A(n18796), .ZN(n18816) );
  AOI22_X1 U21172 ( .A1(n9829), .A2(n18131), .B1(n18125), .B2(n18124), .ZN(
        n18108) );
  OAI221_X1 U21173 ( .B1(n18816), .B2(n18090), .C1(n18816), .C2(n18073), .A(
        n18108), .ZN(n18046) );
  OAI21_X1 U21174 ( .B1(n18048), .B2(n18174), .A(n18071), .ZN(n18049) );
  AOI21_X1 U21175 ( .B1(n18796), .B2(n18050), .A(n18049), .ZN(n18064) );
  INV_X1 U21176 ( .A(n18190), .ZN(n18051) );
  AOI22_X1 U21177 ( .A1(n10076), .A2(n18062), .B1(n18052), .B2(n18051), .ZN(
        n18054) );
  NAND3_X1 U21178 ( .A1(n18064), .A2(n18054), .A3(n18053), .ZN(n18055) );
  OAI211_X1 U21179 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18056), .A(
        n18293), .B(n18055), .ZN(n18057) );
  OAI211_X1 U21180 ( .C1(n18236), .C2(n18059), .A(n18058), .B(n18057), .ZN(
        P3_U2840) );
  INV_X1 U21181 ( .A(n18060), .ZN(n18078) );
  NOR2_X1 U21182 ( .A1(n18078), .A2(n18063), .ZN(n18081) );
  AOI22_X1 U21183 ( .A1(n18296), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18061), 
        .B2(n18081), .ZN(n18068) );
  INV_X1 U21184 ( .A(n18062), .ZN(n18065) );
  NOR2_X1 U21185 ( .A1(n10076), .A2(n18814), .ZN(n18288) );
  AOI221_X1 U21186 ( .B1(n18111), .B2(n18814), .C1(n18063), .C2(n18814), .A(
        n18287), .ZN(n18072) );
  OAI211_X1 U21187 ( .C1(n18065), .C2(n18288), .A(n18072), .B(n18064), .ZN(
        n18066) );
  NAND3_X1 U21188 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n16515), .A3(
        n18066), .ZN(n18067) );
  OAI211_X1 U21189 ( .C1(n18069), .C2(n18223), .A(n18068), .B(n18067), .ZN(
        P3_U2841) );
  AOI22_X1 U21190 ( .A1(n18199), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18194), 
        .B2(n18070), .ZN(n18077) );
  OAI211_X1 U21191 ( .C1(n18073), .C2(n18174), .A(n18072), .B(n18071), .ZN(
        n18074) );
  NOR3_X1 U21192 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18288), .A3(
        n18840), .ZN(n18075) );
  OAI21_X1 U21193 ( .B1(n18082), .B2(n18075), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18076) );
  OAI211_X1 U21194 ( .C1(n18079), .C2(n18078), .A(n18077), .B(n18076), .ZN(
        P3_U2842) );
  AOI22_X1 U21195 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18082), .B1(
        n18081), .B2(n18080), .ZN(n18084) );
  NAND2_X1 U21196 ( .A1(n18199), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18083) );
  OAI211_X1 U21197 ( .C1(n18085), .C2(n18223), .A(n18084), .B(n18083), .ZN(
        P3_U2843) );
  OAI22_X1 U21198 ( .A1(n18809), .A2(n18208), .B1(n18268), .B2(n18269), .ZN(
        n18263) );
  INV_X1 U21199 ( .A(n18263), .ZN(n18088) );
  NOR3_X1 U21200 ( .A1(n18088), .A2(n18087), .A3(n18086), .ZN(n18122) );
  OAI211_X1 U21201 ( .C1(n18089), .C2(n18122), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18293), .ZN(n18102) );
  NOR2_X1 U21202 ( .A1(n18804), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18207) );
  INV_X1 U21203 ( .A(n18207), .ZN(n18272) );
  NAND3_X1 U21204 ( .A1(n18090), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18272), .ZN(n18094) );
  AOI21_X1 U21205 ( .B1(n10007), .B2(n18091), .A(n18809), .ZN(n18093) );
  OAI211_X1 U21206 ( .C1(n10007), .C2(n18174), .A(n18293), .B(n18108), .ZN(
        n18092) );
  AOI211_X1 U21207 ( .C1(n18095), .C2(n18094), .A(n18093), .B(n18092), .ZN(
        n18101) );
  AOI221_X1 U21208 ( .B1(n18271), .B2(n18101), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18101), .A(n18199), .ZN(
        n18097) );
  AOI22_X1 U21209 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18097), .B1(
        n18194), .B2(n18096), .ZN(n18099) );
  NAND2_X1 U21210 ( .A1(n18199), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18098) );
  OAI211_X1 U21211 ( .C1(n18100), .C2(n18102), .A(n18099), .B(n18098), .ZN(
        P3_U2844) );
  NOR2_X1 U21212 ( .A1(n18296), .A2(n18101), .ZN(n18104) );
  INV_X1 U21213 ( .A(n18102), .ZN(n18117) );
  AOI22_X1 U21214 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18104), .B1(
        n18117), .B2(n18103), .ZN(n18106) );
  NAND2_X1 U21215 ( .A1(n18199), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18105) );
  OAI211_X1 U21216 ( .C1(n18107), .C2(n18223), .A(n18106), .B(n18105), .ZN(
        P3_U2845) );
  NAND2_X1 U21217 ( .A1(n18293), .A2(n18108), .ZN(n18115) );
  INV_X1 U21218 ( .A(n18109), .ZN(n18154) );
  NOR2_X1 U21219 ( .A1(n18110), .A2(n18809), .ZN(n18180) );
  AOI21_X1 U21220 ( .B1(n18796), .B2(n18154), .A(n18180), .ZN(n18201) );
  OAI21_X1 U21221 ( .B1(n18112), .B2(n18814), .A(n18111), .ZN(n18113) );
  OAI211_X1 U21222 ( .C1(n18114), .C2(n18190), .A(n18201), .B(n18113), .ZN(
        n18121) );
  OAI221_X1 U21223 ( .B1(n18115), .B2(n18235), .C1(n18115), .C2(n18121), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18120) );
  AOI22_X1 U21224 ( .A1(n18118), .A2(n18194), .B1(n18117), .B2(n18116), .ZN(
        n18119) );
  OAI221_X1 U21225 ( .B1(n18296), .B2(n18120), .C1(n16515), .C2(n18905), .A(
        n18119), .ZN(P3_U2846) );
  NOR2_X1 U21226 ( .A1(n16515), .A2(n18903), .ZN(n18129) );
  OAI21_X1 U21227 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18122), .A(
        n18121), .ZN(n18127) );
  NAND3_X1 U21228 ( .A1(n18125), .A2(n18124), .A3(n18123), .ZN(n18126) );
  AOI21_X1 U21229 ( .B1(n18127), .B2(n18126), .A(n18287), .ZN(n18128) );
  AOI211_X1 U21230 ( .C1(n18289), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18129), .B(n18128), .ZN(n18133) );
  NAND3_X1 U21231 ( .A1(n18277), .A2(n18131), .A3(n18130), .ZN(n18132) );
  OAI211_X1 U21232 ( .C1(n18134), .C2(n18223), .A(n18133), .B(n18132), .ZN(
        P3_U2847) );
  NAND2_X1 U21233 ( .A1(n18293), .A2(n18263), .ZN(n18245) );
  NOR2_X1 U21234 ( .A1(n18211), .A2(n18245), .ZN(n18225) );
  NAND3_X1 U21235 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n18225), .ZN(n18151) );
  NOR2_X1 U21236 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18151), .ZN(
        n18143) );
  NOR2_X1 U21237 ( .A1(n18816), .A2(n18144), .ZN(n18136) );
  OAI211_X1 U21238 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18288), .A(
        n18293), .B(n18201), .ZN(n18135) );
  AOI211_X1 U21239 ( .C1(n10076), .C2(n18137), .A(n18136), .B(n18135), .ZN(
        n18140) );
  INV_X1 U21240 ( .A(n18137), .ZN(n18138) );
  NOR2_X1 U21241 ( .A1(n18984), .A2(n18154), .ZN(n18202) );
  NAND2_X1 U21242 ( .A1(n18138), .A2(n18202), .ZN(n18164) );
  NAND2_X1 U21243 ( .A1(n18814), .A2(n18164), .ZN(n18159) );
  AOI211_X1 U21244 ( .C1(n18140), .C2(n18159), .A(n18199), .B(n18139), .ZN(
        n18142) );
  AOI211_X1 U21245 ( .C1(n18144), .C2(n18143), .A(n18142), .B(n18141), .ZN(
        n18148) );
  AOI22_X1 U21246 ( .A1(n18277), .A2(n18146), .B1(n18194), .B2(n18145), .ZN(
        n18147) );
  OAI211_X1 U21247 ( .C1(n18218), .C2(n18149), .A(n18148), .B(n18147), .ZN(
        P3_U2848) );
  AOI22_X1 U21248 ( .A1(n18177), .A2(n18150), .B1(n18277), .B2(n18175), .ZN(
        n18152) );
  NAND2_X1 U21249 ( .A1(n18152), .A2(n18151), .ZN(n18197) );
  NAND2_X1 U21250 ( .A1(n18155), .A2(n18197), .ZN(n18167) );
  AOI22_X1 U21251 ( .A1(n18296), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18194), 
        .B2(n18153), .ZN(n18162) );
  NAND2_X1 U21252 ( .A1(n18796), .A2(n18154), .ZN(n18188) );
  AOI21_X1 U21253 ( .B1(n18155), .B2(n18188), .A(n18190), .ZN(n18184) );
  OAI22_X1 U21254 ( .A1(n18157), .A2(n18176), .B1(n18156), .B2(n18773), .ZN(
        n18158) );
  NOR3_X1 U21255 ( .A1(n18180), .A2(n18184), .A3(n18158), .ZN(n18165) );
  OAI211_X1 U21256 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18190), .A(
        n18165), .B(n18159), .ZN(n18160) );
  OAI211_X1 U21257 ( .C1(n18287), .C2(n18160), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n16515), .ZN(n18161) );
  OAI211_X1 U21258 ( .C1(n18167), .C2(n18163), .A(n18162), .B(n18161), .ZN(
        P3_U2849) );
  OAI21_X1 U21259 ( .B1(n18814), .B2(n11418), .A(n18164), .ZN(n18166) );
  NAND2_X1 U21260 ( .A1(n18166), .A2(n18165), .ZN(n18169) );
  OAI21_X1 U21261 ( .B1(n18287), .B2(n11418), .A(n18167), .ZN(n18168) );
  AOI22_X1 U21262 ( .A1(n18194), .A2(n18170), .B1(n18169), .B2(n18168), .ZN(
        n18172) );
  OAI211_X1 U21263 ( .C1(n18236), .C2(n11418), .A(n18172), .B(n18171), .ZN(
        P3_U2850) );
  AOI22_X1 U21264 ( .A1(n18296), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18173), 
        .B2(n18197), .ZN(n18186) );
  INV_X1 U21265 ( .A(n18174), .ZN(n18181) );
  OAI22_X1 U21266 ( .A1(n18177), .A2(n18176), .B1(n18773), .B2(n18175), .ZN(
        n18178) );
  NOR2_X1 U21267 ( .A1(n18287), .A2(n18178), .ZN(n18200) );
  OAI221_X1 U21268 ( .B1(n18804), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18804), .C2(n18202), .A(n18200), .ZN(n18179) );
  AOI211_X1 U21269 ( .C1(n18182), .C2(n18181), .A(n18180), .B(n18179), .ZN(
        n18189) );
  OAI21_X1 U21270 ( .B1(n18804), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18189), .ZN(n18183) );
  OAI211_X1 U21271 ( .C1(n18184), .C2(n18183), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16515), .ZN(n18185) );
  OAI211_X1 U21272 ( .C1(n18187), .C2(n18223), .A(n18186), .B(n18185), .ZN(
        P3_U2851) );
  OAI211_X1 U21273 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18190), .A(
        n18189), .B(n18188), .ZN(n18191) );
  NAND2_X1 U21274 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18191), .ZN(
        n18196) );
  NOR2_X1 U21275 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18198), .ZN(
        n18192) );
  AOI22_X1 U21276 ( .A1(n18194), .A2(n18193), .B1(n18192), .B2(n18197), .ZN(
        n18195) );
  OAI221_X1 U21277 ( .B1(n18296), .B2(n18196), .C1(n16515), .C2(n18893), .A(
        n18195), .ZN(P3_U2852) );
  AOI22_X1 U21278 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18199), .B1(n18198), 
        .B2(n18197), .ZN(n18205) );
  OAI211_X1 U21279 ( .C1(n18202), .C2(n18804), .A(n18201), .B(n18200), .ZN(
        n18203) );
  NAND3_X1 U21280 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16515), .A3(
        n18203), .ZN(n18204) );
  OAI211_X1 U21281 ( .C1(n18206), .C2(n18223), .A(n18205), .B(n18204), .ZN(
        P3_U2853) );
  NOR2_X1 U21282 ( .A1(n18268), .A2(n18207), .ZN(n18209) );
  INV_X1 U21283 ( .A(n18208), .ZN(n18267) );
  OAI22_X1 U21284 ( .A1(n18271), .A2(n18209), .B1(n18809), .B2(n18267), .ZN(
        n18250) );
  AOI211_X1 U21285 ( .C1(n18235), .C2(n18211), .A(n18210), .B(n18250), .ZN(
        n18231) );
  OAI21_X1 U21286 ( .B1(n18231), .B2(n18282), .A(n18236), .ZN(n18221) );
  NAND2_X1 U21287 ( .A1(n18213), .A2(n18212), .ZN(n18215) );
  OAI21_X1 U21288 ( .B1(n18245), .B2(n18215), .A(n18214), .ZN(n18220) );
  OAI22_X1 U21289 ( .A1(n18218), .A2(n18217), .B1(n18302), .B2(n18216), .ZN(
        n18219) );
  AOI211_X1 U21290 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n18221), .A(
        n18220), .B(n18219), .ZN(n18222) );
  OAI21_X1 U21291 ( .B1(n18224), .B2(n18223), .A(n18222), .ZN(P3_U2854) );
  AOI21_X1 U21292 ( .B1(n18293), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18225), .ZN(n18230) );
  AOI22_X1 U21293 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18289), .B1(
        n18296), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n18229) );
  INV_X1 U21294 ( .A(n18300), .ZN(n18285) );
  AOI22_X1 U21295 ( .A1(n18285), .A2(n18227), .B1(n18277), .B2(n18226), .ZN(
        n18228) );
  OAI211_X1 U21296 ( .C1(n18231), .C2(n18230), .A(n18229), .B(n18228), .ZN(
        P3_U2855) );
  NOR2_X1 U21297 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18245), .ZN(
        n18232) );
  AOI22_X1 U21298 ( .A1(n18296), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18233), 
        .B2(n18232), .ZN(n18240) );
  INV_X1 U21299 ( .A(n18233), .ZN(n18234) );
  AOI21_X1 U21300 ( .B1(n18235), .B2(n18234), .A(n18250), .ZN(n18237) );
  OAI21_X1 U21301 ( .B1(n18237), .B2(n18287), .A(n18236), .ZN(n18244) );
  AOI22_X1 U21302 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18244), .B1(
        n18285), .B2(n18238), .ZN(n18239) );
  OAI211_X1 U21303 ( .C1(n18241), .C2(n18302), .A(n18240), .B(n18239), .ZN(
        P3_U2856) );
  AOI22_X1 U21304 ( .A1(n18296), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18277), 
        .B2(n18242), .ZN(n18249) );
  AOI22_X1 U21305 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18244), .B1(
        n18285), .B2(n18243), .ZN(n18248) );
  NOR2_X1 U21306 ( .A1(n18251), .A2(n18245), .ZN(n18254) );
  NAND3_X1 U21307 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18254), .A3(
        n18246), .ZN(n18247) );
  NAND3_X1 U21308 ( .A1(n18249), .A2(n18248), .A3(n18247), .ZN(P3_U2857) );
  INV_X1 U21309 ( .A(n18282), .ZN(n18252) );
  OR2_X1 U21310 ( .A1(n18251), .A2(n18250), .ZN(n18262) );
  AOI21_X1 U21311 ( .B1(n18252), .B2(n18262), .A(n18289), .ZN(n18259) );
  AOI22_X1 U21312 ( .A1(n18296), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18285), 
        .B2(n18253), .ZN(n18257) );
  AOI22_X1 U21313 ( .A1(n18255), .A2(n18277), .B1(n18254), .B2(n18258), .ZN(
        n18256) );
  OAI211_X1 U21314 ( .C1(n18259), .C2(n18258), .A(n18257), .B(n18256), .ZN(
        P3_U2858) );
  AOI22_X1 U21315 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18289), .B1(
        n18296), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18266) );
  AOI22_X1 U21316 ( .A1(n18285), .A2(n18261), .B1(n18277), .B2(n18260), .ZN(
        n18265) );
  OAI211_X1 U21317 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18263), .A(
        n18293), .B(n18262), .ZN(n18264) );
  NAND3_X1 U21318 ( .A1(n18266), .A2(n18265), .A3(n18264), .ZN(P3_U2859) );
  OAI21_X1 U21319 ( .B1(n18984), .B2(n18268), .A(n18267), .ZN(n18275) );
  NOR3_X1 U21320 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18968), .A3(
        n18269), .ZN(n18274) );
  AOI211_X1 U21321 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18272), .A(
        n18271), .B(n18270), .ZN(n18273) );
  AOI211_X1 U21322 ( .C1(n10076), .C2(n18275), .A(n18274), .B(n18273), .ZN(
        n18281) );
  AOI22_X1 U21323 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18289), .B1(
        n18296), .B2(P3_REIP_REG_2__SCAN_IN), .ZN(n18280) );
  AOI22_X1 U21324 ( .A1(n18285), .A2(n18278), .B1(n18277), .B2(n18276), .ZN(
        n18279) );
  OAI211_X1 U21325 ( .C1(n18281), .C2(n18287), .A(n18280), .B(n18279), .ZN(
        P3_U2860) );
  NOR2_X1 U21326 ( .A1(n16515), .A2(n18989), .ZN(n18284) );
  AOI211_X1 U21327 ( .C1(n18816), .C2(n18984), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18282), .ZN(n18283) );
  AOI211_X1 U21328 ( .C1(n18286), .C2(n18285), .A(n18284), .B(n18283), .ZN(
        n18291) );
  NOR3_X1 U21329 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18288), .A3(
        n18287), .ZN(n18295) );
  OAI21_X1 U21330 ( .B1(n18289), .B2(n18295), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18290) );
  OAI211_X1 U21331 ( .C1(n18292), .C2(n18302), .A(n18291), .B(n18290), .ZN(
        P3_U2861) );
  AOI21_X1 U21332 ( .B1(n18816), .B2(n18293), .A(n18984), .ZN(n18294) );
  NOR2_X1 U21333 ( .A1(n18295), .A2(n18294), .ZN(n18298) );
  INV_X1 U21334 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18297) );
  MUX2_X1 U21335 ( .A(n18298), .B(n18297), .S(n18296), .Z(n18299) );
  OAI221_X1 U21336 ( .B1(n18303), .B2(n18302), .C1(n18301), .C2(n18300), .A(
        n18299), .ZN(P3_U2862) );
  AOI211_X1 U21337 ( .C1(n18305), .C2(n18304), .A(n18840), .B(n18966), .ZN(
        n18841) );
  OAI21_X1 U21338 ( .B1(n18841), .B2(n18355), .A(n18310), .ZN(n18306) );
  OAI221_X1 U21339 ( .B1(n18819), .B2(n19003), .C1(n18819), .C2(n18310), .A(
        n18306), .ZN(P3_U2863) );
  INV_X1 U21340 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18829) );
  NOR2_X1 U21341 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18829), .ZN(
        n18612) );
  NOR2_X1 U21342 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18826), .ZN(
        n18491) );
  NOR2_X1 U21343 ( .A1(n18612), .A2(n18491), .ZN(n18308) );
  OAI22_X1 U21344 ( .A1(n18309), .A2(n18829), .B1(n18308), .B2(n18307), .ZN(
        P3_U2866) );
  NOR2_X1 U21345 ( .A1(n18830), .A2(n18310), .ZN(P3_U2867) );
  NOR2_X1 U21346 ( .A1(n18829), .A2(n18492), .ZN(n18706) );
  INV_X1 U21347 ( .A(n18706), .ZN(n18709) );
  OR2_X1 U21348 ( .A1(n18819), .A2(n18709), .ZN(n18751) );
  INV_X1 U21349 ( .A(n18751), .ZN(n18764) );
  NAND2_X1 U21350 ( .A1(n18821), .A2(n18819), .ZN(n18822) );
  NAND2_X1 U21351 ( .A1(n18826), .A2(n18829), .ZN(n18401) );
  NOR2_X1 U21352 ( .A1(n18822), .A2(n18401), .ZN(n18419) );
  NOR2_X1 U21353 ( .A1(n18764), .A2(n18415), .ZN(n18375) );
  OAI21_X1 U21354 ( .B1(n18819), .B2(n18954), .A(n18673), .ZN(n18560) );
  NAND2_X1 U21355 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18311) );
  INV_X1 U21356 ( .A(n18311), .ZN(n18639) );
  NAND2_X1 U21357 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18819), .ZN(
        n18559) );
  NAND2_X1 U21358 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18821), .ZN(
        n18446) );
  NAND2_X1 U21359 ( .A1(n18559), .A2(n18446), .ZN(n18611) );
  NAND2_X1 U21360 ( .A1(n18639), .A2(n18611), .ZN(n18669) );
  OAI22_X1 U21361 ( .A1(n18375), .A2(n18560), .B1(n18348), .B2(n18669), .ZN(
        n18353) );
  NOR2_X1 U21362 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18311), .ZN(
        n18707) );
  NAND2_X1 U21363 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18707), .ZN(
        n18671) );
  INV_X1 U21364 ( .A(n18671), .ZN(n18767) );
  NOR2_X2 U21365 ( .A1(n19319), .A2(n18348), .ZN(n18713) );
  AND2_X1 U21366 ( .A1(n18673), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18710) );
  NOR2_X1 U21367 ( .A1(n18849), .A2(n18375), .ZN(n18347) );
  AOI22_X1 U21368 ( .A1(n18767), .A2(n18713), .B1(n18710), .B2(n18347), .ZN(
        n18316) );
  NOR2_X1 U21369 ( .A1(n18311), .A2(n18559), .ZN(n18699) );
  NAND2_X1 U21370 ( .A1(n18708), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18678) );
  INV_X1 U21371 ( .A(n18678), .ZN(n18711) );
  NAND2_X1 U21372 ( .A1(n18313), .A2(n18312), .ZN(n18349) );
  NOR2_X2 U21373 ( .A1(n18314), .A2(n18349), .ZN(n18712) );
  AOI22_X1 U21374 ( .A1(n18675), .A2(n18711), .B1(n18712), .B2(n18415), .ZN(
        n18315) );
  OAI211_X1 U21375 ( .C1(n18317), .C2(n18353), .A(n18316), .B(n18315), .ZN(
        P3_U2868) );
  AND2_X1 U21376 ( .A1(n18708), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18718) );
  AND2_X1 U21377 ( .A1(n18673), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18717) );
  AOI22_X1 U21378 ( .A1(n18675), .A2(n18718), .B1(n18717), .B2(n18347), .ZN(
        n18319) );
  NAND2_X1 U21379 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18708), .ZN(n18681) );
  INV_X1 U21380 ( .A(n18681), .ZN(n18720) );
  NOR2_X1 U21381 ( .A1(n19008), .A2(n18349), .ZN(n18719) );
  AOI22_X1 U21382 ( .A1(n18767), .A2(n18720), .B1(n18719), .B2(n18415), .ZN(
        n18318) );
  OAI211_X1 U21383 ( .C1(n18320), .C2(n18353), .A(n18319), .B(n18318), .ZN(
        P3_U2869) );
  NAND2_X1 U21384 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18708), .ZN(n18684) );
  INV_X1 U21385 ( .A(n18684), .ZN(n18727) );
  NOR2_X2 U21386 ( .A1(n18356), .A2(n18321), .ZN(n18724) );
  AOI22_X1 U21387 ( .A1(n18767), .A2(n18727), .B1(n18724), .B2(n18347), .ZN(
        n18324) );
  NOR2_X1 U21388 ( .A1(n9803), .A2(n18349), .ZN(n18726) );
  AOI22_X1 U21389 ( .A1(n18675), .A2(n18725), .B1(n18726), .B2(n18419), .ZN(
        n18323) );
  OAI211_X1 U21390 ( .C1(n18325), .C2(n18353), .A(n18324), .B(n18323), .ZN(
        P3_U2870) );
  NAND2_X1 U21391 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18708), .ZN(n18687) );
  INV_X1 U21392 ( .A(n18687), .ZN(n18734) );
  NOR2_X2 U21393 ( .A1(n18356), .A2(n18326), .ZN(n18731) );
  AOI22_X1 U21394 ( .A1(n18767), .A2(n18734), .B1(n18731), .B2(n18347), .ZN(
        n18329) );
  AND2_X1 U21395 ( .A1(n18708), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18732) );
  NOR2_X1 U21396 ( .A1(n18327), .A2(n18349), .ZN(n18733) );
  AOI22_X1 U21397 ( .A1(n18675), .A2(n18732), .B1(n18733), .B2(n18419), .ZN(
        n18328) );
  OAI211_X1 U21398 ( .C1(n18330), .C2(n18353), .A(n18329), .B(n18328), .ZN(
        P3_U2871) );
  NOR2_X2 U21399 ( .A1(n18348), .A2(n19345), .ZN(n18739) );
  NOR2_X2 U21400 ( .A1(n18356), .A2(n18331), .ZN(n18738) );
  AOI22_X1 U21401 ( .A1(n18675), .A2(n18739), .B1(n18738), .B2(n18347), .ZN(
        n18334) );
  NAND2_X1 U21402 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18708), .ZN(n18743) );
  INV_X1 U21403 ( .A(n18743), .ZN(n18653) );
  NOR2_X1 U21404 ( .A1(n18332), .A2(n18349), .ZN(n18740) );
  AOI22_X1 U21405 ( .A1(n18767), .A2(n18653), .B1(n18740), .B2(n18419), .ZN(
        n18333) );
  OAI211_X1 U21406 ( .C1(n18335), .C2(n18353), .A(n18334), .B(n18333), .ZN(
        P3_U2872) );
  NOR2_X1 U21407 ( .A1(n18348), .A2(n19351), .ZN(n18746) );
  NOR2_X2 U21408 ( .A1(n18356), .A2(n18336), .ZN(n18745) );
  AOI22_X1 U21409 ( .A1(n18675), .A2(n18746), .B1(n18745), .B2(n18347), .ZN(
        n18339) );
  NOR2_X2 U21410 ( .A1(n19352), .A2(n18348), .ZN(n18747) );
  AOI22_X1 U21411 ( .A1(n18767), .A2(n18747), .B1(n18691), .B2(n18419), .ZN(
        n18338) );
  OAI211_X1 U21412 ( .C1(n18340), .C2(n18353), .A(n18339), .B(n18338), .ZN(
        P3_U2873) );
  NAND2_X1 U21413 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18708), .ZN(n18697) );
  INV_X1 U21414 ( .A(n18697), .ZN(n18754) );
  NOR2_X2 U21415 ( .A1(n18356), .A2(n18341), .ZN(n18753) );
  AOI22_X1 U21416 ( .A1(n18767), .A2(n18754), .B1(n18753), .B2(n18347), .ZN(
        n18344) );
  AND2_X1 U21417 ( .A1(n18708), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18756) );
  NOR2_X1 U21418 ( .A1(n9806), .A2(n18349), .ZN(n18755) );
  AOI22_X1 U21419 ( .A1(n18675), .A2(n18756), .B1(n18755), .B2(n18419), .ZN(
        n18343) );
  OAI211_X1 U21420 ( .C1(n18345), .C2(n18353), .A(n18344), .B(n18343), .ZN(
        P3_U2874) );
  NOR2_X2 U21421 ( .A1(n19362), .A2(n18348), .ZN(n18766) );
  NOR2_X2 U21422 ( .A1(n18346), .A2(n18356), .ZN(n18761) );
  AOI22_X1 U21423 ( .A1(n18675), .A2(n18766), .B1(n18761), .B2(n18347), .ZN(
        n18352) );
  NOR2_X1 U21424 ( .A1(n18348), .A2(n19365), .ZN(n18762) );
  AOI22_X1 U21425 ( .A1(n18767), .A2(n18762), .B1(n18765), .B2(n18419), .ZN(
        n18351) );
  OAI211_X1 U21426 ( .C1(n18354), .C2(n18353), .A(n18352), .B(n18351), .ZN(
        P3_U2875) );
  INV_X1 U21427 ( .A(n18712), .ZN(n18643) );
  INV_X1 U21428 ( .A(n18446), .ZN(n18537) );
  INV_X1 U21429 ( .A(n18401), .ZN(n18399) );
  NAND2_X1 U21430 ( .A1(n18537), .A2(n18399), .ZN(n18444) );
  AOI22_X1 U21431 ( .A1(n18711), .A2(n18764), .B1(n18710), .B2(n18371), .ZN(
        n18358) );
  NOR2_X1 U21432 ( .A1(n18356), .A2(n18355), .ZN(n18705) );
  AND2_X1 U21433 ( .A1(n18821), .A2(n18705), .ZN(n18638) );
  AOI22_X1 U21434 ( .A1(n18708), .A2(n18706), .B1(n18399), .B2(n18638), .ZN(
        n18372) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18372), .B1(
        n18699), .B2(n18713), .ZN(n18357) );
  OAI211_X1 U21436 ( .C1(n18643), .C2(n18444), .A(n18358), .B(n18357), .ZN(
        P3_U2876) );
  INV_X1 U21437 ( .A(n18719), .ZN(n18594) );
  AOI22_X1 U21438 ( .A1(n18675), .A2(n18720), .B1(n18717), .B2(n18371), .ZN(
        n18360) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18372), .B1(
        n18718), .B2(n18764), .ZN(n18359) );
  OAI211_X1 U21440 ( .C1(n18594), .C2(n18444), .A(n18360), .B(n18359), .ZN(
        P3_U2877) );
  INV_X1 U21441 ( .A(n18726), .ZN(n18649) );
  AOI22_X1 U21442 ( .A1(n18725), .A2(n18764), .B1(n18724), .B2(n18371), .ZN(
        n18362) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18372), .B1(
        n18675), .B2(n18727), .ZN(n18361) );
  OAI211_X1 U21444 ( .C1(n18649), .C2(n18444), .A(n18362), .B(n18361), .ZN(
        P3_U2878) );
  INV_X1 U21445 ( .A(n18733), .ZN(n18652) );
  AOI22_X1 U21446 ( .A1(n18675), .A2(n18734), .B1(n18731), .B2(n18371), .ZN(
        n18364) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18372), .B1(
        n18732), .B2(n18764), .ZN(n18363) );
  OAI211_X1 U21448 ( .C1(n18652), .C2(n18444), .A(n18364), .B(n18363), .ZN(
        P3_U2879) );
  AOI22_X1 U21449 ( .A1(n18739), .A2(n18764), .B1(n18738), .B2(n18371), .ZN(
        n18366) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18372), .B1(
        n18675), .B2(n18653), .ZN(n18365) );
  OAI211_X1 U21451 ( .C1(n18656), .C2(n18444), .A(n18366), .B(n18365), .ZN(
        P3_U2880) );
  AOI22_X1 U21452 ( .A1(n18746), .A2(n18764), .B1(n18745), .B2(n18371), .ZN(
        n18368) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18372), .B1(
        n18675), .B2(n18747), .ZN(n18367) );
  OAI211_X1 U21454 ( .C1(n18752), .C2(n18444), .A(n18368), .B(n18367), .ZN(
        P3_U2881) );
  AOI22_X1 U21455 ( .A1(n18675), .A2(n18754), .B1(n18753), .B2(n18371), .ZN(
        n18370) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18372), .B1(
        n18756), .B2(n18764), .ZN(n18369) );
  OAI211_X1 U21457 ( .C1(n18662), .C2(n18444), .A(n18370), .B(n18369), .ZN(
        P3_U2882) );
  INV_X1 U21458 ( .A(n18765), .ZN(n18668) );
  AOI22_X1 U21459 ( .A1(n18761), .A2(n18371), .B1(n18766), .B2(n18764), .ZN(
        n18374) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18372), .B1(
        n18699), .B2(n18762), .ZN(n18373) );
  OAI211_X1 U21461 ( .C1(n18668), .C2(n18444), .A(n18374), .B(n18373), .ZN(
        P3_U2883) );
  NOR2_X2 U21462 ( .A1(n18559), .A2(n18401), .ZN(n18459) );
  NOR2_X1 U21463 ( .A1(n18435), .A2(n18459), .ZN(n18423) );
  INV_X1 U21464 ( .A(n18613), .ZN(n18670) );
  AOI221_X1 U21465 ( .B1(n18375), .B2(n18423), .C1(n18670), .C2(n18423), .A(
        n18560), .ZN(n18398) );
  NOR2_X1 U21466 ( .A1(n18849), .A2(n18423), .ZN(n18394) );
  AOI22_X1 U21467 ( .A1(n18711), .A2(n18415), .B1(n18710), .B2(n18394), .ZN(
        n18377) );
  AOI22_X1 U21468 ( .A1(n18712), .A2(n18459), .B1(n18713), .B2(n18764), .ZN(
        n18376) );
  OAI211_X1 U21469 ( .C1(n18398), .C2(n18378), .A(n18377), .B(n18376), .ZN(
        P3_U2884) );
  INV_X1 U21470 ( .A(n18459), .ZN(n18466) );
  AOI22_X1 U21471 ( .A1(n18720), .A2(n18764), .B1(n18717), .B2(n18394), .ZN(
        n18380) );
  INV_X1 U21472 ( .A(n18398), .ZN(n18391) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18391), .B1(
        n18718), .B2(n18419), .ZN(n18379) );
  OAI211_X1 U21474 ( .C1(n18594), .C2(n18466), .A(n18380), .B(n18379), .ZN(
        P3_U2885) );
  AOI22_X1 U21475 ( .A1(n18725), .A2(n18415), .B1(n18724), .B2(n18394), .ZN(
        n18382) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18391), .B1(
        n18727), .B2(n18764), .ZN(n18381) );
  OAI211_X1 U21477 ( .C1(n18649), .C2(n18466), .A(n18382), .B(n18381), .ZN(
        P3_U2886) );
  AOI22_X1 U21478 ( .A1(n18734), .A2(n18764), .B1(n18731), .B2(n18394), .ZN(
        n18384) );
  AOI22_X1 U21479 ( .A1(n18733), .A2(n18459), .B1(n18732), .B2(n18419), .ZN(
        n18383) );
  OAI211_X1 U21480 ( .C1(n18398), .C2(n18385), .A(n18384), .B(n18383), .ZN(
        P3_U2887) );
  AOI22_X1 U21481 ( .A1(n18653), .A2(n18764), .B1(n18738), .B2(n18394), .ZN(
        n18387) );
  AOI22_X1 U21482 ( .A1(n18740), .A2(n18459), .B1(n18739), .B2(n18419), .ZN(
        n18386) );
  OAI211_X1 U21483 ( .C1(n18398), .C2(n18388), .A(n18387), .B(n18386), .ZN(
        P3_U2888) );
  AOI22_X1 U21484 ( .A1(n18747), .A2(n18764), .B1(n18745), .B2(n18394), .ZN(
        n18390) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18391), .B1(
        n18746), .B2(n18415), .ZN(n18389) );
  OAI211_X1 U21486 ( .C1(n18752), .C2(n18466), .A(n18390), .B(n18389), .ZN(
        P3_U2889) );
  AOI22_X1 U21487 ( .A1(n18756), .A2(n18415), .B1(n18753), .B2(n18394), .ZN(
        n18393) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18391), .B1(
        n18754), .B2(n18764), .ZN(n18392) );
  OAI211_X1 U21489 ( .C1(n18662), .C2(n18466), .A(n18393), .B(n18392), .ZN(
        P3_U2890) );
  AOI22_X1 U21490 ( .A1(n18761), .A2(n18394), .B1(n18766), .B2(n18415), .ZN(
        n18396) );
  AOI22_X1 U21491 ( .A1(n18762), .A2(n18764), .B1(n18765), .B2(n18459), .ZN(
        n18395) );
  OAI211_X1 U21492 ( .C1(n18398), .C2(n18397), .A(n18396), .B(n18395), .ZN(
        P3_U2891) );
  NAND2_X1 U21493 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18399), .ZN(
        n18400) );
  NOR2_X1 U21494 ( .A1(n18849), .A2(n18400), .ZN(n18418) );
  AOI22_X1 U21495 ( .A1(n18713), .A2(n18415), .B1(n18710), .B2(n18418), .ZN(
        n18404) );
  NAND2_X1 U21496 ( .A1(n18821), .A2(n18670), .ZN(n18490) );
  INV_X1 U21497 ( .A(n18400), .ZN(n18445) );
  NAND2_X1 U21498 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18445), .ZN(
        n18489) );
  OAI21_X1 U21499 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18401), .A(n18489), 
        .ZN(n18402) );
  NAND3_X1 U21500 ( .A1(n18673), .A2(n18490), .A3(n18402), .ZN(n18420) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18420), .B1(
        n18712), .B2(n18482), .ZN(n18403) );
  OAI211_X1 U21502 ( .C1(n18678), .C2(n18444), .A(n18404), .B(n18403), .ZN(
        P3_U2892) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18420), .B1(
        n18717), .B2(n18418), .ZN(n18406) );
  AOI22_X1 U21504 ( .A1(n18720), .A2(n18415), .B1(n18718), .B2(n18435), .ZN(
        n18405) );
  OAI211_X1 U21505 ( .C1(n18594), .C2(n18489), .A(n18406), .B(n18405), .ZN(
        P3_U2893) );
  AOI22_X1 U21506 ( .A1(n18725), .A2(n18435), .B1(n18724), .B2(n18418), .ZN(
        n18408) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18420), .B1(
        n18727), .B2(n18415), .ZN(n18407) );
  OAI211_X1 U21508 ( .C1(n18649), .C2(n18489), .A(n18408), .B(n18407), .ZN(
        P3_U2894) );
  AOI22_X1 U21509 ( .A1(n18732), .A2(n18435), .B1(n18731), .B2(n18418), .ZN(
        n18410) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18420), .B1(
        n18734), .B2(n18419), .ZN(n18409) );
  OAI211_X1 U21511 ( .C1(n18652), .C2(n18489), .A(n18410), .B(n18409), .ZN(
        P3_U2895) );
  AOI22_X1 U21512 ( .A1(n18739), .A2(n18435), .B1(n18738), .B2(n18418), .ZN(
        n18412) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18420), .B1(
        n18653), .B2(n18415), .ZN(n18411) );
  OAI211_X1 U21514 ( .C1(n18656), .C2(n18489), .A(n18412), .B(n18411), .ZN(
        P3_U2896) );
  INV_X1 U21515 ( .A(n18746), .ZN(n18694) );
  AOI22_X1 U21516 ( .A1(n18747), .A2(n18415), .B1(n18745), .B2(n18418), .ZN(
        n18414) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18420), .B1(
        n18691), .B2(n18482), .ZN(n18413) );
  OAI211_X1 U21518 ( .C1(n18694), .C2(n18444), .A(n18414), .B(n18413), .ZN(
        P3_U2897) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18420), .B1(
        n18753), .B2(n18418), .ZN(n18417) );
  AOI22_X1 U21520 ( .A1(n18754), .A2(n18415), .B1(n18756), .B2(n18435), .ZN(
        n18416) );
  OAI211_X1 U21521 ( .C1(n18662), .C2(n18489), .A(n18417), .B(n18416), .ZN(
        P3_U2898) );
  AOI22_X1 U21522 ( .A1(n18761), .A2(n18418), .B1(n18766), .B2(n18435), .ZN(
        n18422) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18420), .B1(
        n18762), .B2(n18419), .ZN(n18421) );
  OAI211_X1 U21524 ( .C1(n18668), .C2(n18489), .A(n18422), .B(n18421), .ZN(
        P3_U2899) );
  INV_X1 U21525 ( .A(n18491), .ZN(n18467) );
  NOR2_X1 U21526 ( .A1(n18482), .A2(n9798), .ZN(n18468) );
  NOR2_X1 U21527 ( .A1(n18849), .A2(n18468), .ZN(n18440) );
  AOI22_X1 U21528 ( .A1(n18713), .A2(n18435), .B1(n18710), .B2(n18440), .ZN(
        n18426) );
  OAI21_X1 U21529 ( .B1(n18423), .B2(n18670), .A(n18468), .ZN(n18424) );
  OAI211_X1 U21530 ( .C1(n9798), .C2(n18954), .A(n18673), .B(n18424), .ZN(
        n18441) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18441), .B1(
        n18712), .B2(n9798), .ZN(n18425) );
  OAI211_X1 U21532 ( .C1(n18678), .C2(n18466), .A(n18426), .B(n18425), .ZN(
        P3_U2900) );
  INV_X1 U21533 ( .A(n9798), .ZN(n18504) );
  AOI22_X1 U21534 ( .A1(n18720), .A2(n18435), .B1(n18717), .B2(n18440), .ZN(
        n18428) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18441), .B1(
        n18718), .B2(n18459), .ZN(n18427) );
  OAI211_X1 U21536 ( .C1(n18594), .C2(n18504), .A(n18428), .B(n18427), .ZN(
        P3_U2901) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18441), .B1(
        n18724), .B2(n18440), .ZN(n18430) );
  AOI22_X1 U21538 ( .A1(n18726), .A2(n9798), .B1(n18725), .B2(n18459), .ZN(
        n18429) );
  OAI211_X1 U21539 ( .C1(n18684), .C2(n18444), .A(n18430), .B(n18429), .ZN(
        P3_U2902) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18441), .B1(
        n18731), .B2(n18440), .ZN(n18432) );
  AOI22_X1 U21541 ( .A1(n18733), .A2(n9798), .B1(n18732), .B2(n18459), .ZN(
        n18431) );
  OAI211_X1 U21542 ( .C1(n18687), .C2(n18444), .A(n18432), .B(n18431), .ZN(
        P3_U2903) );
  AOI22_X1 U21543 ( .A1(n18653), .A2(n18435), .B1(n18738), .B2(n18440), .ZN(
        n18434) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18441), .B1(
        n18739), .B2(n18459), .ZN(n18433) );
  OAI211_X1 U21545 ( .C1(n18656), .C2(n18504), .A(n18434), .B(n18433), .ZN(
        P3_U2904) );
  AOI22_X1 U21546 ( .A1(n18747), .A2(n18435), .B1(n18745), .B2(n18440), .ZN(
        n18437) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18441), .B1(
        n18691), .B2(n9798), .ZN(n18436) );
  OAI211_X1 U21548 ( .C1(n18694), .C2(n18466), .A(n18437), .B(n18436), .ZN(
        P3_U2905) );
  AOI22_X1 U21549 ( .A1(n18756), .A2(n18459), .B1(n18753), .B2(n18440), .ZN(
        n18439) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18441), .B1(
        n18755), .B2(n9798), .ZN(n18438) );
  OAI211_X1 U21551 ( .C1(n18697), .C2(n18444), .A(n18439), .B(n18438), .ZN(
        P3_U2906) );
  INV_X1 U21552 ( .A(n18762), .ZN(n18703) );
  AOI22_X1 U21553 ( .A1(n18761), .A2(n18440), .B1(n18766), .B2(n18459), .ZN(
        n18443) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18441), .B1(
        n18765), .B2(n9798), .ZN(n18442) );
  OAI211_X1 U21555 ( .C1(n18703), .C2(n18444), .A(n18443), .B(n18442), .ZN(
        P3_U2907) );
  AOI22_X1 U21556 ( .A1(n18713), .A2(n18459), .B1(n18710), .B2(n18462), .ZN(
        n18448) );
  AOI22_X1 U21557 ( .A1(n18708), .A2(n18445), .B1(n18491), .B2(n18638), .ZN(
        n18463) );
  NOR2_X2 U21558 ( .A1(n18446), .A2(n18467), .ZN(n18529) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18463), .B1(
        n18712), .B2(n18529), .ZN(n18447) );
  OAI211_X1 U21560 ( .C1(n18678), .C2(n18489), .A(n18448), .B(n18447), .ZN(
        P3_U2908) );
  AOI22_X1 U21561 ( .A1(n18717), .A2(n18462), .B1(n18718), .B2(n18482), .ZN(
        n18450) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18463), .B1(
        n18719), .B2(n18529), .ZN(n18449) );
  OAI211_X1 U21563 ( .C1(n18681), .C2(n18466), .A(n18450), .B(n18449), .ZN(
        P3_U2909) );
  INV_X1 U21564 ( .A(n18529), .ZN(n18536) );
  AOI22_X1 U21565 ( .A1(n18727), .A2(n18459), .B1(n18724), .B2(n18462), .ZN(
        n18452) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18463), .B1(
        n18725), .B2(n18482), .ZN(n18451) );
  OAI211_X1 U21567 ( .C1(n18649), .C2(n18536), .A(n18452), .B(n18451), .ZN(
        P3_U2910) );
  AOI22_X1 U21568 ( .A1(n18732), .A2(n18482), .B1(n18731), .B2(n18462), .ZN(
        n18454) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18463), .B1(
        n18733), .B2(n18529), .ZN(n18453) );
  OAI211_X1 U21570 ( .C1(n18687), .C2(n18466), .A(n18454), .B(n18453), .ZN(
        P3_U2911) );
  AOI22_X1 U21571 ( .A1(n18653), .A2(n18459), .B1(n18738), .B2(n18462), .ZN(
        n18456) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18463), .B1(
        n18739), .B2(n18482), .ZN(n18455) );
  OAI211_X1 U21573 ( .C1(n18656), .C2(n18536), .A(n18456), .B(n18455), .ZN(
        P3_U2912) );
  AOI22_X1 U21574 ( .A1(n18747), .A2(n18459), .B1(n18745), .B2(n18462), .ZN(
        n18458) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18463), .B1(
        n18691), .B2(n18529), .ZN(n18457) );
  OAI211_X1 U21576 ( .C1(n18694), .C2(n18489), .A(n18458), .B(n18457), .ZN(
        P3_U2913) );
  AOI22_X1 U21577 ( .A1(n18754), .A2(n18459), .B1(n18753), .B2(n18462), .ZN(
        n18461) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18463), .B1(
        n18756), .B2(n18482), .ZN(n18460) );
  OAI211_X1 U21579 ( .C1(n18662), .C2(n18536), .A(n18461), .B(n18460), .ZN(
        P3_U2914) );
  AOI22_X1 U21580 ( .A1(n18761), .A2(n18462), .B1(n18766), .B2(n18482), .ZN(
        n18465) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18463), .B1(
        n18765), .B2(n18529), .ZN(n18464) );
  OAI211_X1 U21582 ( .C1(n18703), .C2(n18466), .A(n18465), .B(n18464), .ZN(
        P3_U2915) );
  NOR2_X2 U21583 ( .A1(n18559), .A2(n18467), .ZN(n18554) );
  NOR2_X1 U21584 ( .A1(n18529), .A2(n18554), .ZN(n18514) );
  NOR2_X1 U21585 ( .A1(n18849), .A2(n18514), .ZN(n18485) );
  AOI22_X1 U21586 ( .A1(n18713), .A2(n18482), .B1(n18710), .B2(n18485), .ZN(
        n18471) );
  AOI221_X1 U21587 ( .B1(n18514), .B2(n18670), .C1(n18514), .C2(n18468), .A(
        n18560), .ZN(n18469) );
  INV_X1 U21588 ( .A(n18469), .ZN(n18486) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18486), .B1(
        n18712), .B2(n18554), .ZN(n18470) );
  OAI211_X1 U21590 ( .C1(n18678), .C2(n18504), .A(n18471), .B(n18470), .ZN(
        P3_U2916) );
  AOI22_X1 U21591 ( .A1(n18717), .A2(n18485), .B1(n18718), .B2(n9798), .ZN(
        n18473) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18486), .B1(
        n18719), .B2(n18554), .ZN(n18472) );
  OAI211_X1 U21593 ( .C1(n18681), .C2(n18489), .A(n18473), .B(n18472), .ZN(
        P3_U2917) );
  AOI22_X1 U21594 ( .A1(n18725), .A2(n9798), .B1(n18724), .B2(n18485), .ZN(
        n18475) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18486), .B1(
        n18726), .B2(n18554), .ZN(n18474) );
  OAI211_X1 U21596 ( .C1(n18684), .C2(n18489), .A(n18475), .B(n18474), .ZN(
        P3_U2918) );
  INV_X1 U21597 ( .A(n18554), .ZN(n18528) );
  AOI22_X1 U21598 ( .A1(n18734), .A2(n18482), .B1(n18731), .B2(n18485), .ZN(
        n18477) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18486), .B1(
        n18732), .B2(n9798), .ZN(n18476) );
  OAI211_X1 U21600 ( .C1(n18652), .C2(n18528), .A(n18477), .B(n18476), .ZN(
        P3_U2919) );
  AOI22_X1 U21601 ( .A1(n18653), .A2(n18482), .B1(n18738), .B2(n18485), .ZN(
        n18479) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18486), .B1(
        n18739), .B2(n9798), .ZN(n18478) );
  OAI211_X1 U21603 ( .C1(n18656), .C2(n18528), .A(n18479), .B(n18478), .ZN(
        P3_U2920) );
  AOI22_X1 U21604 ( .A1(n18746), .A2(n9798), .B1(n18745), .B2(n18485), .ZN(
        n18481) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18486), .B1(
        n18747), .B2(n18482), .ZN(n18480) );
  OAI211_X1 U21606 ( .C1(n18752), .C2(n18528), .A(n18481), .B(n18480), .ZN(
        P3_U2921) );
  AOI22_X1 U21607 ( .A1(n18754), .A2(n18482), .B1(n18753), .B2(n18485), .ZN(
        n18484) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18486), .B1(
        n18756), .B2(n9798), .ZN(n18483) );
  OAI211_X1 U21609 ( .C1(n18662), .C2(n18528), .A(n18484), .B(n18483), .ZN(
        P3_U2922) );
  AOI22_X1 U21610 ( .A1(n18761), .A2(n18485), .B1(n18766), .B2(n9798), .ZN(
        n18488) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18486), .B1(
        n18765), .B2(n18554), .ZN(n18487) );
  OAI211_X1 U21612 ( .C1(n18703), .C2(n18489), .A(n18488), .B(n18487), .ZN(
        P3_U2923) );
  NAND3_X1 U21613 ( .A1(n18491), .A2(n18705), .A3(n18490), .ZN(n18511) );
  NOR2_X1 U21614 ( .A1(n18492), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18538) );
  INV_X1 U21615 ( .A(n18538), .ZN(n18493) );
  NOR2_X1 U21616 ( .A1(n18849), .A2(n18493), .ZN(n18510) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18511), .B1(
        n18710), .B2(n18510), .ZN(n18495) );
  NOR2_X2 U21618 ( .A1(n18819), .A2(n18493), .ZN(n18579) );
  AOI22_X1 U21619 ( .A1(n18712), .A2(n18579), .B1(n18713), .B2(n9798), .ZN(
        n18494) );
  OAI211_X1 U21620 ( .C1(n18678), .C2(n18536), .A(n18495), .B(n18494), .ZN(
        P3_U2924) );
  INV_X1 U21621 ( .A(n18579), .ZN(n18588) );
  AOI22_X1 U21622 ( .A1(n18720), .A2(n9798), .B1(n18717), .B2(n18510), .ZN(
        n18497) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18511), .B1(
        n18718), .B2(n18529), .ZN(n18496) );
  OAI211_X1 U21624 ( .C1(n18594), .C2(n18588), .A(n18497), .B(n18496), .ZN(
        P3_U2925) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18511), .B1(
        n18724), .B2(n18510), .ZN(n18499) );
  AOI22_X1 U21626 ( .A1(n18726), .A2(n18579), .B1(n18725), .B2(n18529), .ZN(
        n18498) );
  OAI211_X1 U21627 ( .C1(n18684), .C2(n18504), .A(n18499), .B(n18498), .ZN(
        P3_U2926) );
  AOI22_X1 U21628 ( .A1(n18734), .A2(n9798), .B1(n18731), .B2(n18510), .ZN(
        n18501) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18511), .B1(
        n18732), .B2(n18529), .ZN(n18500) );
  OAI211_X1 U21630 ( .C1(n18652), .C2(n18588), .A(n18501), .B(n18500), .ZN(
        P3_U2927) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18511), .B1(
        n18738), .B2(n18510), .ZN(n18503) );
  AOI22_X1 U21632 ( .A1(n18740), .A2(n18579), .B1(n18739), .B2(n18529), .ZN(
        n18502) );
  OAI211_X1 U21633 ( .C1(n18743), .C2(n18504), .A(n18503), .B(n18502), .ZN(
        P3_U2928) );
  AOI22_X1 U21634 ( .A1(n18747), .A2(n9798), .B1(n18745), .B2(n18510), .ZN(
        n18507) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18511), .B1(
        n18691), .B2(n18579), .ZN(n18506) );
  OAI211_X1 U21636 ( .C1(n18694), .C2(n18536), .A(n18507), .B(n18506), .ZN(
        P3_U2929) );
  AOI22_X1 U21637 ( .A1(n18754), .A2(n9798), .B1(n18753), .B2(n18510), .ZN(
        n18509) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18511), .B1(
        n18756), .B2(n18529), .ZN(n18508) );
  OAI211_X1 U21639 ( .C1(n18662), .C2(n18588), .A(n18509), .B(n18508), .ZN(
        P3_U2930) );
  AOI22_X1 U21640 ( .A1(n18762), .A2(n9798), .B1(n18761), .B2(n18510), .ZN(
        n18513) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18511), .B1(
        n18766), .B2(n18529), .ZN(n18512) );
  OAI211_X1 U21642 ( .C1(n18668), .C2(n18588), .A(n18513), .B(n18512), .ZN(
        P3_U2931) );
  INV_X1 U21643 ( .A(n18612), .ZN(n18558) );
  NOR2_X2 U21644 ( .A1(n18822), .A2(n18558), .ZN(n18603) );
  NOR2_X1 U21645 ( .A1(n18579), .A2(n18603), .ZN(n18562) );
  OAI21_X1 U21646 ( .B1(n18514), .B2(n18670), .A(n18562), .ZN(n18515) );
  OAI211_X1 U21647 ( .C1(n18603), .C2(n18954), .A(n18673), .B(n18515), .ZN(
        n18533) );
  NOR2_X1 U21648 ( .A1(n18849), .A2(n18562), .ZN(n18532) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18533), .B1(
        n18710), .B2(n18532), .ZN(n18517) );
  AOI22_X1 U21650 ( .A1(n18712), .A2(n18603), .B1(n18713), .B2(n18529), .ZN(
        n18516) );
  OAI211_X1 U21651 ( .C1(n18678), .C2(n18528), .A(n18517), .B(n18516), .ZN(
        P3_U2932) );
  INV_X1 U21652 ( .A(n18603), .ZN(n18610) );
  AOI22_X1 U21653 ( .A1(n18720), .A2(n18529), .B1(n18717), .B2(n18532), .ZN(
        n18519) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18533), .B1(
        n18718), .B2(n18554), .ZN(n18518) );
  OAI211_X1 U21655 ( .C1(n18594), .C2(n18610), .A(n18519), .B(n18518), .ZN(
        P3_U2933) );
  AOI22_X1 U21656 ( .A1(n18727), .A2(n18529), .B1(n18724), .B2(n18532), .ZN(
        n18521) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18533), .B1(
        n18725), .B2(n18554), .ZN(n18520) );
  OAI211_X1 U21658 ( .C1(n18649), .C2(n18610), .A(n18521), .B(n18520), .ZN(
        P3_U2934) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18533), .B1(
        n18731), .B2(n18532), .ZN(n18523) );
  AOI22_X1 U21660 ( .A1(n18733), .A2(n18603), .B1(n18732), .B2(n18554), .ZN(
        n18522) );
  OAI211_X1 U21661 ( .C1(n18687), .C2(n18536), .A(n18523), .B(n18522), .ZN(
        P3_U2935) );
  AOI22_X1 U21662 ( .A1(n18653), .A2(n18529), .B1(n18738), .B2(n18532), .ZN(
        n18525) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18533), .B1(
        n18739), .B2(n18554), .ZN(n18524) );
  OAI211_X1 U21664 ( .C1(n18656), .C2(n18610), .A(n18525), .B(n18524), .ZN(
        P3_U2936) );
  AOI22_X1 U21665 ( .A1(n18747), .A2(n18529), .B1(n18745), .B2(n18532), .ZN(
        n18527) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18533), .B1(
        n18691), .B2(n18603), .ZN(n18526) );
  OAI211_X1 U21667 ( .C1(n18694), .C2(n18528), .A(n18527), .B(n18526), .ZN(
        P3_U2937) );
  AOI22_X1 U21668 ( .A1(n18754), .A2(n18529), .B1(n18753), .B2(n18532), .ZN(
        n18531) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18533), .B1(
        n18756), .B2(n18554), .ZN(n18530) );
  OAI211_X1 U21670 ( .C1(n18662), .C2(n18610), .A(n18531), .B(n18530), .ZN(
        P3_U2938) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18533), .B1(
        n18761), .B2(n18532), .ZN(n18535) );
  AOI22_X1 U21672 ( .A1(n18765), .A2(n18603), .B1(n18766), .B2(n18554), .ZN(
        n18534) );
  OAI211_X1 U21673 ( .C1(n18703), .C2(n18536), .A(n18535), .B(n18534), .ZN(
        P3_U2939) );
  NAND2_X1 U21674 ( .A1(n18612), .A2(n18537), .ZN(n18631) );
  AOI22_X1 U21675 ( .A1(n18711), .A2(n18579), .B1(n18710), .B2(n18553), .ZN(
        n18540) );
  AOI22_X1 U21676 ( .A1(n18708), .A2(n18538), .B1(n18612), .B2(n18638), .ZN(
        n18555) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18555), .B1(
        n18713), .B2(n18554), .ZN(n18539) );
  OAI211_X1 U21678 ( .C1(n18643), .C2(n18631), .A(n18540), .B(n18539), .ZN(
        P3_U2940) );
  AOI22_X1 U21679 ( .A1(n18717), .A2(n18553), .B1(n18718), .B2(n18579), .ZN(
        n18542) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18555), .B1(
        n18720), .B2(n18554), .ZN(n18541) );
  OAI211_X1 U21681 ( .C1(n18594), .C2(n18631), .A(n18542), .B(n18541), .ZN(
        P3_U2941) );
  AOI22_X1 U21682 ( .A1(n18725), .A2(n18579), .B1(n18724), .B2(n18553), .ZN(
        n18544) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18555), .B1(
        n18727), .B2(n18554), .ZN(n18543) );
  OAI211_X1 U21684 ( .C1(n18649), .C2(n18631), .A(n18544), .B(n18543), .ZN(
        P3_U2942) );
  AOI22_X1 U21685 ( .A1(n18734), .A2(n18554), .B1(n18731), .B2(n18553), .ZN(
        n18546) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18555), .B1(
        n18732), .B2(n18579), .ZN(n18545) );
  OAI211_X1 U21687 ( .C1(n18652), .C2(n18631), .A(n18546), .B(n18545), .ZN(
        P3_U2943) );
  AOI22_X1 U21688 ( .A1(n18653), .A2(n18554), .B1(n18738), .B2(n18553), .ZN(
        n18548) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18555), .B1(
        n18739), .B2(n18579), .ZN(n18547) );
  OAI211_X1 U21690 ( .C1(n18656), .C2(n18631), .A(n18548), .B(n18547), .ZN(
        P3_U2944) );
  AOI22_X1 U21691 ( .A1(n18747), .A2(n18554), .B1(n18745), .B2(n18553), .ZN(
        n18550) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18555), .B1(
        n18746), .B2(n18579), .ZN(n18549) );
  OAI211_X1 U21693 ( .C1(n18752), .C2(n18631), .A(n18550), .B(n18549), .ZN(
        P3_U2945) );
  AOI22_X1 U21694 ( .A1(n18754), .A2(n18554), .B1(n18753), .B2(n18553), .ZN(
        n18552) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18555), .B1(
        n18756), .B2(n18579), .ZN(n18551) );
  OAI211_X1 U21696 ( .C1(n18662), .C2(n18631), .A(n18552), .B(n18551), .ZN(
        P3_U2946) );
  AOI22_X1 U21697 ( .A1(n18761), .A2(n18553), .B1(n18766), .B2(n18579), .ZN(
        n18557) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18555), .B1(
        n18762), .B2(n18554), .ZN(n18556) );
  OAI211_X1 U21699 ( .C1(n18668), .C2(n18631), .A(n18557), .B(n18556), .ZN(
        P3_U2947) );
  INV_X1 U21700 ( .A(n18631), .ZN(n18633) );
  NOR2_X1 U21701 ( .A1(n18559), .A2(n18558), .ZN(n18657) );
  INV_X1 U21702 ( .A(n18657), .ZN(n18646) );
  NOR2_X1 U21703 ( .A1(n18633), .A2(n18664), .ZN(n18561) );
  AOI221_X1 U21704 ( .B1(n18562), .B2(n18561), .C1(n18670), .C2(n18561), .A(
        n18560), .ZN(n18583) );
  AOI21_X1 U21705 ( .B1(n18631), .B2(n18646), .A(n18849), .ZN(n18584) );
  AOI22_X1 U21706 ( .A1(n18711), .A2(n18603), .B1(n18710), .B2(n18584), .ZN(
        n18564) );
  AOI22_X1 U21707 ( .A1(n18712), .A2(n18664), .B1(n18713), .B2(n18579), .ZN(
        n18563) );
  OAI211_X1 U21708 ( .C1(n18583), .C2(n18565), .A(n18564), .B(n18563), .ZN(
        P3_U2948) );
  AOI22_X1 U21709 ( .A1(n18717), .A2(n18584), .B1(n18718), .B2(n18603), .ZN(
        n18567) );
  AOI22_X1 U21710 ( .A1(n18720), .A2(n18579), .B1(n18719), .B2(n18657), .ZN(
        n18566) );
  OAI211_X1 U21711 ( .C1(n18583), .C2(n18568), .A(n18567), .B(n18566), .ZN(
        P3_U2949) );
  AOI22_X1 U21712 ( .A1(n18725), .A2(n18603), .B1(n18724), .B2(n18584), .ZN(
        n18570) );
  INV_X1 U21713 ( .A(n18583), .ZN(n18585) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18585), .B1(
        n18726), .B2(n18664), .ZN(n18569) );
  OAI211_X1 U21715 ( .C1(n18684), .C2(n18588), .A(n18570), .B(n18569), .ZN(
        P3_U2950) );
  AOI22_X1 U21716 ( .A1(n18732), .A2(n18603), .B1(n18731), .B2(n18584), .ZN(
        n18572) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18585), .B1(
        n18733), .B2(n18657), .ZN(n18571) );
  OAI211_X1 U21718 ( .C1(n18687), .C2(n18588), .A(n18572), .B(n18571), .ZN(
        P3_U2951) );
  AOI22_X1 U21719 ( .A1(n18739), .A2(n18603), .B1(n18738), .B2(n18584), .ZN(
        n18574) );
  AOI22_X1 U21720 ( .A1(n18653), .A2(n18579), .B1(n18740), .B2(n18657), .ZN(
        n18573) );
  OAI211_X1 U21721 ( .C1(n18583), .C2(n18575), .A(n18574), .B(n18573), .ZN(
        P3_U2952) );
  AOI22_X1 U21722 ( .A1(n18746), .A2(n18603), .B1(n18745), .B2(n18584), .ZN(
        n18577) );
  AOI22_X1 U21723 ( .A1(n18691), .A2(n18664), .B1(n18747), .B2(n18579), .ZN(
        n18576) );
  OAI211_X1 U21724 ( .C1(n18583), .C2(n18578), .A(n18577), .B(n18576), .ZN(
        P3_U2953) );
  AOI22_X1 U21725 ( .A1(n18754), .A2(n18579), .B1(n18753), .B2(n18584), .ZN(
        n18581) );
  AOI22_X1 U21726 ( .A1(n18755), .A2(n18664), .B1(n18756), .B2(n18603), .ZN(
        n18580) );
  OAI211_X1 U21727 ( .C1(n18583), .C2(n18582), .A(n18581), .B(n18580), .ZN(
        P3_U2954) );
  AOI22_X1 U21728 ( .A1(n18761), .A2(n18584), .B1(n18766), .B2(n18603), .ZN(
        n18587) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18585), .B1(
        n18765), .B2(n18657), .ZN(n18586) );
  OAI211_X1 U21730 ( .C1(n18703), .C2(n18588), .A(n18587), .B(n18586), .ZN(
        P3_U2955) );
  NAND2_X1 U21731 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18612), .ZN(
        n18589) );
  NOR2_X2 U21732 ( .A1(n18819), .A2(n18589), .ZN(n18690) );
  NOR2_X1 U21733 ( .A1(n18849), .A2(n18589), .ZN(n18606) );
  AOI22_X1 U21734 ( .A1(n18711), .A2(n18633), .B1(n18710), .B2(n18606), .ZN(
        n18591) );
  INV_X1 U21735 ( .A(n18589), .ZN(n18640) );
  AOI22_X1 U21736 ( .A1(n18708), .A2(n18612), .B1(n18640), .B2(n18705), .ZN(
        n18607) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18607), .B1(
        n18713), .B2(n18603), .ZN(n18590) );
  OAI211_X1 U21738 ( .C1(n18704), .C2(n18643), .A(n18591), .B(n18590), .ZN(
        P3_U2956) );
  AOI22_X1 U21739 ( .A1(n18720), .A2(n18603), .B1(n18717), .B2(n18606), .ZN(
        n18593) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18607), .B1(
        n18718), .B2(n18633), .ZN(n18592) );
  OAI211_X1 U21741 ( .C1(n18704), .C2(n18594), .A(n18593), .B(n18592), .ZN(
        P3_U2957) );
  AOI22_X1 U21742 ( .A1(n18725), .A2(n18633), .B1(n18724), .B2(n18606), .ZN(
        n18596) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18607), .B1(
        n18690), .B2(n18726), .ZN(n18595) );
  OAI211_X1 U21744 ( .C1(n18684), .C2(n18610), .A(n18596), .B(n18595), .ZN(
        P3_U2958) );
  AOI22_X1 U21745 ( .A1(n18732), .A2(n18633), .B1(n18731), .B2(n18606), .ZN(
        n18598) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18607), .B1(
        n18690), .B2(n18733), .ZN(n18597) );
  OAI211_X1 U21747 ( .C1(n18687), .C2(n18610), .A(n18598), .B(n18597), .ZN(
        P3_U2959) );
  AOI22_X1 U21748 ( .A1(n18653), .A2(n18603), .B1(n18738), .B2(n18606), .ZN(
        n18600) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18607), .B1(
        n18739), .B2(n18633), .ZN(n18599) );
  OAI211_X1 U21750 ( .C1(n18704), .C2(n18656), .A(n18600), .B(n18599), .ZN(
        P3_U2960) );
  AOI22_X1 U21751 ( .A1(n18747), .A2(n18603), .B1(n18745), .B2(n18606), .ZN(
        n18602) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18607), .B1(
        n18690), .B2(n18691), .ZN(n18601) );
  OAI211_X1 U21753 ( .C1(n18694), .C2(n18631), .A(n18602), .B(n18601), .ZN(
        P3_U2961) );
  AOI22_X1 U21754 ( .A1(n18754), .A2(n18603), .B1(n18753), .B2(n18606), .ZN(
        n18605) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18607), .B1(
        n18756), .B2(n18633), .ZN(n18604) );
  OAI211_X1 U21756 ( .C1(n18704), .C2(n18662), .A(n18605), .B(n18604), .ZN(
        P3_U2962) );
  AOI22_X1 U21757 ( .A1(n18761), .A2(n18606), .B1(n18766), .B2(n18633), .ZN(
        n18609) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18607), .B1(
        n18690), .B2(n18765), .ZN(n18608) );
  OAI211_X1 U21759 ( .C1(n18703), .C2(n18610), .A(n18609), .B(n18608), .ZN(
        P3_U2963) );
  NAND2_X1 U21760 ( .A1(n18707), .A2(n18819), .ZN(n18744) );
  NOR2_X1 U21761 ( .A1(n18763), .A2(n18690), .ZN(n18672) );
  NOR2_X1 U21762 ( .A1(n18849), .A2(n18672), .ZN(n18632) );
  AOI22_X1 U21763 ( .A1(n18713), .A2(n18633), .B1(n18710), .B2(n18632), .ZN(
        n18618) );
  INV_X1 U21764 ( .A(n18611), .ZN(n18615) );
  NAND2_X1 U21765 ( .A1(n18613), .A2(n18612), .ZN(n18614) );
  OAI21_X1 U21766 ( .B1(n18615), .B2(n18614), .A(n18672), .ZN(n18616) );
  OAI211_X1 U21767 ( .C1(n18763), .C2(n18954), .A(n18673), .B(n18616), .ZN(
        n18634) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18634), .B1(
        n18763), .B2(n18712), .ZN(n18617) );
  OAI211_X1 U21769 ( .C1(n18678), .C2(n18646), .A(n18618), .B(n18617), .ZN(
        P3_U2964) );
  AOI22_X1 U21770 ( .A1(n18717), .A2(n18632), .B1(n18718), .B2(n18664), .ZN(
        n18620) );
  AOI22_X1 U21771 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18634), .B1(
        n18763), .B2(n18719), .ZN(n18619) );
  OAI211_X1 U21772 ( .C1(n18681), .C2(n18631), .A(n18620), .B(n18619), .ZN(
        P3_U2965) );
  AOI22_X1 U21773 ( .A1(n18725), .A2(n18664), .B1(n18724), .B2(n18632), .ZN(
        n18622) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18634), .B1(
        n18763), .B2(n18726), .ZN(n18621) );
  OAI211_X1 U21775 ( .C1(n18684), .C2(n18631), .A(n18622), .B(n18621), .ZN(
        P3_U2966) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18634), .B1(
        n18731), .B2(n18632), .ZN(n18624) );
  AOI22_X1 U21777 ( .A1(n18763), .A2(n18733), .B1(n18732), .B2(n18657), .ZN(
        n18623) );
  OAI211_X1 U21778 ( .C1(n18687), .C2(n18631), .A(n18624), .B(n18623), .ZN(
        P3_U2967) );
  AOI22_X1 U21779 ( .A1(n18739), .A2(n18664), .B1(n18738), .B2(n18632), .ZN(
        n18626) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18634), .B1(
        n18763), .B2(n18740), .ZN(n18625) );
  OAI211_X1 U21781 ( .C1(n18743), .C2(n18631), .A(n18626), .B(n18625), .ZN(
        P3_U2968) );
  AOI22_X1 U21782 ( .A1(n18746), .A2(n18664), .B1(n18745), .B2(n18632), .ZN(
        n18628) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18634), .B1(
        n18747), .B2(n18633), .ZN(n18627) );
  OAI211_X1 U21784 ( .C1(n18744), .C2(n18752), .A(n18628), .B(n18627), .ZN(
        P3_U2969) );
  AOI22_X1 U21785 ( .A1(n18756), .A2(n18657), .B1(n18753), .B2(n18632), .ZN(
        n18630) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18634), .B1(
        n18763), .B2(n18755), .ZN(n18629) );
  OAI211_X1 U21787 ( .C1(n18697), .C2(n18631), .A(n18630), .B(n18629), .ZN(
        P3_U2970) );
  AOI22_X1 U21788 ( .A1(n18762), .A2(n18633), .B1(n18761), .B2(n18632), .ZN(
        n18636) );
  AOI22_X1 U21789 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18634), .B1(
        n18766), .B2(n18664), .ZN(n18635) );
  OAI211_X1 U21790 ( .C1(n18744), .C2(n18668), .A(n18636), .B(n18635), .ZN(
        P3_U2971) );
  INV_X1 U21791 ( .A(n18707), .ZN(n18637) );
  NOR2_X1 U21792 ( .A1(n18849), .A2(n18637), .ZN(n18663) );
  AOI22_X1 U21793 ( .A1(n18690), .A2(n18711), .B1(n18710), .B2(n18663), .ZN(
        n18642) );
  AOI22_X1 U21794 ( .A1(n18708), .A2(n18640), .B1(n18639), .B2(n18638), .ZN(
        n18665) );
  AOI22_X1 U21795 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18665), .B1(
        n18713), .B2(n18657), .ZN(n18641) );
  OAI211_X1 U21796 ( .C1(n18671), .C2(n18643), .A(n18642), .B(n18641), .ZN(
        P3_U2972) );
  AOI22_X1 U21797 ( .A1(n18690), .A2(n18718), .B1(n18717), .B2(n18663), .ZN(
        n18645) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18665), .B1(
        n18767), .B2(n18719), .ZN(n18644) );
  OAI211_X1 U21799 ( .C1(n18681), .C2(n18646), .A(n18645), .B(n18644), .ZN(
        P3_U2973) );
  AOI22_X1 U21800 ( .A1(n18727), .A2(n18664), .B1(n18724), .B2(n18663), .ZN(
        n18648) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18665), .B1(
        n18690), .B2(n18725), .ZN(n18647) );
  OAI211_X1 U21802 ( .C1(n18671), .C2(n18649), .A(n18648), .B(n18647), .ZN(
        P3_U2974) );
  AOI22_X1 U21803 ( .A1(n18734), .A2(n18664), .B1(n18731), .B2(n18663), .ZN(
        n18651) );
  AOI22_X1 U21804 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18665), .B1(
        n18690), .B2(n18732), .ZN(n18650) );
  OAI211_X1 U21805 ( .C1(n18671), .C2(n18652), .A(n18651), .B(n18650), .ZN(
        P3_U2975) );
  AOI22_X1 U21806 ( .A1(n18653), .A2(n18664), .B1(n18738), .B2(n18663), .ZN(
        n18655) );
  AOI22_X1 U21807 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18665), .B1(
        n18690), .B2(n18739), .ZN(n18654) );
  OAI211_X1 U21808 ( .C1(n18671), .C2(n18656), .A(n18655), .B(n18654), .ZN(
        P3_U2976) );
  AOI22_X1 U21809 ( .A1(n18690), .A2(n18746), .B1(n18745), .B2(n18663), .ZN(
        n18659) );
  AOI22_X1 U21810 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18665), .B1(
        n18747), .B2(n18657), .ZN(n18658) );
  OAI211_X1 U21811 ( .C1(n18671), .C2(n18752), .A(n18659), .B(n18658), .ZN(
        P3_U2977) );
  AOI22_X1 U21812 ( .A1(n18754), .A2(n18664), .B1(n18753), .B2(n18663), .ZN(
        n18661) );
  AOI22_X1 U21813 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18665), .B1(
        n18690), .B2(n18756), .ZN(n18660) );
  OAI211_X1 U21814 ( .C1(n18671), .C2(n18662), .A(n18661), .B(n18660), .ZN(
        P3_U2978) );
  AOI22_X1 U21815 ( .A1(n18762), .A2(n18664), .B1(n18761), .B2(n18663), .ZN(
        n18667) );
  AOI22_X1 U21816 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18665), .B1(
        n18690), .B2(n18766), .ZN(n18666) );
  OAI211_X1 U21817 ( .C1(n18671), .C2(n18668), .A(n18667), .B(n18666), .ZN(
        P3_U2979) );
  NOR2_X1 U21818 ( .A1(n18849), .A2(n18669), .ZN(n18698) );
  AOI22_X1 U21819 ( .A1(n18690), .A2(n18713), .B1(n18710), .B2(n18698), .ZN(
        n18677) );
  AOI221_X1 U21820 ( .B1(n18672), .B2(n18671), .C1(n18670), .C2(n18671), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18674) );
  OAI21_X1 U21821 ( .B1(n18675), .B2(n18674), .A(n18673), .ZN(n18700) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18700), .B1(
        n18699), .B2(n18712), .ZN(n18676) );
  OAI211_X1 U21823 ( .C1(n18744), .C2(n18678), .A(n18677), .B(n18676), .ZN(
        P3_U2980) );
  AOI22_X1 U21824 ( .A1(n18763), .A2(n18718), .B1(n18698), .B2(n18717), .ZN(
        n18680) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18700), .B1(
        n18699), .B2(n18719), .ZN(n18679) );
  OAI211_X1 U21826 ( .C1(n18704), .C2(n18681), .A(n18680), .B(n18679), .ZN(
        P3_U2981) );
  AOI22_X1 U21827 ( .A1(n18763), .A2(n18725), .B1(n18698), .B2(n18724), .ZN(
        n18683) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18700), .B1(
        n18699), .B2(n18726), .ZN(n18682) );
  OAI211_X1 U21829 ( .C1(n18704), .C2(n18684), .A(n18683), .B(n18682), .ZN(
        P3_U2982) );
  AOI22_X1 U21830 ( .A1(n18763), .A2(n18732), .B1(n18698), .B2(n18731), .ZN(
        n18686) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18700), .B1(
        n18699), .B2(n18733), .ZN(n18685) );
  OAI211_X1 U21832 ( .C1(n18704), .C2(n18687), .A(n18686), .B(n18685), .ZN(
        P3_U2983) );
  AOI22_X1 U21833 ( .A1(n18763), .A2(n18739), .B1(n18698), .B2(n18738), .ZN(
        n18689) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18700), .B1(
        n18699), .B2(n18740), .ZN(n18688) );
  OAI211_X1 U21835 ( .C1(n18704), .C2(n18743), .A(n18689), .B(n18688), .ZN(
        P3_U2984) );
  AOI22_X1 U21836 ( .A1(n18690), .A2(n18747), .B1(n18698), .B2(n18745), .ZN(
        n18693) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18700), .B1(
        n18699), .B2(n18691), .ZN(n18692) );
  OAI211_X1 U21838 ( .C1(n18744), .C2(n18694), .A(n18693), .B(n18692), .ZN(
        P3_U2985) );
  AOI22_X1 U21839 ( .A1(n18763), .A2(n18756), .B1(n18698), .B2(n18753), .ZN(
        n18696) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18700), .B1(
        n18699), .B2(n18755), .ZN(n18695) );
  OAI211_X1 U21841 ( .C1(n18704), .C2(n18697), .A(n18696), .B(n18695), .ZN(
        P3_U2986) );
  AOI22_X1 U21842 ( .A1(n18763), .A2(n18766), .B1(n18698), .B2(n18761), .ZN(
        n18702) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18700), .B1(
        n18699), .B2(n18765), .ZN(n18701) );
  OAI211_X1 U21844 ( .C1(n18704), .C2(n18703), .A(n18702), .B(n18701), .ZN(
        P3_U2987) );
  AOI22_X1 U21845 ( .A1(n18708), .A2(n18707), .B1(n18706), .B2(n18705), .ZN(
        n18748) );
  INV_X1 U21846 ( .A(n18748), .ZN(n18770) );
  NOR2_X1 U21847 ( .A1(n18849), .A2(n18709), .ZN(n18760) );
  AOI22_X1 U21848 ( .A1(n18767), .A2(n18711), .B1(n18710), .B2(n18760), .ZN(
        n18715) );
  AOI22_X1 U21849 ( .A1(n18763), .A2(n18713), .B1(n18712), .B2(n18764), .ZN(
        n18714) );
  OAI211_X1 U21850 ( .C1(n18716), .C2(n18770), .A(n18715), .B(n18714), .ZN(
        P3_U2988) );
  AOI22_X1 U21851 ( .A1(n18767), .A2(n18718), .B1(n18717), .B2(n18760), .ZN(
        n18722) );
  AOI22_X1 U21852 ( .A1(n18763), .A2(n18720), .B1(n18719), .B2(n18764), .ZN(
        n18721) );
  OAI211_X1 U21853 ( .C1(n18723), .C2(n18770), .A(n18722), .B(n18721), .ZN(
        P3_U2989) );
  AOI22_X1 U21854 ( .A1(n18767), .A2(n18725), .B1(n18724), .B2(n18760), .ZN(
        n18729) );
  AOI22_X1 U21855 ( .A1(n18763), .A2(n18727), .B1(n18726), .B2(n18764), .ZN(
        n18728) );
  OAI211_X1 U21856 ( .C1(n18730), .C2(n18770), .A(n18729), .B(n18728), .ZN(
        P3_U2990) );
  AOI22_X1 U21857 ( .A1(n18767), .A2(n18732), .B1(n18731), .B2(n18760), .ZN(
        n18736) );
  AOI22_X1 U21858 ( .A1(n18763), .A2(n18734), .B1(n18733), .B2(n18764), .ZN(
        n18735) );
  OAI211_X1 U21859 ( .C1(n18737), .C2(n18770), .A(n18736), .B(n18735), .ZN(
        P3_U2991) );
  AOI22_X1 U21860 ( .A1(n18767), .A2(n18739), .B1(n18738), .B2(n18760), .ZN(
        n18742) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18748), .B1(
        n18740), .B2(n18764), .ZN(n18741) );
  OAI211_X1 U21862 ( .C1(n18744), .C2(n18743), .A(n18742), .B(n18741), .ZN(
        P3_U2992) );
  AOI22_X1 U21863 ( .A1(n18767), .A2(n18746), .B1(n18745), .B2(n18760), .ZN(
        n18750) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18748), .B1(
        n18763), .B2(n18747), .ZN(n18749) );
  OAI211_X1 U21865 ( .C1(n18752), .C2(n18751), .A(n18750), .B(n18749), .ZN(
        P3_U2993) );
  AOI22_X1 U21866 ( .A1(n18763), .A2(n18754), .B1(n18753), .B2(n18760), .ZN(
        n18758) );
  AOI22_X1 U21867 ( .A1(n18767), .A2(n18756), .B1(n18755), .B2(n18764), .ZN(
        n18757) );
  OAI211_X1 U21868 ( .C1(n18759), .C2(n18770), .A(n18758), .B(n18757), .ZN(
        P3_U2994) );
  AOI22_X1 U21869 ( .A1(n18763), .A2(n18762), .B1(n18761), .B2(n18760), .ZN(
        n18769) );
  AOI22_X1 U21870 ( .A1(n18767), .A2(n18766), .B1(n18765), .B2(n18764), .ZN(
        n18768) );
  OAI211_X1 U21871 ( .C1(n18771), .C2(n18770), .A(n18769), .B(n18768), .ZN(
        P3_U2995) );
  AOI21_X1 U21872 ( .B1(n18809), .B2(n18773), .A(n18772), .ZN(n18774) );
  AOI21_X1 U21873 ( .B1(n18776), .B2(n18775), .A(n18774), .ZN(n18777) );
  OAI21_X1 U21874 ( .B1(n18779), .B2(n18778), .A(n18777), .ZN(n19000) );
  OAI21_X1 U21875 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18780), .ZN(n18781) );
  OAI211_X1 U21876 ( .C1(n18783), .C2(n18813), .A(n18782), .B(n18781), .ZN(
        n18835) );
  NOR2_X1 U21877 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18796), .ZN(
        n18817) );
  OAI22_X1 U21878 ( .A1(n18802), .A2(n18817), .B1(n18809), .B2(n18784), .ZN(
        n18785) );
  INV_X1 U21879 ( .A(n18785), .ZN(n18957) );
  NOR2_X1 U21880 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18957), .ZN(
        n18798) );
  INV_X1 U21881 ( .A(n18786), .ZN(n18787) );
  OAI22_X1 U21882 ( .A1(n18790), .A2(n18789), .B1(n18788), .B2(n18787), .ZN(
        n18791) );
  NOR2_X1 U21883 ( .A1(n18792), .A2(n18791), .ZN(n18800) );
  OAI21_X1 U21884 ( .B1(n18794), .B2(n18800), .A(n18793), .ZN(n18795) );
  AOI21_X1 U21885 ( .B1(n18802), .B2(n18796), .A(n18795), .ZN(n18960) );
  NAND2_X1 U21886 ( .A1(n18813), .A2(n18960), .ZN(n18797) );
  AOI22_X1 U21887 ( .A1(n18813), .A2(n18798), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18797), .ZN(n18833) );
  INV_X1 U21888 ( .A(n18813), .ZN(n18824) );
  NOR2_X1 U21889 ( .A1(n18799), .A2(n18972), .ZN(n18812) );
  OAI21_X1 U21890 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18801), .A(
        n18800), .ZN(n18811) );
  OAI211_X1 U21891 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18803), .B(n18802), .ZN(
        n18808) );
  NOR2_X1 U21892 ( .A1(n18804), .A2(n18987), .ZN(n18806) );
  OAI211_X1 U21893 ( .C1(n18806), .C2(n18805), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18972), .ZN(n18807) );
  OAI211_X1 U21894 ( .C1(n18969), .C2(n18809), .A(n18808), .B(n18807), .ZN(
        n18810) );
  AOI21_X1 U21895 ( .B1(n18812), .B2(n18811), .A(n18810), .ZN(n18965) );
  AOI22_X1 U21896 ( .A1(n18824), .A2(n18972), .B1(n18965), .B2(n18813), .ZN(
        n18828) );
  NOR2_X1 U21897 ( .A1(n9824), .A2(n18814), .ZN(n18818) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18816), .B1(
        n18818), .B2(n18987), .ZN(n18982) );
  OAI22_X1 U21899 ( .A1(n18818), .A2(n18973), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18817), .ZN(n18978) );
  OR3_X1 U21900 ( .A1(n18982), .A2(n18821), .A3(n18819), .ZN(n18820) );
  AOI22_X1 U21901 ( .A1(n18982), .A2(n18821), .B1(n18978), .B2(n18820), .ZN(
        n18823) );
  OAI21_X1 U21902 ( .B1(n18824), .B2(n18823), .A(n18822), .ZN(n18827) );
  AND2_X1 U21903 ( .A1(n18828), .A2(n18827), .ZN(n18825) );
  OAI221_X1 U21904 ( .B1(n18828), .B2(n18827), .C1(n18826), .C2(n18825), .A(
        n18830), .ZN(n18832) );
  AOI21_X1 U21905 ( .B1(n18830), .B2(n18829), .A(n18828), .ZN(n18831) );
  AOI222_X1 U21906 ( .A1(n18833), .A2(n18832), .B1(n18833), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18832), .C2(n18831), .ZN(
        n18834) );
  NOR4_X1 U21907 ( .A1(n18836), .A2(n19000), .A3(n18835), .A4(n18834), .ZN(
        n18847) );
  NOR2_X1 U21908 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19011) );
  AOI22_X1 U21909 ( .A1(n18981), .A2(n19011), .B1(n18860), .B2(n19001), .ZN(
        n18837) );
  INV_X1 U21910 ( .A(n18837), .ZN(n18843) );
  OAI211_X1 U21911 ( .C1(n18839), .C2(n18838), .A(n19004), .B(n18847), .ZN(
        n18953) );
  NAND2_X1 U21912 ( .A1(n18860), .A2(n18840), .ZN(n18854) );
  NAND2_X1 U21913 ( .A1(n18953), .A2(n18854), .ZN(n18848) );
  NOR2_X1 U21914 ( .A1(n18841), .A2(n18848), .ZN(n18842) );
  MUX2_X1 U21915 ( .A(n18843), .B(n18842), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18845) );
  OAI211_X1 U21916 ( .C1(n18847), .C2(n18846), .A(n18845), .B(n18844), .ZN(
        P3_U2996) );
  NOR2_X1 U21917 ( .A1(n18849), .A2(n18848), .ZN(n18850) );
  AOI22_X1 U21918 ( .A1(n18851), .A2(n18850), .B1(n18860), .B2(n19001), .ZN(
        n18853) );
  OAI211_X1 U21919 ( .C1(n18854), .C2(n18856), .A(n18853), .B(n18852), .ZN(
        P3_U2997) );
  INV_X1 U21920 ( .A(n18952), .ZN(n18859) );
  AOI221_X1 U21921 ( .B1(n18857), .B2(n19009), .C1(n18856), .C2(n18855), .A(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18858) );
  NOR2_X1 U21922 ( .A1(n18859), .A2(n18858), .ZN(P3_U2998) );
  AND2_X1 U21923 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18948), .ZN(
        P3_U2999) );
  AND2_X1 U21924 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18948), .ZN(
        P3_U3000) );
  AND2_X1 U21925 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18948), .ZN(
        P3_U3001) );
  AND2_X1 U21926 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18948), .ZN(
        P3_U3002) );
  AND2_X1 U21927 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18948), .ZN(
        P3_U3003) );
  AND2_X1 U21928 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18948), .ZN(
        P3_U3004) );
  AND2_X1 U21929 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18948), .ZN(
        P3_U3005) );
  AND2_X1 U21930 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18948), .ZN(
        P3_U3006) );
  AND2_X1 U21931 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18948), .ZN(
        P3_U3007) );
  AND2_X1 U21932 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18948), .ZN(
        P3_U3008) );
  AND2_X1 U21933 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18948), .ZN(
        P3_U3009) );
  AND2_X1 U21934 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18948), .ZN(
        P3_U3010) );
  AND2_X1 U21935 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18948), .ZN(
        P3_U3011) );
  AND2_X1 U21936 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18948), .ZN(
        P3_U3012) );
  AND2_X1 U21937 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18948), .ZN(
        P3_U3013) );
  AND2_X1 U21938 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18948), .ZN(
        P3_U3014) );
  AND2_X1 U21939 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18948), .ZN(
        P3_U3015) );
  AND2_X1 U21940 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18948), .ZN(
        P3_U3016) );
  AND2_X1 U21941 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18948), .ZN(
        P3_U3017) );
  AND2_X1 U21942 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18948), .ZN(
        P3_U3018) );
  AND2_X1 U21943 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18948), .ZN(
        P3_U3019) );
  AND2_X1 U21944 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18948), .ZN(
        P3_U3020) );
  AND2_X1 U21945 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18948), .ZN(P3_U3021) );
  AND2_X1 U21946 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18948), .ZN(P3_U3022) );
  AND2_X1 U21947 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18948), .ZN(P3_U3023) );
  AND2_X1 U21948 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18948), .ZN(P3_U3024) );
  AND2_X1 U21949 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18948), .ZN(P3_U3025) );
  AND2_X1 U21950 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18948), .ZN(P3_U3026) );
  AND2_X1 U21951 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18948), .ZN(P3_U3027) );
  AND2_X1 U21952 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18948), .ZN(P3_U3028) );
  NAND2_X1 U21953 ( .A1(n18860), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18869) );
  OAI21_X1 U21954 ( .B1(n18861), .B2(n20842), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18863) );
  INV_X1 U21955 ( .A(NA), .ZN(n21006) );
  NOR3_X1 U21956 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .A3(n21006), .ZN(n18862) );
  AOI21_X1 U21957 ( .B1(n18997), .B2(n18863), .A(n18862), .ZN(n18864) );
  OAI221_X1 U21958 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(P3_STATE_REG_0__SCAN_IN), .C1(P3_STATE_REG_2__SCAN_IN), .C2(n18869), .A(n18864), .ZN(P3_U3029) );
  NOR2_X1 U21959 ( .A1(n18875), .A2(n20842), .ZN(n18871) );
  NOR2_X1 U21960 ( .A1(n18873), .A2(n18871), .ZN(n18865) );
  INV_X1 U21961 ( .A(n18869), .ZN(n18868) );
  AOI21_X1 U21962 ( .B1(n18865), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n18868), .ZN(n18866) );
  OAI211_X1 U21963 ( .C1(n20842), .C2(n18867), .A(n18866), .B(n19006), .ZN(
        P3_U3030) );
  AOI221_X1 U21964 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18873), .C1(n21006), 
        .C2(n18873), .A(n18868), .ZN(n18874) );
  OAI22_X1 U21965 ( .A1(NA), .A2(n18869), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18870) );
  OAI22_X1 U21966 ( .A1(n18871), .A2(n18870), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18872) );
  OAI22_X1 U21967 ( .A1(n18874), .A2(n18875), .B1(n18873), .B2(n18872), .ZN(
        P3_U3031) );
  INV_X1 U21968 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18877) );
  NAND2_X1 U21969 ( .A1(n18936), .A2(n18875), .ZN(n18933) );
  OAI222_X1 U21970 ( .A1(n18989), .A2(n18939), .B1(n18876), .B2(n18936), .C1(
        n18877), .C2(n18934), .ZN(P3_U3032) );
  OAI222_X1 U21971 ( .A1(n18934), .A2(n18879), .B1(n18878), .B2(n18936), .C1(
        n18877), .C2(n18939), .ZN(P3_U3033) );
  OAI222_X1 U21972 ( .A1(n18933), .A2(n18881), .B1(n18880), .B2(n18936), .C1(
        n18879), .C2(n18939), .ZN(P3_U3034) );
  INV_X1 U21973 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18883) );
  OAI222_X1 U21974 ( .A1(n18933), .A2(n18883), .B1(n18882), .B2(n18936), .C1(
        n18881), .C2(n18939), .ZN(P3_U3035) );
  OAI222_X1 U21975 ( .A1(n18933), .A2(n18885), .B1(n18884), .B2(n18936), .C1(
        n18883), .C2(n18939), .ZN(P3_U3036) );
  OAI222_X1 U21976 ( .A1(n18933), .A2(n18887), .B1(n18886), .B2(n18936), .C1(
        n18885), .C2(n18939), .ZN(P3_U3037) );
  OAI222_X1 U21977 ( .A1(n18933), .A2(n18889), .B1(n18888), .B2(n18936), .C1(
        n18887), .C2(n18939), .ZN(P3_U3038) );
  INV_X1 U21978 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18891) );
  OAI222_X1 U21979 ( .A1(n18934), .A2(n18891), .B1(n18890), .B2(n18936), .C1(
        n18889), .C2(n18939), .ZN(P3_U3039) );
  OAI222_X1 U21980 ( .A1(n18934), .A2(n18893), .B1(n18892), .B2(n18936), .C1(
        n18891), .C2(n18939), .ZN(P3_U3040) );
  INV_X1 U21981 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18895) );
  OAI222_X1 U21982 ( .A1(n18934), .A2(n18895), .B1(n18894), .B2(n18936), .C1(
        n18893), .C2(n18939), .ZN(P3_U3041) );
  OAI222_X1 U21983 ( .A1(n18934), .A2(n18897), .B1(n18896), .B2(n18936), .C1(
        n18895), .C2(n18939), .ZN(P3_U3042) );
  INV_X1 U21984 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18899) );
  OAI222_X1 U21985 ( .A1(n18934), .A2(n18899), .B1(n18898), .B2(n18936), .C1(
        n18897), .C2(n18939), .ZN(P3_U3043) );
  OAI222_X1 U21986 ( .A1(n18934), .A2(n18901), .B1(n18900), .B2(n18936), .C1(
        n18899), .C2(n18939), .ZN(P3_U3044) );
  OAI222_X1 U21987 ( .A1(n18933), .A2(n18903), .B1(n18902), .B2(n18936), .C1(
        n18901), .C2(n18939), .ZN(P3_U3045) );
  OAI222_X1 U21988 ( .A1(n18933), .A2(n18905), .B1(n18904), .B2(n18936), .C1(
        n18903), .C2(n18939), .ZN(P3_U3046) );
  INV_X1 U21989 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18907) );
  OAI222_X1 U21990 ( .A1(n18933), .A2(n18907), .B1(n18906), .B2(n18936), .C1(
        n18905), .C2(n18939), .ZN(P3_U3047) );
  OAI222_X1 U21991 ( .A1(n18933), .A2(n18909), .B1(n18908), .B2(n18936), .C1(
        n18907), .C2(n18939), .ZN(P3_U3048) );
  OAI222_X1 U21992 ( .A1(n18933), .A2(n18912), .B1(n18910), .B2(n18936), .C1(
        n18909), .C2(n18939), .ZN(P3_U3049) );
  OAI222_X1 U21993 ( .A1(n18912), .A2(n18939), .B1(n18911), .B2(n18936), .C1(
        n18913), .C2(n18934), .ZN(P3_U3050) );
  OAI222_X1 U21994 ( .A1(n18934), .A2(n18916), .B1(n18914), .B2(n18936), .C1(
        n18913), .C2(n18939), .ZN(P3_U3051) );
  INV_X1 U21995 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18917) );
  OAI222_X1 U21996 ( .A1(n18916), .A2(n18939), .B1(n18915), .B2(n18936), .C1(
        n18917), .C2(n18934), .ZN(P3_U3052) );
  OAI222_X1 U21997 ( .A1(n18934), .A2(n18920), .B1(n18918), .B2(n18936), .C1(
        n18917), .C2(n18939), .ZN(P3_U3053) );
  OAI222_X1 U21998 ( .A1(n18920), .A2(n18939), .B1(n18919), .B2(n18936), .C1(
        n18921), .C2(n18934), .ZN(P3_U3054) );
  OAI222_X1 U21999 ( .A1(n18933), .A2(n18923), .B1(n18922), .B2(n18936), .C1(
        n18921), .C2(n18939), .ZN(P3_U3055) );
  INV_X1 U22000 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18925) );
  OAI222_X1 U22001 ( .A1(n18934), .A2(n18925), .B1(n18924), .B2(n18936), .C1(
        n18923), .C2(n18939), .ZN(P3_U3056) );
  OAI222_X1 U22002 ( .A1(n18934), .A2(n18927), .B1(n18926), .B2(n18936), .C1(
        n18925), .C2(n18939), .ZN(P3_U3057) );
  OAI222_X1 U22003 ( .A1(n18934), .A2(n18930), .B1(n18928), .B2(n18936), .C1(
        n18927), .C2(n18939), .ZN(P3_U3058) );
  OAI222_X1 U22004 ( .A1(n18930), .A2(n18939), .B1(n18929), .B2(n18936), .C1(
        n18931), .C2(n18934), .ZN(P3_U3059) );
  OAI222_X1 U22005 ( .A1(n18933), .A2(n18938), .B1(n18932), .B2(n18936), .C1(
        n18931), .C2(n18939), .ZN(P3_U3060) );
  INV_X1 U22006 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18937) );
  OAI222_X1 U22007 ( .A1(n18939), .A2(n18938), .B1(n18937), .B2(n18936), .C1(
        n18935), .C2(n18934), .ZN(P3_U3061) );
  INV_X1 U22008 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18940) );
  AOI22_X1 U22009 ( .A1(n18936), .A2(n18941), .B1(n18940), .B2(n18997), .ZN(
        P3_U3274) );
  INV_X1 U22010 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18992) );
  INV_X1 U22011 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18942) );
  AOI22_X1 U22012 ( .A1(n18936), .A2(n18992), .B1(n18942), .B2(n18997), .ZN(
        P3_U3275) );
  INV_X1 U22013 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18943) );
  AOI22_X1 U22014 ( .A1(n18936), .A2(n18944), .B1(n18943), .B2(n18997), .ZN(
        P3_U3276) );
  INV_X1 U22015 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18995) );
  INV_X1 U22016 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18945) );
  AOI22_X1 U22017 ( .A1(n18936), .A2(n18995), .B1(n18945), .B2(n18997), .ZN(
        P3_U3277) );
  INV_X1 U22018 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18947) );
  INV_X1 U22019 ( .A(n18949), .ZN(n18946) );
  AOI21_X1 U22020 ( .B1(n18948), .B2(n18947), .A(n18946), .ZN(P3_U3280) );
  OAI21_X1 U22021 ( .B1(n18951), .B2(n18950), .A(n18949), .ZN(P3_U3281) );
  OAI221_X1 U22022 ( .B1(n18954), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18954), 
        .C2(n18953), .A(n18952), .ZN(P3_U3282) );
  INV_X1 U22023 ( .A(n18955), .ZN(n18959) );
  NOR3_X1 U22024 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18957), .A3(
        n18956), .ZN(n18958) );
  AOI21_X1 U22025 ( .B1(n18959), .B2(n18981), .A(n18958), .ZN(n18964) );
  INV_X1 U22026 ( .A(n18960), .ZN(n18961) );
  AOI21_X1 U22027 ( .B1(n18983), .B2(n18961), .A(n18988), .ZN(n18963) );
  OAI22_X1 U22028 ( .A1(n18988), .A2(n18964), .B1(n18963), .B2(n18962), .ZN(
        P3_U3285) );
  INV_X1 U22029 ( .A(n18965), .ZN(n18970) );
  NOR2_X1 U22030 ( .A1(n18966), .A2(n18984), .ZN(n18975) );
  AOI22_X1 U22031 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18968), .B2(n18967), .ZN(
        n18974) );
  AOI222_X1 U22032 ( .A1(n18970), .A2(n18983), .B1(n18975), .B2(n18974), .C1(
        n18981), .C2(n18969), .ZN(n18971) );
  AOI22_X1 U22033 ( .A1(n18988), .A2(n18972), .B1(n18971), .B2(n18985), .ZN(
        P3_U3288) );
  INV_X1 U22034 ( .A(n18973), .ZN(n18977) );
  INV_X1 U22035 ( .A(n18974), .ZN(n18976) );
  AOI222_X1 U22036 ( .A1(n18978), .A2(n18983), .B1(n18981), .B2(n18977), .C1(
        n18976), .C2(n18975), .ZN(n18979) );
  AOI22_X1 U22037 ( .A1(n18988), .A2(n18980), .B1(n18979), .B2(n18985), .ZN(
        P3_U3289) );
  AOI222_X1 U22038 ( .A1(n18984), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18983), 
        .B2(n18982), .C1(n18987), .C2(n18981), .ZN(n18986) );
  AOI22_X1 U22039 ( .A1(n18988), .A2(n18987), .B1(n18986), .B2(n18985), .ZN(
        P3_U3290) );
  AOI21_X1 U22040 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18990) );
  AOI22_X1 U22041 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18990), .B2(n18989), .ZN(n18993) );
  AOI22_X1 U22042 ( .A1(n18996), .A2(n18993), .B1(n18992), .B2(n18991), .ZN(
        P3_U3292) );
  OAI21_X1 U22043 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18996), .ZN(n18994) );
  OAI21_X1 U22044 ( .B1(n18996), .B2(n18995), .A(n18994), .ZN(P3_U3293) );
  INV_X1 U22045 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18998) );
  AOI22_X1 U22046 ( .A1(n18936), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18998), 
        .B2(n18997), .ZN(P3_U3294) );
  MUX2_X1 U22047 ( .A(P3_MORE_REG_SCAN_IN), .B(n19000), .S(n18999), .Z(
        P3_U3295) );
  AOI21_X1 U22048 ( .B1(n19009), .B2(n19001), .A(n19023), .ZN(n19002) );
  OAI21_X1 U22049 ( .B1(n19004), .B2(n19003), .A(n19002), .ZN(n19005) );
  INV_X1 U22050 ( .A(n19005), .ZN(n19015) );
  AOI21_X1 U22051 ( .B1(n19008), .B2(n19007), .A(n19006), .ZN(n19010) );
  OAI211_X1 U22052 ( .C1(n19016), .C2(n19010), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19009), .ZN(n19012) );
  AOI21_X1 U22053 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19012), .A(n19011), 
        .ZN(n19014) );
  NAND2_X1 U22054 ( .A1(n19015), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19013) );
  OAI21_X1 U22055 ( .B1(n19015), .B2(n19014), .A(n19013), .ZN(P3_U3296) );
  MUX2_X1 U22056 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n18936), .Z(P3_U3297) );
  INV_X1 U22057 ( .A(n19016), .ZN(n19018) );
  OAI21_X1 U22058 ( .B1(n19020), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19019), 
        .ZN(n19017) );
  OAI21_X1 U22059 ( .B1(n19019), .B2(n19018), .A(n19017), .ZN(P3_U3298) );
  NOR2_X1 U22060 ( .A1(n19020), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19022)
         );
  OAI21_X1 U22061 ( .B1(n19023), .B2(n19022), .A(n19021), .ZN(P3_U3299) );
  INV_X1 U22062 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19025) );
  NAND2_X1 U22063 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19913), .ZN(n19905) );
  INV_X1 U22064 ( .A(n19905), .ZN(n19024) );
  NOR2_X1 U22065 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19902) );
  AOI21_X1 U22066 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19024), .A(n19902), 
        .ZN(n19895) );
  INV_X1 U22067 ( .A(n19895), .ZN(n19985) );
  OAI21_X1 U22068 ( .B1(n19029), .B2(n19025), .A(n19896), .ZN(P2_U2815) );
  INV_X1 U22069 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19027) );
  OAI22_X1 U22070 ( .A1(n20052), .A2(n19027), .B1(n20054), .B2(n19026), .ZN(
        P2_U2816) );
  NAND2_X1 U22071 ( .A1(n20068), .A2(n19028), .ZN(n19900) );
  AOI21_X1 U22072 ( .B1(n19029), .B2(n19900), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19030) );
  AOI21_X1 U22073 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n20071), .A(n19030), 
        .ZN(P2_U2817) );
  OAI21_X1 U22074 ( .B1(n19906), .B2(BS16), .A(n19985), .ZN(n19983) );
  OAI21_X1 U22075 ( .B1(n19985), .B2(n20001), .A(n19983), .ZN(P2_U2818) );
  NOR4_X1 U22076 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19034) );
  NOR4_X1 U22077 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19033) );
  NOR4_X1 U22078 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19032) );
  NOR4_X1 U22079 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19031) );
  NAND4_X1 U22080 ( .A1(n19034), .A2(n19033), .A3(n19032), .A4(n19031), .ZN(
        n19040) );
  NOR4_X1 U22081 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19038) );
  AOI211_X1 U22082 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19037) );
  NOR4_X1 U22083 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19036) );
  NOR4_X1 U22084 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19035) );
  NAND4_X1 U22085 ( .A1(n19038), .A2(n19037), .A3(n19036), .A4(n19035), .ZN(
        n19039) );
  NOR2_X1 U22086 ( .A1(n19040), .A2(n19039), .ZN(n19047) );
  INV_X1 U22087 ( .A(n19047), .ZN(n19046) );
  NOR2_X1 U22088 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19046), .ZN(n19041) );
  INV_X1 U22089 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19180) );
  INV_X1 U22090 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U22091 ( .A1(n19041), .A2(n19180), .B1(n19046), .B2(n19981), .ZN(
        P2_U2820) );
  OR3_X1 U22092 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19045) );
  INV_X1 U22093 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19979) );
  AOI22_X1 U22094 ( .A1(n19041), .A2(n19045), .B1(n19046), .B2(n19979), .ZN(
        P2_U2821) );
  INV_X1 U22095 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19984) );
  NAND2_X1 U22096 ( .A1(n19041), .A2(n19984), .ZN(n19044) );
  INV_X1 U22097 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19914) );
  OAI21_X1 U22098 ( .B1(n19180), .B2(n19914), .A(n19047), .ZN(n19042) );
  OAI21_X1 U22099 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19047), .A(n19042), 
        .ZN(n19043) );
  OAI221_X1 U22100 ( .B1(n19044), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19044), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19043), .ZN(P2_U2822) );
  INV_X1 U22101 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19977) );
  OAI221_X1 U22102 ( .B1(n19047), .B2(n19977), .C1(n19046), .C2(n19045), .A(
        n19044), .ZN(P2_U2823) );
  AOI21_X1 U22103 ( .B1(n19050), .B2(n19049), .A(n19048), .ZN(n19052) );
  AOI22_X1 U22104 ( .A1(n19052), .A2(n19190), .B1(n19102), .B2(n19051), .ZN(
        n19059) );
  OAI22_X1 U22105 ( .A1(n19134), .A2(n12593), .B1(n19053), .B2(n19100), .ZN(
        n19056) );
  INV_X1 U22106 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n19054) );
  OAI22_X1 U22107 ( .A1(n19054), .A2(n19163), .B1(n19950), .B2(n19181), .ZN(
        n19055) );
  AOI211_X1 U22108 ( .C1(n19188), .C2(n19057), .A(n19056), .B(n19055), .ZN(
        n19058) );
  OAI211_X1 U22109 ( .C1(n19060), .C2(n19179), .A(n19059), .B(n19058), .ZN(
        P2_U2835) );
  OAI21_X1 U22110 ( .B1(n19946), .B2(n19181), .A(n19150), .ZN(n19064) );
  OAI22_X1 U22111 ( .A1(n19062), .A2(n19186), .B1(n19061), .B2(n19134), .ZN(
        n19063) );
  AOI211_X1 U22112 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19193), .A(
        n19064), .B(n19063), .ZN(n19071) );
  NAND2_X1 U22113 ( .A1(n9807), .A2(n19065), .ZN(n19073) );
  XNOR2_X1 U22114 ( .A(n19066), .B(n19073), .ZN(n19069) );
  INV_X1 U22115 ( .A(n19067), .ZN(n19068) );
  AOI22_X1 U22116 ( .A1(n19069), .A2(n19190), .B1(n19068), .B2(n19188), .ZN(
        n19070) );
  OAI211_X1 U22117 ( .C1(n19072), .C2(n19179), .A(n19071), .B(n19070), .ZN(
        P2_U2837) );
  AOI211_X1 U22118 ( .C1(n19075), .C2(n19074), .A(n19891), .B(n19073), .ZN(
        n19079) );
  AOI22_X1 U22119 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19193), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19166), .ZN(n19076) );
  OAI211_X1 U22120 ( .C1(n19077), .C2(n19186), .A(n19076), .B(n19150), .ZN(
        n19078) );
  AOI211_X1 U22121 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19183), .A(n19079), .B(
        n19078), .ZN(n19083) );
  AOI22_X1 U22122 ( .A1(n19081), .A2(n19188), .B1(n19080), .B2(n19168), .ZN(
        n19082) );
  OAI211_X1 U22123 ( .C1(n19084), .C2(n19100), .A(n19083), .B(n19082), .ZN(
        P2_U2838) );
  AOI22_X1 U22124 ( .A1(n19085), .A2(n19102), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19183), .ZN(n19086) );
  OAI211_X1 U22125 ( .C1(n19942), .C2(n19181), .A(n19086), .B(n19150), .ZN(
        n19087) );
  AOI21_X1 U22126 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19193), .A(
        n19087), .ZN(n19093) );
  NAND2_X1 U22127 ( .A1(n15019), .A2(n19104), .ZN(n19088) );
  XOR2_X1 U22128 ( .A(n19089), .B(n19088), .Z(n19091) );
  AOI22_X1 U22129 ( .A1(n19091), .A2(n19190), .B1(n19090), .B2(n19188), .ZN(
        n19092) );
  OAI211_X1 U22130 ( .C1(n19094), .C2(n19179), .A(n19093), .B(n19092), .ZN(
        P2_U2839) );
  INV_X1 U22131 ( .A(n19095), .ZN(n19103) );
  AOI22_X1 U22132 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19193), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19166), .ZN(n19096) );
  OAI211_X1 U22133 ( .C1(n19134), .C2(n12337), .A(n19096), .B(n19150), .ZN(
        n19097) );
  AOI21_X1 U22134 ( .B1(n19098), .B2(n19188), .A(n19097), .ZN(n19099) );
  OAI21_X1 U22135 ( .B1(n19106), .B2(n19100), .A(n19099), .ZN(n19101) );
  AOI21_X1 U22136 ( .B1(n19103), .B2(n19102), .A(n19101), .ZN(n19109) );
  OAI211_X1 U22137 ( .C1(n19107), .C2(n19106), .A(n19105), .B(n19104), .ZN(
        n19108) );
  OAI211_X1 U22138 ( .C1(n19179), .C2(n19110), .A(n19109), .B(n19108), .ZN(
        P2_U2840) );
  AOI22_X1 U22139 ( .A1(n19183), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19193), .ZN(n19111) );
  OAI21_X1 U22140 ( .B1(n19112), .B2(n19186), .A(n19111), .ZN(n19113) );
  AOI211_X1 U22141 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19166), .A(n19287), 
        .B(n19113), .ZN(n19120) );
  NAND2_X1 U22142 ( .A1(n9807), .A2(n19114), .ZN(n19115) );
  XNOR2_X1 U22143 ( .A(n19116), .B(n19115), .ZN(n19118) );
  AOI22_X1 U22144 ( .A1(n19118), .A2(n19190), .B1(n19117), .B2(n19188), .ZN(
        n19119) );
  OAI211_X1 U22145 ( .C1(n19205), .C2(n19179), .A(n19120), .B(n19119), .ZN(
        P2_U2841) );
  INV_X1 U22146 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n19123) );
  OAI222_X1 U22147 ( .A1(n19163), .A2(n19123), .B1(n19122), .B2(n19134), .C1(
        n19121), .C2(n19186), .ZN(n19124) );
  AOI211_X1 U22148 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19166), .A(n19271), 
        .B(n19124), .ZN(n19131) );
  NAND2_X1 U22149 ( .A1(n9807), .A2(n19125), .ZN(n19126) );
  XNOR2_X1 U22150 ( .A(n19127), .B(n19126), .ZN(n19129) );
  AOI22_X1 U22151 ( .A1(n19129), .A2(n19190), .B1(n19128), .B2(n19188), .ZN(
        n19130) );
  OAI211_X1 U22152 ( .C1(n19132), .C2(n19179), .A(n19131), .B(n19130), .ZN(
        P2_U2843) );
  OAI22_X1 U22153 ( .A1(n19135), .A2(n19186), .B1(n19134), .B2(n19133), .ZN(
        n19136) );
  INV_X1 U22154 ( .A(n19136), .ZN(n19137) );
  OAI211_X1 U22155 ( .C1(n19927), .C2(n19181), .A(n19137), .B(n19150), .ZN(
        n19138) );
  AOI21_X1 U22156 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19193), .A(
        n19138), .ZN(n19145) );
  NAND2_X1 U22157 ( .A1(n9807), .A2(n19139), .ZN(n19140) );
  XNOR2_X1 U22158 ( .A(n19141), .B(n19140), .ZN(n19143) );
  AOI22_X1 U22159 ( .A1(n19143), .A2(n19190), .B1(n19142), .B2(n19188), .ZN(
        n19144) );
  OAI211_X1 U22160 ( .C1(n19146), .C2(n19179), .A(n19145), .B(n19144), .ZN(
        P2_U2847) );
  NAND2_X1 U22161 ( .A1(n9807), .A2(n19147), .ZN(n19148) );
  XOR2_X1 U22162 ( .A(n19149), .B(n19148), .Z(n19162) );
  OAI21_X1 U22163 ( .B1(n19924), .B2(n19181), .A(n19150), .ZN(n19154) );
  OAI22_X1 U22164 ( .A1(n19152), .A2(n19186), .B1(n19151), .B2(n19163), .ZN(
        n19153) );
  AOI211_X1 U22165 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19183), .A(n19154), .B(
        n19153), .ZN(n19161) );
  INV_X1 U22166 ( .A(n19155), .ZN(n19156) );
  OAI22_X1 U22167 ( .A1(n19158), .A2(n19179), .B1(n19157), .B2(n19156), .ZN(
        n19159) );
  INV_X1 U22168 ( .A(n19159), .ZN(n19160) );
  OAI211_X1 U22169 ( .C1(n19891), .C2(n19162), .A(n19161), .B(n19160), .ZN(
        P2_U2849) );
  OAI22_X1 U22170 ( .A1(n19164), .A2(n19186), .B1(n19286), .B2(n19163), .ZN(
        n19165) );
  AOI211_X1 U22171 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19166), .A(n19287), .B(
        n19165), .ZN(n19176) );
  AOI22_X1 U22172 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19183), .B1(n19168), .B2(
        n19167), .ZN(n19175) );
  AOI22_X1 U22173 ( .A1(n19169), .A2(n19189), .B1(n19188), .B2(n19281), .ZN(
        n19174) );
  AND2_X1 U22174 ( .A1(n15019), .A2(n19170), .ZN(n19172) );
  AOI21_X1 U22175 ( .B1(n19269), .B2(n19172), .A(n19891), .ZN(n19171) );
  OAI21_X1 U22176 ( .B1(n19269), .B2(n19172), .A(n19171), .ZN(n19173) );
  NAND4_X1 U22177 ( .A1(n19176), .A2(n19175), .A3(n19174), .A4(n19173), .ZN(
        P2_U2851) );
  INV_X1 U22178 ( .A(n19177), .ZN(n19185) );
  OAI22_X1 U22179 ( .A1(n19181), .A2(n19180), .B1(n19179), .B2(n19178), .ZN(
        n19182) );
  AOI21_X1 U22180 ( .B1(n19183), .B2(P2_EBX_REG_0__SCAN_IN), .A(n19182), .ZN(
        n19184) );
  OAI21_X1 U22181 ( .B1(n19186), .B2(n19185), .A(n19184), .ZN(n19187) );
  AOI21_X1 U22182 ( .B1(n12974), .B2(n19188), .A(n19187), .ZN(n19196) );
  AOI22_X1 U22183 ( .A1(n19191), .A2(n19190), .B1(n19586), .B2(n19189), .ZN(
        n19195) );
  OAI21_X1 U22184 ( .B1(n19193), .B2(n19192), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19194) );
  NAND3_X1 U22185 ( .A1(n19196), .A2(n19195), .A3(n19194), .ZN(P2_U2855) );
  AOI22_X1 U22186 ( .A1(n19199), .A2(n19198), .B1(n19197), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19202) );
  AOI22_X1 U22187 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19200), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19203), .ZN(n19201) );
  NAND2_X1 U22188 ( .A1(n19202), .A2(n19201), .ZN(P2_U2888) );
  AOI22_X1 U22189 ( .A1(n19213), .A2(n19260), .B1(n19203), .B2(
        P2_EAX_REG_14__SCAN_IN), .ZN(n19204) );
  OAI21_X1 U22190 ( .B1(n19206), .B2(n19205), .A(n19204), .ZN(P2_U2905) );
  INV_X1 U22191 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19231) );
  INV_X1 U22192 ( .A(n19206), .ZN(n19215) );
  AOI22_X1 U22193 ( .A1(n19215), .A2(n19207), .B1(n19213), .B2(n19258), .ZN(
        n19208) );
  OAI21_X1 U22194 ( .B1(n19217), .B2(n19231), .A(n19208), .ZN(P2_U2906) );
  AOI22_X1 U22195 ( .A1(n19215), .A2(n19210), .B1(n19213), .B2(n19209), .ZN(
        n19211) );
  OAI21_X1 U22196 ( .B1(n19217), .B2(n19235), .A(n19211), .ZN(P2_U2908) );
  AOI22_X1 U22197 ( .A1(n19215), .A2(n19214), .B1(n19213), .B2(n19212), .ZN(
        n19216) );
  OAI21_X1 U22198 ( .B1(n19217), .B2(n19239), .A(n19216), .ZN(P2_U2910) );
  NOR2_X1 U22199 ( .A1(n19225), .A2(n19218), .ZN(P2_U2920) );
  INV_X1 U22200 ( .A(n19219), .ZN(n19222) );
  AOI22_X1 U22201 ( .A1(n19222), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19227), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19220) );
  OAI21_X1 U22202 ( .B1(n19221), .B2(n19225), .A(n19220), .ZN(P2_U2921) );
  AOI22_X1 U22203 ( .A1(n19222), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n19227), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19223) );
  OAI21_X1 U22204 ( .B1(n19225), .B2(n19224), .A(n19223), .ZN(P2_U2922) );
  AOI22_X1 U22205 ( .A1(n19227), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19226) );
  OAI21_X1 U22206 ( .B1(n13357), .B2(n19256), .A(n19226), .ZN(P2_U2936) );
  INV_X1 U22207 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19229) );
  AOI22_X1 U22208 ( .A1(n19227), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19228) );
  OAI21_X1 U22209 ( .B1(n19229), .B2(n19256), .A(n19228), .ZN(P2_U2937) );
  AOI22_X1 U22210 ( .A1(n19227), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19230) );
  OAI21_X1 U22211 ( .B1(n19231), .B2(n19256), .A(n19230), .ZN(P2_U2938) );
  AOI22_X1 U22212 ( .A1(n19227), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19232) );
  OAI21_X1 U22213 ( .B1(n19233), .B2(n19256), .A(n19232), .ZN(P2_U2939) );
  AOI22_X1 U22214 ( .A1(n19227), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19234) );
  OAI21_X1 U22215 ( .B1(n19235), .B2(n19256), .A(n19234), .ZN(P2_U2940) );
  INV_X1 U22216 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19237) );
  AOI22_X1 U22217 ( .A1(n19227), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19236) );
  OAI21_X1 U22218 ( .B1(n19237), .B2(n19256), .A(n19236), .ZN(P2_U2941) );
  AOI22_X1 U22219 ( .A1(n19227), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19238) );
  OAI21_X1 U22220 ( .B1(n19239), .B2(n19256), .A(n19238), .ZN(P2_U2942) );
  AOI22_X1 U22221 ( .A1(n19227), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19240) );
  OAI21_X1 U22222 ( .B1(n19241), .B2(n19256), .A(n19240), .ZN(P2_U2943) );
  AOI22_X1 U22223 ( .A1(n19227), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19242) );
  OAI21_X1 U22224 ( .B1(n13556), .B2(n19256), .A(n19242), .ZN(P2_U2944) );
  AOI22_X1 U22225 ( .A1(n19227), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19243) );
  OAI21_X1 U22226 ( .B1(n13505), .B2(n19256), .A(n19243), .ZN(P2_U2945) );
  INV_X1 U22227 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19245) );
  AOI22_X1 U22228 ( .A1(n19227), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19244) );
  OAI21_X1 U22229 ( .B1(n19245), .B2(n19256), .A(n19244), .ZN(P2_U2946) );
  INV_X1 U22230 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19247) );
  AOI22_X1 U22231 ( .A1(n19227), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19246) );
  OAI21_X1 U22232 ( .B1(n19247), .B2(n19256), .A(n19246), .ZN(P2_U2947) );
  INV_X1 U22233 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19249) );
  AOI22_X1 U22234 ( .A1(n19227), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19248) );
  OAI21_X1 U22235 ( .B1(n19249), .B2(n19256), .A(n19248), .ZN(P2_U2948) );
  INV_X1 U22236 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19251) );
  AOI22_X1 U22237 ( .A1(n19227), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19250) );
  OAI21_X1 U22238 ( .B1(n19251), .B2(n19256), .A(n19250), .ZN(P2_U2949) );
  INV_X1 U22239 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19253) );
  AOI22_X1 U22240 ( .A1(n19227), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19252) );
  OAI21_X1 U22241 ( .B1(n19253), .B2(n19256), .A(n19252), .ZN(P2_U2950) );
  INV_X1 U22242 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19257) );
  AOI22_X1 U22243 ( .A1(n19227), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19254), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19255) );
  OAI21_X1 U22244 ( .B1(n19257), .B2(n19256), .A(n19255), .ZN(P2_U2951) );
  AOI22_X1 U22245 ( .A1(n19263), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19266), .ZN(n19259) );
  NAND2_X1 U22246 ( .A1(n19261), .A2(n19258), .ZN(n19264) );
  NAND2_X1 U22247 ( .A1(n19259), .A2(n19264), .ZN(P2_U2965) );
  AOI22_X1 U22248 ( .A1(n19263), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19266), .ZN(n19262) );
  NAND2_X1 U22249 ( .A1(n19261), .A2(n19260), .ZN(n19267) );
  NAND2_X1 U22250 ( .A1(n19262), .A2(n19267), .ZN(P2_U2966) );
  AOI22_X1 U22251 ( .A1(n19263), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19266), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n19265) );
  NAND2_X1 U22252 ( .A1(n19265), .A2(n19264), .ZN(P2_U2980) );
  AOI22_X1 U22253 ( .A1(n19263), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19266), .ZN(n19268) );
  NAND2_X1 U22254 ( .A1(n19268), .A2(n19267), .ZN(P2_U2981) );
  AOI22_X1 U22255 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19271), .B1(n19270), 
        .B2(n19269), .ZN(n19284) );
  XOR2_X1 U22256 ( .A(n9813), .B(n19272), .Z(n19297) );
  INV_X1 U22257 ( .A(n19297), .ZN(n19279) );
  XNOR2_X1 U22258 ( .A(n19274), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19275) );
  XNOR2_X1 U22259 ( .A(n19276), .B(n19275), .ZN(n19299) );
  OAI22_X1 U22260 ( .A1(n19279), .A2(n19278), .B1(n19277), .B2(n19299), .ZN(
        n19280) );
  AOI21_X1 U22261 ( .B1(n19282), .B2(n19281), .A(n19280), .ZN(n19283) );
  OAI211_X1 U22262 ( .C1(n19286), .C2(n19285), .A(n19284), .B(n19283), .ZN(
        P2_U3010) );
  NAND2_X1 U22263 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19287), .ZN(n19288) );
  OAI221_X1 U22264 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19291), .C1(
        n19290), .C2(n19289), .A(n19288), .ZN(n19295) );
  OAI22_X1 U22265 ( .A1(n19293), .A2(n19301), .B1(n19308), .B2(n19292), .ZN(
        n19294) );
  AOI211_X1 U22266 ( .C1(n19297), .C2(n19296), .A(n19295), .B(n19294), .ZN(
        n19298) );
  OAI21_X1 U22267 ( .B1(n19303), .B2(n19299), .A(n19298), .ZN(P2_U3042) );
  OAI22_X1 U22268 ( .A1(n19303), .A2(n19302), .B1(n19301), .B2(n19300), .ZN(
        n19310) );
  OAI211_X1 U22269 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n19305), .B(n19304), .ZN(n19306) );
  OAI21_X1 U22270 ( .B1(n19308), .B2(n19307), .A(n19306), .ZN(n19309) );
  AOI211_X1 U22271 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n19311), .A(
        n19310), .B(n19309), .ZN(n19313) );
  OAI211_X1 U22272 ( .C1(n19315), .C2(n19314), .A(n19313), .B(n19312), .ZN(
        P2_U3045) );
  AOI22_X1 U22273 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19357), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19356), .ZN(n19665) );
  OAI22_X2 U22274 ( .A1(n14567), .A2(n19366), .B1(n19319), .B2(n19364), .ZN(
        n19796) );
  NOR2_X2 U22275 ( .A1(n11815), .A2(n19368), .ZN(n19830) );
  NAND2_X1 U22276 ( .A1(n20012), .A2(n20019), .ZN(n19435) );
  OR2_X1 U22277 ( .A1(n19435), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19381) );
  NOR2_X1 U22278 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19381), .ZN(
        n19370) );
  AOI22_X1 U22279 ( .A1(n19796), .A2(n19881), .B1(n19830), .B2(n19370), .ZN(
        n19330) );
  OAI21_X1 U22280 ( .B1(n19881), .B2(n19401), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19320) );
  NAND2_X1 U22281 ( .A1(n19320), .A2(n20007), .ZN(n19328) );
  INV_X1 U22282 ( .A(n19834), .ZN(n19877) );
  NOR2_X1 U22283 ( .A1(n19328), .A2(n19877), .ZN(n19321) );
  AOI211_X1 U22284 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n12064), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19321), .ZN(n19322) );
  OAI21_X1 U22285 ( .B1(n19322), .B2(n19370), .A(n19836), .ZN(n19373) );
  NOR2_X1 U22286 ( .A1(n19877), .A2(n19370), .ZN(n19327) );
  INV_X1 U22287 ( .A(n12064), .ZN(n19325) );
  OAI21_X1 U22288 ( .B1(n19325), .B2(n19370), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19326) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19373), .B1(
        n19324), .B2(n19372), .ZN(n19329) );
  OAI211_X1 U22290 ( .C1(n19665), .C2(n19398), .A(n19330), .B(n19329), .ZN(
        P2_U3048) );
  AOI22_X1 U22291 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19357), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19356), .ZN(n19804) );
  NOR2_X2 U22292 ( .A1(n9802), .A2(n19368), .ZN(n19842) );
  AOI22_X1 U22293 ( .A1(n19800), .A2(n19881), .B1(n19842), .B2(n19370), .ZN(
        n19335) );
  AOI22_X1 U22294 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19373), .B1(
        n19333), .B2(n19372), .ZN(n19334) );
  OAI211_X1 U22295 ( .C1(n19804), .C2(n19398), .A(n19335), .B(n19334), .ZN(
        P2_U3049) );
  AOI22_X1 U22296 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19357), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19356), .ZN(n19763) );
  NOR2_X2 U22297 ( .A1(n9948), .A2(n19368), .ZN(n19847) );
  AOI22_X1 U22298 ( .A1(n19760), .A2(n19881), .B1(n19847), .B2(n19370), .ZN(
        n19339) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19373), .B1(
        n19337), .B2(n19372), .ZN(n19338) );
  OAI211_X1 U22300 ( .C1(n19763), .C2(n19398), .A(n19339), .B(n19338), .ZN(
        P2_U3050) );
  AOI22_X1 U22301 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19357), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19356), .ZN(n19767) );
  NOR2_X2 U22302 ( .A1(n19341), .A2(n19368), .ZN(n19852) );
  AOI22_X1 U22303 ( .A1(n19764), .A2(n19881), .B1(n19852), .B2(n19370), .ZN(
        n19344) );
  NOR2_X2 U22304 ( .A1(n19342), .A2(n19786), .ZN(n19853) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19373), .B1(
        n19853), .B2(n19372), .ZN(n19343) );
  OAI211_X1 U22306 ( .C1(n19767), .C2(n19398), .A(n19344), .B(n19343), .ZN(
        P2_U3051) );
  OAI22_X2 U22307 ( .A1(n19346), .A2(n19366), .B1(n19345), .B2(n19364), .ZN(
        n19860) );
  INV_X1 U22308 ( .A(n19860), .ZN(n19674) );
  AOI22_X1 U22309 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19356), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19357), .ZN(n19863) );
  INV_X1 U22310 ( .A(n19863), .ZN(n19768) );
  NOR2_X2 U22311 ( .A1(n19347), .A2(n19368), .ZN(n19858) );
  AOI22_X1 U22312 ( .A1(n19768), .A2(n19881), .B1(n19858), .B2(n19370), .ZN(
        n19350) );
  NOR2_X2 U22313 ( .A1(n19348), .A2(n19786), .ZN(n19859) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19373), .B1(
        n19859), .B2(n19372), .ZN(n19349) );
  OAI211_X1 U22315 ( .C1(n19674), .C2(n19398), .A(n19350), .B(n19349), .ZN(
        P2_U3052) );
  NOR2_X2 U22316 ( .A1(n12785), .A2(n19368), .ZN(n19864) );
  AOI22_X1 U22317 ( .A1(n19811), .A2(n19881), .B1(n19864), .B2(n19370), .ZN(
        n19355) );
  NOR2_X2 U22318 ( .A1(n19353), .A2(n19786), .ZN(n19865) );
  AOI22_X1 U22319 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19373), .B1(
        n19865), .B2(n19372), .ZN(n19354) );
  OAI211_X1 U22320 ( .C1(n19814), .C2(n19398), .A(n19355), .B(n19354), .ZN(
        P2_U3053) );
  AOI22_X1 U22321 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19357), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19356), .ZN(n19679) );
  NOR2_X2 U22322 ( .A1(n12957), .A2(n19368), .ZN(n19870) );
  AOI22_X1 U22323 ( .A1(n19774), .A2(n19881), .B1(n19870), .B2(n19370), .ZN(
        n19361) );
  NOR2_X2 U22324 ( .A1(n19359), .A2(n19786), .ZN(n19871) );
  AOI22_X1 U22325 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19373), .B1(
        n19871), .B2(n19372), .ZN(n19360) );
  OAI211_X1 U22326 ( .C1(n19679), .C2(n19398), .A(n19361), .B(n19360), .ZN(
        P2_U3054) );
  OAI22_X2 U22327 ( .A1(n19367), .A2(n19366), .B1(n19365), .B2(n19364), .ZN(
        n19821) );
  NOR2_X2 U22328 ( .A1(n19369), .A2(n19368), .ZN(n19876) );
  AOI22_X1 U22329 ( .A1(n19821), .A2(n19881), .B1(n19876), .B2(n19370), .ZN(
        n19375) );
  NOR2_X2 U22330 ( .A1(n19371), .A2(n19786), .ZN(n19878) );
  AOI22_X1 U22331 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19373), .B1(
        n19878), .B2(n19372), .ZN(n19374) );
  OAI211_X1 U22332 ( .C1(n19826), .C2(n19398), .A(n19375), .B(n19374), .ZN(
        P2_U3055) );
  NOR2_X2 U22333 ( .A1(n19624), .A2(n19559), .ZN(n19431) );
  INV_X1 U22334 ( .A(n19431), .ZN(n19405) );
  INV_X1 U22335 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19533) );
  INV_X1 U22336 ( .A(n19887), .ZN(n19377) );
  INV_X1 U22337 ( .A(n12044), .ZN(n19376) );
  NOR2_X1 U22338 ( .A1(n19620), .A2(n19435), .ZN(n19399) );
  NOR3_X1 U22339 ( .A1(n19376), .A2(n19399), .A3(n19533), .ZN(n19380) );
  AOI211_X2 U22340 ( .C1(n19381), .C2(n19533), .A(n19377), .B(n19380), .ZN(
        n19400) );
  AOI22_X1 U22341 ( .A1(n19400), .A2(n19324), .B1(n19830), .B2(n19399), .ZN(
        n19385) );
  NAND2_X1 U22342 ( .A1(n19987), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19563) );
  INV_X1 U22343 ( .A(n19563), .ZN(n19379) );
  INV_X1 U22344 ( .A(n19624), .ZN(n19378) );
  NAND2_X1 U22345 ( .A1(n19379), .A2(n19378), .ZN(n19382) );
  AOI21_X1 U22346 ( .B1(n19382), .B2(n19381), .A(n19380), .ZN(n19383) );
  OAI211_X1 U22347 ( .C1(n19399), .C2(n12958), .A(n19383), .B(n19836), .ZN(
        n19402) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19796), .ZN(n19384) );
  OAI211_X1 U22349 ( .C1(n19665), .C2(n19405), .A(n19385), .B(n19384), .ZN(
        P2_U3056) );
  AOI22_X1 U22350 ( .A1(n19400), .A2(n19333), .B1(n19842), .B2(n19399), .ZN(
        n19387) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19800), .ZN(n19386) );
  OAI211_X1 U22352 ( .C1(n19804), .C2(n19405), .A(n19387), .B(n19386), .ZN(
        P2_U3057) );
  INV_X1 U22353 ( .A(n19760), .ZN(n19851) );
  AOI22_X1 U22354 ( .A1(n19400), .A2(n19337), .B1(n19847), .B2(n19399), .ZN(
        n19389) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19402), .B1(
        n19431), .B2(n19848), .ZN(n19388) );
  OAI211_X1 U22356 ( .C1(n19851), .C2(n19398), .A(n19389), .B(n19388), .ZN(
        P2_U3058) );
  INV_X1 U22357 ( .A(n19764), .ZN(n19857) );
  AOI22_X1 U22358 ( .A1(n19400), .A2(n19853), .B1(n19852), .B2(n19399), .ZN(
        n19391) );
  INV_X1 U22359 ( .A(n19767), .ZN(n19854) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19402), .B1(
        n19431), .B2(n19854), .ZN(n19390) );
  OAI211_X1 U22361 ( .C1(n19857), .C2(n19398), .A(n19391), .B(n19390), .ZN(
        P2_U3059) );
  AOI22_X1 U22362 ( .A1(n19400), .A2(n19859), .B1(n19858), .B2(n19399), .ZN(
        n19393) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19402), .B1(
        n19431), .B2(n19860), .ZN(n19392) );
  OAI211_X1 U22364 ( .C1(n19863), .C2(n19398), .A(n19393), .B(n19392), .ZN(
        P2_U3060) );
  INV_X1 U22365 ( .A(n19811), .ZN(n19869) );
  AOI22_X1 U22366 ( .A1(n19400), .A2(n19865), .B1(n19864), .B2(n19399), .ZN(
        n19395) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19402), .B1(
        n19431), .B2(n19866), .ZN(n19394) );
  OAI211_X1 U22368 ( .C1(n19869), .C2(n19398), .A(n19395), .B(n19394), .ZN(
        P2_U3061) );
  AOI22_X1 U22369 ( .A1(n19400), .A2(n19871), .B1(n19870), .B2(n19399), .ZN(
        n19397) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19402), .B1(
        n19431), .B2(n19872), .ZN(n19396) );
  OAI211_X1 U22371 ( .C1(n19875), .C2(n19398), .A(n19397), .B(n19396), .ZN(
        P2_U3062) );
  AOI22_X1 U22372 ( .A1(n19400), .A2(n19878), .B1(n19876), .B2(n19399), .ZN(
        n19404) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19821), .ZN(n19403) );
  OAI211_X1 U22374 ( .C1(n19826), .C2(n19405), .A(n19404), .B(n19403), .ZN(
        P2_U3063) );
  INV_X1 U22375 ( .A(n12061), .ZN(n19406) );
  NOR2_X1 U22376 ( .A1(n19653), .A2(n19435), .ZN(n19429) );
  OAI21_X1 U22377 ( .B1(n19406), .B2(n19429), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19408) );
  INV_X1 U22378 ( .A(n19435), .ZN(n19407) );
  NAND2_X1 U22379 ( .A1(n19652), .A2(n19407), .ZN(n19409) );
  NAND2_X1 U22380 ( .A1(n19408), .A2(n19409), .ZN(n19430) );
  AOI22_X1 U22381 ( .A1(n19430), .A2(n19324), .B1(n19830), .B2(n19429), .ZN(
        n19416) );
  INV_X1 U22382 ( .A(n19462), .ZN(n19452) );
  OAI21_X1 U22383 ( .B1(n19452), .B2(n19431), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19410) );
  NAND2_X1 U22384 ( .A1(n19410), .A2(n19409), .ZN(n19413) );
  INV_X1 U22385 ( .A(n19429), .ZN(n19411) );
  OAI21_X1 U22386 ( .B1(n12061), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19411), 
        .ZN(n19412) );
  MUX2_X1 U22387 ( .A(n19413), .B(n19412), .S(n20002), .Z(n19414) );
  NAND2_X1 U22388 ( .A1(n19414), .A2(n19836), .ZN(n19432) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19796), .ZN(n19415) );
  OAI211_X1 U22390 ( .C1(n19665), .C2(n19462), .A(n19416), .B(n19415), .ZN(
        P2_U3064) );
  AOI22_X1 U22391 ( .A1(n19430), .A2(n19333), .B1(n19842), .B2(n19429), .ZN(
        n19418) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19800), .ZN(n19417) );
  OAI211_X1 U22393 ( .C1(n19804), .C2(n19462), .A(n19418), .B(n19417), .ZN(
        P2_U3065) );
  AOI22_X1 U22394 ( .A1(n19430), .A2(n19337), .B1(n19847), .B2(n19429), .ZN(
        n19420) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19760), .ZN(n19419) );
  OAI211_X1 U22396 ( .C1(n19763), .C2(n19462), .A(n19420), .B(n19419), .ZN(
        P2_U3066) );
  AOI22_X1 U22397 ( .A1(n19430), .A2(n19853), .B1(n19852), .B2(n19429), .ZN(
        n19422) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19764), .ZN(n19421) );
  OAI211_X1 U22399 ( .C1(n19767), .C2(n19462), .A(n19422), .B(n19421), .ZN(
        P2_U3067) );
  AOI22_X1 U22400 ( .A1(n19430), .A2(n19859), .B1(n19858), .B2(n19429), .ZN(
        n19424) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19768), .ZN(n19423) );
  OAI211_X1 U22402 ( .C1(n19674), .C2(n19462), .A(n19424), .B(n19423), .ZN(
        P2_U3068) );
  AOI22_X1 U22403 ( .A1(n19430), .A2(n19865), .B1(n19864), .B2(n19429), .ZN(
        n19426) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19811), .ZN(n19425) );
  OAI211_X1 U22405 ( .C1(n19814), .C2(n19462), .A(n19426), .B(n19425), .ZN(
        P2_U3069) );
  AOI22_X1 U22406 ( .A1(n19430), .A2(n19871), .B1(n19870), .B2(n19429), .ZN(
        n19428) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19774), .ZN(n19427) );
  OAI211_X1 U22408 ( .C1(n19679), .C2(n19462), .A(n19428), .B(n19427), .ZN(
        P2_U3070) );
  AOI22_X1 U22409 ( .A1(n19430), .A2(n19878), .B1(n19876), .B2(n19429), .ZN(
        n19434) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19821), .ZN(n19433) );
  OAI211_X1 U22411 ( .C1(n19826), .C2(n19462), .A(n19434), .B(n19433), .ZN(
        P2_U3071) );
  INV_X1 U22412 ( .A(n19796), .ZN(n19841) );
  NOR2_X1 U22413 ( .A1(n19686), .A2(n19435), .ZN(n19457) );
  AOI22_X1 U22414 ( .A1(n19494), .A2(n19838), .B1(n19457), .B2(n19830), .ZN(
        n19443) );
  OAI21_X1 U22415 ( .B1(n19563), .B2(n19698), .A(n20007), .ZN(n19441) );
  NOR2_X1 U22416 ( .A1(n20028), .A2(n19435), .ZN(n19438) );
  INV_X1 U22417 ( .A(n19457), .ZN(n19436) );
  OAI211_X1 U22418 ( .C1(n12065), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20002), 
        .B(n19436), .ZN(n19437) );
  OAI211_X1 U22419 ( .C1(n19441), .C2(n19438), .A(n19836), .B(n19437), .ZN(
        n19459) );
  INV_X1 U22420 ( .A(n19438), .ZN(n19440) );
  OAI21_X1 U22421 ( .B1(n11988), .B2(n19457), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19439) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19459), .B1(
        n19324), .B2(n19458), .ZN(n19442) );
  OAI211_X1 U22423 ( .C1(n19841), .C2(n19462), .A(n19443), .B(n19442), .ZN(
        P2_U3072) );
  INV_X1 U22424 ( .A(n19804), .ZN(n19843) );
  AOI22_X1 U22425 ( .A1(n19494), .A2(n19843), .B1(n19457), .B2(n19842), .ZN(
        n19445) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19459), .B1(
        n19333), .B2(n19458), .ZN(n19444) );
  OAI211_X1 U22427 ( .C1(n19846), .C2(n19462), .A(n19445), .B(n19444), .ZN(
        P2_U3073) );
  AOI22_X1 U22428 ( .A1(n19494), .A2(n19848), .B1(n19457), .B2(n19847), .ZN(
        n19447) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19459), .B1(
        n19337), .B2(n19458), .ZN(n19446) );
  OAI211_X1 U22430 ( .C1(n19851), .C2(n19462), .A(n19447), .B(n19446), .ZN(
        P2_U3074) );
  AOI22_X1 U22431 ( .A1(n19764), .A2(n19452), .B1(n19457), .B2(n19852), .ZN(
        n19449) );
  AOI22_X1 U22432 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19459), .B1(
        n19853), .B2(n19458), .ZN(n19448) );
  OAI211_X1 U22433 ( .C1(n19767), .C2(n19491), .A(n19449), .B(n19448), .ZN(
        P2_U3075) );
  AOI22_X1 U22434 ( .A1(n19860), .A2(n19494), .B1(n19457), .B2(n19858), .ZN(
        n19451) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19459), .B1(
        n19859), .B2(n19458), .ZN(n19450) );
  OAI211_X1 U22436 ( .C1(n19863), .C2(n19462), .A(n19451), .B(n19450), .ZN(
        P2_U3076) );
  AOI22_X1 U22437 ( .A1(n19811), .A2(n19452), .B1(n19457), .B2(n19864), .ZN(
        n19454) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19459), .B1(
        n19865), .B2(n19458), .ZN(n19453) );
  OAI211_X1 U22439 ( .C1(n19814), .C2(n19491), .A(n19454), .B(n19453), .ZN(
        P2_U3077) );
  AOI22_X1 U22440 ( .A1(n19494), .A2(n19872), .B1(n19457), .B2(n19870), .ZN(
        n19456) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19459), .B1(
        n19871), .B2(n19458), .ZN(n19455) );
  OAI211_X1 U22442 ( .C1(n19875), .C2(n19462), .A(n19456), .B(n19455), .ZN(
        P2_U3078) );
  INV_X1 U22443 ( .A(n19821), .ZN(n19886) );
  AOI22_X1 U22444 ( .A1(n19880), .A2(n19494), .B1(n19457), .B2(n19876), .ZN(
        n19461) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19459), .B1(
        n19878), .B2(n19458), .ZN(n19460) );
  OAI211_X1 U22446 ( .C1(n19886), .C2(n19462), .A(n19461), .B(n19460), .ZN(
        P2_U3079) );
  NAND3_X1 U22447 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20012), .A3(
        n20028), .ZN(n19504) );
  NOR2_X1 U22448 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19504), .ZN(
        n19492) );
  NOR2_X1 U22449 ( .A1(n20007), .A2(n19492), .ZN(n19463) );
  OAI21_X1 U22450 ( .B1(n19471), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19463), 
        .ZN(n19470) );
  NOR2_X1 U22451 ( .A1(n19465), .A2(n19464), .ZN(n19719) );
  NAND2_X1 U22452 ( .A1(n19719), .A2(n20012), .ZN(n19474) );
  OAI21_X1 U22453 ( .B1(n19494), .B2(n19521), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19467) );
  NAND2_X1 U22454 ( .A1(n19474), .A2(n19467), .ZN(n19468) );
  AND2_X1 U22455 ( .A1(n19836), .A2(n19468), .ZN(n19469) );
  INV_X1 U22456 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19477) );
  INV_X1 U22457 ( .A(n19471), .ZN(n19472) );
  OAI21_X1 U22458 ( .B1(n19472), .B2(n19492), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19473) );
  OAI21_X1 U22459 ( .B1(n19474), .B2(n20002), .A(n19473), .ZN(n19493) );
  AOI22_X1 U22460 ( .A1(n19493), .A2(n19324), .B1(n19830), .B2(n19492), .ZN(
        n19476) );
  AOI22_X1 U22461 ( .A1(n19494), .A2(n19796), .B1(n19521), .B2(n19838), .ZN(
        n19475) );
  OAI211_X1 U22462 ( .C1(n19478), .C2(n19477), .A(n19476), .B(n19475), .ZN(
        P2_U3080) );
  AOI22_X1 U22463 ( .A1(n19493), .A2(n19333), .B1(n19842), .B2(n19492), .ZN(
        n19480) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19495), .B1(
        n19521), .B2(n19843), .ZN(n19479) );
  OAI211_X1 U22465 ( .C1(n19846), .C2(n19491), .A(n19480), .B(n19479), .ZN(
        P2_U3081) );
  AOI22_X1 U22466 ( .A1(n19493), .A2(n19337), .B1(n19847), .B2(n19492), .ZN(
        n19482) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19495), .B1(
        n19521), .B2(n19848), .ZN(n19481) );
  OAI211_X1 U22468 ( .C1(n19851), .C2(n19491), .A(n19482), .B(n19481), .ZN(
        P2_U3082) );
  AOI22_X1 U22469 ( .A1(n19493), .A2(n19853), .B1(n19852), .B2(n19492), .ZN(
        n19484) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19495), .B1(
        n19521), .B2(n19854), .ZN(n19483) );
  OAI211_X1 U22471 ( .C1(n19857), .C2(n19491), .A(n19484), .B(n19483), .ZN(
        P2_U3083) );
  AOI22_X1 U22472 ( .A1(n19493), .A2(n19859), .B1(n19858), .B2(n19492), .ZN(
        n19486) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19495), .B1(
        n19521), .B2(n19860), .ZN(n19485) );
  OAI211_X1 U22474 ( .C1(n19863), .C2(n19491), .A(n19486), .B(n19485), .ZN(
        P2_U3084) );
  AOI22_X1 U22475 ( .A1(n19493), .A2(n19865), .B1(n19864), .B2(n19492), .ZN(
        n19488) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19495), .B1(
        n19494), .B2(n19811), .ZN(n19487) );
  OAI211_X1 U22477 ( .C1(n19814), .C2(n19518), .A(n19488), .B(n19487), .ZN(
        P2_U3085) );
  AOI22_X1 U22478 ( .A1(n19493), .A2(n19871), .B1(n19870), .B2(n19492), .ZN(
        n19490) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19495), .B1(
        n19521), .B2(n19872), .ZN(n19489) );
  OAI211_X1 U22480 ( .C1(n19875), .C2(n19491), .A(n19490), .B(n19489), .ZN(
        P2_U3086) );
  AOI22_X1 U22481 ( .A1(n19493), .A2(n19878), .B1(n19876), .B2(n19492), .ZN(
        n19497) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19495), .B1(
        n19494), .B2(n19821), .ZN(n19496) );
  OAI211_X1 U22483 ( .C1(n19826), .C2(n19518), .A(n19497), .B(n19496), .ZN(
        P2_U3087) );
  NOR2_X1 U22484 ( .A1(n20036), .A2(n19504), .ZN(n19532) );
  AOI22_X1 U22485 ( .A1(n19555), .A2(n19838), .B1(n19830), .B2(n19532), .ZN(
        n19507) );
  OAI21_X1 U22486 ( .B1(n19563), .B2(n19754), .A(n20007), .ZN(n19505) );
  INV_X1 U22487 ( .A(n19504), .ZN(n19501) );
  INV_X1 U22488 ( .A(n12054), .ZN(n19502) );
  OAI21_X1 U22489 ( .B1(n19502), .B2(n19533), .A(n12958), .ZN(n19499) );
  INV_X1 U22490 ( .A(n19532), .ZN(n19498) );
  AOI21_X1 U22491 ( .B1(n19499), .B2(n19498), .A(n19786), .ZN(n19500) );
  OAI21_X1 U22492 ( .B1(n19502), .B2(n19532), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19503) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19523), .B1(
        n19324), .B2(n19522), .ZN(n19506) );
  OAI211_X1 U22494 ( .C1(n19841), .C2(n19518), .A(n19507), .B(n19506), .ZN(
        P2_U3088) );
  AOI22_X1 U22495 ( .A1(n19555), .A2(n19843), .B1(n19842), .B2(n19532), .ZN(
        n19509) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19523), .B1(
        n19333), .B2(n19522), .ZN(n19508) );
  OAI211_X1 U22497 ( .C1(n19846), .C2(n19518), .A(n19509), .B(n19508), .ZN(
        P2_U3089) );
  AOI22_X1 U22498 ( .A1(n19555), .A2(n19848), .B1(n19847), .B2(n19532), .ZN(
        n19511) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19523), .B1(
        n19337), .B2(n19522), .ZN(n19510) );
  OAI211_X1 U22500 ( .C1(n19851), .C2(n19518), .A(n19511), .B(n19510), .ZN(
        P2_U3090) );
  AOI22_X1 U22501 ( .A1(n19764), .A2(n19521), .B1(n19852), .B2(n19532), .ZN(
        n19513) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19523), .B1(
        n19853), .B2(n19522), .ZN(n19512) );
  OAI211_X1 U22503 ( .C1(n19767), .C2(n19552), .A(n19513), .B(n19512), .ZN(
        P2_U3091) );
  AOI22_X1 U22504 ( .A1(n19768), .A2(n19521), .B1(n19858), .B2(n19532), .ZN(
        n19515) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19523), .B1(
        n19859), .B2(n19522), .ZN(n19514) );
  OAI211_X1 U22506 ( .C1(n19674), .C2(n19552), .A(n19515), .B(n19514), .ZN(
        P2_U3092) );
  AOI22_X1 U22507 ( .A1(n19866), .A2(n19555), .B1(n19864), .B2(n19532), .ZN(
        n19517) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19523), .B1(
        n19865), .B2(n19522), .ZN(n19516) );
  OAI211_X1 U22509 ( .C1(n19869), .C2(n19518), .A(n19517), .B(n19516), .ZN(
        P2_U3093) );
  AOI22_X1 U22510 ( .A1(n19774), .A2(n19521), .B1(n19870), .B2(n19532), .ZN(
        n19520) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19523), .B1(
        n19871), .B2(n19522), .ZN(n19519) );
  OAI211_X1 U22512 ( .C1(n19679), .C2(n19552), .A(n19520), .B(n19519), .ZN(
        P2_U3094) );
  AOI22_X1 U22513 ( .A1(n19821), .A2(n19521), .B1(n19876), .B2(n19532), .ZN(
        n19525) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19523), .B1(
        n19878), .B2(n19522), .ZN(n19524) );
  OAI211_X1 U22515 ( .C1(n19826), .C2(n19552), .A(n19525), .B(n19524), .ZN(
        P2_U3095) );
  AOI21_X1 U22516 ( .B1(n19552), .B2(n19580), .A(n20001), .ZN(n19527) );
  NOR2_X1 U22517 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19831), .ZN(
        n19565) );
  INV_X1 U22518 ( .A(n19565), .ZN(n19562) );
  NOR2_X1 U22519 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19562), .ZN(
        n19553) );
  AOI221_X1 U22520 ( .B1(n19532), .B2(n12958), .C1(n19527), .C2(n12958), .A(
        n19553), .ZN(n19531) );
  INV_X1 U22521 ( .A(n19553), .ZN(n19528) );
  AND2_X1 U22522 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19528), .ZN(n19529) );
  NAND2_X1 U22523 ( .A1(n12059), .A2(n19529), .ZN(n19536) );
  NAND2_X1 U22524 ( .A1(n19536), .A2(n19836), .ZN(n19530) );
  INV_X1 U22525 ( .A(n19556), .ZN(n19539) );
  NOR2_X1 U22526 ( .A1(n19532), .A2(n19553), .ZN(n19534) );
  OAI21_X1 U22527 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19534), .A(n19533), 
        .ZN(n19535) );
  AND2_X1 U22528 ( .A1(n19536), .A2(n19535), .ZN(n19554) );
  AOI22_X1 U22529 ( .A1(n19554), .A2(n19324), .B1(n19830), .B2(n19553), .ZN(
        n19538) );
  AOI22_X1 U22530 ( .A1(n19555), .A2(n19796), .B1(n19582), .B2(n19838), .ZN(
        n19537) );
  OAI211_X1 U22531 ( .C1(n19539), .C2(n13078), .A(n19538), .B(n19537), .ZN(
        P2_U3096) );
  AOI22_X1 U22532 ( .A1(n19554), .A2(n19333), .B1(n19842), .B2(n19553), .ZN(
        n19541) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19556), .B1(
        n19555), .B2(n19800), .ZN(n19540) );
  OAI211_X1 U22534 ( .C1(n19804), .C2(n19580), .A(n19541), .B(n19540), .ZN(
        P2_U3097) );
  AOI22_X1 U22535 ( .A1(n19554), .A2(n19337), .B1(n19847), .B2(n19553), .ZN(
        n19543) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19556), .B1(
        n19582), .B2(n19848), .ZN(n19542) );
  OAI211_X1 U22537 ( .C1(n19851), .C2(n19552), .A(n19543), .B(n19542), .ZN(
        P2_U3098) );
  AOI22_X1 U22538 ( .A1(n19554), .A2(n19853), .B1(n19852), .B2(n19553), .ZN(
        n19545) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19556), .B1(
        n19555), .B2(n19764), .ZN(n19544) );
  OAI211_X1 U22540 ( .C1(n19767), .C2(n19580), .A(n19545), .B(n19544), .ZN(
        P2_U3099) );
  AOI22_X1 U22541 ( .A1(n19554), .A2(n19859), .B1(n19858), .B2(n19553), .ZN(
        n19547) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19556), .B1(
        n19582), .B2(n19860), .ZN(n19546) );
  OAI211_X1 U22543 ( .C1(n19863), .C2(n19552), .A(n19547), .B(n19546), .ZN(
        P2_U3100) );
  AOI22_X1 U22544 ( .A1(n19554), .A2(n19865), .B1(n19864), .B2(n19553), .ZN(
        n19549) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19556), .B1(
        n19555), .B2(n19811), .ZN(n19548) );
  OAI211_X1 U22546 ( .C1(n19814), .C2(n19580), .A(n19549), .B(n19548), .ZN(
        P2_U3101) );
  AOI22_X1 U22547 ( .A1(n19554), .A2(n19871), .B1(n19870), .B2(n19553), .ZN(
        n19551) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19556), .B1(
        n19582), .B2(n19872), .ZN(n19550) );
  OAI211_X1 U22549 ( .C1(n19875), .C2(n19552), .A(n19551), .B(n19550), .ZN(
        P2_U3102) );
  AOI22_X1 U22550 ( .A1(n19554), .A2(n19878), .B1(n19876), .B2(n19553), .ZN(
        n19558) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19556), .B1(
        n19555), .B2(n19821), .ZN(n19557) );
  OAI211_X1 U22552 ( .C1(n19826), .C2(n19580), .A(n19558), .B(n19557), .ZN(
        P2_U3103) );
  INV_X1 U22553 ( .A(n12058), .ZN(n19560) );
  NOR2_X1 U22554 ( .A1(n20036), .A2(n19562), .ZN(n19593) );
  OAI21_X1 U22555 ( .B1(n19560), .B2(n19593), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19561) );
  OAI21_X1 U22556 ( .B1(n19562), .B2(n20002), .A(n19561), .ZN(n19581) );
  AOI22_X1 U22557 ( .A1(n19581), .A2(n19324), .B1(n19830), .B2(n19593), .ZN(
        n19567) );
  NOR2_X1 U22558 ( .A1(n19563), .A2(n19832), .ZN(n20006) );
  INV_X1 U22559 ( .A(n19593), .ZN(n19590) );
  OAI211_X1 U22560 ( .C1(n12058), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20002), 
        .B(n19590), .ZN(n19564) );
  OAI211_X1 U22561 ( .C1(n20006), .C2(n19565), .A(n19836), .B(n19564), .ZN(
        n19583) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19583), .B1(
        n19582), .B2(n19796), .ZN(n19566) );
  OAI211_X1 U22563 ( .C1(n19665), .C2(n19617), .A(n19567), .B(n19566), .ZN(
        P2_U3104) );
  AOI22_X1 U22564 ( .A1(n19581), .A2(n19333), .B1(n19842), .B2(n19593), .ZN(
        n19569) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19583), .B1(
        n19609), .B2(n19843), .ZN(n19568) );
  OAI211_X1 U22566 ( .C1(n19846), .C2(n19580), .A(n19569), .B(n19568), .ZN(
        P2_U3105) );
  AOI22_X1 U22567 ( .A1(n19581), .A2(n19337), .B1(n19847), .B2(n19593), .ZN(
        n19571) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19583), .B1(
        n19609), .B2(n19848), .ZN(n19570) );
  OAI211_X1 U22569 ( .C1(n19851), .C2(n19580), .A(n19571), .B(n19570), .ZN(
        P2_U3106) );
  AOI22_X1 U22570 ( .A1(n19581), .A2(n19853), .B1(n19852), .B2(n19593), .ZN(
        n19573) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19583), .B1(
        n19582), .B2(n19764), .ZN(n19572) );
  OAI211_X1 U22572 ( .C1(n19767), .C2(n19617), .A(n19573), .B(n19572), .ZN(
        P2_U3107) );
  AOI22_X1 U22573 ( .A1(n19581), .A2(n19859), .B1(n19858), .B2(n19593), .ZN(
        n19575) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19583), .B1(
        n19609), .B2(n19860), .ZN(n19574) );
  OAI211_X1 U22575 ( .C1(n19863), .C2(n19580), .A(n19575), .B(n19574), .ZN(
        P2_U3108) );
  AOI22_X1 U22576 ( .A1(n19581), .A2(n19865), .B1(n19864), .B2(n19593), .ZN(
        n19577) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19583), .B1(
        n19609), .B2(n19866), .ZN(n19576) );
  OAI211_X1 U22578 ( .C1(n19869), .C2(n19580), .A(n19577), .B(n19576), .ZN(
        P2_U3109) );
  AOI22_X1 U22579 ( .A1(n19581), .A2(n19871), .B1(n19870), .B2(n19593), .ZN(
        n19579) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19583), .B1(
        n19609), .B2(n19872), .ZN(n19578) );
  OAI211_X1 U22581 ( .C1(n19875), .C2(n19580), .A(n19579), .B(n19578), .ZN(
        P2_U3110) );
  AOI22_X1 U22582 ( .A1(n19581), .A2(n19878), .B1(n19876), .B2(n19593), .ZN(
        n19585) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19583), .B1(
        n19582), .B2(n19821), .ZN(n19584) );
  OAI211_X1 U22584 ( .C1(n19826), .C2(n19617), .A(n19585), .B(n19584), .ZN(
        P2_U3111) );
  NAND2_X1 U22585 ( .A1(n20019), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19689) );
  OR2_X1 U22586 ( .A1(n19689), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19627) );
  NOR2_X1 U22587 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19627), .ZN(
        n19612) );
  AOI22_X1 U22588 ( .A1(n19796), .A2(n19609), .B1(n19830), .B2(n19612), .ZN(
        n19598) );
  NAND2_X1 U22589 ( .A1(n19645), .A2(n19617), .ZN(n19587) );
  AOI21_X1 U22590 ( .B1(n19587), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20002), 
        .ZN(n19592) );
  INV_X1 U22591 ( .A(n19588), .ZN(n19594) );
  OAI21_X1 U22592 ( .B1(n19594), .B2(n19533), .A(n12958), .ZN(n19589) );
  AOI21_X1 U22593 ( .B1(n19592), .B2(n19590), .A(n19589), .ZN(n19591) );
  OAI21_X1 U22594 ( .B1(n19612), .B2(n19591), .A(n19836), .ZN(n19614) );
  OAI21_X1 U22595 ( .B1(n19612), .B2(n19593), .A(n19592), .ZN(n19596) );
  OAI21_X1 U22596 ( .B1(n19594), .B2(n19612), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19595) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19614), .B1(
        n19324), .B2(n19613), .ZN(n19597) );
  OAI211_X1 U22598 ( .C1(n19665), .C2(n19645), .A(n19598), .B(n19597), .ZN(
        P2_U3112) );
  AOI22_X1 U22599 ( .A1(n19800), .A2(n19609), .B1(n19612), .B2(n19842), .ZN(
        n19600) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19614), .B1(
        n19613), .B2(n19333), .ZN(n19599) );
  OAI211_X1 U22601 ( .C1(n19804), .C2(n19645), .A(n19600), .B(n19599), .ZN(
        P2_U3113) );
  AOI22_X1 U22602 ( .A1(n19760), .A2(n19609), .B1(n19847), .B2(n19612), .ZN(
        n19602) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19614), .B1(
        n19613), .B2(n19337), .ZN(n19601) );
  OAI211_X1 U22604 ( .C1(n19763), .C2(n19645), .A(n19602), .B(n19601), .ZN(
        P2_U3114) );
  AOI22_X1 U22605 ( .A1(n19764), .A2(n19609), .B1(n19852), .B2(n19612), .ZN(
        n19604) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19614), .B1(
        n19613), .B2(n19853), .ZN(n19603) );
  OAI211_X1 U22607 ( .C1(n19767), .C2(n19645), .A(n19604), .B(n19603), .ZN(
        P2_U3115) );
  INV_X1 U22608 ( .A(n19645), .ZN(n19647) );
  AOI22_X1 U22609 ( .A1(n19860), .A2(n19647), .B1(n19858), .B2(n19612), .ZN(
        n19606) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19614), .B1(
        n19613), .B2(n19859), .ZN(n19605) );
  OAI211_X1 U22611 ( .C1(n19863), .C2(n19617), .A(n19606), .B(n19605), .ZN(
        P2_U3116) );
  AOI22_X1 U22612 ( .A1(n19811), .A2(n19609), .B1(n19612), .B2(n19864), .ZN(
        n19608) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19614), .B1(
        n19613), .B2(n19865), .ZN(n19607) );
  OAI211_X1 U22614 ( .C1(n19814), .C2(n19645), .A(n19608), .B(n19607), .ZN(
        P2_U3117) );
  AOI22_X1 U22615 ( .A1(n19774), .A2(n19609), .B1(n19870), .B2(n19612), .ZN(
        n19611) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19614), .B1(
        n19613), .B2(n19871), .ZN(n19610) );
  OAI211_X1 U22617 ( .C1(n19679), .C2(n19645), .A(n19611), .B(n19610), .ZN(
        P2_U3118) );
  AOI22_X1 U22618 ( .A1(n19880), .A2(n19647), .B1(n19612), .B2(n19876), .ZN(
        n19616) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19614), .B1(
        n19613), .B2(n19878), .ZN(n19615) );
  OAI211_X1 U22620 ( .C1(n19886), .C2(n19617), .A(n19616), .B(n19615), .ZN(
        P2_U3119) );
  OR2_X1 U22621 ( .A1(n19987), .A2(n20001), .ZN(n19833) );
  OAI21_X1 U22622 ( .B1(n19833), .B2(n19624), .A(n20007), .ZN(n19628) );
  INV_X1 U22623 ( .A(n19627), .ZN(n19618) );
  OR2_X1 U22624 ( .A1(n19628), .A2(n19618), .ZN(n19623) );
  NAND2_X1 U22625 ( .A1(n12046), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19619) );
  NAND2_X1 U22626 ( .A1(n19619), .A2(n12958), .ZN(n19621) );
  NOR2_X1 U22627 ( .A1(n19620), .A2(n19689), .ZN(n19646) );
  INV_X1 U22628 ( .A(n19646), .ZN(n19659) );
  AOI21_X1 U22629 ( .B1(n19621), .B2(n19659), .A(n19786), .ZN(n19622) );
  AOI22_X1 U22630 ( .A1(n19682), .A2(n19838), .B1(n19830), .B2(n19646), .ZN(
        n19630) );
  INV_X1 U22631 ( .A(n12046), .ZN(n19625) );
  OAI21_X1 U22632 ( .B1(n19625), .B2(n19646), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19626) );
  AOI22_X1 U22633 ( .A1(n19324), .A2(n19648), .B1(n19647), .B2(n19796), .ZN(
        n19629) );
  OAI211_X1 U22634 ( .C1(n19632), .C2(n19631), .A(n19630), .B(n19629), .ZN(
        P2_U3120) );
  AOI22_X1 U22635 ( .A1(n19682), .A2(n19843), .B1(n19646), .B2(n19842), .ZN(
        n19634) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19649), .B1(
        n19333), .B2(n19648), .ZN(n19633) );
  OAI211_X1 U22637 ( .C1(n19846), .C2(n19645), .A(n19634), .B(n19633), .ZN(
        P2_U3121) );
  AOI22_X1 U22638 ( .A1(n19760), .A2(n19647), .B1(n19847), .B2(n19646), .ZN(
        n19636) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19649), .B1(
        n19337), .B2(n19648), .ZN(n19635) );
  OAI211_X1 U22640 ( .C1(n19763), .C2(n19660), .A(n19636), .B(n19635), .ZN(
        P2_U3122) );
  AOI22_X1 U22641 ( .A1(n19854), .A2(n19682), .B1(n19852), .B2(n19646), .ZN(
        n19638) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19649), .B1(
        n19853), .B2(n19648), .ZN(n19637) );
  OAI211_X1 U22643 ( .C1(n19857), .C2(n19645), .A(n19638), .B(n19637), .ZN(
        P2_U3123) );
  AOI22_X1 U22644 ( .A1(n19768), .A2(n19647), .B1(n19858), .B2(n19646), .ZN(
        n19640) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19649), .B1(
        n19859), .B2(n19648), .ZN(n19639) );
  OAI211_X1 U22646 ( .C1(n19674), .C2(n19660), .A(n19640), .B(n19639), .ZN(
        P2_U3124) );
  AOI22_X1 U22647 ( .A1(n19866), .A2(n19682), .B1(n19646), .B2(n19864), .ZN(
        n19642) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19649), .B1(
        n19865), .B2(n19648), .ZN(n19641) );
  OAI211_X1 U22649 ( .C1(n19869), .C2(n19645), .A(n19642), .B(n19641), .ZN(
        P2_U3125) );
  AOI22_X1 U22650 ( .A1(n19682), .A2(n19872), .B1(n19870), .B2(n19646), .ZN(
        n19644) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19649), .B1(
        n19871), .B2(n19648), .ZN(n19643) );
  OAI211_X1 U22652 ( .C1(n19875), .C2(n19645), .A(n19644), .B(n19643), .ZN(
        P2_U3126) );
  AOI22_X1 U22653 ( .A1(n19821), .A2(n19647), .B1(n19876), .B2(n19646), .ZN(
        n19651) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19649), .B1(
        n19878), .B2(n19648), .ZN(n19650) );
  OAI211_X1 U22655 ( .C1(n19826), .C2(n19660), .A(n19651), .B(n19650), .ZN(
        P2_U3127) );
  INV_X1 U22656 ( .A(n19652), .ZN(n19655) );
  INV_X1 U22657 ( .A(n12045), .ZN(n19656) );
  NOR2_X1 U22658 ( .A1(n19653), .A2(n19689), .ZN(n19680) );
  OAI21_X1 U22659 ( .B1(n19656), .B2(n19680), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19654) );
  OAI21_X1 U22660 ( .B1(n19689), .B2(n19655), .A(n19654), .ZN(n19681) );
  AOI22_X1 U22661 ( .A1(n19681), .A2(n19324), .B1(n19830), .B2(n19680), .ZN(
        n19664) );
  NAND3_X1 U22662 ( .A1(n19656), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n12958), 
        .ZN(n19658) );
  INV_X1 U22663 ( .A(n19680), .ZN(n19657) );
  NAND2_X1 U22664 ( .A1(n19658), .A2(n19657), .ZN(n19662) );
  OAI221_X1 U22665 ( .B1(n20001), .B2(n19718), .C1(n20001), .C2(n19660), .A(
        n19659), .ZN(n19661) );
  OAI221_X1 U22666 ( .B1(n19662), .B2(n20007), .C1(n19662), .C2(n19661), .A(
        n19836), .ZN(n19683) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19796), .ZN(n19663) );
  OAI211_X1 U22668 ( .C1(n19665), .C2(n19718), .A(n19664), .B(n19663), .ZN(
        P2_U3128) );
  AOI22_X1 U22669 ( .A1(n19681), .A2(n19333), .B1(n19842), .B2(n19680), .ZN(
        n19667) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19800), .ZN(n19666) );
  OAI211_X1 U22671 ( .C1(n19804), .C2(n19718), .A(n19667), .B(n19666), .ZN(
        P2_U3129) );
  AOI22_X1 U22672 ( .A1(n19681), .A2(n19337), .B1(n19847), .B2(n19680), .ZN(
        n19669) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19760), .ZN(n19668) );
  OAI211_X1 U22674 ( .C1(n19763), .C2(n19718), .A(n19669), .B(n19668), .ZN(
        P2_U3130) );
  AOI22_X1 U22675 ( .A1(n19681), .A2(n19853), .B1(n19852), .B2(n19680), .ZN(
        n19671) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19764), .ZN(n19670) );
  OAI211_X1 U22677 ( .C1(n19767), .C2(n19718), .A(n19671), .B(n19670), .ZN(
        P2_U3131) );
  AOI22_X1 U22678 ( .A1(n19681), .A2(n19859), .B1(n19858), .B2(n19680), .ZN(
        n19673) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19768), .ZN(n19672) );
  OAI211_X1 U22680 ( .C1(n19674), .C2(n19718), .A(n19673), .B(n19672), .ZN(
        P2_U3132) );
  AOI22_X1 U22681 ( .A1(n19681), .A2(n19865), .B1(n19864), .B2(n19680), .ZN(
        n19676) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19811), .ZN(n19675) );
  OAI211_X1 U22683 ( .C1(n19814), .C2(n19718), .A(n19676), .B(n19675), .ZN(
        P2_U3133) );
  AOI22_X1 U22684 ( .A1(n19681), .A2(n19871), .B1(n19870), .B2(n19680), .ZN(
        n19678) );
  AOI22_X1 U22685 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19774), .ZN(n19677) );
  OAI211_X1 U22686 ( .C1(n19679), .C2(n19718), .A(n19678), .B(n19677), .ZN(
        P2_U3134) );
  AOI22_X1 U22687 ( .A1(n19681), .A2(n19878), .B1(n19876), .B2(n19680), .ZN(
        n19685) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19821), .ZN(n19684) );
  OAI211_X1 U22689 ( .C1(n19826), .C2(n19718), .A(n19685), .B(n19684), .ZN(
        P2_U3135) );
  INV_X1 U22690 ( .A(n19686), .ZN(n19688) );
  INV_X1 U22691 ( .A(n19689), .ZN(n19687) );
  NAND2_X1 U22692 ( .A1(n19688), .A2(n19687), .ZN(n19694) );
  NAND3_X1 U22693 ( .A1(n12051), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19694), 
        .ZN(n19692) );
  NOR2_X1 U22694 ( .A1(n20028), .A2(n19689), .ZN(n19697) );
  INV_X1 U22695 ( .A(n19697), .ZN(n19690) );
  OAI21_X1 U22696 ( .B1(n19690), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19533), 
        .ZN(n19691) );
  INV_X1 U22697 ( .A(n19694), .ZN(n19713) );
  AOI22_X1 U22698 ( .A1(n19714), .A2(n19324), .B1(n19830), .B2(n19713), .ZN(
        n19700) );
  INV_X1 U22699 ( .A(n19833), .ZN(n19696) );
  INV_X1 U22700 ( .A(n19692), .ZN(n19693) );
  AOI211_X1 U22701 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19694), .A(n19786), 
        .B(n19693), .ZN(n19695) );
  OAI221_X1 U22702 ( .B1(n19697), .B2(n20003), .C1(n19697), .C2(n19696), .A(
        n19695), .ZN(n19715) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19715), .B1(
        n19722), .B2(n19838), .ZN(n19699) );
  OAI211_X1 U22704 ( .C1(n19841), .C2(n19718), .A(n19700), .B(n19699), .ZN(
        P2_U3136) );
  AOI22_X1 U22705 ( .A1(n19714), .A2(n19333), .B1(n19842), .B2(n19713), .ZN(
        n19702) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19715), .B1(
        n19722), .B2(n19843), .ZN(n19701) );
  OAI211_X1 U22707 ( .C1(n19846), .C2(n19718), .A(n19702), .B(n19701), .ZN(
        P2_U3137) );
  AOI22_X1 U22708 ( .A1(n19714), .A2(n19337), .B1(n19847), .B2(n19713), .ZN(
        n19704) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19715), .B1(
        n19722), .B2(n19848), .ZN(n19703) );
  OAI211_X1 U22710 ( .C1(n19851), .C2(n19718), .A(n19704), .B(n19703), .ZN(
        P2_U3138) );
  AOI22_X1 U22711 ( .A1(n19714), .A2(n19853), .B1(n19852), .B2(n19713), .ZN(
        n19706) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19715), .B1(
        n19722), .B2(n19854), .ZN(n19705) );
  OAI211_X1 U22713 ( .C1(n19857), .C2(n19718), .A(n19706), .B(n19705), .ZN(
        P2_U3139) );
  AOI22_X1 U22714 ( .A1(n19714), .A2(n19859), .B1(n19858), .B2(n19713), .ZN(
        n19708) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19715), .B1(
        n19722), .B2(n19860), .ZN(n19707) );
  OAI211_X1 U22716 ( .C1(n19863), .C2(n19718), .A(n19708), .B(n19707), .ZN(
        P2_U3140) );
  AOI22_X1 U22717 ( .A1(n19714), .A2(n19865), .B1(n19864), .B2(n19713), .ZN(
        n19710) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19715), .B1(
        n19722), .B2(n19866), .ZN(n19709) );
  OAI211_X1 U22719 ( .C1(n19869), .C2(n19718), .A(n19710), .B(n19709), .ZN(
        P2_U3141) );
  AOI22_X1 U22720 ( .A1(n19714), .A2(n19871), .B1(n19870), .B2(n19713), .ZN(
        n19712) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19715), .B1(
        n19722), .B2(n19872), .ZN(n19711) );
  OAI211_X1 U22722 ( .C1(n19875), .C2(n19718), .A(n19712), .B(n19711), .ZN(
        P2_U3142) );
  AOI22_X1 U22723 ( .A1(n19714), .A2(n19878), .B1(n19876), .B2(n19713), .ZN(
        n19717) );
  AOI22_X1 U22724 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19715), .B1(
        n19722), .B2(n19880), .ZN(n19716) );
  OAI211_X1 U22725 ( .C1(n19886), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P2_U3143) );
  NAND2_X1 U22726 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19719), .ZN(
        n19724) );
  OR2_X1 U22727 ( .A1(n19724), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19721) );
  INV_X1 U22728 ( .A(n12050), .ZN(n19720) );
  NAND3_X1 U22729 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20028), .ZN(n19753) );
  NOR2_X1 U22730 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19753), .ZN(
        n19741) );
  NOR3_X1 U22731 ( .A1(n19720), .A2(n19741), .A3(n19533), .ZN(n19723) );
  AOI21_X1 U22732 ( .B1(n19533), .B2(n19721), .A(n19723), .ZN(n19742) );
  AOI22_X1 U22733 ( .A1(n19742), .A2(n19324), .B1(n19830), .B2(n19741), .ZN(
        n19728) );
  NOR2_X2 U22734 ( .A1(n19783), .A2(n19754), .ZN(n19778) );
  OAI21_X1 U22735 ( .B1(n19722), .B2(n19778), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19725) );
  AOI211_X1 U22736 ( .C1(n19725), .C2(n19724), .A(n19786), .B(n19723), .ZN(
        n19726) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19743), .B1(
        n19778), .B2(n19838), .ZN(n19727) );
  OAI211_X1 U22738 ( .C1(n19841), .C2(n19746), .A(n19728), .B(n19727), .ZN(
        P2_U3144) );
  AOI22_X1 U22739 ( .A1(n19742), .A2(n19333), .B1(n19842), .B2(n19741), .ZN(
        n19730) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19743), .B1(
        n19778), .B2(n19843), .ZN(n19729) );
  OAI211_X1 U22741 ( .C1(n19846), .C2(n19746), .A(n19730), .B(n19729), .ZN(
        P2_U3145) );
  AOI22_X1 U22742 ( .A1(n19742), .A2(n19337), .B1(n19847), .B2(n19741), .ZN(
        n19732) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19743), .B1(
        n19778), .B2(n19848), .ZN(n19731) );
  OAI211_X1 U22744 ( .C1(n19851), .C2(n19746), .A(n19732), .B(n19731), .ZN(
        P2_U3146) );
  AOI22_X1 U22745 ( .A1(n19742), .A2(n19853), .B1(n19852), .B2(n19741), .ZN(
        n19734) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19743), .B1(
        n19778), .B2(n19854), .ZN(n19733) );
  OAI211_X1 U22747 ( .C1(n19857), .C2(n19746), .A(n19734), .B(n19733), .ZN(
        P2_U3147) );
  AOI22_X1 U22748 ( .A1(n19742), .A2(n19859), .B1(n19858), .B2(n19741), .ZN(
        n19736) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19743), .B1(
        n19778), .B2(n19860), .ZN(n19735) );
  OAI211_X1 U22750 ( .C1(n19863), .C2(n19746), .A(n19736), .B(n19735), .ZN(
        P2_U3148) );
  AOI22_X1 U22751 ( .A1(n19742), .A2(n19865), .B1(n19864), .B2(n19741), .ZN(
        n19738) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19743), .B1(
        n19778), .B2(n19866), .ZN(n19737) );
  OAI211_X1 U22753 ( .C1(n19869), .C2(n19746), .A(n19738), .B(n19737), .ZN(
        P2_U3149) );
  AOI22_X1 U22754 ( .A1(n19742), .A2(n19871), .B1(n19870), .B2(n19741), .ZN(
        n19740) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19743), .B1(
        n19778), .B2(n19872), .ZN(n19739) );
  OAI211_X1 U22756 ( .C1(n19875), .C2(n19746), .A(n19740), .B(n19739), .ZN(
        P2_U3150) );
  AOI22_X1 U22757 ( .A1(n19742), .A2(n19878), .B1(n19876), .B2(n19741), .ZN(
        n19745) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19743), .B1(
        n19778), .B2(n19880), .ZN(n19744) );
  OAI211_X1 U22759 ( .C1(n19886), .C2(n19746), .A(n19745), .B(n19744), .ZN(
        P2_U3151) );
  OAI21_X1 U22760 ( .B1(n19833), .B2(n19754), .A(n19753), .ZN(n19750) );
  OR2_X1 U22761 ( .A1(n12055), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19748) );
  NOR2_X1 U22762 ( .A1(n20036), .A2(n19753), .ZN(n19785) );
  NOR2_X1 U22763 ( .A1(n20007), .A2(n19785), .ZN(n19747) );
  AOI21_X1 U22764 ( .B1(n19748), .B2(n19747), .A(n19786), .ZN(n19749) );
  INV_X1 U22765 ( .A(n12055), .ZN(n19751) );
  OAI21_X1 U22766 ( .B1(n19751), .B2(n19785), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19752) );
  OAI21_X1 U22767 ( .B1(n19753), .B2(n20002), .A(n19752), .ZN(n19777) );
  AOI22_X1 U22768 ( .A1(n19777), .A2(n19324), .B1(n19830), .B2(n19785), .ZN(
        n19757) );
  AOI22_X1 U22769 ( .A1(n19778), .A2(n19796), .B1(n19820), .B2(n19838), .ZN(
        n19756) );
  OAI211_X1 U22770 ( .C1(n19782), .C2(n13088), .A(n19757), .B(n19756), .ZN(
        P2_U3152) );
  AOI22_X1 U22771 ( .A1(n19777), .A2(n19333), .B1(n19842), .B2(n19785), .ZN(
        n19759) );
  INV_X1 U22772 ( .A(n19782), .ZN(n19771) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19771), .B1(
        n19778), .B2(n19800), .ZN(n19758) );
  OAI211_X1 U22774 ( .C1(n19804), .C2(n19818), .A(n19759), .B(n19758), .ZN(
        P2_U3153) );
  AOI22_X1 U22775 ( .A1(n19777), .A2(n19337), .B1(n19847), .B2(n19785), .ZN(
        n19762) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19771), .B1(
        n19778), .B2(n19760), .ZN(n19761) );
  OAI211_X1 U22777 ( .C1(n19763), .C2(n19818), .A(n19762), .B(n19761), .ZN(
        P2_U3154) );
  AOI22_X1 U22778 ( .A1(n19777), .A2(n19853), .B1(n19852), .B2(n19785), .ZN(
        n19766) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19771), .B1(
        n19778), .B2(n19764), .ZN(n19765) );
  OAI211_X1 U22780 ( .C1(n19767), .C2(n19818), .A(n19766), .B(n19765), .ZN(
        P2_U3155) );
  AOI22_X1 U22781 ( .A1(n19777), .A2(n19859), .B1(n19858), .B2(n19785), .ZN(
        n19770) );
  AOI22_X1 U22782 ( .A1(n19820), .A2(n19860), .B1(n19778), .B2(n19768), .ZN(
        n19769) );
  OAI211_X1 U22783 ( .C1(n19782), .C2(n13205), .A(n19770), .B(n19769), .ZN(
        P2_U3156) );
  AOI22_X1 U22784 ( .A1(n19777), .A2(n19865), .B1(n19864), .B2(n19785), .ZN(
        n19773) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19771), .B1(
        n19778), .B2(n19811), .ZN(n19772) );
  OAI211_X1 U22786 ( .C1(n19814), .C2(n19818), .A(n19773), .B(n19772), .ZN(
        P2_U3157) );
  AOI22_X1 U22787 ( .A1(n19777), .A2(n19871), .B1(n19870), .B2(n19785), .ZN(
        n19776) );
  AOI22_X1 U22788 ( .A1(n19778), .A2(n19774), .B1(n19820), .B2(n19872), .ZN(
        n19775) );
  OAI211_X1 U22789 ( .C1(n19782), .C2(n12101), .A(n19776), .B(n19775), .ZN(
        P2_U3158) );
  INV_X1 U22790 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n19781) );
  AOI22_X1 U22791 ( .A1(n19777), .A2(n19878), .B1(n19876), .B2(n19785), .ZN(
        n19780) );
  AOI22_X1 U22792 ( .A1(n19820), .A2(n19880), .B1(n19778), .B2(n19821), .ZN(
        n19779) );
  OAI211_X1 U22793 ( .C1(n19782), .C2(n19781), .A(n19780), .B(n19779), .ZN(
        P2_U3159) );
  NAND2_X1 U22794 ( .A1(n19818), .A2(n19885), .ZN(n19784) );
  AOI21_X1 U22795 ( .B1(n19784), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20002), 
        .ZN(n19791) );
  NOR3_X2 U22796 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20012), .A3(
        n19831), .ZN(n19819) );
  NOR2_X1 U22797 ( .A1(n19819), .A2(n19785), .ZN(n19794) );
  NAND2_X1 U22798 ( .A1(n19791), .A2(n19794), .ZN(n19790) );
  OR2_X1 U22799 ( .A1(n12047), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19788) );
  NOR2_X1 U22800 ( .A1(n20007), .A2(n19819), .ZN(n19787) );
  AOI21_X1 U22801 ( .B1(n19788), .B2(n19787), .A(n19786), .ZN(n19789) );
  INV_X1 U22802 ( .A(n19885), .ZN(n19815) );
  AOI22_X1 U22803 ( .A1(n19815), .A2(n19838), .B1(n19830), .B2(n19819), .ZN(
        n19798) );
  INV_X1 U22804 ( .A(n19791), .ZN(n19795) );
  INV_X1 U22805 ( .A(n12047), .ZN(n19792) );
  OAI21_X1 U22806 ( .B1(n19792), .B2(n19819), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19793) );
  AOI22_X1 U22807 ( .A1(n19324), .A2(n19822), .B1(n19820), .B2(n19796), .ZN(
        n19797) );
  OAI211_X1 U22808 ( .C1(n19801), .C2(n19799), .A(n19798), .B(n19797), .ZN(
        P2_U3160) );
  AOI22_X1 U22809 ( .A1(n19800), .A2(n19820), .B1(n19819), .B2(n19842), .ZN(
        n19803) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19823), .B1(
        n19333), .B2(n19822), .ZN(n19802) );
  OAI211_X1 U22811 ( .C1(n19804), .C2(n19885), .A(n19803), .B(n19802), .ZN(
        P2_U3161) );
  AOI22_X1 U22812 ( .A1(n19815), .A2(n19848), .B1(n19819), .B2(n19847), .ZN(
        n19806) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19823), .B1(
        n19337), .B2(n19822), .ZN(n19805) );
  OAI211_X1 U22814 ( .C1(n19851), .C2(n19818), .A(n19806), .B(n19805), .ZN(
        P2_U3162) );
  AOI22_X1 U22815 ( .A1(n19854), .A2(n19815), .B1(n19819), .B2(n19852), .ZN(
        n19808) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19823), .B1(
        n19853), .B2(n19822), .ZN(n19807) );
  OAI211_X1 U22817 ( .C1(n19857), .C2(n19818), .A(n19808), .B(n19807), .ZN(
        P2_U3163) );
  AOI22_X1 U22818 ( .A1(n19860), .A2(n19815), .B1(n19819), .B2(n19858), .ZN(
        n19810) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19823), .B1(
        n19859), .B2(n19822), .ZN(n19809) );
  OAI211_X1 U22820 ( .C1(n19863), .C2(n19818), .A(n19810), .B(n19809), .ZN(
        P2_U3164) );
  AOI22_X1 U22821 ( .A1(n19811), .A2(n19820), .B1(n19819), .B2(n19864), .ZN(
        n19813) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19823), .B1(
        n19865), .B2(n19822), .ZN(n19812) );
  OAI211_X1 U22823 ( .C1(n19814), .C2(n19885), .A(n19813), .B(n19812), .ZN(
        P2_U3165) );
  AOI22_X1 U22824 ( .A1(n19815), .A2(n19872), .B1(n19819), .B2(n19870), .ZN(
        n19817) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19823), .B1(
        n19871), .B2(n19822), .ZN(n19816) );
  OAI211_X1 U22826 ( .C1(n19875), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        P2_U3166) );
  AOI22_X1 U22827 ( .A1(n19821), .A2(n19820), .B1(n19819), .B2(n19876), .ZN(
        n19825) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19823), .B1(
        n19878), .B2(n19822), .ZN(n19824) );
  OAI211_X1 U22829 ( .C1(n19826), .C2(n19885), .A(n19825), .B(n19824), .ZN(
        P2_U3167) );
  OR2_X1 U22830 ( .A1(n20012), .A2(n19831), .ZN(n19829) );
  INV_X1 U22831 ( .A(n12067), .ZN(n19827) );
  OAI21_X1 U22832 ( .B1(n19827), .B2(n19877), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19828) );
  OAI21_X1 U22833 ( .B1(n19829), .B2(n20002), .A(n19828), .ZN(n19879) );
  AOI22_X1 U22834 ( .A1(n19879), .A2(n19324), .B1(n19877), .B2(n19830), .ZN(
        n19840) );
  OAI22_X1 U22835 ( .A1(n19833), .A2(n19832), .B1(n19831), .B2(n20012), .ZN(
        n19837) );
  OAI211_X1 U22836 ( .C1(n12067), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20002), 
        .B(n19834), .ZN(n19835) );
  NAND3_X1 U22837 ( .A1(n19837), .A2(n19836), .A3(n19835), .ZN(n19882) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19882), .B1(
        n19881), .B2(n19838), .ZN(n19839) );
  OAI211_X1 U22839 ( .C1(n19841), .C2(n19885), .A(n19840), .B(n19839), .ZN(
        P2_U3168) );
  AOI22_X1 U22840 ( .A1(n19879), .A2(n19333), .B1(n19877), .B2(n19842), .ZN(
        n19845) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19882), .B1(
        n19881), .B2(n19843), .ZN(n19844) );
  OAI211_X1 U22842 ( .C1(n19846), .C2(n19885), .A(n19845), .B(n19844), .ZN(
        P2_U3169) );
  AOI22_X1 U22843 ( .A1(n19879), .A2(n19337), .B1(n19877), .B2(n19847), .ZN(
        n19850) );
  AOI22_X1 U22844 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19882), .B1(
        n19881), .B2(n19848), .ZN(n19849) );
  OAI211_X1 U22845 ( .C1(n19851), .C2(n19885), .A(n19850), .B(n19849), .ZN(
        P2_U3170) );
  AOI22_X1 U22846 ( .A1(n19879), .A2(n19853), .B1(n19877), .B2(n19852), .ZN(
        n19856) );
  AOI22_X1 U22847 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19882), .B1(
        n19881), .B2(n19854), .ZN(n19855) );
  OAI211_X1 U22848 ( .C1(n19857), .C2(n19885), .A(n19856), .B(n19855), .ZN(
        P2_U3171) );
  AOI22_X1 U22849 ( .A1(n19879), .A2(n19859), .B1(n19877), .B2(n19858), .ZN(
        n19862) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19882), .B1(
        n19881), .B2(n19860), .ZN(n19861) );
  OAI211_X1 U22851 ( .C1(n19863), .C2(n19885), .A(n19862), .B(n19861), .ZN(
        P2_U3172) );
  AOI22_X1 U22852 ( .A1(n19879), .A2(n19865), .B1(n19877), .B2(n19864), .ZN(
        n19868) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19882), .B1(
        n19881), .B2(n19866), .ZN(n19867) );
  OAI211_X1 U22854 ( .C1(n19869), .C2(n19885), .A(n19868), .B(n19867), .ZN(
        P2_U3173) );
  AOI22_X1 U22855 ( .A1(n19879), .A2(n19871), .B1(n19877), .B2(n19870), .ZN(
        n19874) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19882), .B1(
        n19881), .B2(n19872), .ZN(n19873) );
  OAI211_X1 U22857 ( .C1(n19875), .C2(n19885), .A(n19874), .B(n19873), .ZN(
        P2_U3174) );
  AOI22_X1 U22858 ( .A1(n19879), .A2(n19878), .B1(n19877), .B2(n19876), .ZN(
        n19884) );
  AOI22_X1 U22859 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19882), .B1(
        n19881), .B2(n19880), .ZN(n19883) );
  OAI211_X1 U22860 ( .C1(n19886), .C2(n19885), .A(n19884), .B(n19883), .ZN(
        P2_U3175) );
  OAI211_X1 U22861 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20057), .A(n19888), 
        .B(n19887), .ZN(n19893) );
  NOR2_X1 U22862 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20054), .ZN(n19889) );
  OAI211_X1 U22863 ( .C1(n19890), .C2(n19889), .A(n19897), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19892) );
  OAI211_X1 U22864 ( .C1(n19894), .C2(n19893), .A(n19892), .B(n19891), .ZN(
        P2_U3177) );
  AND2_X1 U22865 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19896), .ZN(
        P2_U3179) );
  AND2_X1 U22866 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19896), .ZN(
        P2_U3180) );
  AND2_X1 U22867 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19896), .ZN(
        P2_U3181) );
  AND2_X1 U22868 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19896), .ZN(
        P2_U3182) );
  AND2_X1 U22869 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19896), .ZN(
        P2_U3183) );
  AND2_X1 U22870 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19896), .ZN(
        P2_U3184) );
  AND2_X1 U22871 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19896), .ZN(
        P2_U3185) );
  AND2_X1 U22872 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19896), .ZN(
        P2_U3186) );
  AND2_X1 U22873 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19896), .ZN(
        P2_U3187) );
  AND2_X1 U22874 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19896), .ZN(
        P2_U3188) );
  AND2_X1 U22875 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19896), .ZN(
        P2_U3189) );
  AND2_X1 U22876 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19896), .ZN(
        P2_U3190) );
  AND2_X1 U22877 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19896), .ZN(
        P2_U3191) );
  AND2_X1 U22878 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19896), .ZN(
        P2_U3192) );
  AND2_X1 U22879 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19896), .ZN(
        P2_U3193) );
  AND2_X1 U22880 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19895), .ZN(
        P2_U3194) );
  AND2_X1 U22881 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19895), .ZN(
        P2_U3195) );
  AND2_X1 U22882 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19895), .ZN(
        P2_U3196) );
  AND2_X1 U22883 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19895), .ZN(
        P2_U3197) );
  AND2_X1 U22884 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19895), .ZN(
        P2_U3198) );
  AND2_X1 U22885 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19895), .ZN(
        P2_U3199) );
  AND2_X1 U22886 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19895), .ZN(
        P2_U3200) );
  AND2_X1 U22887 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19895), .ZN(P2_U3201) );
  AND2_X1 U22888 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19895), .ZN(P2_U3202) );
  AND2_X1 U22889 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19895), .ZN(P2_U3203) );
  AND2_X1 U22890 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19895), .ZN(P2_U3204) );
  AND2_X1 U22891 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19895), .ZN(P2_U3205) );
  AND2_X1 U22892 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19896), .ZN(P2_U3206) );
  AND2_X1 U22893 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19896), .ZN(P2_U3207) );
  AND2_X1 U22894 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19896), .ZN(P2_U3208) );
  INV_X1 U22895 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20067) );
  NOR2_X1 U22896 ( .A1(HOLD), .A2(n20067), .ZN(n19901) );
  NAND2_X1 U22897 ( .A1(NA), .A2(n19902), .ZN(n19907) );
  AND2_X1 U22898 ( .A1(n19897), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19909) );
  NAND2_X1 U22899 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19898) );
  OAI21_X1 U22900 ( .B1(n19909), .B2(n19898), .A(n19913), .ZN(n19899) );
  OAI211_X1 U22901 ( .C1(n19901), .C2(n19900), .A(n19907), .B(n19899), .ZN(
        P2_U3209) );
  NAND2_X1 U22902 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20842), .ZN(n19908) );
  AOI211_X1 U22903 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n19908), .A(n19902), 
        .B(n20067), .ZN(n19903) );
  NOR3_X1 U22904 ( .A1(n20062), .A2(n19909), .A3(n19903), .ZN(n19904) );
  OAI21_X1 U22905 ( .B1(n20842), .B2(n19905), .A(n19904), .ZN(P2_U3210) );
  AOI22_X1 U22906 ( .A1(n19906), .A2(n20067), .B1(n19909), .B2(n21006), .ZN(
        n19912) );
  OAI21_X1 U22907 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19911) );
  OAI211_X1 U22908 ( .C1(n19909), .C2(n19908), .A(P2_STATE_REG_2__SCAN_IN), 
        .B(n19907), .ZN(n19910) );
  OAI21_X1 U22909 ( .B1(n19912), .B2(n19911), .A(n19910), .ZN(P2_U3211) );
  NAND2_X1 U22910 ( .A1(n20071), .A2(n19913), .ZN(n19975) );
  CLKBUF_X1 U22911 ( .A(n19975), .Z(n19970) );
  OAI222_X1 U22912 ( .A1(n19970), .A2(n19917), .B1(n19915), .B2(n20071), .C1(
        n19914), .C2(n19971), .ZN(P2_U3212) );
  OAI222_X1 U22913 ( .A1(n19971), .A2(n19917), .B1(n19916), .B2(n20071), .C1(
        n19919), .C2(n19970), .ZN(P2_U3213) );
  INV_X1 U22914 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19920) );
  OAI222_X1 U22915 ( .A1(n19971), .A2(n19919), .B1(n19918), .B2(n20071), .C1(
        n19920), .C2(n19970), .ZN(P2_U3214) );
  OAI222_X1 U22916 ( .A1(n19975), .A2(n19922), .B1(n19921), .B2(n20071), .C1(
        n19920), .C2(n19971), .ZN(P2_U3215) );
  OAI222_X1 U22917 ( .A1(n19975), .A2(n19924), .B1(n19923), .B2(n20071), .C1(
        n19922), .C2(n19971), .ZN(P2_U3216) );
  OAI222_X1 U22918 ( .A1(n19975), .A2(n15089), .B1(n19925), .B2(n20071), .C1(
        n19924), .C2(n19971), .ZN(P2_U3217) );
  OAI222_X1 U22919 ( .A1(n19975), .A2(n19927), .B1(n19926), .B2(n20071), .C1(
        n15089), .C2(n19971), .ZN(P2_U3218) );
  OAI222_X1 U22920 ( .A1(n19975), .A2(n19929), .B1(n19928), .B2(n20071), .C1(
        n19927), .C2(n19971), .ZN(P2_U3219) );
  OAI222_X1 U22921 ( .A1(n19970), .A2(n15068), .B1(n19930), .B2(n20071), .C1(
        n19929), .C2(n19971), .ZN(P2_U3220) );
  OAI222_X1 U22922 ( .A1(n19970), .A2(n19932), .B1(n19931), .B2(n20071), .C1(
        n15068), .C2(n19971), .ZN(P2_U3221) );
  OAI222_X1 U22923 ( .A1(n19970), .A2(n19934), .B1(n19933), .B2(n20071), .C1(
        n19932), .C2(n19971), .ZN(P2_U3222) );
  OAI222_X1 U22924 ( .A1(n19970), .A2(n19936), .B1(n19935), .B2(n20071), .C1(
        n19934), .C2(n19971), .ZN(P2_U3223) );
  OAI222_X1 U22925 ( .A1(n19970), .A2(n19938), .B1(n19937), .B2(n20071), .C1(
        n19936), .C2(n19971), .ZN(P2_U3224) );
  OAI222_X1 U22926 ( .A1(n19970), .A2(n19940), .B1(n19939), .B2(n20071), .C1(
        n19938), .C2(n19971), .ZN(P2_U3225) );
  OAI222_X1 U22927 ( .A1(n19975), .A2(n19942), .B1(n19941), .B2(n20071), .C1(
        n19940), .C2(n19971), .ZN(P2_U3226) );
  OAI222_X1 U22928 ( .A1(n19975), .A2(n19944), .B1(n19943), .B2(n20071), .C1(
        n19942), .C2(n19971), .ZN(P2_U3227) );
  OAI222_X1 U22929 ( .A1(n19975), .A2(n19946), .B1(n19945), .B2(n20071), .C1(
        n19944), .C2(n19971), .ZN(P2_U3228) );
  INV_X1 U22930 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19948) );
  OAI222_X1 U22931 ( .A1(n19975), .A2(n19948), .B1(n19947), .B2(n20071), .C1(
        n19946), .C2(n19971), .ZN(P2_U3229) );
  OAI222_X1 U22932 ( .A1(n19975), .A2(n19950), .B1(n19949), .B2(n20071), .C1(
        n19948), .C2(n19971), .ZN(P2_U3230) );
  OAI222_X1 U22933 ( .A1(n19975), .A2(n19952), .B1(n19951), .B2(n20071), .C1(
        n19950), .C2(n19971), .ZN(P2_U3231) );
  OAI222_X1 U22934 ( .A1(n19970), .A2(n19954), .B1(n19953), .B2(n20071), .C1(
        n19952), .C2(n19971), .ZN(P2_U3232) );
  INV_X1 U22935 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19956) );
  OAI222_X1 U22936 ( .A1(n19970), .A2(n19956), .B1(n19955), .B2(n20071), .C1(
        n19954), .C2(n19971), .ZN(P2_U3233) );
  OAI222_X1 U22937 ( .A1(n19970), .A2(n19958), .B1(n19957), .B2(n20071), .C1(
        n19956), .C2(n19971), .ZN(P2_U3234) );
  OAI222_X1 U22938 ( .A1(n19970), .A2(n19960), .B1(n19959), .B2(n20071), .C1(
        n19958), .C2(n19971), .ZN(P2_U3235) );
  OAI222_X1 U22939 ( .A1(n19970), .A2(n19962), .B1(n19961), .B2(n20071), .C1(
        n19960), .C2(n19971), .ZN(P2_U3236) );
  OAI222_X1 U22940 ( .A1(n19970), .A2(n19965), .B1(n19963), .B2(n20071), .C1(
        n19962), .C2(n19971), .ZN(P2_U3237) );
  OAI222_X1 U22941 ( .A1(n19971), .A2(n19965), .B1(n19964), .B2(n20071), .C1(
        n19966), .C2(n19970), .ZN(P2_U3238) );
  OAI222_X1 U22942 ( .A1(n19970), .A2(n19968), .B1(n19967), .B2(n20071), .C1(
        n19966), .C2(n19971), .ZN(P2_U3239) );
  INV_X1 U22943 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19972) );
  OAI222_X1 U22944 ( .A1(n19970), .A2(n19972), .B1(n19969), .B2(n20071), .C1(
        n19968), .C2(n19971), .ZN(P2_U3240) );
  INV_X1 U22945 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19973) );
  OAI222_X1 U22946 ( .A1(n19975), .A2(n19974), .B1(n19973), .B2(n20071), .C1(
        n19972), .C2(n19971), .ZN(P2_U3241) );
  INV_X1 U22947 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19976) );
  AOI22_X1 U22948 ( .A1(n20071), .A2(n19977), .B1(n19976), .B2(n20068), .ZN(
        P2_U3585) );
  MUX2_X1 U22949 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20071), .Z(P2_U3586) );
  INV_X1 U22950 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19978) );
  AOI22_X1 U22951 ( .A1(n20071), .A2(n19979), .B1(n19978), .B2(n20068), .ZN(
        P2_U3587) );
  INV_X1 U22952 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19980) );
  AOI22_X1 U22953 ( .A1(n20071), .A2(n19981), .B1(n19980), .B2(n20068), .ZN(
        P2_U3588) );
  OAI21_X1 U22954 ( .B1(n19985), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19983), 
        .ZN(n19982) );
  INV_X1 U22955 ( .A(n19982), .ZN(P2_U3591) );
  OAI21_X1 U22956 ( .B1(n19985), .B2(n19984), .A(n19983), .ZN(P2_U3592) );
  OAI22_X1 U22957 ( .A1(n19987), .A2(n19995), .B1(n19986), .B2(n20004), .ZN(
        n19988) );
  OAI22_X1 U22958 ( .A1(n19999), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19988), .B2(n19996), .ZN(n19989) );
  INV_X1 U22959 ( .A(n19989), .ZN(P2_U3596) );
  INV_X1 U22960 ( .A(n19990), .ZN(n19992) );
  OAI222_X1 U22961 ( .A1(n19995), .A2(n19994), .B1(n20004), .B2(n19993), .C1(
        n19992), .C2(n19991), .ZN(n19997) );
  OAI22_X1 U22962 ( .A1(n19999), .A2(n19998), .B1(n19997), .B2(n19996), .ZN(
        n20000) );
  INV_X1 U22963 ( .A(n20000), .ZN(P2_U3600) );
  NOR2_X1 U22964 ( .A1(n20002), .A2(n20001), .ZN(n20024) );
  NAND2_X1 U22965 ( .A1(n20003), .A2(n20024), .ZN(n20013) );
  NAND3_X1 U22966 ( .A1(n20022), .A2(n20004), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20005) );
  NAND2_X1 U22967 ( .A1(n20005), .A2(n20020), .ZN(n20014) );
  NAND2_X1 U22968 ( .A1(n20013), .A2(n20014), .ZN(n20010) );
  AOI222_X1 U22969 ( .A1(n20010), .A2(n20009), .B1(n20008), .B2(
        P2_STATE2_REG_3__SCAN_IN), .C1(n20007), .C2(n20006), .ZN(n20011) );
  AOI22_X1 U22970 ( .A1(n20034), .A2(n20012), .B1(n20011), .B2(n20035), .ZN(
        P2_U3602) );
  OAI21_X1 U22971 ( .B1(n20015), .B2(n20014), .A(n20013), .ZN(n20016) );
  AOI21_X1 U22972 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20017), .A(n20016), 
        .ZN(n20018) );
  AOI22_X1 U22973 ( .A1(n20034), .A2(n20019), .B1(n20018), .B2(n20035), .ZN(
        P2_U3603) );
  INV_X1 U22974 ( .A(n20020), .ZN(n20030) );
  AND2_X1 U22975 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20021) );
  NOR2_X1 U22976 ( .A1(n20030), .A2(n20021), .ZN(n20023) );
  MUX2_X1 U22977 ( .A(n20024), .B(n20023), .S(n20022), .Z(n20025) );
  AOI21_X1 U22978 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20026), .A(n20025), 
        .ZN(n20027) );
  AOI22_X1 U22979 ( .A1(n20034), .A2(n20028), .B1(n20027), .B2(n20035), .ZN(
        P2_U3604) );
  OAI21_X1 U22980 ( .B1(n20031), .B2(n20030), .A(n20029), .ZN(n20032) );
  AOI21_X1 U22981 ( .B1(n20036), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20032), 
        .ZN(n20033) );
  OAI22_X1 U22982 ( .A1(n20036), .A2(n20035), .B1(n20034), .B2(n20033), .ZN(
        P2_U3605) );
  INV_X1 U22983 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20037) );
  AOI22_X1 U22984 ( .A1(n20071), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20037), 
        .B2(n20068), .ZN(P2_U3608) );
  INV_X1 U22985 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n20050) );
  INV_X1 U22986 ( .A(n20038), .ZN(n20049) );
  INV_X1 U22987 ( .A(n20039), .ZN(n20043) );
  INV_X1 U22988 ( .A(n20040), .ZN(n20041) );
  OAI22_X1 U22989 ( .A1(n20044), .A2(n20043), .B1(n20042), .B2(n20041), .ZN(
        n20045) );
  INV_X1 U22990 ( .A(n20045), .ZN(n20048) );
  NOR2_X1 U22991 ( .A1(n20049), .A2(n20046), .ZN(n20047) );
  AOI22_X1 U22992 ( .A1(n20050), .A2(n20049), .B1(n20048), .B2(n20047), .ZN(
        P2_U3609) );
  AOI21_X1 U22993 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20051), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20053) );
  AOI211_X1 U22994 ( .C1(n20057), .C2(n19227), .A(n20053), .B(n20052), .ZN(
        n20066) );
  NOR4_X1 U22995 ( .A1(n20062), .A2(n12173), .A3(n20055), .A4(n20054), .ZN(
        n20059) );
  AOI21_X1 U22996 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20057), .A(n20056), 
        .ZN(n20058) );
  NOR2_X1 U22997 ( .A1(n20059), .A2(n20058), .ZN(n20065) );
  AOI211_X1 U22998 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n20062), .A(n20061), 
        .B(n12584), .ZN(n20063) );
  NOR2_X1 U22999 ( .A1(n20066), .A2(n20063), .ZN(n20064) );
  AOI22_X1 U23000 ( .A1(n20067), .A2(n20066), .B1(n20065), .B2(n20064), .ZN(
        P2_U3610) );
  INV_X1 U23001 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20069) );
  AOI22_X1 U23002 ( .A1(n20071), .A2(n20070), .B1(n20069), .B2(n20068), .ZN(
        P2_U3611) );
  AND2_X1 U23003 ( .A1(n20845), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20073) );
  INV_X1 U23004 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20072) );
  INV_X2 U23005 ( .A(n20944), .ZN(n20890) );
  AOI21_X1 U23006 ( .B1(n20073), .B2(n20072), .A(n20890), .ZN(P1_U2802) );
  OAI21_X1 U23007 ( .B1(n20075), .B2(n20074), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20076) );
  OAI21_X1 U23008 ( .B1(n20077), .B2(n20936), .A(n20076), .ZN(P1_U2803) );
  NOR2_X1 U23009 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20079) );
  OAI21_X1 U23010 ( .B1(n20079), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20944), .ZN(
        n20078) );
  OAI21_X1 U23011 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20944), .A(n20078), 
        .ZN(P1_U2804) );
  AOI21_X1 U23012 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20845), .A(n20890), 
        .ZN(n20903) );
  OAI21_X1 U23013 ( .B1(BS16), .B2(n20079), .A(n20903), .ZN(n20901) );
  OAI21_X1 U23014 ( .B1(n20903), .B2(n21137), .A(n20901), .ZN(P1_U2805) );
  OAI21_X1 U23015 ( .B1(n20081), .B2(n21151), .A(n20080), .ZN(P1_U2806) );
  NOR4_X1 U23016 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20085) );
  NOR4_X1 U23017 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20084) );
  NOR4_X1 U23018 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20083) );
  NOR4_X1 U23019 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20082) );
  NAND4_X1 U23020 ( .A1(n20085), .A2(n20084), .A3(n20083), .A4(n20082), .ZN(
        n20091) );
  NOR4_X1 U23021 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20089) );
  AOI211_X1 U23022 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20088) );
  NOR4_X1 U23023 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20087) );
  NOR4_X1 U23024 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20086) );
  NAND4_X1 U23025 ( .A1(n20089), .A2(n20088), .A3(n20087), .A4(n20086), .ZN(
        n20090) );
  NOR2_X1 U23026 ( .A1(n20091), .A2(n20090), .ZN(n20926) );
  INV_X1 U23027 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20896) );
  NOR3_X1 U23028 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20093) );
  OAI21_X1 U23029 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20093), .A(n20926), .ZN(
        n20092) );
  OAI21_X1 U23030 ( .B1(n20926), .B2(n20896), .A(n20092), .ZN(P1_U2807) );
  INV_X1 U23031 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20902) );
  AOI21_X1 U23032 ( .B1(n21275), .B2(n20902), .A(n20093), .ZN(n20094) );
  INV_X1 U23033 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21074) );
  INV_X1 U23034 ( .A(n20926), .ZN(n20928) );
  AOI22_X1 U23035 ( .A1(n20926), .A2(n20094), .B1(n21074), .B2(n20928), .ZN(
        P1_U2808) );
  NOR2_X1 U23036 ( .A1(n20095), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n20104) );
  AOI22_X1 U23037 ( .A1(n20161), .A2(n20130), .B1(n20127), .B2(n20096), .ZN(
        n20103) );
  OAI21_X1 U23038 ( .B1(n20098), .B2(n20097), .A(n20134), .ZN(n20101) );
  NOR2_X1 U23039 ( .A1(n20163), .A2(n20099), .ZN(n20100) );
  AOI211_X1 U23040 ( .C1(n20152), .C2(P1_EBX_REG_9__SCAN_IN), .A(n20101), .B(
        n20100), .ZN(n20102) );
  OAI211_X1 U23041 ( .C1(n20105), .C2(n20104), .A(n20103), .B(n20102), .ZN(
        P1_U2831) );
  OR2_X1 U23042 ( .A1(n20112), .A2(n20106), .ZN(n20118) );
  NOR2_X1 U23043 ( .A1(n20107), .A2(n20168), .ZN(n20108) );
  AOI211_X1 U23044 ( .C1(n20139), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20138), .B(n20108), .ZN(n20109) );
  OAI21_X1 U23045 ( .B1(n20110), .B2(n20142), .A(n20109), .ZN(n20111) );
  AOI21_X1 U23046 ( .B1(n20130), .B2(n9917), .A(n20111), .ZN(n20114) );
  AOI22_X1 U23047 ( .A1(n20166), .A2(n20123), .B1(n21261), .B2(n20112), .ZN(
        n20113) );
  OAI211_X1 U23048 ( .C1(n21261), .C2(n20118), .A(n20114), .B(n20113), .ZN(
        P1_U2833) );
  AOI22_X1 U23049 ( .A1(n20152), .A2(P1_EBX_REG_6__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20139), .ZN(n20126) );
  OAI21_X1 U23050 ( .B1(n20117), .B2(n20116), .A(n20115), .ZN(n20149) );
  NAND2_X1 U23051 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20149), .ZN(n20132) );
  AOI21_X1 U23052 ( .B1(n21255), .B2(n20132), .A(n20118), .ZN(n20122) );
  OAI22_X1 U23053 ( .A1(n20120), .A2(n20142), .B1(n20119), .B2(n20155), .ZN(
        n20121) );
  AOI211_X1 U23054 ( .C1(n20124), .C2(n20123), .A(n20122), .B(n20121), .ZN(
        n20125) );
  NAND3_X1 U23055 ( .A1(n20126), .A2(n20125), .A3(n20134), .ZN(P1_U2834) );
  AOI22_X1 U23056 ( .A1(n20128), .A2(n20127), .B1(n20152), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n20137) );
  INV_X1 U23057 ( .A(n20169), .ZN(n20129) );
  AOI22_X1 U23058 ( .A1(n20130), .A2(n20129), .B1(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20139), .ZN(n20136) );
  INV_X1 U23059 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21121) );
  NAND2_X1 U23060 ( .A1(n20131), .A2(n21121), .ZN(n20133) );
  AOI22_X1 U23061 ( .A1(n20171), .A2(n20157), .B1(n20133), .B2(n20132), .ZN(
        n20135) );
  NAND4_X1 U23062 ( .A1(n20137), .A2(n20136), .A3(n20135), .A4(n20134), .ZN(
        P1_U2835) );
  AOI21_X1 U23063 ( .B1(n20139), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20138), .ZN(n20140) );
  OAI21_X1 U23064 ( .B1(n20142), .B2(n20141), .A(n20140), .ZN(n20143) );
  AOI21_X1 U23065 ( .B1(n20145), .B2(n20144), .A(n20143), .ZN(n20160) );
  NOR3_X1 U23066 ( .A1(n20148), .A2(n20147), .A3(n20146), .ZN(n20151) );
  NOR2_X1 U23067 ( .A1(n20149), .A2(n21299), .ZN(n20150) );
  AOI211_X1 U23068 ( .C1(n20152), .C2(P1_EBX_REG_4__SCAN_IN), .A(n20151), .B(
        n20150), .ZN(n20153) );
  OAI21_X1 U23069 ( .B1(n20155), .B2(n20154), .A(n20153), .ZN(n20156) );
  AOI21_X1 U23070 ( .B1(n20158), .B2(n20157), .A(n20156), .ZN(n20159) );
  NAND2_X1 U23071 ( .A1(n20160), .A2(n20159), .ZN(P1_U2836) );
  INV_X1 U23072 ( .A(n20161), .ZN(n20162) );
  OAI22_X1 U23073 ( .A1(n20163), .A2(n14532), .B1(n14521), .B2(n20162), .ZN(
        n20164) );
  INV_X1 U23074 ( .A(n20164), .ZN(n20165) );
  OAI21_X1 U23075 ( .B1(n20179), .B2(n21307), .A(n20165), .ZN(P1_U2863) );
  AOI22_X1 U23076 ( .A1(n20166), .A2(n20176), .B1(n20175), .B2(n9917), .ZN(
        n20167) );
  OAI21_X1 U23077 ( .B1(n20179), .B2(n20168), .A(n20167), .ZN(P1_U2865) );
  NOR2_X1 U23078 ( .A1(n20169), .A2(n14521), .ZN(n20170) );
  AOI21_X1 U23079 ( .B1(n20171), .B2(n20176), .A(n20170), .ZN(n20172) );
  OAI21_X1 U23080 ( .B1(n20179), .B2(n20173), .A(n20172), .ZN(P1_U2867) );
  AOI22_X1 U23081 ( .A1(n20177), .A2(n20176), .B1(n20175), .B2(n20174), .ZN(
        n20178) );
  OAI21_X1 U23082 ( .B1(n20179), .B2(n21284), .A(n20178), .ZN(P1_U2869) );
  AOI22_X1 U23083 ( .A1(n20941), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20181) );
  OAI21_X1 U23084 ( .B1(n20182), .B2(n20210), .A(n20181), .ZN(P1_U2921) );
  INV_X1 U23085 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20184) );
  AOI22_X1 U23086 ( .A1(n20941), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20183) );
  OAI21_X1 U23087 ( .B1(n20184), .B2(n20210), .A(n20183), .ZN(P1_U2922) );
  INV_X1 U23088 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20186) );
  AOI22_X1 U23089 ( .A1(n20941), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20185) );
  OAI21_X1 U23090 ( .B1(n20186), .B2(n20210), .A(n20185), .ZN(P1_U2923) );
  INV_X1 U23091 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20188) );
  AOI22_X1 U23092 ( .A1(n20941), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20187) );
  OAI21_X1 U23093 ( .B1(n20188), .B2(n20210), .A(n20187), .ZN(P1_U2924) );
  INV_X1 U23094 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20190) );
  AOI22_X1 U23095 ( .A1(n20941), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20189) );
  OAI21_X1 U23096 ( .B1(n20190), .B2(n20210), .A(n20189), .ZN(P1_U2925) );
  INV_X1 U23097 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20192) );
  AOI22_X1 U23098 ( .A1(n20941), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20191) );
  OAI21_X1 U23099 ( .B1(n20192), .B2(n20210), .A(n20191), .ZN(P1_U2926) );
  INV_X1 U23100 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20194) );
  AOI22_X1 U23101 ( .A1(n20941), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20193) );
  OAI21_X1 U23102 ( .B1(n20194), .B2(n20210), .A(n20193), .ZN(P1_U2927) );
  AOI22_X1 U23103 ( .A1(n20941), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20196) );
  OAI21_X1 U23104 ( .B1(n20197), .B2(n20210), .A(n20196), .ZN(P1_U2928) );
  AOI22_X1 U23105 ( .A1(n20941), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20198) );
  OAI21_X1 U23106 ( .B1(n10706), .B2(n20210), .A(n20198), .ZN(P1_U2929) );
  AOI22_X1 U23107 ( .A1(n20941), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20199) );
  OAI21_X1 U23108 ( .B1(n10696), .B2(n20210), .A(n20199), .ZN(P1_U2930) );
  AOI22_X1 U23109 ( .A1(n20941), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20200) );
  OAI21_X1 U23110 ( .B1(n10675), .B2(n20210), .A(n20200), .ZN(P1_U2931) );
  AOI22_X1 U23111 ( .A1(n20941), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20201) );
  OAI21_X1 U23112 ( .B1(n20202), .B2(n20210), .A(n20201), .ZN(P1_U2932) );
  AOI22_X1 U23113 ( .A1(n20941), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20203) );
  OAI21_X1 U23114 ( .B1(n20204), .B2(n20210), .A(n20203), .ZN(P1_U2933) );
  AOI22_X1 U23115 ( .A1(n20941), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20205) );
  OAI21_X1 U23116 ( .B1(n20206), .B2(n20210), .A(n20205), .ZN(P1_U2934) );
  AOI22_X1 U23117 ( .A1(n20941), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20207) );
  OAI21_X1 U23118 ( .B1(n20208), .B2(n20210), .A(n20207), .ZN(P1_U2935) );
  AOI22_X1 U23119 ( .A1(n20941), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20195), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20209) );
  OAI21_X1 U23120 ( .B1(n20211), .B2(n20210), .A(n20209), .ZN(P1_U2936) );
  AOI22_X1 U23121 ( .A1(n20251), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20223), .ZN(n20213) );
  OAI21_X1 U23122 ( .B1(n20267), .B2(n20253), .A(n20213), .ZN(P1_U2937) );
  AOI22_X1 U23123 ( .A1(n20251), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20223), .ZN(n20214) );
  OAI21_X1 U23124 ( .B1(n20276), .B2(n20253), .A(n20214), .ZN(P1_U2938) );
  AOI22_X1 U23125 ( .A1(n20251), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20223), .ZN(n20215) );
  OAI21_X1 U23126 ( .B1(n20283), .B2(n20253), .A(n20215), .ZN(P1_U2939) );
  AOI22_X1 U23127 ( .A1(n20251), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20223), .ZN(n20216) );
  OAI21_X1 U23128 ( .B1(n20288), .B2(n20253), .A(n20216), .ZN(P1_U2940) );
  AOI22_X1 U23129 ( .A1(n20251), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20223), .ZN(n20217) );
  OAI21_X1 U23130 ( .B1(n20227), .B2(n20253), .A(n20217), .ZN(P1_U2941) );
  AOI22_X1 U23131 ( .A1(n20251), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20223), .ZN(n20218) );
  OAI21_X1 U23132 ( .B1(n20295), .B2(n20253), .A(n20218), .ZN(P1_U2942) );
  AOI22_X1 U23133 ( .A1(n20251), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20223), .ZN(n20219) );
  OAI21_X1 U23134 ( .B1(n20303), .B2(n20253), .A(n20219), .ZN(P1_U2943) );
  AOI22_X1 U23135 ( .A1(n20251), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20223), .ZN(n20220) );
  OAI21_X1 U23136 ( .B1(n20231), .B2(n20253), .A(n20220), .ZN(P1_U2944) );
  AOI22_X1 U23137 ( .A1(n20251), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20223), .ZN(n20221) );
  OAI21_X1 U23138 ( .B1(n20267), .B2(n20253), .A(n20221), .ZN(P1_U2952) );
  AOI22_X1 U23139 ( .A1(n20251), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20223), .ZN(n20222) );
  OAI21_X1 U23140 ( .B1(n20276), .B2(n20253), .A(n20222), .ZN(P1_U2953) );
  AOI22_X1 U23141 ( .A1(n20251), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20223), .ZN(n20224) );
  OAI21_X1 U23142 ( .B1(n20283), .B2(n20253), .A(n20224), .ZN(P1_U2954) );
  AOI22_X1 U23143 ( .A1(n20251), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20223), .ZN(n20225) );
  OAI21_X1 U23144 ( .B1(n20288), .B2(n20253), .A(n20225), .ZN(P1_U2955) );
  AOI22_X1 U23145 ( .A1(n20251), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20223), .ZN(n20226) );
  OAI21_X1 U23146 ( .B1(n20227), .B2(n20253), .A(n20226), .ZN(P1_U2956) );
  AOI22_X1 U23147 ( .A1(n20251), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20223), .ZN(n20228) );
  OAI21_X1 U23148 ( .B1(n20295), .B2(n20253), .A(n20228), .ZN(P1_U2957) );
  AOI22_X1 U23149 ( .A1(n20251), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20223), .ZN(n20229) );
  OAI21_X1 U23150 ( .B1(n20303), .B2(n20253), .A(n20229), .ZN(P1_U2958) );
  AOI22_X1 U23151 ( .A1(n20251), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20223), .ZN(n20230) );
  OAI21_X1 U23152 ( .B1(n20231), .B2(n20253), .A(n20230), .ZN(P1_U2959) );
  AOI22_X1 U23153 ( .A1(n20251), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20223), .ZN(n20234) );
  NAND2_X1 U23154 ( .A1(n20248), .A2(n20232), .ZN(n20233) );
  NAND2_X1 U23155 ( .A1(n20234), .A2(n20233), .ZN(P1_U2961) );
  AOI22_X1 U23156 ( .A1(n20251), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20223), .ZN(n20237) );
  NAND2_X1 U23157 ( .A1(n20248), .A2(n20235), .ZN(n20236) );
  NAND2_X1 U23158 ( .A1(n20237), .A2(n20236), .ZN(P1_U2962) );
  AOI22_X1 U23159 ( .A1(n20251), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20223), .ZN(n20240) );
  NAND2_X1 U23160 ( .A1(n20248), .A2(n20238), .ZN(n20239) );
  NAND2_X1 U23161 ( .A1(n20240), .A2(n20239), .ZN(P1_U2963) );
  AOI22_X1 U23162 ( .A1(n20251), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20223), .ZN(n20243) );
  NAND2_X1 U23163 ( .A1(n20248), .A2(n20241), .ZN(n20242) );
  NAND2_X1 U23164 ( .A1(n20243), .A2(n20242), .ZN(P1_U2964) );
  AOI22_X1 U23165 ( .A1(n20251), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20223), .ZN(n20246) );
  NAND2_X1 U23166 ( .A1(n20248), .A2(n20244), .ZN(n20245) );
  NAND2_X1 U23167 ( .A1(n20246), .A2(n20245), .ZN(P1_U2965) );
  AOI22_X1 U23168 ( .A1(n20251), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20223), .ZN(n20250) );
  NAND2_X1 U23169 ( .A1(n20248), .A2(n20247), .ZN(n20249) );
  NAND2_X1 U23170 ( .A1(n20250), .A2(n20249), .ZN(P1_U2966) );
  AOI22_X1 U23171 ( .A1(n20251), .A2(P1_EAX_REG_15__SCAN_IN), .B1(
        P1_LWORD_REG_15__SCAN_IN), .B2(n20223), .ZN(n20252) );
  OAI21_X1 U23172 ( .B1(n20254), .B2(n20253), .A(n20252), .ZN(P1_U2967) );
  OAI211_X1 U23173 ( .C1(n20258), .C2(n20257), .A(n20256), .B(n20255), .ZN(
        n20259) );
  AOI21_X1 U23174 ( .B1(n20261), .B2(n20260), .A(n20259), .ZN(n20262) );
  OAI221_X1 U23175 ( .B1(n20265), .B2(n20264), .C1(n20265), .C2(n20263), .A(
        n20262), .ZN(P1_U3031) );
  NOR2_X1 U23176 ( .A1(n11147), .A2(n20923), .ZN(P1_U3032) );
  INV_X1 U23177 ( .A(DATAI_24_), .ZN(n21262) );
  OAI22_X2 U23178 ( .A1(n14567), .A2(n20306), .B1(n21262), .B2(n20304), .ZN(
        n20738) );
  NOR2_X2 U23179 ( .A1(n20273), .A2(n20266), .ZN(n20774) );
  AOI22_X1 U23180 ( .A1(n20828), .A2(n20738), .B1(n20294), .B2(n20774), .ZN(
        n20270) );
  INV_X1 U23181 ( .A(DATAI_16_), .ZN(n21073) );
  AOI22_X1 U23182 ( .A1(n20773), .A2(n20307), .B1(n20334), .B2(n20781), .ZN(
        n20269) );
  OAI211_X1 U23183 ( .C1(n20311), .C2(n20271), .A(n20270), .B(n20269), .ZN(
        P1_U3033) );
  INV_X1 U23184 ( .A(DATAI_25_), .ZN(n20272) );
  INV_X1 U23185 ( .A(n20787), .ZN(n20709) );
  INV_X1 U23186 ( .A(n20294), .ZN(n20301) );
  NAND2_X1 U23187 ( .A1(n20300), .A2(n20274), .ZN(n20665) );
  OAI22_X1 U23188 ( .A1(n20803), .A2(n20709), .B1(n20301), .B2(n20665), .ZN(
        n20275) );
  INV_X1 U23189 ( .A(n20275), .ZN(n20280) );
  INV_X1 U23190 ( .A(DATAI_17_), .ZN(n20278) );
  OAI22_X1 U23191 ( .A1(n20278), .A2(n20304), .B1(n20277), .B2(n20306), .ZN(
        n20706) );
  AOI22_X1 U23192 ( .A1(n20785), .A2(n20307), .B1(n20334), .B2(n20706), .ZN(
        n20279) );
  OAI211_X1 U23193 ( .C1(n20311), .C2(n10525), .A(n20280), .B(n20279), .ZN(
        P1_U3034) );
  INV_X1 U23194 ( .A(DATAI_26_), .ZN(n21156) );
  OAI22_X1 U23195 ( .A1(n15260), .A2(n20306), .B1(n21156), .B2(n20304), .ZN(
        n20744) );
  INV_X1 U23196 ( .A(n20744), .ZN(n20796) );
  NAND2_X1 U23197 ( .A1(n20300), .A2(n20281), .ZN(n20353) );
  OAI22_X1 U23198 ( .A1(n20803), .A2(n20796), .B1(n20301), .B2(n20353), .ZN(
        n20282) );
  INV_X1 U23199 ( .A(n20282), .ZN(n20285) );
  INV_X1 U23200 ( .A(DATAI_18_), .ZN(n21140) );
  OAI22_X2 U23201 ( .A1(n21140), .A2(n20304), .B1(n15322), .B2(n20306), .ZN(
        n20793) );
  AOI22_X1 U23202 ( .A1(n20791), .A2(n20307), .B1(n20334), .B2(n20793), .ZN(
        n20284) );
  OAI211_X1 U23203 ( .C1(n20311), .C2(n20286), .A(n20285), .B(n20284), .ZN(
        P1_U3035) );
  INV_X1 U23204 ( .A(DATAI_27_), .ZN(n21169) );
  OAI22_X2 U23205 ( .A1(n14551), .A2(n20306), .B1(n21169), .B2(n20304), .ZN(
        n20799) );
  NAND2_X1 U23206 ( .A1(n20300), .A2(n20287), .ZN(n20596) );
  AOI22_X1 U23207 ( .A1(n20828), .A2(n20799), .B1(n20294), .B2(n20798), .ZN(
        n20291) );
  INV_X1 U23208 ( .A(DATAI_19_), .ZN(n20289) );
  OAI22_X1 U23209 ( .A1(n20289), .A2(n20304), .B1(n14593), .B2(n20306), .ZN(
        n20712) );
  AOI22_X1 U23210 ( .A1(n20797), .A2(n20307), .B1(n20334), .B2(n20712), .ZN(
        n20290) );
  OAI211_X1 U23211 ( .C1(n20311), .C2(n20292), .A(n20291), .B(n20290), .ZN(
        P1_U3036) );
  INV_X1 U23212 ( .A(DATAI_29_), .ZN(n20293) );
  NAND2_X1 U23213 ( .A1(n20300), .A2(n10450), .ZN(n20364) );
  AOI22_X1 U23214 ( .A1(n20828), .A2(n20754), .B1(n20294), .B2(n20812), .ZN(
        n20298) );
  INV_X1 U23215 ( .A(DATAI_21_), .ZN(n21277) );
  OAI22_X2 U23216 ( .A1(n20296), .A2(n20306), .B1(n21277), .B2(n20304), .ZN(
        n20813) );
  AOI22_X1 U23217 ( .A1(n20811), .A2(n20307), .B1(n20334), .B2(n20813), .ZN(
        n20297) );
  OAI211_X1 U23218 ( .C1(n20311), .C2(n20299), .A(n20298), .B(n20297), .ZN(
        P1_U3038) );
  INV_X1 U23219 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20310) );
  INV_X1 U23220 ( .A(DATAI_30_), .ZN(n21128) );
  OAI22_X1 U23221 ( .A1(n14535), .A2(n20306), .B1(n21128), .B2(n20304), .ZN(
        n20758) );
  INV_X1 U23222 ( .A(n20758), .ZN(n20822) );
  NAND2_X1 U23223 ( .A1(n20300), .A2(n10574), .ZN(n20683) );
  OAI22_X1 U23224 ( .A1(n20803), .A2(n20822), .B1(n20301), .B2(n20683), .ZN(
        n20302) );
  INV_X1 U23225 ( .A(n20302), .ZN(n20309) );
  INV_X1 U23226 ( .A(DATAI_22_), .ZN(n20305) );
  OAI22_X1 U23227 ( .A1(n14579), .A2(n20306), .B1(n20305), .B2(n20304), .ZN(
        n20819) );
  AOI22_X1 U23228 ( .A1(n20817), .A2(n20307), .B1(n20334), .B2(n20819), .ZN(
        n20308) );
  OAI211_X1 U23229 ( .C1(n20311), .C2(n20310), .A(n20309), .B(n20308), .ZN(
        P1_U3039) );
  INV_X1 U23230 ( .A(n20781), .ZN(n20741) );
  INV_X1 U23231 ( .A(n20703), .ZN(n20444) );
  INV_X1 U23232 ( .A(n20380), .ZN(n20313) );
  INV_X1 U23233 ( .A(n20312), .ZN(n20551) );
  NOR2_X1 U23234 ( .A1(n20696), .A2(n20314), .ZN(n20332) );
  AOI21_X1 U23235 ( .B1(n20313), .B2(n20551), .A(n20332), .ZN(n20315) );
  OAI22_X1 U23236 ( .A1(n20315), .A2(n20920), .B1(n20314), .B2(n10577), .ZN(
        n20333) );
  AOI22_X1 U23237 ( .A1(n20773), .A2(n20333), .B1(n20774), .B2(n20332), .ZN(
        n20319) );
  INV_X1 U23238 ( .A(n20314), .ZN(n20317) );
  OR2_X1 U23239 ( .A1(n20339), .A2(n21137), .ZN(n20701) );
  OAI21_X1 U23240 ( .B1(n20383), .B2(n20701), .A(n20315), .ZN(n20316) );
  OAI221_X1 U23241 ( .B1(n20698), .B2(n20317), .C1(n20920), .C2(n20316), .A(
        n20779), .ZN(n20335) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20738), .ZN(n20318) );
  OAI211_X1 U23243 ( .C1(n20741), .C2(n20372), .A(n20319), .B(n20318), .ZN(
        P1_U3041) );
  AOI22_X1 U23244 ( .A1(n20786), .A2(n20332), .B1(n20333), .B2(n20785), .ZN(
        n20321) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20787), .ZN(n20320) );
  OAI211_X1 U23246 ( .C1(n20790), .C2(n20372), .A(n20321), .B(n20320), .ZN(
        P1_U3042) );
  INV_X1 U23247 ( .A(n20793), .ZN(n20747) );
  AOI22_X1 U23248 ( .A1(n20792), .A2(n20332), .B1(n20333), .B2(n20791), .ZN(
        n20323) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20744), .ZN(n20322) );
  OAI211_X1 U23250 ( .C1(n20747), .C2(n20372), .A(n20323), .B(n20322), .ZN(
        P1_U3043) );
  INV_X1 U23251 ( .A(n20712), .ZN(n20804) );
  AOI22_X1 U23252 ( .A1(n20798), .A2(n20332), .B1(n20333), .B2(n20797), .ZN(
        n20325) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20799), .ZN(n20324) );
  OAI211_X1 U23254 ( .C1(n20804), .C2(n20372), .A(n20325), .B(n20324), .ZN(
        P1_U3044) );
  INV_X1 U23255 ( .A(n20807), .ZN(n20753) );
  AOI22_X1 U23256 ( .A1(n20806), .A2(n20333), .B1(n20805), .B2(n20332), .ZN(
        n20327) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20750), .ZN(n20326) );
  OAI211_X1 U23258 ( .C1(n20753), .C2(n20372), .A(n20327), .B(n20326), .ZN(
        P1_U3045) );
  INV_X1 U23259 ( .A(n20813), .ZN(n20757) );
  AOI22_X1 U23260 ( .A1(n20812), .A2(n20332), .B1(n20811), .B2(n20333), .ZN(
        n20329) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20754), .ZN(n20328) );
  OAI211_X1 U23262 ( .C1(n20757), .C2(n20372), .A(n20329), .B(n20328), .ZN(
        P1_U3046) );
  INV_X1 U23263 ( .A(n20819), .ZN(n20761) );
  AOI22_X1 U23264 ( .A1(n20818), .A2(n20332), .B1(n20817), .B2(n20333), .ZN(
        n20331) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20758), .ZN(n20330) );
  OAI211_X1 U23266 ( .C1(n20761), .C2(n20372), .A(n20331), .B(n20330), .ZN(
        P1_U3047) );
  INV_X1 U23267 ( .A(n20827), .ZN(n20769) );
  AOI22_X1 U23268 ( .A1(n20826), .A2(n20333), .B1(n20824), .B2(n20332), .ZN(
        n20337) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20335), .B1(
        n20334), .B2(n20764), .ZN(n20336) );
  OAI211_X1 U23270 ( .C1(n20769), .C2(n20372), .A(n20337), .B(n20336), .ZN(
        P1_U3048) );
  NAND2_X1 U23271 ( .A1(n20372), .A2(n20698), .ZN(n20340) );
  INV_X1 U23272 ( .A(n20915), .ZN(n20650) );
  OAI21_X1 U23273 ( .B1(n20405), .B2(n20340), .A(n20650), .ZN(n20342) );
  NOR2_X1 U23274 ( .A1(n20380), .A2(n13559), .ZN(n20345) );
  INV_X1 U23275 ( .A(n20773), .ZN(n20664) );
  NOR3_X1 U23276 ( .A1(n20655), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20385) );
  NAND2_X1 U23277 ( .A1(n20696), .A2(n20385), .ZN(n20371) );
  INV_X1 U23278 ( .A(n20371), .ZN(n20341) );
  AOI22_X1 U23279 ( .A1(n20405), .A2(n20781), .B1(n20774), .B2(n20341), .ZN(
        n20349) );
  INV_X1 U23280 ( .A(n20342), .ZN(n20346) );
  NOR2_X1 U23281 ( .A1(n10347), .A2(n10577), .ZN(n20469) );
  AOI211_X1 U23282 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20371), .A(n20469), 
        .B(n20343), .ZN(n20344) );
  INV_X1 U23283 ( .A(n20372), .ZN(n20347) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20374), .B1(
        n20347), .B2(n20738), .ZN(n20348) );
  OAI211_X1 U23285 ( .C1(n20377), .C2(n20664), .A(n20349), .B(n20348), .ZN(
        P1_U3049) );
  OAI22_X1 U23286 ( .A1(n20372), .A2(n20709), .B1(n20665), .B2(n20371), .ZN(
        n20350) );
  INV_X1 U23287 ( .A(n20350), .ZN(n20352) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20706), .ZN(n20351) );
  OAI211_X1 U23289 ( .C1(n20377), .C2(n20669), .A(n20352), .B(n20351), .ZN(
        P1_U3050) );
  INV_X1 U23290 ( .A(n20791), .ZN(n20672) );
  OAI22_X1 U23291 ( .A1(n20372), .A2(n20796), .B1(n20353), .B2(n20371), .ZN(
        n20354) );
  INV_X1 U23292 ( .A(n20354), .ZN(n20356) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20793), .ZN(n20355) );
  OAI211_X1 U23294 ( .C1(n20377), .C2(n20672), .A(n20356), .B(n20355), .ZN(
        P1_U3051) );
  INV_X1 U23295 ( .A(n20797), .ZN(n20675) );
  INV_X1 U23296 ( .A(n20799), .ZN(n20715) );
  OAI22_X1 U23297 ( .A1(n20372), .A2(n20715), .B1(n20596), .B2(n20371), .ZN(
        n20357) );
  INV_X1 U23298 ( .A(n20357), .ZN(n20359) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20712), .ZN(n20358) );
  OAI211_X1 U23300 ( .C1(n20377), .C2(n20675), .A(n20359), .B(n20358), .ZN(
        P1_U3052) );
  INV_X1 U23301 ( .A(n20806), .ZN(n20678) );
  INV_X1 U23302 ( .A(n20805), .ZN(n20360) );
  OAI22_X1 U23303 ( .A1(n20372), .A2(n20810), .B1(n20360), .B2(n20371), .ZN(
        n20361) );
  INV_X1 U23304 ( .A(n20361), .ZN(n20363) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20807), .ZN(n20362) );
  OAI211_X1 U23306 ( .C1(n20377), .C2(n20678), .A(n20363), .B(n20362), .ZN(
        P1_U3053) );
  INV_X1 U23307 ( .A(n20811), .ZN(n20681) );
  INV_X1 U23308 ( .A(n20754), .ZN(n20816) );
  OAI22_X1 U23309 ( .A1(n20372), .A2(n20816), .B1(n20364), .B2(n20371), .ZN(
        n20365) );
  INV_X1 U23310 ( .A(n20365), .ZN(n20367) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20813), .ZN(n20366) );
  OAI211_X1 U23312 ( .C1(n20377), .C2(n20681), .A(n20367), .B(n20366), .ZN(
        P1_U3054) );
  OAI22_X1 U23313 ( .A1(n20372), .A2(n20822), .B1(n20683), .B2(n20371), .ZN(
        n20368) );
  INV_X1 U23314 ( .A(n20368), .ZN(n20370) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20819), .ZN(n20369) );
  OAI211_X1 U23316 ( .C1(n20377), .C2(n20687), .A(n20370), .B(n20369), .ZN(
        P1_U3055) );
  INV_X1 U23317 ( .A(n20826), .ZN(n20694) );
  INV_X1 U23318 ( .A(n20824), .ZN(n20610) );
  OAI22_X1 U23319 ( .A1(n20372), .A2(n20833), .B1(n20610), .B2(n20371), .ZN(
        n20373) );
  INV_X1 U23320 ( .A(n20373), .ZN(n20376) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20827), .ZN(n20375) );
  OAI211_X1 U23322 ( .C1(n20377), .C2(n20694), .A(n20376), .B(n20375), .ZN(
        P1_U3056) );
  AND2_X1 U23323 ( .A1(n20378), .A2(n10591), .ZN(n20619) );
  INV_X1 U23324 ( .A(n20619), .ZN(n20771) );
  NOR2_X1 U23325 ( .A1(n20618), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20404) );
  INV_X1 U23326 ( .A(n20404), .ZN(n20379) );
  OAI21_X1 U23327 ( .B1(n20380), .B2(n20771), .A(n20379), .ZN(n20388) );
  INV_X1 U23328 ( .A(n20623), .ZN(n20381) );
  AOI21_X1 U23329 ( .B1(n20382), .B2(n20381), .A(n20920), .ZN(n20384) );
  AOI22_X1 U23330 ( .A1(n20435), .A2(n20781), .B1(n20774), .B2(n20404), .ZN(
        n20391) );
  INV_X1 U23331 ( .A(n20384), .ZN(n20389) );
  OAI21_X1 U23332 ( .B1(n20698), .B2(n20385), .A(n20779), .ZN(n20386) );
  INV_X1 U23333 ( .A(n20386), .ZN(n20387) );
  OAI21_X1 U23334 ( .B1(n20389), .B2(n20388), .A(n20387), .ZN(n20406) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20738), .ZN(n20390) );
  OAI211_X1 U23336 ( .C1(n20409), .C2(n20664), .A(n20391), .B(n20390), .ZN(
        P1_U3057) );
  AOI22_X1 U23337 ( .A1(n20405), .A2(n20787), .B1(n20786), .B2(n20404), .ZN(
        n20393) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20406), .B1(
        n20435), .B2(n20706), .ZN(n20392) );
  OAI211_X1 U23339 ( .C1(n20409), .C2(n20669), .A(n20393), .B(n20392), .ZN(
        P1_U3058) );
  AOI22_X1 U23340 ( .A1(n20405), .A2(n20744), .B1(n20792), .B2(n20404), .ZN(
        n20395) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20406), .B1(
        n20435), .B2(n20793), .ZN(n20394) );
  OAI211_X1 U23342 ( .C1(n20409), .C2(n20672), .A(n20395), .B(n20394), .ZN(
        P1_U3059) );
  AOI22_X1 U23343 ( .A1(n20435), .A2(n20712), .B1(n20798), .B2(n20404), .ZN(
        n20397) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20799), .ZN(n20396) );
  OAI211_X1 U23345 ( .C1(n20409), .C2(n20675), .A(n20397), .B(n20396), .ZN(
        P1_U3060) );
  AOI22_X1 U23346 ( .A1(n20435), .A2(n20807), .B1(n20805), .B2(n20404), .ZN(
        n20399) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20750), .ZN(n20398) );
  OAI211_X1 U23348 ( .C1(n20409), .C2(n20678), .A(n20399), .B(n20398), .ZN(
        P1_U3061) );
  AOI22_X1 U23349 ( .A1(n20405), .A2(n20754), .B1(n20812), .B2(n20404), .ZN(
        n20401) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20406), .B1(
        n20435), .B2(n20813), .ZN(n20400) );
  OAI211_X1 U23351 ( .C1(n20409), .C2(n20681), .A(n20401), .B(n20400), .ZN(
        P1_U3062) );
  AOI22_X1 U23352 ( .A1(n20405), .A2(n20758), .B1(n20818), .B2(n20404), .ZN(
        n20403) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20406), .B1(
        n20435), .B2(n20819), .ZN(n20402) );
  OAI211_X1 U23354 ( .C1(n20409), .C2(n20687), .A(n20403), .B(n20402), .ZN(
        P1_U3063) );
  AOI22_X1 U23355 ( .A1(n20405), .A2(n20764), .B1(n20824), .B2(n20404), .ZN(
        n20408) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20406), .B1(
        n20435), .B2(n20827), .ZN(n20407) );
  OAI211_X1 U23357 ( .C1(n20409), .C2(n20694), .A(n20408), .B(n20407), .ZN(
        P1_U3064) );
  NAND3_X1 U23358 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20617), .A3(
        n20655), .ZN(n20439) );
  NOR2_X1 U23359 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20439), .ZN(
        n20433) );
  INV_X1 U23360 ( .A(n20654), .ZN(n20730) );
  NOR2_X1 U23361 ( .A1(n13609), .A2(n20411), .ZN(n20495) );
  NAND3_X1 U23362 ( .A1(n20495), .A2(n20698), .A3(n13559), .ZN(n20412) );
  OAI21_X1 U23363 ( .B1(n20730), .B2(n20413), .A(n20412), .ZN(n20434) );
  AOI22_X1 U23364 ( .A1(n20774), .A2(n20433), .B1(n20773), .B2(n20434), .ZN(
        n20420) );
  INV_X1 U23365 ( .A(n20435), .ZN(n20414) );
  AOI21_X1 U23366 ( .B1(n20414), .B2(n20464), .A(n21137), .ZN(n20415) );
  AOI21_X1 U23367 ( .B1(n20495), .B2(n13559), .A(n20415), .ZN(n20416) );
  NOR2_X1 U23368 ( .A1(n20416), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20418) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20738), .ZN(n20419) );
  OAI211_X1 U23370 ( .C1(n20741), .C2(n20464), .A(n20420), .B(n20419), .ZN(
        P1_U3065) );
  AOI22_X1 U23371 ( .A1(n20786), .A2(n20433), .B1(n20785), .B2(n20434), .ZN(
        n20422) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20787), .ZN(n20421) );
  OAI211_X1 U23373 ( .C1(n20790), .C2(n20464), .A(n20422), .B(n20421), .ZN(
        P1_U3066) );
  AOI22_X1 U23374 ( .A1(n20792), .A2(n20433), .B1(n20791), .B2(n20434), .ZN(
        n20424) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20744), .ZN(n20423) );
  OAI211_X1 U23376 ( .C1(n20747), .C2(n20464), .A(n20424), .B(n20423), .ZN(
        P1_U3067) );
  AOI22_X1 U23377 ( .A1(n20798), .A2(n20433), .B1(n20797), .B2(n20434), .ZN(
        n20426) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20799), .ZN(n20425) );
  OAI211_X1 U23379 ( .C1(n20804), .C2(n20464), .A(n20426), .B(n20425), .ZN(
        P1_U3068) );
  AOI22_X1 U23380 ( .A1(n20806), .A2(n20434), .B1(n20805), .B2(n20433), .ZN(
        n20428) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20750), .ZN(n20427) );
  OAI211_X1 U23382 ( .C1(n20753), .C2(n20464), .A(n20428), .B(n20427), .ZN(
        P1_U3069) );
  AOI22_X1 U23383 ( .A1(n20812), .A2(n20433), .B1(n20811), .B2(n20434), .ZN(
        n20430) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20754), .ZN(n20429) );
  OAI211_X1 U23385 ( .C1(n20757), .C2(n20464), .A(n20430), .B(n20429), .ZN(
        P1_U3070) );
  AOI22_X1 U23386 ( .A1(n20818), .A2(n20433), .B1(n20817), .B2(n20434), .ZN(
        n20432) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20758), .ZN(n20431) );
  OAI211_X1 U23388 ( .C1(n20761), .C2(n20464), .A(n20432), .B(n20431), .ZN(
        P1_U3071) );
  AOI22_X1 U23389 ( .A1(n20826), .A2(n20434), .B1(n20824), .B2(n20433), .ZN(
        n20438) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20436), .B1(
        n20435), .B2(n20764), .ZN(n20437) );
  OAI211_X1 U23391 ( .C1(n20769), .C2(n20464), .A(n20438), .B(n20437), .ZN(
        P1_U3072) );
  INV_X1 U23392 ( .A(n20738), .ZN(n20784) );
  NOR2_X1 U23393 ( .A1(n20696), .A2(n20439), .ZN(n20459) );
  AOI21_X1 U23394 ( .B1(n20495), .B2(n20551), .A(n20459), .ZN(n20440) );
  OAI22_X1 U23395 ( .A1(n20440), .A2(n20920), .B1(n20439), .B2(n10577), .ZN(
        n20460) );
  AOI22_X1 U23396 ( .A1(n20774), .A2(n20459), .B1(n20773), .B2(n20460), .ZN(
        n20446) );
  INV_X1 U23397 ( .A(n20439), .ZN(n20443) );
  INV_X1 U23398 ( .A(n20498), .ZN(n20441) );
  OAI21_X1 U23399 ( .B1(n20441), .B2(n20701), .A(n20440), .ZN(n20442) );
  OAI221_X1 U23400 ( .B1(n20698), .B2(n20443), .C1(n20920), .C2(n20442), .A(
        n20779), .ZN(n20461) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20461), .B1(
        n20488), .B2(n20781), .ZN(n20445) );
  OAI211_X1 U23402 ( .C1(n20784), .C2(n20464), .A(n20446), .B(n20445), .ZN(
        P1_U3073) );
  AOI22_X1 U23403 ( .A1(n20786), .A2(n20459), .B1(n20785), .B2(n20460), .ZN(
        n20448) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20461), .B1(
        n20488), .B2(n20706), .ZN(n20447) );
  OAI211_X1 U23405 ( .C1(n20709), .C2(n20464), .A(n20448), .B(n20447), .ZN(
        P1_U3074) );
  AOI22_X1 U23406 ( .A1(n20792), .A2(n20459), .B1(n20791), .B2(n20460), .ZN(
        n20450) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20461), .B1(
        n20488), .B2(n20793), .ZN(n20449) );
  OAI211_X1 U23408 ( .C1(n20796), .C2(n20464), .A(n20450), .B(n20449), .ZN(
        P1_U3075) );
  AOI22_X1 U23409 ( .A1(n20798), .A2(n20459), .B1(n20797), .B2(n20460), .ZN(
        n20452) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20461), .B1(
        n20488), .B2(n20712), .ZN(n20451) );
  OAI211_X1 U23411 ( .C1(n20715), .C2(n20464), .A(n20452), .B(n20451), .ZN(
        P1_U3076) );
  AOI22_X1 U23412 ( .A1(n20806), .A2(n20460), .B1(n20805), .B2(n20459), .ZN(
        n20454) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20461), .B1(
        n20488), .B2(n20807), .ZN(n20453) );
  OAI211_X1 U23414 ( .C1(n20810), .C2(n20464), .A(n20454), .B(n20453), .ZN(
        P1_U3077) );
  AOI22_X1 U23415 ( .A1(n20812), .A2(n20459), .B1(n20811), .B2(n20460), .ZN(
        n20456) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20461), .B1(
        n20488), .B2(n20813), .ZN(n20455) );
  OAI211_X1 U23417 ( .C1(n20816), .C2(n20464), .A(n20456), .B(n20455), .ZN(
        P1_U3078) );
  AOI22_X1 U23418 ( .A1(n20818), .A2(n20459), .B1(n20817), .B2(n20460), .ZN(
        n20458) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20461), .B1(
        n20488), .B2(n20819), .ZN(n20457) );
  OAI211_X1 U23420 ( .C1(n20822), .C2(n20464), .A(n20458), .B(n20457), .ZN(
        P1_U3079) );
  AOI22_X1 U23421 ( .A1(n20826), .A2(n20460), .B1(n20824), .B2(n20459), .ZN(
        n20463) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20461), .B1(
        n20488), .B2(n20827), .ZN(n20462) );
  OAI211_X1 U23423 ( .C1(n20833), .C2(n20464), .A(n20463), .B(n20462), .ZN(
        P1_U3080) );
  INV_X1 U23424 ( .A(n20488), .ZN(n20465) );
  NAND2_X1 U23425 ( .A1(n20465), .A2(n20698), .ZN(n20467) );
  INV_X1 U23426 ( .A(n20728), .ZN(n20466) );
  OAI21_X1 U23427 ( .B1(n20467), .B2(n20516), .A(n20650), .ZN(n20471) );
  AND2_X1 U23428 ( .A1(n20495), .A2(n20731), .ZN(n20468) );
  INV_X1 U23429 ( .A(n20499), .ZN(n20496) );
  NOR2_X1 U23430 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20496), .ZN(
        n20487) );
  AOI22_X1 U23431 ( .A1(n20516), .A2(n20781), .B1(n20487), .B2(n20774), .ZN(
        n20474) );
  INV_X1 U23432 ( .A(n20468), .ZN(n20470) );
  AOI21_X1 U23433 ( .B1(n20471), .B2(n20470), .A(n20469), .ZN(n20472) );
  OAI211_X1 U23434 ( .C1(n20487), .C2(n20661), .A(n20736), .B(n20472), .ZN(
        n20489) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20489), .B1(
        n20488), .B2(n20738), .ZN(n20473) );
  OAI211_X1 U23436 ( .C1(n20492), .C2(n20664), .A(n20474), .B(n20473), .ZN(
        P1_U3081) );
  AOI22_X1 U23437 ( .A1(n20516), .A2(n20706), .B1(n20487), .B2(n20786), .ZN(
        n20476) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20489), .B1(
        n20488), .B2(n20787), .ZN(n20475) );
  OAI211_X1 U23439 ( .C1(n20492), .C2(n20669), .A(n20476), .B(n20475), .ZN(
        P1_U3082) );
  AOI22_X1 U23440 ( .A1(n20516), .A2(n20793), .B1(n20487), .B2(n20792), .ZN(
        n20478) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20489), .B1(
        n20488), .B2(n20744), .ZN(n20477) );
  OAI211_X1 U23442 ( .C1(n20492), .C2(n20672), .A(n20478), .B(n20477), .ZN(
        P1_U3083) );
  AOI22_X1 U23443 ( .A1(n20488), .A2(n20799), .B1(n20798), .B2(n20487), .ZN(
        n20480) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20489), .B1(
        n20516), .B2(n20712), .ZN(n20479) );
  OAI211_X1 U23445 ( .C1(n20492), .C2(n20675), .A(n20480), .B(n20479), .ZN(
        P1_U3084) );
  AOI22_X1 U23446 ( .A1(n20516), .A2(n20807), .B1(n20805), .B2(n20487), .ZN(
        n20482) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20489), .B1(
        n20488), .B2(n20750), .ZN(n20481) );
  OAI211_X1 U23448 ( .C1(n20492), .C2(n20678), .A(n20482), .B(n20481), .ZN(
        P1_U3085) );
  AOI22_X1 U23449 ( .A1(n20488), .A2(n20754), .B1(n20487), .B2(n20812), .ZN(
        n20484) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20489), .B1(
        n20516), .B2(n20813), .ZN(n20483) );
  OAI211_X1 U23451 ( .C1(n20492), .C2(n20681), .A(n20484), .B(n20483), .ZN(
        P1_U3086) );
  AOI22_X1 U23452 ( .A1(n20516), .A2(n20819), .B1(n20487), .B2(n20818), .ZN(
        n20486) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20489), .B1(
        n20488), .B2(n20758), .ZN(n20485) );
  OAI211_X1 U23454 ( .C1(n20492), .C2(n20687), .A(n20486), .B(n20485), .ZN(
        P1_U3087) );
  AOI22_X1 U23455 ( .A1(n20516), .A2(n20827), .B1(n20824), .B2(n20487), .ZN(
        n20491) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20489), .B1(
        n20488), .B2(n20764), .ZN(n20490) );
  OAI211_X1 U23457 ( .C1(n20492), .C2(n20694), .A(n20491), .B(n20490), .ZN(
        P1_U3088) );
  INV_X1 U23458 ( .A(n20626), .ZN(n20493) );
  INV_X1 U23459 ( .A(n20494), .ZN(n20514) );
  AOI21_X1 U23460 ( .B1(n20495), .B2(n20619), .A(n20514), .ZN(n20497) );
  OAI22_X1 U23461 ( .A1(n20497), .A2(n20920), .B1(n10577), .B2(n20496), .ZN(
        n20515) );
  AOI22_X1 U23462 ( .A1(n20774), .A2(n20514), .B1(n20773), .B2(n20515), .ZN(
        n20501) );
  NOR2_X1 U23463 ( .A1(n20623), .A2(n20920), .ZN(n20775) );
  AND2_X1 U23464 ( .A1(n20498), .A2(n20775), .ZN(n20912) );
  OAI21_X1 U23465 ( .B1(n20499), .B2(n20912), .A(n20779), .ZN(n20517) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20738), .ZN(n20500) );
  OAI211_X1 U23467 ( .C1(n20741), .C2(n20526), .A(n20501), .B(n20500), .ZN(
        P1_U3089) );
  AOI22_X1 U23468 ( .A1(n20786), .A2(n20514), .B1(n20785), .B2(n20515), .ZN(
        n20503) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20787), .ZN(n20502) );
  OAI211_X1 U23470 ( .C1(n20790), .C2(n20526), .A(n20503), .B(n20502), .ZN(
        P1_U3090) );
  AOI22_X1 U23471 ( .A1(n20792), .A2(n20514), .B1(n20791), .B2(n20515), .ZN(
        n20505) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20744), .ZN(n20504) );
  OAI211_X1 U23473 ( .C1(n20747), .C2(n20526), .A(n20505), .B(n20504), .ZN(
        P1_U3091) );
  AOI22_X1 U23474 ( .A1(n20798), .A2(n20514), .B1(n20797), .B2(n20515), .ZN(
        n20507) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20799), .ZN(n20506) );
  OAI211_X1 U23476 ( .C1(n20804), .C2(n20526), .A(n20507), .B(n20506), .ZN(
        P1_U3092) );
  AOI22_X1 U23477 ( .A1(n20806), .A2(n20515), .B1(n20805), .B2(n20514), .ZN(
        n20509) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20750), .ZN(n20508) );
  OAI211_X1 U23479 ( .C1(n20753), .C2(n20526), .A(n20509), .B(n20508), .ZN(
        P1_U3093) );
  AOI22_X1 U23480 ( .A1(n20514), .A2(n20812), .B1(n20811), .B2(n20515), .ZN(
        n20511) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20754), .ZN(n20510) );
  OAI211_X1 U23482 ( .C1(n20757), .C2(n20526), .A(n20511), .B(n20510), .ZN(
        P1_U3094) );
  AOI22_X1 U23483 ( .A1(n20514), .A2(n20818), .B1(n20817), .B2(n20515), .ZN(
        n20513) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20758), .ZN(n20512) );
  OAI211_X1 U23485 ( .C1(n20761), .C2(n20526), .A(n20513), .B(n20512), .ZN(
        P1_U3095) );
  AOI22_X1 U23486 ( .A1(n20826), .A2(n20515), .B1(n20824), .B2(n20514), .ZN(
        n20519) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20764), .ZN(n20518) );
  OAI211_X1 U23488 ( .C1(n20769), .C2(n20526), .A(n20519), .B(n20518), .ZN(
        P1_U3096) );
  INV_X1 U23489 ( .A(n9818), .ZN(n20916) );
  INV_X1 U23490 ( .A(n20919), .ZN(n20522) );
  NAND3_X1 U23491 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11143), .A3(
        n20655), .ZN(n20552) );
  NOR2_X1 U23492 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20552), .ZN(
        n20545) );
  AND2_X1 U23493 ( .A1(n20913), .A2(n13609), .ZN(n20620) );
  AOI21_X1 U23494 ( .B1(n20620), .B2(n13559), .A(n20545), .ZN(n20528) );
  INV_X1 U23495 ( .A(n20578), .ZN(n20524) );
  NOR2_X1 U23496 ( .A1(n20524), .A2(n20523), .ZN(n20653) );
  INV_X1 U23497 ( .A(n20653), .ZN(n20657) );
  OAI22_X1 U23498 ( .A1(n20528), .A2(n20920), .B1(n20525), .B2(n20657), .ZN(
        n20546) );
  AOI22_X1 U23499 ( .A1(n20774), .A2(n20545), .B1(n20546), .B2(n20773), .ZN(
        n20532) );
  INV_X1 U23500 ( .A(n20575), .ZN(n20527) );
  OAI21_X1 U23501 ( .B1(n20527), .B2(n20547), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20529) );
  NAND2_X1 U23502 ( .A1(n20529), .A2(n20528), .ZN(n20530) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20738), .ZN(n20531) );
  OAI211_X1 U23504 ( .C1(n20741), .C2(n20575), .A(n20532), .B(n20531), .ZN(
        P1_U3097) );
  AOI22_X1 U23505 ( .A1(n20786), .A2(n20545), .B1(n20785), .B2(n20546), .ZN(
        n20534) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20787), .ZN(n20533) );
  OAI211_X1 U23507 ( .C1(n20790), .C2(n20575), .A(n20534), .B(n20533), .ZN(
        P1_U3098) );
  AOI22_X1 U23508 ( .A1(n20792), .A2(n20545), .B1(n20791), .B2(n20546), .ZN(
        n20536) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20744), .ZN(n20535) );
  OAI211_X1 U23510 ( .C1(n20747), .C2(n20575), .A(n20536), .B(n20535), .ZN(
        P1_U3099) );
  AOI22_X1 U23511 ( .A1(n20798), .A2(n20545), .B1(n20797), .B2(n20546), .ZN(
        n20538) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20799), .ZN(n20537) );
  OAI211_X1 U23513 ( .C1(n20804), .C2(n20575), .A(n20538), .B(n20537), .ZN(
        P1_U3100) );
  AOI22_X1 U23514 ( .A1(n20806), .A2(n20546), .B1(n20805), .B2(n20545), .ZN(
        n20540) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20750), .ZN(n20539) );
  OAI211_X1 U23516 ( .C1(n20753), .C2(n20575), .A(n20540), .B(n20539), .ZN(
        P1_U3101) );
  AOI22_X1 U23517 ( .A1(n20812), .A2(n20545), .B1(n20811), .B2(n20546), .ZN(
        n20542) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20754), .ZN(n20541) );
  OAI211_X1 U23519 ( .C1(n20757), .C2(n20575), .A(n20542), .B(n20541), .ZN(
        P1_U3102) );
  AOI22_X1 U23520 ( .A1(n20818), .A2(n20545), .B1(n20817), .B2(n20546), .ZN(
        n20544) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20758), .ZN(n20543) );
  OAI211_X1 U23522 ( .C1(n20761), .C2(n20575), .A(n20544), .B(n20543), .ZN(
        P1_U3103) );
  AOI22_X1 U23523 ( .A1(n20826), .A2(n20546), .B1(n20824), .B2(n20545), .ZN(
        n20550) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20764), .ZN(n20549) );
  OAI211_X1 U23525 ( .C1(n20769), .C2(n20575), .A(n20550), .B(n20549), .ZN(
        P1_U3104) );
  NOR2_X1 U23526 ( .A1(n20696), .A2(n20552), .ZN(n20570) );
  AOI21_X1 U23527 ( .B1(n20620), .B2(n20551), .A(n20570), .ZN(n20553) );
  OAI22_X1 U23528 ( .A1(n20553), .A2(n20920), .B1(n20552), .B2(n10577), .ZN(
        n20571) );
  AOI22_X1 U23529 ( .A1(n20774), .A2(n20570), .B1(n20571), .B2(n20773), .ZN(
        n20557) );
  INV_X1 U23530 ( .A(n20552), .ZN(n20555) );
  OAI21_X1 U23531 ( .B1(n20919), .B2(n20701), .A(n20553), .ZN(n20554) );
  OAI221_X1 U23532 ( .B1(n20698), .B2(n20555), .C1(n20920), .C2(n20554), .A(
        n20779), .ZN(n20572) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20572), .B1(
        n20612), .B2(n20781), .ZN(n20556) );
  OAI211_X1 U23534 ( .C1(n20784), .C2(n20575), .A(n20557), .B(n20556), .ZN(
        P1_U3105) );
  AOI22_X1 U23535 ( .A1(n20786), .A2(n20570), .B1(n20785), .B2(n20571), .ZN(
        n20559) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20572), .B1(
        n20612), .B2(n20706), .ZN(n20558) );
  OAI211_X1 U23537 ( .C1(n20709), .C2(n20575), .A(n20559), .B(n20558), .ZN(
        P1_U3106) );
  AOI22_X1 U23538 ( .A1(n20792), .A2(n20570), .B1(n20791), .B2(n20571), .ZN(
        n20561) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20572), .B1(
        n20612), .B2(n20793), .ZN(n20560) );
  OAI211_X1 U23540 ( .C1(n20796), .C2(n20575), .A(n20561), .B(n20560), .ZN(
        P1_U3107) );
  AOI22_X1 U23541 ( .A1(n20798), .A2(n20570), .B1(n20797), .B2(n20571), .ZN(
        n20563) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20572), .B1(
        n20612), .B2(n20712), .ZN(n20562) );
  OAI211_X1 U23543 ( .C1(n20715), .C2(n20575), .A(n20563), .B(n20562), .ZN(
        P1_U3108) );
  AOI22_X1 U23544 ( .A1(n20806), .A2(n20571), .B1(n20805), .B2(n20570), .ZN(
        n20565) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20572), .B1(
        n20612), .B2(n20807), .ZN(n20564) );
  OAI211_X1 U23546 ( .C1(n20810), .C2(n20575), .A(n20565), .B(n20564), .ZN(
        P1_U3109) );
  AOI22_X1 U23547 ( .A1(n20812), .A2(n20570), .B1(n20811), .B2(n20571), .ZN(
        n20567) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20572), .B1(
        n20612), .B2(n20813), .ZN(n20566) );
  OAI211_X1 U23549 ( .C1(n20816), .C2(n20575), .A(n20567), .B(n20566), .ZN(
        P1_U3110) );
  AOI22_X1 U23550 ( .A1(n20818), .A2(n20570), .B1(n20817), .B2(n20571), .ZN(
        n20569) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20572), .B1(
        n20612), .B2(n20819), .ZN(n20568) );
  OAI211_X1 U23552 ( .C1(n20822), .C2(n20575), .A(n20569), .B(n20568), .ZN(
        P1_U3111) );
  AOI22_X1 U23553 ( .A1(n20826), .A2(n20571), .B1(n20824), .B2(n20570), .ZN(
        n20574) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20572), .B1(
        n20612), .B2(n20827), .ZN(n20573) );
  OAI211_X1 U23555 ( .C1(n20833), .C2(n20575), .A(n20574), .B(n20573), .ZN(
        P1_U3112) );
  NAND3_X1 U23556 ( .A1(n20646), .A2(n20576), .A3(n20698), .ZN(n20577) );
  NAND2_X1 U23557 ( .A1(n20577), .A2(n20650), .ZN(n20587) );
  AND2_X1 U23558 ( .A1(n20620), .A2(n20731), .ZN(n20583) );
  OR2_X1 U23559 ( .A1(n20578), .A2(n20617), .ZN(n20729) );
  INV_X1 U23560 ( .A(n20729), .ZN(n20579) );
  INV_X1 U23561 ( .A(n20774), .ZN(n20581) );
  NAND3_X1 U23562 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n11143), .ZN(n20621) );
  NOR2_X1 U23563 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20621), .ZN(
        n20602) );
  INV_X1 U23564 ( .A(n20602), .ZN(n20609) );
  OAI22_X1 U23565 ( .A1(n20646), .A2(n20741), .B1(n20581), .B2(n20609), .ZN(
        n20582) );
  INV_X1 U23566 ( .A(n20582), .ZN(n20590) );
  INV_X1 U23567 ( .A(n20583), .ZN(n20586) );
  NAND2_X1 U23568 ( .A1(n20729), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20735) );
  OAI211_X1 U23569 ( .C1(n20661), .C2(n20602), .A(n20735), .B(n20584), .ZN(
        n20585) );
  AOI21_X1 U23570 ( .B1(n20587), .B2(n20586), .A(n20585), .ZN(n20588) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20738), .ZN(n20589) );
  OAI211_X1 U23572 ( .C1(n20616), .C2(n20664), .A(n20590), .B(n20589), .ZN(
        P1_U3113) );
  OAI22_X1 U23573 ( .A1(n20646), .A2(n20790), .B1(n20665), .B2(n20609), .ZN(
        n20591) );
  INV_X1 U23574 ( .A(n20591), .ZN(n20593) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20787), .ZN(n20592) );
  OAI211_X1 U23576 ( .C1(n20616), .C2(n20669), .A(n20593), .B(n20592), .ZN(
        P1_U3114) );
  AOI22_X1 U23577 ( .A1(n20612), .A2(n20744), .B1(n20792), .B2(n20602), .ZN(
        n20595) );
  INV_X1 U23578 ( .A(n20646), .ZN(n20603) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20613), .B1(
        n20603), .B2(n20793), .ZN(n20594) );
  OAI211_X1 U23580 ( .C1(n20616), .C2(n20672), .A(n20595), .B(n20594), .ZN(
        P1_U3115) );
  OAI22_X1 U23581 ( .A1(n20646), .A2(n20804), .B1(n20596), .B2(n20609), .ZN(
        n20597) );
  INV_X1 U23582 ( .A(n20597), .ZN(n20599) );
  AOI22_X1 U23583 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20799), .ZN(n20598) );
  OAI211_X1 U23584 ( .C1(n20616), .C2(n20675), .A(n20599), .B(n20598), .ZN(
        P1_U3116) );
  AOI22_X1 U23585 ( .A1(n20612), .A2(n20750), .B1(n20805), .B2(n20602), .ZN(
        n20601) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20613), .B1(
        n20603), .B2(n20807), .ZN(n20600) );
  OAI211_X1 U23587 ( .C1(n20616), .C2(n20678), .A(n20601), .B(n20600), .ZN(
        P1_U3117) );
  AOI22_X1 U23588 ( .A1(n20603), .A2(n20813), .B1(n20812), .B2(n20602), .ZN(
        n20605) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20754), .ZN(n20604) );
  OAI211_X1 U23590 ( .C1(n20616), .C2(n20681), .A(n20605), .B(n20604), .ZN(
        P1_U3118) );
  OAI22_X1 U23591 ( .A1(n20646), .A2(n20761), .B1(n20683), .B2(n20609), .ZN(
        n20606) );
  INV_X1 U23592 ( .A(n20606), .ZN(n20608) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20758), .ZN(n20607) );
  OAI211_X1 U23594 ( .C1(n20616), .C2(n20687), .A(n20608), .B(n20607), .ZN(
        P1_U3119) );
  OAI22_X1 U23595 ( .A1(n20646), .A2(n20769), .B1(n20610), .B2(n20609), .ZN(
        n20611) );
  INV_X1 U23596 ( .A(n20611), .ZN(n20615) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20764), .ZN(n20614) );
  OAI211_X1 U23598 ( .C1(n20616), .C2(n20694), .A(n20615), .B(n20614), .ZN(
        P1_U3120) );
  NOR2_X1 U23599 ( .A1(n20618), .A2(n20617), .ZN(n20641) );
  AOI21_X1 U23600 ( .B1(n20620), .B2(n20619), .A(n20641), .ZN(n20622) );
  OAI22_X1 U23601 ( .A1(n20622), .A2(n20920), .B1(n20621), .B2(n10577), .ZN(
        n20642) );
  AOI22_X1 U23602 ( .A1(n20774), .A2(n20641), .B1(n20642), .B2(n20773), .ZN(
        n20628) );
  INV_X1 U23603 ( .A(n20621), .ZN(n20625) );
  OAI21_X1 U23604 ( .B1(n20919), .B2(n20623), .A(n20622), .ZN(n20624) );
  OAI221_X1 U23605 ( .B1(n20698), .B2(n20625), .C1(n20920), .C2(n20624), .A(
        n20779), .ZN(n20643) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20643), .B1(
        n20690), .B2(n20781), .ZN(n20627) );
  OAI211_X1 U23607 ( .C1(n20784), .C2(n20646), .A(n20628), .B(n20627), .ZN(
        P1_U3121) );
  AOI22_X1 U23608 ( .A1(n20786), .A2(n20641), .B1(n20785), .B2(n20642), .ZN(
        n20630) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20643), .B1(
        n20690), .B2(n20706), .ZN(n20629) );
  OAI211_X1 U23610 ( .C1(n20709), .C2(n20646), .A(n20630), .B(n20629), .ZN(
        P1_U3122) );
  AOI22_X1 U23611 ( .A1(n20792), .A2(n20641), .B1(n20791), .B2(n20642), .ZN(
        n20632) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20643), .B1(
        n20690), .B2(n20793), .ZN(n20631) );
  OAI211_X1 U23613 ( .C1(n20796), .C2(n20646), .A(n20632), .B(n20631), .ZN(
        P1_U3123) );
  AOI22_X1 U23614 ( .A1(n20798), .A2(n20641), .B1(n20797), .B2(n20642), .ZN(
        n20634) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20643), .B1(
        n20690), .B2(n20712), .ZN(n20633) );
  OAI211_X1 U23616 ( .C1(n20715), .C2(n20646), .A(n20634), .B(n20633), .ZN(
        P1_U3124) );
  AOI22_X1 U23617 ( .A1(n20806), .A2(n20642), .B1(n20805), .B2(n20641), .ZN(
        n20636) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20643), .B1(
        n20690), .B2(n20807), .ZN(n20635) );
  OAI211_X1 U23619 ( .C1(n20810), .C2(n20646), .A(n20636), .B(n20635), .ZN(
        P1_U3125) );
  AOI22_X1 U23620 ( .A1(n20812), .A2(n20641), .B1(n20811), .B2(n20642), .ZN(
        n20638) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20643), .B1(
        n20690), .B2(n20813), .ZN(n20637) );
  OAI211_X1 U23622 ( .C1(n20816), .C2(n20646), .A(n20638), .B(n20637), .ZN(
        P1_U3126) );
  AOI22_X1 U23623 ( .A1(n20818), .A2(n20641), .B1(n20817), .B2(n20642), .ZN(
        n20640) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20643), .B1(
        n20690), .B2(n20819), .ZN(n20639) );
  OAI211_X1 U23625 ( .C1(n20822), .C2(n20646), .A(n20640), .B(n20639), .ZN(
        P1_U3127) );
  AOI22_X1 U23626 ( .A1(n20826), .A2(n20642), .B1(n20824), .B2(n20641), .ZN(
        n20645) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20643), .B1(
        n20690), .B2(n20827), .ZN(n20644) );
  OAI211_X1 U23628 ( .C1(n20833), .C2(n20646), .A(n20645), .B(n20644), .ZN(
        P1_U3128) );
  INV_X1 U23629 ( .A(n20647), .ZN(n20648) );
  NAND3_X1 U23630 ( .A1(n20649), .A2(n20698), .A3(n20727), .ZN(n20651) );
  NAND2_X1 U23631 ( .A1(n20651), .A2(n20650), .ZN(n20659) );
  OR2_X1 U23632 ( .A1(n13609), .A2(n20652), .ZN(n20697) );
  NOR2_X1 U23633 ( .A1(n20697), .A2(n20731), .ZN(n20656) );
  AOI22_X1 U23634 ( .A1(n20659), .A2(n20656), .B1(n20654), .B2(n20653), .ZN(
        n20695) );
  NAND3_X1 U23635 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20655), .ZN(n20700) );
  NOR2_X1 U23636 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20700), .ZN(
        n20688) );
  AOI22_X1 U23637 ( .A1(n20689), .A2(n20781), .B1(n20774), .B2(n20688), .ZN(
        n20663) );
  INV_X1 U23638 ( .A(n20656), .ZN(n20658) );
  AOI22_X1 U23639 ( .A1(n20659), .A2(n20658), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20657), .ZN(n20660) );
  OAI211_X1 U23640 ( .C1(n20688), .C2(n20661), .A(n20736), .B(n20660), .ZN(
        n20691) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20738), .ZN(n20662) );
  OAI211_X1 U23642 ( .C1(n20695), .C2(n20664), .A(n20663), .B(n20662), .ZN(
        P1_U3129) );
  INV_X1 U23643 ( .A(n20688), .ZN(n20682) );
  OAI22_X1 U23644 ( .A1(n20727), .A2(n20790), .B1(n20665), .B2(n20682), .ZN(
        n20666) );
  INV_X1 U23645 ( .A(n20666), .ZN(n20668) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20787), .ZN(n20667) );
  OAI211_X1 U23647 ( .C1(n20695), .C2(n20669), .A(n20668), .B(n20667), .ZN(
        P1_U3130) );
  AOI22_X1 U23648 ( .A1(n20689), .A2(n20793), .B1(n20792), .B2(n20688), .ZN(
        n20671) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20744), .ZN(n20670) );
  OAI211_X1 U23650 ( .C1(n20695), .C2(n20672), .A(n20671), .B(n20670), .ZN(
        P1_U3131) );
  AOI22_X1 U23651 ( .A1(n20689), .A2(n20712), .B1(n20798), .B2(n20688), .ZN(
        n20674) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20799), .ZN(n20673) );
  OAI211_X1 U23653 ( .C1(n20695), .C2(n20675), .A(n20674), .B(n20673), .ZN(
        P1_U3132) );
  AOI22_X1 U23654 ( .A1(n20689), .A2(n20807), .B1(n20805), .B2(n20688), .ZN(
        n20677) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20750), .ZN(n20676) );
  OAI211_X1 U23656 ( .C1(n20695), .C2(n20678), .A(n20677), .B(n20676), .ZN(
        P1_U3133) );
  AOI22_X1 U23657 ( .A1(n20689), .A2(n20813), .B1(n20812), .B2(n20688), .ZN(
        n20680) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20754), .ZN(n20679) );
  OAI211_X1 U23659 ( .C1(n20695), .C2(n20681), .A(n20680), .B(n20679), .ZN(
        P1_U3134) );
  OAI22_X1 U23660 ( .A1(n20727), .A2(n20761), .B1(n20683), .B2(n20682), .ZN(
        n20684) );
  INV_X1 U23661 ( .A(n20684), .ZN(n20686) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20758), .ZN(n20685) );
  OAI211_X1 U23663 ( .C1(n20695), .C2(n20687), .A(n20686), .B(n20685), .ZN(
        P1_U3135) );
  AOI22_X1 U23664 ( .A1(n20689), .A2(n20827), .B1(n20824), .B2(n20688), .ZN(
        n20693) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20691), .B1(
        n20690), .B2(n20764), .ZN(n20692) );
  OAI211_X1 U23666 ( .C1(n20695), .C2(n20694), .A(n20693), .B(n20692), .ZN(
        P1_U3136) );
  NOR2_X1 U23667 ( .A1(n20696), .A2(n20700), .ZN(n20722) );
  INV_X1 U23668 ( .A(n20722), .ZN(n20699) );
  INV_X1 U23669 ( .A(n20697), .ZN(n20732) );
  NAND2_X1 U23670 ( .A1(n20732), .A2(n20698), .ZN(n20772) );
  OAI222_X1 U23671 ( .A1(n20699), .A2(n20920), .B1(n10577), .B2(n20700), .C1(
        n20312), .C2(n20772), .ZN(n20723) );
  AOI22_X1 U23672 ( .A1(n20774), .A2(n20722), .B1(n20723), .B2(n20773), .ZN(
        n20705) );
  INV_X1 U23673 ( .A(n20700), .ZN(n20702) );
  NOR3_X1 U23674 ( .A1(n20777), .A2(n20920), .A3(n20701), .ZN(n20911) );
  OAI21_X1 U23675 ( .B1(n20702), .B2(n20911), .A(n20779), .ZN(n20724) );
  AOI22_X1 U23676 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20724), .B1(
        n20765), .B2(n20781), .ZN(n20704) );
  OAI211_X1 U23677 ( .C1(n20784), .C2(n20727), .A(n20705), .B(n20704), .ZN(
        P1_U3137) );
  AOI22_X1 U23678 ( .A1(n20786), .A2(n20722), .B1(n20785), .B2(n20723), .ZN(
        n20708) );
  AOI22_X1 U23679 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20724), .B1(
        n20765), .B2(n20706), .ZN(n20707) );
  OAI211_X1 U23680 ( .C1(n20709), .C2(n20727), .A(n20708), .B(n20707), .ZN(
        P1_U3138) );
  AOI22_X1 U23681 ( .A1(n20792), .A2(n20722), .B1(n20791), .B2(n20723), .ZN(
        n20711) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20724), .B1(
        n20765), .B2(n20793), .ZN(n20710) );
  OAI211_X1 U23683 ( .C1(n20796), .C2(n20727), .A(n20711), .B(n20710), .ZN(
        P1_U3139) );
  AOI22_X1 U23684 ( .A1(n20798), .A2(n20722), .B1(n20797), .B2(n20723), .ZN(
        n20714) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20724), .B1(
        n20765), .B2(n20712), .ZN(n20713) );
  OAI211_X1 U23686 ( .C1(n20715), .C2(n20727), .A(n20714), .B(n20713), .ZN(
        P1_U3140) );
  AOI22_X1 U23687 ( .A1(n20806), .A2(n20723), .B1(n20805), .B2(n20722), .ZN(
        n20717) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20724), .B1(
        n20765), .B2(n20807), .ZN(n20716) );
  OAI211_X1 U23689 ( .C1(n20810), .C2(n20727), .A(n20717), .B(n20716), .ZN(
        P1_U3141) );
  AOI22_X1 U23690 ( .A1(n20812), .A2(n20722), .B1(n20811), .B2(n20723), .ZN(
        n20719) );
  AOI22_X1 U23691 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20724), .B1(
        n20765), .B2(n20813), .ZN(n20718) );
  OAI211_X1 U23692 ( .C1(n20816), .C2(n20727), .A(n20719), .B(n20718), .ZN(
        P1_U3142) );
  AOI22_X1 U23693 ( .A1(n20818), .A2(n20722), .B1(n20817), .B2(n20723), .ZN(
        n20721) );
  AOI22_X1 U23694 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20724), .B1(
        n20765), .B2(n20819), .ZN(n20720) );
  OAI211_X1 U23695 ( .C1(n20822), .C2(n20727), .A(n20721), .B(n20720), .ZN(
        P1_U3143) );
  AOI22_X1 U23696 ( .A1(n20826), .A2(n20723), .B1(n20824), .B2(n20722), .ZN(
        n20726) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20724), .B1(
        n20765), .B2(n20827), .ZN(n20725) );
  OAI211_X1 U23698 ( .C1(n20833), .C2(n20727), .A(n20726), .B(n20725), .ZN(
        P1_U3144) );
  NOR2_X1 U23699 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20776), .ZN(
        n20762) );
  OAI22_X1 U23700 ( .A1(n20772), .A2(n13559), .B1(n20730), .B2(n20729), .ZN(
        n20763) );
  AOI22_X1 U23701 ( .A1(n20774), .A2(n20762), .B1(n20773), .B2(n20763), .ZN(
        n20740) );
  INV_X1 U23702 ( .A(n20832), .ZN(n20800) );
  OAI21_X1 U23703 ( .B1(n20765), .B2(n20800), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20734) );
  NAND2_X1 U23704 ( .A1(n20732), .A2(n20731), .ZN(n20733) );
  AOI21_X1 U23705 ( .B1(n20734), .B2(n20733), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20737) );
  AOI22_X1 U23706 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20766), .B1(
        n20765), .B2(n20738), .ZN(n20739) );
  OAI211_X1 U23707 ( .C1(n20741), .C2(n20832), .A(n20740), .B(n20739), .ZN(
        P1_U3145) );
  AOI22_X1 U23708 ( .A1(n20786), .A2(n20762), .B1(n20785), .B2(n20763), .ZN(
        n20743) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20766), .B1(
        n20765), .B2(n20787), .ZN(n20742) );
  OAI211_X1 U23710 ( .C1(n20790), .C2(n20832), .A(n20743), .B(n20742), .ZN(
        P1_U3146) );
  AOI22_X1 U23711 ( .A1(n20792), .A2(n20762), .B1(n20791), .B2(n20763), .ZN(
        n20746) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20766), .B1(
        n20765), .B2(n20744), .ZN(n20745) );
  OAI211_X1 U23713 ( .C1(n20747), .C2(n20832), .A(n20746), .B(n20745), .ZN(
        P1_U3147) );
  AOI22_X1 U23714 ( .A1(n20798), .A2(n20762), .B1(n20797), .B2(n20763), .ZN(
        n20749) );
  AOI22_X1 U23715 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20766), .B1(
        n20765), .B2(n20799), .ZN(n20748) );
  OAI211_X1 U23716 ( .C1(n20804), .C2(n20832), .A(n20749), .B(n20748), .ZN(
        P1_U3148) );
  AOI22_X1 U23717 ( .A1(n20806), .A2(n20763), .B1(n20805), .B2(n20762), .ZN(
        n20752) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20766), .B1(
        n20765), .B2(n20750), .ZN(n20751) );
  OAI211_X1 U23719 ( .C1(n20753), .C2(n20832), .A(n20752), .B(n20751), .ZN(
        P1_U3149) );
  AOI22_X1 U23720 ( .A1(n20812), .A2(n20762), .B1(n20811), .B2(n20763), .ZN(
        n20756) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20766), .B1(
        n20765), .B2(n20754), .ZN(n20755) );
  OAI211_X1 U23722 ( .C1(n20757), .C2(n20832), .A(n20756), .B(n20755), .ZN(
        P1_U3150) );
  AOI22_X1 U23723 ( .A1(n20818), .A2(n20762), .B1(n20817), .B2(n20763), .ZN(
        n20760) );
  AOI22_X1 U23724 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20766), .B1(
        n20765), .B2(n20758), .ZN(n20759) );
  OAI211_X1 U23725 ( .C1(n20761), .C2(n20832), .A(n20760), .B(n20759), .ZN(
        P1_U3151) );
  AOI22_X1 U23726 ( .A1(n20826), .A2(n20763), .B1(n20824), .B2(n20762), .ZN(
        n20768) );
  AOI22_X1 U23727 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20766), .B1(
        n20765), .B2(n20764), .ZN(n20767) );
  OAI211_X1 U23728 ( .C1(n20769), .C2(n20832), .A(n20768), .B(n20767), .ZN(
        P1_U3152) );
  INV_X1 U23729 ( .A(n20770), .ZN(n20823) );
  OAI222_X1 U23730 ( .A1(n20772), .A2(n20771), .B1(n10577), .B2(n20776), .C1(
        n20920), .C2(n20770), .ZN(n20825) );
  AOI22_X1 U23731 ( .A1(n20774), .A2(n20823), .B1(n20773), .B2(n20825), .ZN(
        n20783) );
  INV_X1 U23732 ( .A(n20775), .ZN(n20778) );
  OAI21_X1 U23733 ( .B1(n20778), .B2(n20777), .A(n20776), .ZN(n20780) );
  NAND2_X1 U23734 ( .A1(n20780), .A2(n20779), .ZN(n20829) );
  AOI22_X1 U23735 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20829), .B1(
        n20828), .B2(n20781), .ZN(n20782) );
  OAI211_X1 U23736 ( .C1(n20784), .C2(n20832), .A(n20783), .B(n20782), .ZN(
        P1_U3153) );
  AOI22_X1 U23737 ( .A1(n20786), .A2(n20823), .B1(n20785), .B2(n20825), .ZN(
        n20789) );
  AOI22_X1 U23738 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20829), .B1(
        n20800), .B2(n20787), .ZN(n20788) );
  OAI211_X1 U23739 ( .C1(n20790), .C2(n20803), .A(n20789), .B(n20788), .ZN(
        P1_U3154) );
  AOI22_X1 U23740 ( .A1(n20792), .A2(n20823), .B1(n20791), .B2(n20825), .ZN(
        n20795) );
  AOI22_X1 U23741 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20829), .B1(
        n20828), .B2(n20793), .ZN(n20794) );
  OAI211_X1 U23742 ( .C1(n20796), .C2(n20832), .A(n20795), .B(n20794), .ZN(
        P1_U3155) );
  AOI22_X1 U23743 ( .A1(n20798), .A2(n20823), .B1(n20797), .B2(n20825), .ZN(
        n20802) );
  AOI22_X1 U23744 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20829), .B1(
        n20800), .B2(n20799), .ZN(n20801) );
  OAI211_X1 U23745 ( .C1(n20804), .C2(n20803), .A(n20802), .B(n20801), .ZN(
        P1_U3156) );
  AOI22_X1 U23746 ( .A1(n20806), .A2(n20825), .B1(n20805), .B2(n20823), .ZN(
        n20809) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20829), .B1(
        n20828), .B2(n20807), .ZN(n20808) );
  OAI211_X1 U23748 ( .C1(n20810), .C2(n20832), .A(n20809), .B(n20808), .ZN(
        P1_U3157) );
  AOI22_X1 U23749 ( .A1(n20823), .A2(n20812), .B1(n20811), .B2(n20825), .ZN(
        n20815) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20829), .B1(
        n20828), .B2(n20813), .ZN(n20814) );
  OAI211_X1 U23751 ( .C1(n20816), .C2(n20832), .A(n20815), .B(n20814), .ZN(
        P1_U3158) );
  AOI22_X1 U23752 ( .A1(n20823), .A2(n20818), .B1(n20817), .B2(n20825), .ZN(
        n20821) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20829), .B1(
        n20828), .B2(n20819), .ZN(n20820) );
  OAI211_X1 U23754 ( .C1(n20822), .C2(n20832), .A(n20821), .B(n20820), .ZN(
        P1_U3159) );
  AOI22_X1 U23755 ( .A1(n20826), .A2(n20825), .B1(n20824), .B2(n20823), .ZN(
        n20831) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20829), .B1(
        n20828), .B2(n20827), .ZN(n20830) );
  OAI211_X1 U23757 ( .C1(n20833), .C2(n20832), .A(n20831), .B(n20830), .ZN(
        P1_U3160) );
  NOR2_X1 U23758 ( .A1(n20936), .A2(n20834), .ZN(n20836) );
  AOI22_X1 U23759 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20836), .B1(n20835), 
        .B2(n10577), .ZN(P1_U3163) );
  AND2_X1 U23760 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20899), .ZN(
        P1_U3164) );
  AND2_X1 U23761 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20899), .ZN(
        P1_U3165) );
  AND2_X1 U23762 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20899), .ZN(
        P1_U3166) );
  AND2_X1 U23763 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20899), .ZN(
        P1_U3167) );
  AND2_X1 U23764 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20899), .ZN(
        P1_U3168) );
  AND2_X1 U23765 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20899), .ZN(
        P1_U3169) );
  AND2_X1 U23766 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20899), .ZN(
        P1_U3170) );
  AND2_X1 U23767 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20899), .ZN(
        P1_U3171) );
  AND2_X1 U23768 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20899), .ZN(
        P1_U3172) );
  AND2_X1 U23769 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20899), .ZN(
        P1_U3173) );
  AND2_X1 U23770 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20899), .ZN(
        P1_U3174) );
  AND2_X1 U23771 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20899), .ZN(
        P1_U3175) );
  AND2_X1 U23772 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20899), .ZN(
        P1_U3176) );
  AND2_X1 U23773 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20899), .ZN(
        P1_U3177) );
  AND2_X1 U23774 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20899), .ZN(
        P1_U3178) );
  AND2_X1 U23775 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20899), .ZN(
        P1_U3179) );
  AND2_X1 U23776 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20899), .ZN(
        P1_U3180) );
  AND2_X1 U23777 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20899), .ZN(
        P1_U3181) );
  AND2_X1 U23778 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20899), .ZN(
        P1_U3182) );
  AND2_X1 U23779 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20899), .ZN(
        P1_U3183) );
  AND2_X1 U23780 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20899), .ZN(
        P1_U3184) );
  AND2_X1 U23781 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20899), .ZN(
        P1_U3185) );
  AND2_X1 U23782 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20899), .ZN(P1_U3186) );
  AND2_X1 U23783 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20899), .ZN(P1_U3187) );
  AND2_X1 U23784 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20899), .ZN(P1_U3188) );
  AND2_X1 U23785 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20899), .ZN(P1_U3189) );
  AND2_X1 U23786 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20899), .ZN(P1_U3190) );
  AND2_X1 U23787 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20899), .ZN(P1_U3191) );
  AND2_X1 U23788 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20899), .ZN(P1_U3192) );
  AND2_X1 U23789 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20899), .ZN(P1_U3193) );
  NOR2_X1 U23790 ( .A1(n20837), .A2(n20843), .ZN(n20847) );
  NOR2_X1 U23791 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20838) );
  OAI22_X1 U23792 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21006), .B1(n20838), 
        .B2(n20842), .ZN(n20839) );
  NOR2_X1 U23793 ( .A1(n20840), .A2(n20839), .ZN(n20841) );
  OAI22_X1 U23794 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20847), .B1(n20890), 
        .B2(n20841), .ZN(P1_U3194) );
  AOI21_X1 U23795 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20852), .A(n20842), .ZN(n20844) );
  OAI221_X1 U23796 ( .B1(n20844), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20844), .C2(n20843), .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20851) );
  AOI21_X1 U23797 ( .B1(n20846), .B2(n21006), .A(n20845), .ZN(n20850) );
  INV_X1 U23798 ( .A(n20847), .ZN(n20848) );
  OAI211_X1 U23799 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21006), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20848), .ZN(n20849) );
  OAI21_X1 U23800 ( .B1(n20851), .B2(n20850), .A(n20849), .ZN(P1_U3196) );
  NAND2_X1 U23801 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20890), .ZN(n20892) );
  INV_X1 U23802 ( .A(n20892), .ZN(n20866) );
  INV_X1 U23803 ( .A(n20866), .ZN(n20887) );
  INV_X1 U23804 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20853) );
  INV_X1 U23805 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21054) );
  NAND2_X1 U23806 ( .A1(n20890), .A2(n20852), .ZN(n20889) );
  INV_X1 U23807 ( .A(n20889), .ZN(n20864) );
  OAI222_X1 U23808 ( .A1(n20887), .A2(n21275), .B1(n20853), .B2(n20890), .C1(
        n21054), .C2(n20881), .ZN(P1_U3197) );
  INV_X1 U23809 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20854) );
  OAI222_X1 U23810 ( .A1(n20892), .A2(n21054), .B1(n20854), .B2(n20890), .C1(
        n14063), .C2(n20881), .ZN(P1_U3198) );
  OAI222_X1 U23811 ( .A1(n20887), .A2(n14063), .B1(n20855), .B2(n20890), .C1(
        n21299), .C2(n20881), .ZN(P1_U3199) );
  INV_X1 U23812 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20856) );
  OAI222_X1 U23813 ( .A1(n20889), .A2(n21121), .B1(n20856), .B2(n20890), .C1(
        n21299), .C2(n20892), .ZN(P1_U3200) );
  INV_X1 U23814 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20857) );
  OAI222_X1 U23815 ( .A1(n20892), .A2(n21121), .B1(n20857), .B2(n20890), .C1(
        n21255), .C2(n20881), .ZN(P1_U3201) );
  INV_X1 U23816 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20858) );
  OAI222_X1 U23817 ( .A1(n20892), .A2(n21255), .B1(n20858), .B2(n20890), .C1(
        n21261), .C2(n20881), .ZN(P1_U3202) );
  INV_X1 U23818 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20859) );
  OAI222_X1 U23819 ( .A1(n20892), .A2(n21261), .B1(n20859), .B2(n20890), .C1(
        n20860), .C2(n20881), .ZN(P1_U3203) );
  INV_X1 U23820 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20861) );
  OAI222_X1 U23821 ( .A1(n20881), .A2(n14191), .B1(n20861), .B2(n20890), .C1(
        n20860), .C2(n20892), .ZN(P1_U3204) );
  INV_X1 U23822 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21278) );
  INV_X1 U23823 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20862) );
  OAI222_X1 U23824 ( .A1(n20889), .A2(n21278), .B1(n20862), .B2(n20890), .C1(
        n14191), .C2(n20892), .ZN(P1_U3205) );
  INV_X1 U23825 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21143) );
  INV_X1 U23826 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20863) );
  OAI222_X1 U23827 ( .A1(n20881), .A2(n21143), .B1(n20863), .B2(n20890), .C1(
        n21278), .C2(n20887), .ZN(P1_U3206) );
  AOI22_X1 U23828 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20944), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20864), .ZN(n20865) );
  OAI21_X1 U23829 ( .B1(n21143), .B2(n20887), .A(n20865), .ZN(P1_U3207) );
  AOI22_X1 U23830 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20944), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20866), .ZN(n20867) );
  OAI21_X1 U23831 ( .B1(n14773), .B2(n20881), .A(n20867), .ZN(P1_U3208) );
  INV_X1 U23832 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20868) );
  OAI222_X1 U23833 ( .A1(n20889), .A2(n21300), .B1(n20868), .B2(n20890), .C1(
        n14773), .C2(n20887), .ZN(P1_U3209) );
  INV_X1 U23834 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20869) );
  OAI222_X1 U23835 ( .A1(n20889), .A2(n21122), .B1(n20869), .B2(n20890), .C1(
        n21300), .C2(n20887), .ZN(P1_U3210) );
  INV_X1 U23836 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20870) );
  OAI222_X1 U23837 ( .A1(n20892), .A2(n21122), .B1(n20870), .B2(n20890), .C1(
        n21042), .C2(n20881), .ZN(P1_U3211) );
  INV_X1 U23838 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20871) );
  OAI222_X1 U23839 ( .A1(n20892), .A2(n21042), .B1(n20871), .B2(n20890), .C1(
        n14755), .C2(n20881), .ZN(P1_U3212) );
  INV_X1 U23840 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20872) );
  OAI222_X1 U23841 ( .A1(n20889), .A2(n21039), .B1(n20872), .B2(n20890), .C1(
        n14755), .C2(n20887), .ZN(P1_U3213) );
  INV_X1 U23842 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20873) );
  OAI222_X1 U23843 ( .A1(n20892), .A2(n21039), .B1(n20873), .B2(n20890), .C1(
        n21041), .C2(n20881), .ZN(P1_U3214) );
  INV_X1 U23844 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20874) );
  OAI222_X1 U23845 ( .A1(n20889), .A2(n21131), .B1(n20874), .B2(n20890), .C1(
        n21041), .C2(n20887), .ZN(P1_U3215) );
  INV_X1 U23846 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20875) );
  OAI222_X1 U23847 ( .A1(n20892), .A2(n21131), .B1(n20875), .B2(n20890), .C1(
        n21018), .C2(n20889), .ZN(P1_U3216) );
  INV_X1 U23848 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20876) );
  INV_X1 U23849 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21069) );
  OAI222_X1 U23850 ( .A1(n20892), .A2(n21018), .B1(n20876), .B2(n20890), .C1(
        n21069), .C2(n20889), .ZN(P1_U3217) );
  INV_X1 U23851 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20877) );
  INV_X1 U23852 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21243) );
  OAI222_X1 U23853 ( .A1(n20892), .A2(n21069), .B1(n20877), .B2(n20890), .C1(
        n21243), .C2(n20881), .ZN(P1_U3218) );
  INV_X1 U23854 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20878) );
  OAI222_X1 U23855 ( .A1(n20889), .A2(n20879), .B1(n20878), .B2(n20890), .C1(
        n21243), .C2(n20887), .ZN(P1_U3219) );
  INV_X1 U23856 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20880) );
  OAI222_X1 U23857 ( .A1(n20889), .A2(n20883), .B1(n20880), .B2(n20890), .C1(
        n20879), .C2(n20887), .ZN(P1_U3220) );
  INV_X1 U23858 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20882) );
  OAI222_X1 U23859 ( .A1(n20892), .A2(n20883), .B1(n20882), .B2(n20890), .C1(
        n21272), .C2(n20881), .ZN(P1_U3221) );
  INV_X1 U23860 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20884) );
  OAI222_X1 U23861 ( .A1(n20889), .A2(n21103), .B1(n20884), .B2(n20890), .C1(
        n21272), .C2(n20887), .ZN(P1_U3222) );
  INV_X1 U23862 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20885) );
  OAI222_X1 U23863 ( .A1(n20889), .A2(n21268), .B1(n20885), .B2(n20890), .C1(
        n21103), .C2(n20887), .ZN(P1_U3223) );
  INV_X1 U23864 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20886) );
  OAI222_X1 U23865 ( .A1(n20889), .A2(n21044), .B1(n20886), .B2(n20890), .C1(
        n21268), .C2(n20887), .ZN(P1_U3224) );
  INV_X1 U23866 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20888) );
  OAI222_X1 U23867 ( .A1(n20889), .A2(n14626), .B1(n20888), .B2(n20890), .C1(
        n21044), .C2(n20887), .ZN(P1_U3225) );
  INV_X1 U23868 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20891) );
  OAI222_X1 U23869 ( .A1(n20892), .A2(n14626), .B1(n20891), .B2(n20890), .C1(
        n21028), .C2(n20889), .ZN(P1_U3226) );
  INV_X1 U23870 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U23871 ( .A1(n20890), .A2(n21074), .B1(n20893), .B2(n20944), .ZN(
        P1_U3458) );
  INV_X1 U23872 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21161) );
  INV_X1 U23873 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20894) );
  AOI22_X1 U23874 ( .A1(n20890), .A2(n21161), .B1(n20894), .B2(n20944), .ZN(
        P1_U3459) );
  INV_X1 U23875 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20895) );
  AOI22_X1 U23876 ( .A1(n20890), .A2(n20896), .B1(n20895), .B2(n20944), .ZN(
        P1_U3460) );
  INV_X1 U23877 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21102) );
  INV_X1 U23878 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20897) );
  AOI22_X1 U23879 ( .A1(n20890), .A2(n21102), .B1(n20897), .B2(n20944), .ZN(
        P1_U3461) );
  INV_X1 U23880 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20900) );
  INV_X1 U23881 ( .A(n20901), .ZN(n20898) );
  AOI21_X1 U23882 ( .B1(n20900), .B2(n20899), .A(n20898), .ZN(P1_U3464) );
  OAI21_X1 U23883 ( .B1(n20903), .B2(n20902), .A(n20901), .ZN(P1_U3465) );
  AOI22_X1 U23884 ( .A1(n20907), .A2(n20906), .B1(n20905), .B2(n20904), .ZN(
        n20908) );
  INV_X1 U23885 ( .A(n20908), .ZN(n20910) );
  MUX2_X1 U23886 ( .A(n20910), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20909), .Z(P1_U3469) );
  NOR2_X1 U23887 ( .A1(n20912), .A2(n20911), .ZN(n20918) );
  AOI22_X1 U23888 ( .A1(n20916), .A2(n20915), .B1(n20914), .B2(n20913), .ZN(
        n20917) );
  OAI211_X1 U23889 ( .C1(n20920), .C2(n20919), .A(n20918), .B(n20917), .ZN(
        n20921) );
  NAND2_X1 U23890 ( .A1(n20923), .A2(n20921), .ZN(n20922) );
  OAI21_X1 U23891 ( .B1(n20923), .B2(n20617), .A(n20922), .ZN(P1_U3475) );
  AOI21_X1 U23892 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20924) );
  AOI22_X1 U23893 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20924), .B2(n21275), .ZN(n20925) );
  AOI22_X1 U23894 ( .A1(n20926), .A2(n20925), .B1(n21161), .B2(n20928), .ZN(
        P1_U3481) );
  NOR2_X1 U23895 ( .A1(n20928), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20927) );
  AOI22_X1 U23896 ( .A1(n21102), .A2(n20928), .B1(n13727), .B2(n20927), .ZN(
        P1_U3482) );
  AOI22_X1 U23897 ( .A1(n20890), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21130), 
        .B2(n20944), .ZN(P1_U3483) );
  INV_X1 U23898 ( .A(n20929), .ZN(n20930) );
  AOI21_X1 U23899 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20931), .A(n20930), 
        .ZN(n20932) );
  AOI211_X1 U23900 ( .C1(n20934), .C2(n20933), .A(n10577), .B(n20932), .ZN(
        n20937) );
  OAI21_X1 U23901 ( .B1(n20937), .B2(n20936), .A(n20935), .ZN(n20943) );
  AOI211_X1 U23902 ( .C1(n20941), .C2(n20940), .A(n20939), .B(n20938), .ZN(
        n20942) );
  MUX2_X1 U23903 ( .A(n20943), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20942), 
        .Z(P1_U3485) );
  AOI22_X1 U23904 ( .A1(n20890), .A2(n21302), .B1(n21289), .B2(n20944), .ZN(
        P1_U3486) );
  XNOR2_X1 U23905 ( .A(keyinput_g79), .B(n21299), .ZN(n20951) );
  AOI22_X1 U23906 ( .A1(DATAI_10_), .A2(keyinput_g22), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(keyinput_g74), .ZN(n20945) );
  OAI221_X1 U23907 ( .B1(DATAI_10_), .B2(keyinput_g22), .C1(
        P1_REIP_REG_9__SCAN_IN), .C2(keyinput_g74), .A(n20945), .ZN(n20950) );
  AOI22_X1 U23908 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(keyinput_g105), .B1(
        P1_EBX_REG_6__SCAN_IN), .B2(keyinput_g109), .ZN(n20946) );
  OAI221_X1 U23909 ( .B1(P1_EBX_REG_10__SCAN_IN), .B2(keyinput_g105), .C1(
        P1_EBX_REG_6__SCAN_IN), .C2(keyinput_g109), .A(n20946), .ZN(n20949) );
  AOI22_X1 U23910 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(keyinput_g83), .B1(
        DATAI_25_), .B2(keyinput_g7), .ZN(n20947) );
  OAI221_X1 U23911 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(keyinput_g83), .C1(
        DATAI_25_), .C2(keyinput_g7), .A(n20947), .ZN(n20948) );
  NOR4_X1 U23912 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n20979) );
  AOI22_X1 U23913 ( .A1(DATAI_6_), .A2(keyinput_g26), .B1(
        P1_EBX_REG_3__SCAN_IN), .B2(keyinput_g112), .ZN(n20952) );
  OAI221_X1 U23914 ( .B1(DATAI_6_), .B2(keyinput_g26), .C1(
        P1_EBX_REG_3__SCAN_IN), .C2(keyinput_g112), .A(n20952), .ZN(n20959) );
  AOI22_X1 U23915 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g50), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(keyinput_g71), .ZN(n20953) );
  OAI221_X1 U23916 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g50), 
        .C1(P1_REIP_REG_12__SCAN_IN), .C2(keyinput_g71), .A(n20953), .ZN(
        n20958) );
  AOI22_X1 U23917 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g43), 
        .B1(DATAI_15_), .B2(keyinput_g17), .ZN(n20954) );
  OAI221_X1 U23918 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g43), 
        .C1(DATAI_15_), .C2(keyinput_g17), .A(n20954), .ZN(n20957) );
  AOI22_X1 U23919 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_g42), .B1(BS16), 
        .B2(keyinput_g35), .ZN(n20955) );
  OAI221_X1 U23920 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .C1(BS16), 
        .C2(keyinput_g35), .A(n20955), .ZN(n20956) );
  NOR4_X1 U23921 ( .A1(n20959), .A2(n20958), .A3(n20957), .A4(n20956), .ZN(
        n20978) );
  AOI22_X1 U23922 ( .A1(HOLD), .A2(keyinput_g33), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(keyinput_g99), .ZN(n20960) );
  OAI221_X1 U23923 ( .B1(HOLD), .B2(keyinput_g33), .C1(P1_EBX_REG_16__SCAN_IN), 
        .C2(keyinput_g99), .A(n20960), .ZN(n20967) );
  AOI22_X1 U23924 ( .A1(DATAI_17_), .A2(keyinput_g15), .B1(
        P1_EBX_REG_28__SCAN_IN), .B2(keyinput_g87), .ZN(n20961) );
  OAI221_X1 U23925 ( .B1(DATAI_17_), .B2(keyinput_g15), .C1(
        P1_EBX_REG_28__SCAN_IN), .C2(keyinput_g87), .A(n20961), .ZN(n20966) );
  AOI22_X1 U23926 ( .A1(DATAI_26_), .A2(keyinput_g6), .B1(DATAI_13_), .B2(
        keyinput_g19), .ZN(n20962) );
  OAI221_X1 U23927 ( .B1(DATAI_26_), .B2(keyinput_g6), .C1(DATAI_13_), .C2(
        keyinput_g19), .A(n20962), .ZN(n20965) );
  AOI22_X1 U23928 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(keyinput_g68), .B1(
        DATAI_31_), .B2(keyinput_g1), .ZN(n20963) );
  OAI221_X1 U23929 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(keyinput_g68), .C1(
        DATAI_31_), .C2(keyinput_g1), .A(n20963), .ZN(n20964) );
  NOR4_X1 U23930 ( .A1(n20967), .A2(n20966), .A3(n20965), .A4(n20964), .ZN(
        n20977) );
  AOI22_X1 U23931 ( .A1(DATAI_21_), .A2(keyinput_g11), .B1(DATAI_9_), .B2(
        keyinput_g23), .ZN(n20968) );
  OAI221_X1 U23932 ( .B1(DATAI_21_), .B2(keyinput_g11), .C1(DATAI_9_), .C2(
        keyinput_g23), .A(n20968), .ZN(n20975) );
  AOI22_X1 U23933 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_g45), .B1(
        P1_EBX_REG_7__SCAN_IN), .B2(keyinput_g108), .ZN(n20969) );
  OAI221_X1 U23934 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_g45), .C1(
        P1_EBX_REG_7__SCAN_IN), .C2(keyinput_g108), .A(n20969), .ZN(n20974) );
  AOI22_X1 U23935 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_g39), .B1(
        DATAI_22_), .B2(keyinput_g10), .ZN(n20970) );
  OAI221_X1 U23936 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        DATAI_22_), .C2(keyinput_g10), .A(n20970), .ZN(n20973) );
  AOI22_X1 U23937 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g49), .B1(
        P1_EBX_REG_0__SCAN_IN), .B2(keyinput_g115), .ZN(n20971) );
  OAI221_X1 U23938 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g49), 
        .C1(P1_EBX_REG_0__SCAN_IN), .C2(keyinput_g115), .A(n20971), .ZN(n20972) );
  NOR4_X1 U23939 ( .A1(n20975), .A2(n20974), .A3(n20973), .A4(n20972), .ZN(
        n20976) );
  NAND4_X1 U23940 ( .A1(n20979), .A2(n20978), .A3(n20977), .A4(n20976), .ZN(
        n21119) );
  AOI22_X1 U23941 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(keyinput_g122), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_g44), .ZN(n20980) );
  OAI221_X1 U23942 ( .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_g122), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_g44), .A(n20980), .ZN(n20987)
         );
  AOI22_X1 U23943 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_g75), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(keyinput_g103), .ZN(n20981) );
  OAI221_X1 U23944 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_g75), .C1(
        P1_EBX_REG_12__SCAN_IN), .C2(keyinput_g103), .A(n20981), .ZN(n20986)
         );
  AOI22_X1 U23945 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_g55), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_g58), .ZN(n20982) );
  OAI221_X1 U23946 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_g58), .A(n20982), .ZN(n20985)
         );
  AOI22_X1 U23947 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_g59), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(keyinput_g125), .ZN(n20983) );
  OAI221_X1 U23948 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .C1(
        P1_EAX_REG_22__SCAN_IN), .C2(keyinput_g125), .A(n20983), .ZN(n20984)
         );
  NOR4_X1 U23949 ( .A1(n20987), .A2(n20986), .A3(n20985), .A4(n20984), .ZN(
        n21016) );
  AOI22_X1 U23950 ( .A1(DATAI_3_), .A2(keyinput_g29), .B1(DATAI_30_), .B2(
        keyinput_g2), .ZN(n20988) );
  OAI221_X1 U23951 ( .B1(DATAI_3_), .B2(keyinput_g29), .C1(DATAI_30_), .C2(
        keyinput_g2), .A(n20988), .ZN(n20995) );
  AOI22_X1 U23952 ( .A1(DATAI_19_), .A2(keyinput_g13), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(keyinput_g127), .ZN(n20989) );
  OAI221_X1 U23953 ( .B1(DATAI_19_), .B2(keyinput_g13), .C1(
        P1_EAX_REG_20__SCAN_IN), .C2(keyinput_g127), .A(n20989), .ZN(n20994)
         );
  AOI22_X1 U23954 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(keyinput_g94), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(keyinput_g121), .ZN(n20990) );
  OAI221_X1 U23955 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput_g94), .C1(
        P1_EAX_REG_26__SCAN_IN), .C2(keyinput_g121), .A(n20990), .ZN(n20993)
         );
  AOI22_X1 U23956 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_g104), .B1(
        P1_EBX_REG_1__SCAN_IN), .B2(keyinput_g114), .ZN(n20991) );
  OAI221_X1 U23957 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_g104), .C1(
        P1_EBX_REG_1__SCAN_IN), .C2(keyinput_g114), .A(n20991), .ZN(n20992) );
  NOR4_X1 U23958 ( .A1(n20995), .A2(n20994), .A3(n20993), .A4(n20992), .ZN(
        n21015) );
  AOI22_X1 U23959 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_g40), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput_g85), .ZN(n20996) );
  OAI221_X1 U23960 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_g40), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput_g85), .A(n20996), .ZN(n21003) );
  AOI22_X1 U23961 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_g60), .B1(
        P1_EBX_REG_15__SCAN_IN), .B2(keyinput_g100), .ZN(n20997) );
  OAI221_X1 U23962 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .C1(
        P1_EBX_REG_15__SCAN_IN), .C2(keyinput_g100), .A(n20997), .ZN(n21002)
         );
  AOI22_X1 U23963 ( .A1(DATAI_4_), .A2(keyinput_g28), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(keyinput_g126), .ZN(n20998) );
  OAI221_X1 U23964 ( .B1(DATAI_4_), .B2(keyinput_g28), .C1(
        P1_EAX_REG_21__SCAN_IN), .C2(keyinput_g126), .A(n20998), .ZN(n21001)
         );
  AOI22_X1 U23965 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(keyinput_g69), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(keyinput_g116), .ZN(n20999) );
  OAI221_X1 U23966 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(keyinput_g69), .C1(
        P1_EAX_REG_31__SCAN_IN), .C2(keyinput_g116), .A(n20999), .ZN(n21000)
         );
  NOR4_X1 U23967 ( .A1(n21003), .A2(n21002), .A3(n21001), .A4(n21000), .ZN(
        n21014) );
  AOI22_X1 U23968 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(keyinput_g80), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(keyinput_g110), .ZN(n21004) );
  OAI221_X1 U23969 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(keyinput_g80), .C1(
        P1_EBX_REG_5__SCAN_IN), .C2(keyinput_g110), .A(n21004), .ZN(n21012) );
  AOI22_X1 U23970 ( .A1(DATAI_29_), .A2(keyinput_g3), .B1(n21006), .B2(
        keyinput_g34), .ZN(n21005) );
  OAI221_X1 U23971 ( .B1(DATAI_29_), .B2(keyinput_g3), .C1(n21006), .C2(
        keyinput_g34), .A(n21005), .ZN(n21011) );
  AOI22_X1 U23972 ( .A1(n21130), .A2(keyinput_g47), .B1(n21289), .B2(
        keyinput_g41), .ZN(n21007) );
  OAI221_X1 U23973 ( .B1(n21130), .B2(keyinput_g47), .C1(n21289), .C2(
        keyinput_g41), .A(n21007), .ZN(n21010) );
  INV_X1 U23974 ( .A(DATAI_7_), .ZN(n21259) );
  AOI22_X1 U23975 ( .A1(n11076), .A2(keyinput_g119), .B1(keyinput_g25), .B2(
        n21259), .ZN(n21008) );
  OAI221_X1 U23976 ( .B1(n11076), .B2(keyinput_g119), .C1(n21259), .C2(
        keyinput_g25), .A(n21008), .ZN(n21009) );
  NOR4_X1 U23977 ( .A1(n21012), .A2(n21011), .A3(n21010), .A4(n21009), .ZN(
        n21013) );
  NAND4_X1 U23978 ( .A1(n21016), .A2(n21015), .A3(n21014), .A4(n21013), .ZN(
        n21118) );
  AOI22_X1 U23979 ( .A1(n21018), .A2(keyinput_g62), .B1(keyinput_g5), .B2(
        n21169), .ZN(n21017) );
  OAI221_X1 U23980 ( .B1(n21018), .B2(keyinput_g62), .C1(n21169), .C2(
        keyinput_g5), .A(n21017), .ZN(n21026) );
  AOI22_X1 U23981 ( .A1(n21255), .A2(keyinput_g77), .B1(keyinput_g73), .B2(
        n21278), .ZN(n21019) );
  OAI221_X1 U23982 ( .B1(n21255), .B2(keyinput_g77), .C1(n21278), .C2(
        keyinput_g73), .A(n21019), .ZN(n21025) );
  AOI22_X1 U23983 ( .A1(n21021), .A2(keyinput_g9), .B1(n21286), .B2(
        keyinput_g4), .ZN(n21020) );
  OAI221_X1 U23984 ( .B1(n21021), .B2(keyinput_g9), .C1(n21286), .C2(
        keyinput_g4), .A(n21020), .ZN(n21024) );
  AOI22_X1 U23985 ( .A1(n11100), .A2(keyinput_g118), .B1(keyinput_g70), .B2(
        n14773), .ZN(n21022) );
  OAI221_X1 U23986 ( .B1(n11100), .B2(keyinput_g118), .C1(n14773), .C2(
        keyinput_g70), .A(n21022), .ZN(n21023) );
  NOR4_X1 U23987 ( .A1(n21026), .A2(n21025), .A3(n21024), .A4(n21023), .ZN(
        n21067) );
  AOI22_X1 U23988 ( .A1(n21028), .A2(keyinput_g52), .B1(keyinput_g97), .B2(
        n21308), .ZN(n21027) );
  OAI221_X1 U23989 ( .B1(n21028), .B2(keyinput_g52), .C1(n21308), .C2(
        keyinput_g97), .A(n21027), .ZN(n21036) );
  AOI22_X1 U23990 ( .A1(n14626), .A2(keyinput_g53), .B1(n21269), .B2(
        keyinput_g86), .ZN(n21029) );
  OAI221_X1 U23991 ( .B1(n14626), .B2(keyinput_g53), .C1(n21269), .C2(
        keyinput_g86), .A(n21029), .ZN(n21035) );
  INV_X1 U23992 ( .A(READY2), .ZN(n21305) );
  AOI22_X1 U23993 ( .A1(n21287), .A2(keyinput_g93), .B1(keyinput_g37), .B2(
        n21305), .ZN(n21030) );
  OAI221_X1 U23994 ( .B1(n21287), .B2(keyinput_g93), .C1(n21305), .C2(
        keyinput_g37), .A(n21030), .ZN(n21034) );
  AOI22_X1 U23995 ( .A1(n10976), .A2(keyinput_g124), .B1(keyinput_g12), .B2(
        n21032), .ZN(n21031) );
  OAI221_X1 U23996 ( .B1(n10976), .B2(keyinput_g124), .C1(n21032), .C2(
        keyinput_g12), .A(n21031), .ZN(n21033) );
  NOR4_X1 U23997 ( .A1(n21036), .A2(n21035), .A3(n21034), .A4(n21033), .ZN(
        n21066) );
  AOI22_X1 U23998 ( .A1(n21039), .A2(keyinput_g65), .B1(n21038), .B2(
        keyinput_g101), .ZN(n21037) );
  OAI221_X1 U23999 ( .B1(n21039), .B2(keyinput_g65), .C1(n21038), .C2(
        keyinput_g101), .A(n21037), .ZN(n21050) );
  AOI22_X1 U24000 ( .A1(n21042), .A2(keyinput_g67), .B1(keyinput_g64), .B2(
        n21041), .ZN(n21040) );
  OAI221_X1 U24001 ( .B1(n21042), .B2(keyinput_g67), .C1(n21041), .C2(
        keyinput_g64), .A(n21040), .ZN(n21049) );
  INV_X1 U24002 ( .A(DATAI_0_), .ZN(n21045) );
  AOI22_X1 U24003 ( .A1(n21045), .A2(keyinput_g32), .B1(n21044), .B2(
        keyinput_g54), .ZN(n21043) );
  OAI221_X1 U24004 ( .B1(n21045), .B2(keyinput_g32), .C1(n21044), .C2(
        keyinput_g54), .A(n21043), .ZN(n21048) );
  AOI22_X1 U24005 ( .A1(n21302), .A2(keyinput_g0), .B1(n21272), .B2(
        keyinput_g57), .ZN(n21046) );
  OAI221_X1 U24006 ( .B1(n21302), .B2(keyinput_g0), .C1(n21272), .C2(
        keyinput_g57), .A(n21046), .ZN(n21047) );
  NOR4_X1 U24007 ( .A1(n21050), .A2(n21049), .A3(n21048), .A4(n21047), .ZN(
        n21065) );
  AOI22_X1 U24008 ( .A1(n21290), .A2(keyinput_g113), .B1(keyinput_g21), .B2(
        n21052), .ZN(n21051) );
  OAI221_X1 U24009 ( .B1(n21290), .B2(keyinput_g113), .C1(n21052), .C2(
        keyinput_g21), .A(n21051), .ZN(n21063) );
  AOI22_X1 U24010 ( .A1(n21054), .A2(keyinput_g81), .B1(n21307), .B2(
        keyinput_g106), .ZN(n21053) );
  OAI221_X1 U24011 ( .B1(n21054), .B2(keyinput_g81), .C1(n21307), .C2(
        keyinput_g106), .A(n21053), .ZN(n21062) );
  INV_X1 U24012 ( .A(DATAI_5_), .ZN(n21056) );
  AOI22_X1 U24013 ( .A1(n21057), .A2(keyinput_g20), .B1(keyinput_g27), .B2(
        n21056), .ZN(n21055) );
  OAI221_X1 U24014 ( .B1(n21057), .B2(keyinput_g20), .C1(n21056), .C2(
        keyinput_g27), .A(n21055), .ZN(n21061) );
  AOI22_X1 U24015 ( .A1(n21059), .A2(keyinput_g18), .B1(n21293), .B2(
        keyinput_g91), .ZN(n21058) );
  OAI221_X1 U24016 ( .B1(n21059), .B2(keyinput_g18), .C1(n21293), .C2(
        keyinput_g91), .A(n21058), .ZN(n21060) );
  NOR4_X1 U24017 ( .A1(n21063), .A2(n21062), .A3(n21061), .A4(n21060), .ZN(
        n21064) );
  NAND4_X1 U24018 ( .A1(n21067), .A2(n21066), .A3(n21065), .A4(n21064), .ZN(
        n21117) );
  AOI22_X1 U24019 ( .A1(n21143), .A2(keyinput_g72), .B1(keyinput_g61), .B2(
        n21069), .ZN(n21068) );
  OAI221_X1 U24020 ( .B1(n21143), .B2(keyinput_g72), .C1(n21069), .C2(
        keyinput_g61), .A(n21068), .ZN(n21079) );
  INV_X1 U24021 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21071) );
  AOI22_X1 U24022 ( .A1(n21292), .A2(keyinput_g117), .B1(keyinput_g96), .B2(
        n21071), .ZN(n21070) );
  OAI221_X1 U24023 ( .B1(n21292), .B2(keyinput_g117), .C1(n21071), .C2(
        keyinput_g96), .A(n21070), .ZN(n21078) );
  AOI22_X1 U24024 ( .A1(n21074), .A2(keyinput_g51), .B1(n21073), .B2(
        keyinput_g16), .ZN(n21072) );
  OAI221_X1 U24025 ( .B1(n21074), .B2(keyinput_g51), .C1(n21073), .C2(
        keyinput_g16), .A(n21072), .ZN(n21077) );
  AOI22_X1 U24026 ( .A1(n21131), .A2(keyinput_g63), .B1(keyinput_g24), .B2(
        n21172), .ZN(n21075) );
  OAI221_X1 U24027 ( .B1(n21131), .B2(keyinput_g63), .C1(n21172), .C2(
        keyinput_g24), .A(n21075), .ZN(n21076) );
  NOR4_X1 U24028 ( .A1(n21079), .A2(n21078), .A3(n21077), .A4(n21076), .ZN(
        n21115) );
  AOI22_X1 U24029 ( .A1(n21166), .A2(keyinput_g84), .B1(n21138), .B2(
        keyinput_g102), .ZN(n21080) );
  OAI221_X1 U24030 ( .B1(n21166), .B2(keyinput_g84), .C1(n21138), .C2(
        keyinput_g102), .A(n21080), .ZN(n21090) );
  AOI22_X1 U24031 ( .A1(n21082), .A2(keyinput_g95), .B1(keyinput_g98), .B2(
        n14513), .ZN(n21081) );
  OAI221_X1 U24032 ( .B1(n21082), .B2(keyinput_g95), .C1(n14513), .C2(
        keyinput_g98), .A(n21081), .ZN(n21089) );
  INV_X1 U24033 ( .A(DATAI_1_), .ZN(n21163) );
  AOI22_X1 U24034 ( .A1(n21121), .A2(keyinput_g78), .B1(keyinput_g31), .B2(
        n21163), .ZN(n21083) );
  OAI221_X1 U24035 ( .B1(n21121), .B2(keyinput_g78), .C1(n21163), .C2(
        keyinput_g31), .A(n21083), .ZN(n21088) );
  INV_X1 U24036 ( .A(DATAI_2_), .ZN(n21085) );
  AOI22_X1 U24037 ( .A1(n21086), .A2(keyinput_g89), .B1(keyinput_g30), .B2(
        n21085), .ZN(n21084) );
  OAI221_X1 U24038 ( .B1(n21086), .B2(keyinput_g89), .C1(n21085), .C2(
        keyinput_g30), .A(n21084), .ZN(n21087) );
  NOR4_X1 U24039 ( .A1(n21090), .A2(n21089), .A3(n21088), .A4(n21087), .ZN(
        n21114) );
  AOI22_X1 U24040 ( .A1(n21125), .A2(keyinput_g88), .B1(keyinput_g76), .B2(
        n21261), .ZN(n21091) );
  OAI221_X1 U24041 ( .B1(n21125), .B2(keyinput_g88), .C1(n21261), .C2(
        keyinput_g76), .A(n21091), .ZN(n21099) );
  AOI22_X1 U24042 ( .A1(n21275), .A2(keyinput_g82), .B1(n21271), .B2(
        keyinput_g107), .ZN(n21092) );
  OAI221_X1 U24043 ( .B1(n21275), .B2(keyinput_g82), .C1(n21271), .C2(
        keyinput_g107), .A(n21092), .ZN(n21098) );
  INV_X1 U24044 ( .A(READY1), .ZN(n21157) );
  AOI22_X1 U24045 ( .A1(n21151), .A2(keyinput_g46), .B1(n21157), .B2(
        keyinput_g36), .ZN(n21093) );
  OAI221_X1 U24046 ( .B1(n21151), .B2(keyinput_g46), .C1(n21157), .C2(
        keyinput_g36), .A(n21093), .ZN(n21097) );
  AOI22_X1 U24047 ( .A1(n21095), .A2(keyinput_g111), .B1(keyinput_g38), .B2(
        n21256), .ZN(n21094) );
  OAI221_X1 U24048 ( .B1(n21095), .B2(keyinput_g111), .C1(n21256), .C2(
        keyinput_g38), .A(n21094), .ZN(n21096) );
  NOR4_X1 U24049 ( .A1(n21099), .A2(n21098), .A3(n21097), .A4(n21096), .ZN(
        n21113) );
  AOI22_X1 U24050 ( .A1(n21140), .A2(keyinput_g14), .B1(n10995), .B2(
        keyinput_g123), .ZN(n21100) );
  OAI221_X1 U24051 ( .B1(n21140), .B2(keyinput_g14), .C1(n10995), .C2(
        keyinput_g123), .A(n21100), .ZN(n21111) );
  AOI22_X1 U24052 ( .A1(n21103), .A2(keyinput_g56), .B1(keyinput_g48), .B2(
        n21102), .ZN(n21101) );
  OAI221_X1 U24053 ( .B1(n21103), .B2(keyinput_g56), .C1(n21102), .C2(
        keyinput_g48), .A(n21101), .ZN(n21110) );
  AOI22_X1 U24054 ( .A1(n21105), .A2(keyinput_g120), .B1(keyinput_g8), .B2(
        n21262), .ZN(n21104) );
  OAI221_X1 U24055 ( .B1(n21105), .B2(keyinput_g120), .C1(n21262), .C2(
        keyinput_g8), .A(n21104), .ZN(n21109) );
  AOI22_X1 U24056 ( .A1(n14755), .A2(keyinput_g66), .B1(n21107), .B2(
        keyinput_g90), .ZN(n21106) );
  OAI221_X1 U24057 ( .B1(n14755), .B2(keyinput_g66), .C1(n21107), .C2(
        keyinput_g90), .A(n21106), .ZN(n21108) );
  NOR4_X1 U24058 ( .A1(n21111), .A2(n21110), .A3(n21109), .A4(n21108), .ZN(
        n21112) );
  NAND4_X1 U24059 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21116) );
  NOR4_X1 U24060 ( .A1(n21119), .A2(n21118), .A3(n21117), .A4(n21116), .ZN(
        n21329) );
  INV_X1 U24061 ( .A(keyinput_f92), .ZN(n21326) );
  AOI22_X1 U24062 ( .A1(n21122), .A2(keyinput_f68), .B1(n21121), .B2(
        keyinput_f78), .ZN(n21120) );
  OAI221_X1 U24063 ( .B1(n21122), .B2(keyinput_f68), .C1(n21121), .C2(
        keyinput_f78), .A(n21120), .ZN(n21135) );
  INV_X1 U24064 ( .A(keyinput_f48), .ZN(n21124) );
  AOI22_X1 U24065 ( .A1(n21125), .A2(keyinput_f88), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(n21124), .ZN(n21123) );
  OAI221_X1 U24066 ( .B1(n21125), .B2(keyinput_f88), .C1(n21124), .C2(
        P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21123), .ZN(n21134) );
  INV_X1 U24067 ( .A(keyinput_f42), .ZN(n21127) );
  AOI22_X1 U24068 ( .A1(n21128), .A2(keyinput_f2), .B1(P1_D_C_N_REG_SCAN_IN), 
        .B2(n21127), .ZN(n21126) );
  OAI221_X1 U24069 ( .B1(n21128), .B2(keyinput_f2), .C1(n21127), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n21126), .ZN(n21133) );
  AOI22_X1 U24070 ( .A1(n21131), .A2(keyinput_f63), .B1(keyinput_f47), .B2(
        n21130), .ZN(n21129) );
  OAI221_X1 U24071 ( .B1(n21131), .B2(keyinput_f63), .C1(n21130), .C2(
        keyinput_f47), .A(n21129), .ZN(n21132) );
  NOR4_X1 U24072 ( .A1(n21135), .A2(n21134), .A3(n21133), .A4(n21132), .ZN(
        n21324) );
  AOI22_X1 U24073 ( .A1(n21138), .A2(keyinput_f102), .B1(n21137), .B2(
        keyinput_f44), .ZN(n21136) );
  OAI221_X1 U24074 ( .B1(n21138), .B2(keyinput_f102), .C1(n21137), .C2(
        keyinput_f44), .A(n21136), .ZN(n21149) );
  AOI22_X1 U24075 ( .A1(n21141), .A2(keyinput_f115), .B1(keyinput_f14), .B2(
        n21140), .ZN(n21139) );
  OAI221_X1 U24076 ( .B1(n21141), .B2(keyinput_f115), .C1(n21140), .C2(
        keyinput_f14), .A(n21139), .ZN(n21148) );
  AOI22_X1 U24077 ( .A1(n10916), .A2(keyinput_f127), .B1(keyinput_f72), .B2(
        n21143), .ZN(n21142) );
  OAI221_X1 U24078 ( .B1(n10916), .B2(keyinput_f127), .C1(n21143), .C2(
        keyinput_f72), .A(n21142), .ZN(n21147) );
  INV_X1 U24079 ( .A(DATAI_4_), .ZN(n21145) );
  AOI22_X1 U24080 ( .A1(n21145), .A2(keyinput_f28), .B1(keyinput_f17), .B2(
        n14606), .ZN(n21144) );
  OAI221_X1 U24081 ( .B1(n21145), .B2(keyinput_f28), .C1(n14606), .C2(
        keyinput_f17), .A(n21144), .ZN(n21146) );
  NOR4_X1 U24082 ( .A1(n21149), .A2(n21148), .A3(n21147), .A4(n21146), .ZN(
        n21323) );
  AOI22_X1 U24083 ( .A1(n21151), .A2(keyinput_f46), .B1(n11076), .B2(
        keyinput_f119), .ZN(n21150) );
  OAI221_X1 U24084 ( .B1(n21151), .B2(keyinput_f46), .C1(n11076), .C2(
        keyinput_f119), .A(n21150), .ZN(n21180) );
  AOI22_X1 U24085 ( .A1(n21154), .A2(keyinput_f105), .B1(n21153), .B2(
        keyinput_f87), .ZN(n21152) );
  OAI221_X1 U24086 ( .B1(n21154), .B2(keyinput_f105), .C1(n21153), .C2(
        keyinput_f87), .A(n21152), .ZN(n21179) );
  OAI22_X1 U24087 ( .A1(n21157), .A2(keyinput_f36), .B1(n21156), .B2(
        keyinput_f6), .ZN(n21155) );
  AOI221_X1 U24088 ( .B1(n21157), .B2(keyinput_f36), .C1(keyinput_f6), .C2(
        n21156), .A(n21155), .ZN(n21160) );
  XOR2_X1 U24089 ( .A(keyinput_f49), .B(P1_BYTEENABLE_REG_1__SCAN_IN), .Z(
        n21158) );
  AOI21_X1 U24090 ( .B1(keyinput_f50), .B2(n21161), .A(n21158), .ZN(n21159) );
  OAI211_X1 U24091 ( .C1(keyinput_f50), .C2(n21161), .A(n21160), .B(n21159), 
        .ZN(n21178) );
  OAI22_X1 U24092 ( .A1(n21164), .A2(keyinput_f94), .B1(n21163), .B2(
        keyinput_f31), .ZN(n21162) );
  AOI221_X1 U24093 ( .B1(n21164), .B2(keyinput_f94), .C1(keyinput_f31), .C2(
        n21163), .A(n21162), .ZN(n21176) );
  OAI22_X1 U24094 ( .A1(n21167), .A2(keyinput_f126), .B1(n21166), .B2(
        keyinput_f84), .ZN(n21165) );
  AOI221_X1 U24095 ( .B1(n21167), .B2(keyinput_f126), .C1(keyinput_f84), .C2(
        n21166), .A(n21165), .ZN(n21175) );
  OAI22_X1 U24096 ( .A1(n21170), .A2(keyinput_f99), .B1(n21169), .B2(
        keyinput_f5), .ZN(n21168) );
  AOI221_X1 U24097 ( .B1(n21170), .B2(keyinput_f99), .C1(keyinput_f5), .C2(
        n21169), .A(n21168), .ZN(n21174) );
  OAI22_X1 U24098 ( .A1(n14755), .A2(keyinput_f66), .B1(n21172), .B2(
        keyinput_f24), .ZN(n21171) );
  AOI221_X1 U24099 ( .B1(n14755), .B2(keyinput_f66), .C1(keyinput_f24), .C2(
        n21172), .A(n21171), .ZN(n21173) );
  NAND4_X1 U24100 ( .A1(n21176), .A2(n21175), .A3(n21174), .A4(n21173), .ZN(
        n21177) );
  NOR4_X1 U24101 ( .A1(n21180), .A2(n21179), .A3(n21178), .A4(n21177), .ZN(
        n21322) );
  OAI22_X1 U24102 ( .A1(P1_EBX_REG_26__SCAN_IN), .A2(keyinput_f89), .B1(
        keyinput_f109), .B2(P1_EBX_REG_6__SCAN_IN), .ZN(n21181) );
  AOI221_X1 U24103 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(keyinput_f89), .C1(
        P1_EBX_REG_6__SCAN_IN), .C2(keyinput_f109), .A(n21181), .ZN(n21188) );
  OAI22_X1 U24104 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_f123), .B1(
        DATAI_31_), .B2(keyinput_f1), .ZN(n21182) );
  AOI221_X1 U24105 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_f123), .C1(
        keyinput_f1), .C2(DATAI_31_), .A(n21182), .ZN(n21187) );
  OAI22_X1 U24106 ( .A1(P1_EBX_REG_25__SCAN_IN), .A2(keyinput_f90), .B1(
        keyinput_f64), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n21183) );
  AOI221_X1 U24107 ( .B1(P1_EBX_REG_25__SCAN_IN), .B2(keyinput_f90), .C1(
        P1_REIP_REG_19__SCAN_IN), .C2(keyinput_f64), .A(n21183), .ZN(n21186)
         );
  OAI22_X1 U24108 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_f52), .B1(
        DATAI_2_), .B2(keyinput_f30), .ZN(n21184) );
  AOI221_X1 U24109 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .C1(
        keyinput_f30), .C2(DATAI_2_), .A(n21184), .ZN(n21185) );
  NAND4_X1 U24110 ( .A1(n21188), .A2(n21187), .A3(n21186), .A4(n21185), .ZN(
        n21320) );
  OAI22_X1 U24111 ( .A1(DATAI_29_), .A2(keyinput_f3), .B1(keyinput_f29), .B2(
        DATAI_3_), .ZN(n21189) );
  AOI221_X1 U24112 ( .B1(DATAI_29_), .B2(keyinput_f3), .C1(DATAI_3_), .C2(
        keyinput_f29), .A(n21189), .ZN(n21214) );
  OAI22_X1 U24113 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_f67), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_f56), .ZN(n21190) );
  AOI221_X1 U24114 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(keyinput_f67), .C1(
        keyinput_f56), .C2(P1_REIP_REG_27__SCAN_IN), .A(n21190), .ZN(n21193)
         );
  OAI22_X1 U24115 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(
        keyinput_f62), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n21191) );
  AOI221_X1 U24116 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_f62), .A(n21191), .ZN(n21192)
         );
  OAI211_X1 U24117 ( .C1(n11100), .C2(keyinput_f118), .A(n21193), .B(n21192), 
        .ZN(n21194) );
  AOI21_X1 U24118 ( .B1(n11100), .B2(keyinput_f118), .A(n21194), .ZN(n21213)
         );
  AOI22_X1 U24119 ( .A1(DATAI_13_), .A2(keyinput_f19), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_f59), .ZN(n21195) );
  OAI221_X1 U24120 ( .B1(DATAI_13_), .B2(keyinput_f19), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_f59), .A(n21195), .ZN(n21202)
         );
  AOI22_X1 U24121 ( .A1(DATAI_20_), .A2(keyinput_f12), .B1(DATAI_25_), .B2(
        keyinput_f7), .ZN(n21196) );
  OAI221_X1 U24122 ( .B1(DATAI_20_), .B2(keyinput_f12), .C1(DATAI_25_), .C2(
        keyinput_f7), .A(n21196), .ZN(n21201) );
  AOI22_X1 U24123 ( .A1(DATAI_14_), .A2(keyinput_f18), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(keyinput_f71), .ZN(n21197) );
  OAI221_X1 U24124 ( .B1(DATAI_14_), .B2(keyinput_f18), .C1(
        P1_REIP_REG_12__SCAN_IN), .C2(keyinput_f71), .A(n21197), .ZN(n21200)
         );
  AOI22_X1 U24125 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_f65), .B1(
        P1_EBX_REG_1__SCAN_IN), .B2(keyinput_f114), .ZN(n21198) );
  OAI221_X1 U24126 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_f65), .C1(
        P1_EBX_REG_1__SCAN_IN), .C2(keyinput_f114), .A(n21198), .ZN(n21199) );
  NOR4_X1 U24127 ( .A1(n21202), .A2(n21201), .A3(n21200), .A4(n21199), .ZN(
        n21212) );
  AOI22_X1 U24128 ( .A1(DATAI_19_), .A2(keyinput_f13), .B1(DATAI_23_), .B2(
        keyinput_f9), .ZN(n21203) );
  OAI221_X1 U24129 ( .B1(DATAI_19_), .B2(keyinput_f13), .C1(DATAI_23_), .C2(
        keyinput_f9), .A(n21203), .ZN(n21210) );
  AOI22_X1 U24130 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_f75), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(keyinput_f120), .ZN(n21204) );
  OAI221_X1 U24131 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_f75), .C1(
        P1_EAX_REG_27__SCAN_IN), .C2(keyinput_f120), .A(n21204), .ZN(n21209)
         );
  AOI22_X1 U24132 ( .A1(keyinput_f33), .A2(HOLD), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(keyinput_f122), .ZN(n21205) );
  OAI221_X1 U24133 ( .B1(keyinput_f33), .B2(HOLD), .C1(P1_EAX_REG_25__SCAN_IN), 
        .C2(keyinput_f122), .A(n21205), .ZN(n21208) );
  AOI22_X1 U24134 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(keyinput_f83), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput_f85), .ZN(n21206) );
  OAI221_X1 U24135 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(keyinput_f83), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput_f85), .A(n21206), .ZN(n21207) );
  NOR4_X1 U24136 ( .A1(n21210), .A2(n21209), .A3(n21208), .A4(n21207), .ZN(
        n21211) );
  NAND4_X1 U24137 ( .A1(n21214), .A2(n21213), .A3(n21212), .A4(n21211), .ZN(
        n21319) );
  AOI22_X1 U24138 ( .A1(keyinput_f51), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        keyinput_f35), .B2(BS16), .ZN(n21215) );
  OAI221_X1 U24139 ( .B1(keyinput_f51), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), 
        .C1(keyinput_f35), .C2(BS16), .A(n21215), .ZN(n21222) );
  AOI22_X1 U24140 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_f61), .B1(
        P1_EBX_REG_7__SCAN_IN), .B2(keyinput_f108), .ZN(n21216) );
  OAI221_X1 U24141 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .C1(
        P1_EBX_REG_7__SCAN_IN), .C2(keyinput_f108), .A(n21216), .ZN(n21221) );
  AOI22_X1 U24142 ( .A1(DATAI_5_), .A2(keyinput_f27), .B1(DATAI_12_), .B2(
        keyinput_f20), .ZN(n21217) );
  OAI221_X1 U24143 ( .B1(DATAI_5_), .B2(keyinput_f27), .C1(DATAI_12_), .C2(
        keyinput_f20), .A(n21217), .ZN(n21220) );
  AOI22_X1 U24144 ( .A1(DATAI_6_), .A2(keyinput_f26), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_f54), .ZN(n21218) );
  OAI221_X1 U24145 ( .B1(DATAI_6_), .B2(keyinput_f26), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_f54), .A(n21218), .ZN(n21219)
         );
  NOR4_X1 U24146 ( .A1(n21222), .A2(n21221), .A3(n21220), .A4(n21219), .ZN(
        n21251) );
  AOI22_X1 U24147 ( .A1(DATAI_11_), .A2(keyinput_f21), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(keyinput_f81), .ZN(n21223) );
  OAI221_X1 U24148 ( .B1(DATAI_11_), .B2(keyinput_f21), .C1(
        P1_REIP_REG_2__SCAN_IN), .C2(keyinput_f81), .A(n21223), .ZN(n21230) );
  AOI22_X1 U24149 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_f104), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(keyinput_f103), .ZN(n21224) );
  OAI221_X1 U24150 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_f104), .C1(
        P1_EBX_REG_12__SCAN_IN), .C2(keyinput_f103), .A(n21224), .ZN(n21229)
         );
  AOI22_X1 U24151 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(keyinput_f111), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(keyinput_f116), .ZN(n21225) );
  OAI221_X1 U24152 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(keyinput_f111), .C1(
        P1_EAX_REG_31__SCAN_IN), .C2(keyinput_f116), .A(n21225), .ZN(n21228)
         );
  AOI22_X1 U24153 ( .A1(DATAI_22_), .A2(keyinput_f10), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(keyinput_f110), .ZN(n21226) );
  OAI221_X1 U24154 ( .B1(DATAI_22_), .B2(keyinput_f10), .C1(
        P1_EBX_REG_5__SCAN_IN), .C2(keyinput_f110), .A(n21226), .ZN(n21227) );
  NOR4_X1 U24155 ( .A1(n21230), .A2(n21229), .A3(n21228), .A4(n21227), .ZN(
        n21250) );
  AOI22_X1 U24156 ( .A1(keyinput_f34), .A2(NA), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(keyinput_f70), .ZN(n21231) );
  OAI221_X1 U24157 ( .B1(keyinput_f34), .B2(NA), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(keyinput_f70), .A(n21231), .ZN(n21238) );
  AOI22_X1 U24158 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_f45), .B1(DATAI_17_), .B2(keyinput_f15), .ZN(n21232) );
  OAI221_X1 U24159 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_f45), .C1(
        DATAI_17_), .C2(keyinput_f15), .A(n21232), .ZN(n21237) );
  AOI22_X1 U24160 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_f58), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(keyinput_f95), .ZN(n21233) );
  OAI221_X1 U24161 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .C1(
        P1_EBX_REG_20__SCAN_IN), .C2(keyinput_f95), .A(n21233), .ZN(n21236) );
  AOI22_X1 U24162 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_f43), 
        .B1(DATAI_0_), .B2(keyinput_f32), .ZN(n21234) );
  OAI221_X1 U24163 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f43), 
        .C1(DATAI_0_), .C2(keyinput_f32), .A(n21234), .ZN(n21235) );
  NOR4_X1 U24164 ( .A1(n21238), .A2(n21237), .A3(n21236), .A4(n21235), .ZN(
        n21249) );
  AOI22_X1 U24165 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_f53), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(keyinput_f124), .ZN(n21239) );
  OAI221_X1 U24166 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .C1(
        P1_EAX_REG_23__SCAN_IN), .C2(keyinput_f124), .A(n21239), .ZN(n21247)
         );
  AOI22_X1 U24167 ( .A1(DATAI_16_), .A2(keyinput_f16), .B1(
        P1_EBX_REG_19__SCAN_IN), .B2(keyinput_f96), .ZN(n21240) );
  OAI221_X1 U24168 ( .B1(DATAI_16_), .B2(keyinput_f16), .C1(
        P1_EBX_REG_19__SCAN_IN), .C2(keyinput_f96), .A(n21240), .ZN(n21246) );
  AOI22_X1 U24169 ( .A1(keyinput_f39), .A2(P1_ADS_N_REG_SCAN_IN), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(keyinput_f74), .ZN(n21241) );
  OAI221_X1 U24170 ( .B1(keyinput_f39), .B2(P1_ADS_N_REG_SCAN_IN), .C1(
        P1_REIP_REG_9__SCAN_IN), .C2(keyinput_f74), .A(n21241), .ZN(n21245) );
  AOI22_X1 U24171 ( .A1(DATAI_9_), .A2(keyinput_f23), .B1(n21243), .B2(
        keyinput_f60), .ZN(n21242) );
  OAI221_X1 U24172 ( .B1(DATAI_9_), .B2(keyinput_f23), .C1(n21243), .C2(
        keyinput_f60), .A(n21242), .ZN(n21244) );
  NOR4_X1 U24173 ( .A1(n21247), .A2(n21246), .A3(n21245), .A4(n21244), .ZN(
        n21248) );
  NAND4_X1 U24174 ( .A1(n21251), .A2(n21250), .A3(n21249), .A4(n21248), .ZN(
        n21318) );
  AOI22_X1 U24175 ( .A1(n14513), .A2(keyinput_f98), .B1(keyinput_f22), .B2(
        n21253), .ZN(n21252) );
  OAI221_X1 U24176 ( .B1(n14513), .B2(keyinput_f98), .C1(n21253), .C2(
        keyinput_f22), .A(n21252), .ZN(n21266) );
  AOI22_X1 U24177 ( .A1(n21256), .A2(keyinput_f38), .B1(n21255), .B2(
        keyinput_f77), .ZN(n21254) );
  OAI221_X1 U24178 ( .B1(n21256), .B2(keyinput_f38), .C1(n21255), .C2(
        keyinput_f77), .A(n21254), .ZN(n21265) );
  AOI22_X1 U24179 ( .A1(n21259), .A2(keyinput_f25), .B1(n21258), .B2(
        keyinput_f121), .ZN(n21257) );
  OAI221_X1 U24180 ( .B1(n21259), .B2(keyinput_f25), .C1(n21258), .C2(
        keyinput_f121), .A(n21257), .ZN(n21264) );
  AOI22_X1 U24181 ( .A1(n21262), .A2(keyinput_f8), .B1(n21261), .B2(
        keyinput_f76), .ZN(n21260) );
  OAI221_X1 U24182 ( .B1(n21262), .B2(keyinput_f8), .C1(n21261), .C2(
        keyinput_f76), .A(n21260), .ZN(n21263) );
  NOR4_X1 U24183 ( .A1(n21266), .A2(n21265), .A3(n21264), .A4(n21263), .ZN(
        n21316) );
  AOI22_X1 U24184 ( .A1(n21269), .A2(keyinput_f86), .B1(keyinput_f55), .B2(
        n21268), .ZN(n21267) );
  OAI221_X1 U24185 ( .B1(n21269), .B2(keyinput_f86), .C1(n21268), .C2(
        keyinput_f55), .A(n21267), .ZN(n21282) );
  AOI22_X1 U24186 ( .A1(n21272), .A2(keyinput_f57), .B1(n21271), .B2(
        keyinput_f107), .ZN(n21270) );
  OAI221_X1 U24187 ( .B1(n21272), .B2(keyinput_f57), .C1(n21271), .C2(
        keyinput_f107), .A(n21270), .ZN(n21281) );
  AOI22_X1 U24188 ( .A1(n21275), .A2(keyinput_f82), .B1(n21274), .B2(
        keyinput_f125), .ZN(n21273) );
  OAI221_X1 U24189 ( .B1(n21275), .B2(keyinput_f82), .C1(n21274), .C2(
        keyinput_f125), .A(n21273), .ZN(n21280) );
  AOI22_X1 U24190 ( .A1(n21278), .A2(keyinput_f73), .B1(keyinput_f11), .B2(
        n21277), .ZN(n21276) );
  OAI221_X1 U24191 ( .B1(n21278), .B2(keyinput_f73), .C1(n21277), .C2(
        keyinput_f11), .A(n21276), .ZN(n21279) );
  NOR4_X1 U24192 ( .A1(n21282), .A2(n21281), .A3(n21280), .A4(n21279), .ZN(
        n21315) );
  AOI22_X1 U24193 ( .A1(n21284), .A2(keyinput_f112), .B1(keyinput_f80), .B2(
        n14063), .ZN(n21283) );
  OAI221_X1 U24194 ( .B1(n21284), .B2(keyinput_f112), .C1(n14063), .C2(
        keyinput_f80), .A(n21283), .ZN(n21297) );
  AOI22_X1 U24195 ( .A1(n21287), .A2(keyinput_f93), .B1(keyinput_f4), .B2(
        n21286), .ZN(n21285) );
  OAI221_X1 U24196 ( .B1(n21287), .B2(keyinput_f93), .C1(n21286), .C2(
        keyinput_f4), .A(n21285), .ZN(n21296) );
  AOI22_X1 U24197 ( .A1(n21290), .A2(keyinput_f113), .B1(keyinput_f41), .B2(
        n21289), .ZN(n21288) );
  OAI221_X1 U24198 ( .B1(n21290), .B2(keyinput_f113), .C1(n21289), .C2(
        keyinput_f41), .A(n21288), .ZN(n21295) );
  AOI22_X1 U24199 ( .A1(n21293), .A2(keyinput_f91), .B1(n21292), .B2(
        keyinput_f117), .ZN(n21291) );
  OAI221_X1 U24200 ( .B1(n21293), .B2(keyinput_f91), .C1(n21292), .C2(
        keyinput_f117), .A(n21291), .ZN(n21294) );
  NOR4_X1 U24201 ( .A1(n21297), .A2(n21296), .A3(n21295), .A4(n21294), .ZN(
        n21314) );
  AOI22_X1 U24202 ( .A1(n21300), .A2(keyinput_f69), .B1(n21299), .B2(
        keyinput_f79), .ZN(n21298) );
  OAI221_X1 U24203 ( .B1(n21300), .B2(keyinput_f69), .C1(n21299), .C2(
        keyinput_f79), .A(n21298), .ZN(n21312) );
  INV_X1 U24204 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21303) );
  AOI22_X1 U24205 ( .A1(n21303), .A2(keyinput_f40), .B1(keyinput_f0), .B2(
        n21302), .ZN(n21301) );
  OAI221_X1 U24206 ( .B1(n21303), .B2(keyinput_f40), .C1(n21302), .C2(
        keyinput_f0), .A(n21301), .ZN(n21311) );
  AOI22_X1 U24207 ( .A1(n14514), .A2(keyinput_f100), .B1(keyinput_f37), .B2(
        n21305), .ZN(n21304) );
  OAI221_X1 U24208 ( .B1(n14514), .B2(keyinput_f100), .C1(n21305), .C2(
        keyinput_f37), .A(n21304), .ZN(n21310) );
  AOI22_X1 U24209 ( .A1(n21308), .A2(keyinput_f97), .B1(keyinput_f106), .B2(
        n21307), .ZN(n21306) );
  OAI221_X1 U24210 ( .B1(n21308), .B2(keyinput_f97), .C1(n21307), .C2(
        keyinput_f106), .A(n21306), .ZN(n21309) );
  NOR4_X1 U24211 ( .A1(n21312), .A2(n21311), .A3(n21310), .A4(n21309), .ZN(
        n21313) );
  NAND4_X1 U24212 ( .A1(n21316), .A2(n21315), .A3(n21314), .A4(n21313), .ZN(
        n21317) );
  NOR4_X1 U24213 ( .A1(n21320), .A2(n21319), .A3(n21318), .A4(n21317), .ZN(
        n21321) );
  NAND4_X1 U24214 ( .A1(n21324), .A2(n21323), .A3(n21322), .A4(n21321), .ZN(
        n21325) );
  OAI221_X1 U24215 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(keyinput_f92), .C1(
        n21330), .C2(n21326), .A(n21325), .ZN(n21327) );
  OAI21_X1 U24216 ( .B1(n21330), .B2(keyinput_g92), .A(n21327), .ZN(n21328) );
  AOI211_X1 U24217 ( .C1(n21330), .C2(keyinput_g92), .A(n21329), .B(n21328), 
        .ZN(n21332) );
  AOI22_X1 U24218 ( .A1(n16619), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16621), .ZN(n21331) );
  XNOR2_X1 U24219 ( .A(n21332), .B(n21331), .ZN(U355) );
  AND2_X1 U12986 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13612) );
  INV_X1 U11259 ( .A(n20274), .ZN(n12878) );
  NAND2_X1 U12889 ( .A1(n10047), .A2(n12159), .ZN(n10049) );
  INV_X2 U12571 ( .A(n20055), .ZN(n11815) );
  OR2_X1 U11255 ( .A1(n11163), .A2(n11162), .ZN(n11165) );
  AOI21_X1 U11270 ( .B1(n11988), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n11987), .ZN(n11989) );
  CLKBUF_X1 U11313 ( .A(n11068), .Z(n11118) );
  CLKBUF_X1 U11314 ( .A(n10452), .Z(n13680) );
  CLKBUF_X1 U11316 ( .A(n11813), .Z(n11808) );
  NAND2_X1 U11319 ( .A1(n14431), .A2(n12872), .ZN(n14393) );
  CLKBUF_X1 U11341 ( .A(n12672), .Z(n14328) );
  INV_X1 U11367 ( .A(n10155), .ZN(n20266) );
  CLKBUF_X1 U11547 ( .A(n11949), .Z(n11959) );
  INV_X2 U11563 ( .A(n11489), .ZN(n9809) );
  CLKBUF_X1 U11620 ( .A(n18322), .Z(n9803) );
  CLKBUF_X2 U12390 ( .A(n18342), .Z(n9806) );
  NAND3_X1 U12507 ( .A1(n10040), .A2(n10041), .A3(n10043), .ZN(n15480) );
  CLKBUF_X1 U12905 ( .A(n19271), .Z(n19287) );
  CLKBUF_X1 U13115 ( .A(n18815), .Z(n9824) );
  CLKBUF_X1 U15048 ( .A(n17598), .Z(n17606) );
endmodule

