

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453;

  INV_X4 U7246 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OR2_X1 U7247 ( .A1(n14851), .A2(n7136), .ZN(n7131) );
  OAI22_X1 U7248 ( .A1(n12269), .A2(n12268), .B1(n12245), .B2(n10126), .ZN(
        n12639) );
  AOI21_X1 U7249 ( .B1(n10437), .B2(n10436), .A(n10124), .ZN(n12269) );
  OR2_X1 U7250 ( .A1(n8086), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8100) );
  INV_X1 U7251 ( .A(n11287), .ZN(n14994) );
  INV_X2 U7252 ( .A(n12589), .ZN(n10372) );
  INV_X2 U7253 ( .A(n10299), .ZN(n10254) );
  CLKBUF_X1 U7254 ( .A(n8616), .Z(n6910) );
  CLKBUF_X3 U7256 ( .A(n9798), .Z(n6544) );
  BUF_X2 U7257 ( .A(n7755), .Z(n12363) );
  CLKBUF_X2 U7258 ( .A(n6547), .Z(n12360) );
  CLKBUF_X2 U7259 ( .A(n8333), .Z(n8770) );
  NAND2_X1 U7260 ( .A1(n7683), .A2(n8945), .ZN(n8008) );
  XNOR2_X1 U7261 ( .A(n8970), .B(P1_IR_REG_20__SCAN_IN), .ZN(n10681) );
  AND2_X1 U7262 ( .A1(n8967), .A2(n8969), .ZN(n14415) );
  AND2_X1 U7263 ( .A1(n13913), .A2(n13917), .ZN(n8616) );
  INV_X1 U7264 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8519) );
  INV_X1 U7265 ( .A(n9798), .ZN(n9656) );
  OR2_X1 U7266 ( .A1(n6536), .A2(n7612), .ZN(n6535) );
  NAND2_X1 U7267 ( .A1(n13707), .A2(n13710), .ZN(n9881) );
  NAND2_X1 U7268 ( .A1(n8111), .A2(n11208), .ZN(n8109) );
  OAI21_X1 U7269 ( .B1(n8172), .B2(n15388), .A(n6905), .ZN(n6904) );
  NAND2_X1 U7270 ( .A1(n12555), .A2(n12414), .ZN(n12547) );
  AND2_X1 U7271 ( .A1(n15319), .A2(n8126), .ZN(n15308) );
  NAND2_X1 U7272 ( .A1(n8170), .A2(n8169), .ZN(n7683) );
  INV_X1 U7273 ( .A(n13547), .ZN(n10913) );
  INV_X2 U7275 ( .A(n10254), .ZN(n12591) );
  INV_X1 U7276 ( .A(n8983), .ZN(n9266) );
  INV_X1 U7277 ( .A(n10097), .ZN(n10109) );
  INV_X1 U7278 ( .A(n12547), .ZN(n12530) );
  INV_X1 U7279 ( .A(n8008), .ZN(n12370) );
  XNOR2_X1 U7280 ( .A(n6529), .B(n7676), .ZN(n8170) );
  NAND2_X1 U7281 ( .A1(n8746), .A2(n8745), .ZN(n8762) );
  INV_X1 U7282 ( .A(n9767), .ZN(n8359) );
  INV_X1 U7283 ( .A(n10196), .ZN(n10374) );
  INV_X1 U7284 ( .A(n9015), .ZN(n9439) );
  INV_X1 U7285 ( .A(n9417), .ZN(n9014) );
  NAND2_X2 U7286 ( .A1(n9524), .A2(n14545), .ZN(n8983) );
  NAND2_X2 U7287 ( .A1(n10026), .A2(n10180), .ZN(n12589) );
  INV_X1 U7288 ( .A(n11043), .ZN(n11206) );
  INV_X1 U7289 ( .A(n11684), .ZN(n15199) );
  INV_X1 U7290 ( .A(n13668), .ZN(n13815) );
  INV_X2 U7291 ( .A(n11852), .ZN(n13742) );
  OAI21_X2 U7292 ( .B1(n10519), .B2(n8359), .A(n8461), .ZN(n11443) );
  NAND2_X1 U7293 ( .A1(n9246), .A2(n9245), .ZN(n14510) );
  BUF_X1 U7294 ( .A(n11489), .Z(n6543) );
  OR2_X1 U7295 ( .A1(n11825), .A2(n11829), .ZN(n6498) );
  OAI21_X2 U7296 ( .B1(n8007), .B2(n6741), .A(n6739), .ZN(n7441) );
  NAND2_X2 U7297 ( .A1(n10028), .A2(n9479), .ZN(n9960) );
  NAND2_X1 U7298 ( .A1(n8986), .A2(n8985), .ZN(n10028) );
  AND2_X2 U7299 ( .A1(n11766), .A2(n8271), .ZN(n9585) );
  OAI21_X2 U7300 ( .B1(n9881), .B2(n7376), .A(n7374), .ZN(n13676) );
  XNOR2_X1 U7301 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7702) );
  NOR2_X2 U7302 ( .A1(n8059), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8074) );
  NAND2_X2 U7303 ( .A1(n12932), .A2(n8148), .ZN(n12918) );
  OR2_X1 U7304 ( .A1(n6776), .A2(n9686), .ZN(n6773) );
  OAI21_X2 U7305 ( .B1(n9577), .B2(n15388), .A(n9576), .ZN(n12892) );
  XNOR2_X1 U7306 ( .A(n11259), .B(n10913), .ZN(n9905) );
  AOI21_X2 U7307 ( .B1(n14662), .B2(n14601), .A(n14659), .ZN(n15449) );
  NAND2_X2 U7308 ( .A1(n14602), .A2(n14603), .ZN(n14562) );
  XNOR2_X2 U7309 ( .A(n14561), .B(n14560), .ZN(n14602) );
  OR2_X2 U7310 ( .A1(n9324), .A2(n6868), .ZN(n8769) );
  OR2_X2 U7311 ( .A1(n11351), .A2(n11443), .ZN(n11496) );
  BUF_X2 U7312 ( .A(n9742), .Z(n14537) );
  AOI21_X2 U7313 ( .B1(n10065), .B2(n14937), .A(n10064), .ZN(n14444) );
  OAI22_X2 U7314 ( .A1(n14849), .A2(P2_ADDR_REG_12__SCAN_IN), .B1(n6743), .B2(
        n14634), .ZN(n6814) );
  XNOR2_X2 U7315 ( .A(n6744), .B(n7114), .ZN(n14849) );
  NAND2_X2 U7316 ( .A1(n8107), .A2(n8106), .ZN(n12921) );
  XNOR2_X2 U7317 ( .A(n11299), .B(n11033), .ZN(n11034) );
  AND2_X2 U7318 ( .A1(n12726), .A2(n11032), .ZN(n11299) );
  XNOR2_X2 U7319 ( .A(n7362), .B(n7361), .ZN(n14851) );
  OAI21_X2 U7320 ( .B1(n12193), .B2(n9864), .A(n9866), .ZN(n13781) );
  NAND2_X2 U7321 ( .A1(n6844), .A2(n9863), .ZN(n12193) );
  INV_X2 U7322 ( .A(n10681), .ZN(n11764) );
  NAND4_X2 U7323 ( .A1(n8294), .A2(n8295), .A3(n8296), .A4(n8293), .ZN(n13549)
         );
  NOR2_X2 U7324 ( .A1(n14646), .A2(n14645), .ZN(n14647) );
  XNOR2_X2 U7325 ( .A(n12046), .B(n12045), .ZN(n15285) );
  AND2_X2 U7326 ( .A1(n12044), .A2(n12043), .ZN(n12046) );
  OAI22_X2 U7327 ( .A1(n14847), .A2(n6742), .B1(n14846), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n6744) );
  AND2_X2 U7328 ( .A1(n7116), .A2(n7115), .ZN(n14847) );
  OR2_X1 U7329 ( .A1(n13366), .A2(n9580), .ZN(n6525) );
  NAND2_X1 U7330 ( .A1(n6906), .A2(n6903), .ZN(n12905) );
  INV_X1 U7331 ( .A(n10383), .ZN(n6499) );
  CLKBUF_X1 U7332 ( .A(n13968), .Z(n14065) );
  NAND2_X1 U7333 ( .A1(n6528), .A2(n6500), .ZN(n6527) );
  XNOR2_X1 U7334 ( .A(n14638), .B(n14637), .ZN(n6745) );
  INV_X1 U7335 ( .A(n12395), .ZN(n6502) );
  NAND2_X1 U7336 ( .A1(n8562), .A2(n8561), .ZN(n11926) );
  OAI21_X1 U7337 ( .B1(n7801), .B2(n6505), .A(n6515), .ZN(n15306) );
  AOI21_X1 U7338 ( .B1(n12476), .B2(n6524), .A(n6503), .ZN(n6523) );
  NAND2_X1 U7339 ( .A1(n10233), .A2(n6842), .ZN(n11652) );
  NAND2_X1 U7340 ( .A1(n6504), .A2(n14725), .ZN(n6520) );
  NAND2_X1 U7341 ( .A1(n8411), .A2(n8410), .ZN(n15146) );
  NOR2_X2 U7342 ( .A1(n10885), .A2(n10884), .ZN(n10883) );
  NAND2_X1 U7343 ( .A1(n10086), .A2(n10085), .ZN(n10097) );
  OAI21_X1 U7344 ( .B1(n12455), .B2(n6505), .A(n12459), .ZN(n6516) );
  INV_X1 U7345 ( .A(n15322), .ZN(n6505) );
  NAND2_X1 U7346 ( .A1(n12421), .A2(n8109), .ZN(n10087) );
  INV_X1 U7347 ( .A(n14138), .ZN(n8938) );
  INV_X1 U7348 ( .A(n12717), .ZN(n11454) );
  AND2_X1 U7349 ( .A1(n6506), .A2(n8110), .ZN(n12416) );
  INV_X1 U7350 ( .A(n15391), .ZN(n10877) );
  NAND4_X1 U7351 ( .A1(n7693), .A2(n7695), .A3(n7696), .A4(n7694), .ZN(n10839)
         );
  INV_X1 U7352 ( .A(n9799), .ZN(n9798) );
  INV_X1 U7353 ( .A(n11720), .ZN(n11380) );
  CLKBUF_X2 U7354 ( .A(n7729), .Z(n12358) );
  BUF_X1 U7355 ( .A(n7739), .Z(n6547) );
  NAND4_X2 U7356 ( .A1(n8270), .A2(n8269), .A3(n8268), .A4(n8267), .ZN(n13551)
         );
  NAND2_X1 U7357 ( .A1(n8983), .A2(n8945), .ZN(n9118) );
  INV_X1 U7358 ( .A(n14415), .ZN(n14218) );
  CLKBUF_X3 U7359 ( .A(n7683), .Z(n6507) );
  CLKBUF_X2 U7360 ( .A(n8314), .Z(n6545) );
  NOR2_X2 U7361 ( .A1(n13913), .A2(n13917), .ZN(n8314) );
  INV_X2 U7362 ( .A(n12334), .ZN(n8924) );
  NOR2_X1 U7363 ( .A1(n7864), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7881) );
  INV_X2 U7364 ( .A(n8945), .ZN(n9323) );
  AND3_X1 U7365 ( .A1(n8857), .A2(n8518), .A3(n8242), .ZN(n7631) );
  NAND4_X1 U7366 ( .A1(n8220), .A2(n8604), .A3(n8364), .A4(n8363), .ZN(n8237)
         );
  NOR2_X1 U7367 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6831) );
  NAND2_X1 U7368 ( .A1(n7113), .A2(n9803), .ZN(n9833) );
  NAND2_X1 U7369 ( .A1(n6525), .A2(n6886), .ZN(P3_U3454) );
  OR2_X1 U7370 ( .A1(n13366), .A2(n15439), .ZN(n8218) );
  NOR2_X1 U7371 ( .A1(n12905), .A2(n6526), .ZN(n13366) );
  MUX2_X1 U7372 ( .A(n9560), .B(P3_REG1_REG_28__SCAN_IN), .S(n15439), .Z(n9561) );
  NOR2_X1 U7373 ( .A1(n6748), .A2(n6639), .ZN(n6892) );
  OAI21_X1 U7374 ( .B1(n13881), .B2(n15240), .A(n6911), .ZN(n6894) );
  NAND2_X1 U7375 ( .A1(n6846), .A2(n9897), .ZN(n13623) );
  AND2_X1 U7376 ( .A1(n9545), .A2(n9544), .ZN(n12904) );
  NAND2_X1 U7377 ( .A1(n14276), .A2(n14275), .ZN(n14274) );
  XNOR2_X1 U7378 ( .A(n12352), .B(n6757), .ZN(n6508) );
  NAND2_X1 U7379 ( .A1(n9536), .A2(n12399), .ZN(n9563) );
  OR2_X1 U7380 ( .A1(n12568), .A2(n12567), .ZN(n14077) );
  NAND2_X1 U7381 ( .A1(n6534), .A2(n6535), .ZN(n9536) );
  OR2_X1 U7382 ( .A1(n9790), .A2(n9761), .ZN(n9794) );
  NAND2_X1 U7383 ( .A1(n9579), .A2(n9578), .ZN(n12352) );
  AND2_X1 U7384 ( .A1(n12564), .A2(n12563), .ZN(n12566) );
  AND2_X1 U7385 ( .A1(n12909), .A2(n15426), .ZN(n6526) );
  OR2_X1 U7386 ( .A1(n6499), .A2(n10384), .ZN(n12564) );
  OAI21_X1 U7387 ( .B1(n7639), .B2(n8152), .A(n9546), .ZN(n12909) );
  OAI21_X1 U7388 ( .B1(n12912), .B2(n7242), .A(n7238), .ZN(n9547) );
  OAI21_X1 U7389 ( .B1(n8763), .B2(n7527), .A(n8784), .ZN(n7525) );
  AND2_X1 U7390 ( .A1(n12563), .A2(n10380), .ZN(n10383) );
  NAND2_X1 U7391 ( .A1(n8146), .A2(n8145), .ZN(n12946) );
  NOR2_X1 U7392 ( .A1(n13643), .A2(n7373), .ZN(n7372) );
  AND2_X1 U7393 ( .A1(n12915), .A2(n12402), .ZN(n7639) );
  AND2_X1 U7394 ( .A1(n9769), .A2(n9768), .ZN(n13880) );
  NAND2_X1 U7395 ( .A1(n12912), .A2(n8094), .ZN(n12915) );
  NAND2_X1 U7396 ( .A1(n9412), .A2(n9411), .ZN(n14446) );
  CLKBUF_X1 U7397 ( .A(n12995), .Z(n6839) );
  XNOR2_X1 U7398 ( .A(n7360), .B(n6673), .ZN(n14689) );
  NAND2_X1 U7399 ( .A1(n6957), .A2(n6627), .ZN(n8744) );
  NAND2_X1 U7400 ( .A1(n12947), .A2(n12525), .ZN(n12939) );
  OAI21_X1 U7401 ( .B1(n12948), .B2(n6514), .A(n6512), .ZN(n12912) );
  XNOR2_X1 U7402 ( .A(n9426), .B(n9425), .ZN(n12290) );
  NAND2_X1 U7403 ( .A1(n12948), .A2(n7070), .ZN(n12947) );
  NAND2_X1 U7404 ( .A1(n9381), .A2(n9380), .ZN(n14455) );
  AND2_X1 U7405 ( .A1(n8811), .A2(n8810), .ZN(n13668) );
  INV_X1 U7406 ( .A(n6513), .ZN(n6512) );
  AOI21_X1 U7407 ( .B1(n12959), .B2(n12397), .A(n8053), .ZN(n12948) );
  OAI21_X1 U7408 ( .B1(n7070), .B2(n6514), .A(n12938), .ZN(n6513) );
  NAND2_X1 U7409 ( .A1(n8794), .A2(n8793), .ZN(n13682) );
  AND2_X1 U7410 ( .A1(n12527), .A2(n12913), .ZN(n12938) );
  OAI21_X1 U7411 ( .B1(n8827), .B2(n12076), .A(n8826), .ZN(n8829) );
  OAI21_X1 U7412 ( .B1(n8017), .B2(n12516), .A(n6713), .ZN(n12959) );
  XNOR2_X1 U7413 ( .A(n8807), .B(n8806), .ZN(n12175) );
  NAND2_X1 U7414 ( .A1(n12990), .A2(n12506), .ZN(n8017) );
  NAND2_X1 U7415 ( .A1(n9348), .A2(n9347), .ZN(n14314) );
  INV_X1 U7416 ( .A(n12525), .ZN(n6514) );
  NAND2_X1 U7417 ( .A1(n7131), .A2(n7130), .ZN(n14852) );
  AND2_X1 U7418 ( .A1(n8772), .A2(n8771), .ZN(n13891) );
  NAND2_X1 U7419 ( .A1(n8072), .A2(n8071), .ZN(n13375) );
  OAI21_X1 U7420 ( .B1(n13002), .B2(n12996), .A(n6527), .ZN(n12990) );
  NAND2_X1 U7421 ( .A1(n6715), .A2(n12499), .ZN(n13002) );
  XNOR2_X1 U7422 ( .A(n8750), .B(n8749), .ZN(n12070) );
  NAND2_X1 U7423 ( .A1(n6518), .A2(n7222), .ZN(n13288) );
  NAND2_X1 U7424 ( .A1(n6518), .A2(n6517), .ZN(n13286) );
  NAND2_X1 U7425 ( .A1(n6738), .A2(n8069), .ZN(n8081) );
  NAND2_X1 U7426 ( .A1(n6940), .A2(n6939), .ZN(n12317) );
  NAND2_X1 U7427 ( .A1(n12281), .A2(n7224), .ZN(n6518) );
  OAI21_X1 U7428 ( .B1(n6716), .B2(n12408), .A(n6523), .ZN(n12264) );
  NAND2_X1 U7429 ( .A1(n6716), .A2(n7888), .ZN(n12246) );
  NAND2_X1 U7430 ( .A1(n8533), .A2(n11635), .ZN(n11641) );
  INV_X1 U7431 ( .A(n13396), .ZN(n6500) );
  AND2_X1 U7432 ( .A1(n7222), .A2(n12395), .ZN(n6517) );
  NAND2_X1 U7433 ( .A1(n8584), .A2(n8583), .ZN(n12109) );
  NAND2_X1 U7434 ( .A1(n9209), .A2(n9208), .ZN(n14104) );
  OAI21_X1 U7435 ( .B1(n6522), .B2(n6521), .A(n6519), .ZN(n12214) );
  INV_X1 U7436 ( .A(n12086), .ZN(n6501) );
  NAND2_X1 U7437 ( .A1(n6522), .A2(n12469), .ZN(n14724) );
  NAND2_X1 U7438 ( .A1(n15308), .A2(n8127), .ZN(n15307) );
  NAND2_X1 U7439 ( .A1(n15306), .A2(n12463), .ZN(n7838) );
  AOI21_X1 U7440 ( .B1(n7484), .B2(n7477), .A(n7476), .ZN(n7475) );
  NAND2_X1 U7441 ( .A1(n9193), .A2(n9192), .ZN(n14827) );
  NAND2_X1 U7442 ( .A1(n7801), .A2(n12455), .ZN(n15318) );
  NAND2_X1 U7443 ( .A1(n6717), .A2(n12445), .ZN(n11698) );
  NAND2_X1 U7444 ( .A1(n11697), .A2(n12450), .ZN(n15335) );
  NAND2_X1 U7445 ( .A1(n8526), .A2(n8525), .ZN(n11855) );
  AND2_X1 U7446 ( .A1(n6727), .A2(n6726), .ZN(n14668) );
  OAI21_X1 U7447 ( .B1(n11458), .B2(n6511), .A(n6509), .ZN(n11697) );
  NAND2_X1 U7448 ( .A1(n8499), .A2(n8498), .ZN(n11887) );
  INV_X1 U7449 ( .A(n7888), .ZN(n6524) );
  INV_X1 U7450 ( .A(n12412), .ZN(n6503) );
  NAND2_X1 U7451 ( .A1(n11458), .A2(n12385), .ZN(n6717) );
  NAND2_X1 U7452 ( .A1(n8066), .A2(n8065), .ZN(n12960) );
  NAND2_X1 U7453 ( .A1(n9123), .A2(n9122), .ZN(n15022) );
  AND2_X1 U7454 ( .A1(n6520), .A2(n12473), .ZN(n6519) );
  INV_X1 U7455 ( .A(n12615), .ZN(n6528) );
  NAND2_X1 U7456 ( .A1(n9090), .A2(n9089), .ZN(n11878) );
  INV_X1 U7457 ( .A(n14725), .ZN(n6521) );
  NAND2_X1 U7458 ( .A1(n9075), .A2(n9074), .ZN(n15006) );
  NAND2_X1 U7459 ( .A1(n7364), .A2(n14615), .ZN(n14617) );
  INV_X1 U7460 ( .A(n6510), .ZN(n6509) );
  INV_X1 U7461 ( .A(n6516), .ZN(n6515) );
  OAI21_X1 U7462 ( .B1(n12385), .B2(n6511), .A(n12454), .ZN(n6510) );
  NAND2_X1 U7463 ( .A1(n8391), .A2(n8390), .ZN(n11689) );
  INV_X1 U7464 ( .A(n12469), .ZN(n6504) );
  AND2_X1 U7465 ( .A1(n7735), .A2(n12431), .ZN(n8114) );
  NAND2_X1 U7466 ( .A1(n10088), .A2(n8109), .ZN(n15380) );
  AND2_X1 U7467 ( .A1(n10030), .A2(n8994), .ZN(n11324) );
  AOI21_X1 U7468 ( .B1(n7236), .B2(n11035), .A(n7234), .ZN(n7233) );
  INV_X1 U7469 ( .A(n12445), .ZN(n6511) );
  AND2_X1 U7470 ( .A1(n7143), .A2(n7142), .ZN(n14571) );
  NAND2_X1 U7471 ( .A1(n12421), .A2(n12416), .ZN(n10088) );
  AND2_X1 U7472 ( .A1(n12428), .A2(n12427), .ZN(n15379) );
  OR2_X1 U7473 ( .A1(n14612), .A2(n14613), .ZN(n7143) );
  CLKBUF_X1 U7474 ( .A(n8116), .Z(n12719) );
  NAND2_X1 U7475 ( .A1(n6598), .A2(n7741), .ZN(n12718) );
  INV_X1 U7476 ( .A(n8110), .ZN(n12328) );
  NAND4_X1 U7477 ( .A1(n8929), .A2(n8928), .A3(n8927), .A4(n8926), .ZN(n14138)
         );
  NOR2_X1 U7478 ( .A1(n14607), .A2(n14608), .ZN(n14610) );
  NAND2_X2 U7479 ( .A1(n6575), .A2(n8260), .ZN(n15171) );
  NAND4_X1 U7480 ( .A1(n7672), .A2(n7671), .A3(n7670), .A4(n7669), .ZN(n12717)
         );
  AND3_X1 U7481 ( .A1(n7692), .A2(n7691), .A3(n7690), .ZN(n15358) );
  BUF_X4 U7482 ( .A(n9799), .Z(n6542) );
  OR2_X1 U7483 ( .A1(n12724), .A2(n12725), .ZN(n12726) );
  INV_X1 U7484 ( .A(n10839), .ZN(n6506) );
  OAI211_X1 U7485 ( .C1(n7729), .C2(n10450), .A(n7699), .B(n7700), .ZN(n8110)
         );
  NAND2_X1 U7486 ( .A1(n7814), .A2(n7813), .ZN(n7830) );
  AND3_X1 U7487 ( .A1(n7719), .A2(n7718), .A3(n7717), .ZN(n15391) );
  INV_X2 U7488 ( .A(n8000), .ZN(n7981) );
  NAND2_X2 U7489 ( .A1(n11250), .A2(n9586), .ZN(n9799) );
  AND3_X1 U7490 ( .A1(n7734), .A2(n7733), .A3(n7732), .ZN(n15373) );
  CLKBUF_X1 U7491 ( .A(n9417), .Z(n9443) );
  INV_X2 U7492 ( .A(n9118), .ZN(n9466) );
  OAI22_X1 U7493 ( .A1(n7794), .A2(n7793), .B1(P2_DATAO_REG_7__SCAN_IN), .B2(
        n10500), .ZN(n7811) );
  INV_X1 U7494 ( .A(n8008), .ZN(n7746) );
  NAND2_X1 U7495 ( .A1(n14541), .A2(n12334), .ZN(n9017) );
  AND2_X2 U7496 ( .A1(n7663), .A2(n12288), .ZN(n7721) );
  OAI21_X1 U7497 ( .B1(n8303), .B2(n7201), .A(n7198), .ZN(n8331) );
  XNOR2_X1 U7498 ( .A(n9512), .B(n9511), .ZN(n12180) );
  NAND2_X1 U7499 ( .A1(n9520), .A2(n11764), .ZN(n10180) );
  XNOR2_X1 U7500 ( .A(n7246), .B(n11047), .ZN(n11131) );
  INV_X2 U7501 ( .A(n12553), .ZN(n15255) );
  BUF_X2 U7502 ( .A(n8315), .Z(n8369) );
  NAND2_X1 U7503 ( .A1(n8934), .A2(n8933), .ZN(n14545) );
  XNOR2_X1 U7504 ( .A(n7662), .B(P3_IR_REG_29__SCAN_IN), .ZN(n7667) );
  OAI21_X1 U7505 ( .B1(n9513), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9512) );
  AND2_X1 U7506 ( .A1(n9586), .A2(n11820), .ZN(n10766) );
  NOR2_X1 U7507 ( .A1(n13913), .A2(n8266), .ZN(n8315) );
  AOI21_X1 U7508 ( .B1(n8307), .B2(n7200), .A(n7199), .ZN(n7198) );
  MUX2_X1 U7509 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8932), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n8934) );
  NAND2_X1 U7510 ( .A1(n13412), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7662) );
  MUX2_X1 U7511 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8228), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8229) );
  OR2_X1 U7512 ( .A1(n9505), .A2(n8935), .ZN(n7144) );
  NAND2_X1 U7513 ( .A1(n14563), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n7126) );
  INV_X2 U7514 ( .A(n14536), .ZN(n14544) );
  NAND2_X1 U7515 ( .A1(n6777), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U7516 ( .A1(n6530), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6529) );
  XNOR2_X1 U7517 ( .A(n6721), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7663) );
  MUX2_X1 U7518 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7674), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7675) );
  OR2_X1 U7519 ( .A1(n8262), .A2(n6978), .ZN(n6969) );
  NAND2_X1 U7520 ( .A1(n8182), .A2(n6668), .ZN(n6530) );
  NAND2_X2 U7521 ( .A1(n10476), .A2(P2_U3088), .ZN(n13920) );
  OR2_X1 U7522 ( .A1(n8231), .A2(n8519), .ZN(n8226) );
  AOI22_X1 U7523 ( .A1(n11206), .A2(P3_REG2_REG_2__SCAN_IN), .B1(n11006), .B2(
        n11043), .ZN(n11190) );
  NAND2_X2 U7524 ( .A1(n10476), .A2(P3_U3151), .ZN(n13423) );
  AND3_X1 U7525 ( .A1(n8243), .A2(n7631), .A3(n6976), .ZN(n8262) );
  OAI21_X1 U7526 ( .B1(n8247), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n6896), .ZN(
        n7497) );
  AND2_X1 U7527 ( .A1(n6895), .A2(n7857), .ZN(n8182) );
  CLKBUF_X1 U7528 ( .A(n8630), .Z(n8631) );
  AND3_X1 U7529 ( .A1(n6660), .A2(n6820), .A3(n6818), .ZN(n15065) );
  INV_X1 U7530 ( .A(n8237), .ZN(n8243) );
  NOR2_X1 U7531 ( .A1(n7769), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U7532 ( .A1(n6800), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7716) );
  NAND4_X1 U7533 ( .A1(n9200), .A2(n8909), .A3(n8908), .A4(n6831), .ZN(n8912)
         );
  AND2_X2 U7534 ( .A1(n7092), .A2(n7090), .ZN(n8247) );
  NOR2_X1 U7535 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  NAND2_X1 U7536 ( .A1(n8257), .A2(n8256), .ZN(n10553) );
  AND2_X1 U7537 ( .A1(n8248), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7701) );
  AND4_X1 U7538 ( .A1(n8241), .A2(n8240), .A3(n8239), .A4(n8238), .ZN(n8857)
         );
  AND2_X1 U7539 ( .A1(n7660), .A2(n7611), .ZN(n7610) );
  AND2_X1 U7540 ( .A1(n6833), .A2(n6832), .ZN(n9200) );
  AND3_X1 U7541 ( .A1(n8223), .A2(n8222), .A3(n8221), .ZN(n8518) );
  AND2_X1 U7542 ( .A1(n7307), .A2(n7605), .ZN(n7603) );
  NOR2_X1 U7543 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7405) );
  NOR2_X1 U7544 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n8239) );
  XNOR2_X1 U7545 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14596) );
  NOR2_X1 U7546 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8240) );
  NOR2_X1 U7547 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n7406) );
  NOR2_X1 U7548 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8908) );
  NOR2_X1 U7549 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n8909) );
  NOR2_X2 U7550 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8948) );
  INV_X4 U7551 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7552 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6833) );
  INV_X1 U7553 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8238) );
  INV_X1 U7554 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7908) );
  INV_X1 U7555 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7654) );
  INV_X4 U7556 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X2 U7557 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8364) );
  INV_X1 U7558 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7030) );
  INV_X1 U7559 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7358) );
  NOR2_X1 U7560 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7604) );
  INV_X1 U7561 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7686) );
  NOR2_X1 U7562 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7738) );
  AND2_X1 U7563 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7308) );
  NOR2_X1 U7564 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n6531) );
  NOR2_X1 U7565 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n6532) );
  NOR2_X1 U7566 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n6533) );
  NOR2_X1 U7567 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n8363) );
  NOR2_X1 U7568 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n8362) );
  INV_X1 U7569 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7659) );
  NOR2_X1 U7570 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8221) );
  NOR2_X1 U7571 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8222) );
  NOR2_X1 U7572 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n7251) );
  INV_X1 U7573 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7660) );
  NOR2_X1 U7574 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7652) );
  INV_X1 U7575 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7307) );
  AOI21_X1 U7576 ( .B1(n6508), .B2(n15411), .A(n12892), .ZN(n10407) );
  AOI21_X1 U7577 ( .B1(n6508), .B2(n13306), .A(n12895), .ZN(n12896) );
  NAND2_X1 U7578 ( .A1(n14735), .A2(n14737), .ZN(n6522) );
  NAND2_X1 U7579 ( .A1(n12264), .A2(n12482), .ZN(n7920) );
  NAND4_X1 U7580 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n7686), .ZN(n6722)
         );
  NAND2_X1 U7581 ( .A1(n8383), .A2(n8382), .ZN(n8387) );
  NAND2_X1 U7582 ( .A1(n12918), .A2(n6537), .ZN(n6534) );
  INV_X1 U7583 ( .A(n9528), .ZN(n6536) );
  AND2_X1 U7584 ( .A1(n8149), .A2(n9528), .ZN(n6537) );
  NAND2_X1 U7585 ( .A1(n11699), .A2(n6541), .ZN(n6538) );
  AND2_X1 U7586 ( .A1(n6538), .A2(n6539), .ZN(n15319) );
  OR2_X1 U7587 ( .A1(n6540), .A2(n8123), .ZN(n6539) );
  INV_X1 U7588 ( .A(n6566), .ZN(n6540) );
  AND2_X1 U7589 ( .A1(n8122), .A2(n6566), .ZN(n6541) );
  NAND2_X1 U7590 ( .A1(n6718), .A2(n7661), .ZN(n13412) );
  OAI222_X1 U7591 ( .A1(P3_U3151), .A2(n12288), .B1(n13419), .B2(n12287), .C1(
        n12286), .C2(n13423), .ZN(P3_U3266) );
  OAI21_X2 U7592 ( .B1(n9993), .B2(n6795), .A(n6793), .ZN(n14349) );
  XNOR2_X2 U7593 ( .A(n8762), .B(n8760), .ZN(n13432) );
  NAND2_X1 U7594 ( .A1(n6546), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7708) );
  OAI211_X2 U7595 ( .C1(n7117), .C2(n6725), .A(n14559), .B(n6723), .ZN(n14561)
         );
  NAND2_X4 U7596 ( .A1(n9175), .A2(n9174), .ZN(n14820) );
  OAI21_X1 U7597 ( .B1(n7673), .B2(n6719), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n6721) );
  XNOR2_X2 U7598 ( .A(n6732), .B(n6592), .ZN(n14688) );
  NAND2_X2 U7599 ( .A1(n6734), .A2(n6733), .ZN(n6732) );
  AOI21_X2 U7600 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11812), .A(n11798), .ZN(
        n11825) );
  OAI21_X2 U7601 ( .B1(n15266), .B2(n7244), .A(n7243), .ZN(n11798) );
  XNOR2_X2 U7602 ( .A(n7129), .B(n6596), .ZN(n14850) );
  OAI21_X2 U7603 ( .B1(n6745), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n6597), .ZN(
        n7129) );
  OAI22_X1 U7604 ( .A1(n12946), .A2(n8147), .B1(n12655), .B2(n12960), .ZN(
        n12930) );
  INV_X2 U7605 ( .A(n12721), .ZN(n8111) );
  NAND4_X1 U7606 ( .A1(n7705), .A2(n7707), .A3(n7706), .A4(n7708), .ZN(n12721)
         );
  AND2_X1 U7607 ( .A1(n7663), .A2(n12288), .ZN(n6546) );
  NAND2_X1 U7608 ( .A1(n12562), .A2(n7667), .ZN(n7755) );
  NOR2_X1 U7609 ( .A1(n7663), .A2(n7667), .ZN(n7739) );
  NOR2_X1 U7610 ( .A1(n15268), .A2(n11607), .ZN(n11610) );
  NOR2_X1 U7611 ( .A1(n7565), .A2(n6791), .ZN(n6790) );
  INV_X1 U7612 ( .A(n10000), .ZN(n6791) );
  NAND2_X1 U7613 ( .A1(n7521), .A2(n9313), .ZN(n7520) );
  INV_X1 U7614 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U7615 ( .A1(n7295), .A2(n6572), .ZN(n7294) );
  INV_X1 U7616 ( .A(n8142), .ZN(n7608) );
  NAND2_X1 U7617 ( .A1(n12522), .A2(n8052), .ZN(n12519) );
  OR2_X1 U7618 ( .A1(n12979), .A2(n12625), .ZN(n12514) );
  NAND2_X1 U7619 ( .A1(n7351), .A2(n7350), .ZN(n10428) );
  OAI21_X1 U7620 ( .B1(n6551), .B2(n6687), .A(n7353), .ZN(n7350) );
  AND2_X1 U7621 ( .A1(n7354), .A2(n7353), .ZN(n7352) );
  INV_X1 U7622 ( .A(n12360), .ZN(n8167) );
  INV_X1 U7624 ( .A(n7303), .ZN(n7297) );
  NAND2_X1 U7625 ( .A1(n14349), .A2(n9996), .ZN(n9998) );
  INV_X1 U7626 ( .A(n14628), .ZN(n6726) );
  OAI21_X1 U7627 ( .B1(n9592), .B2(n15166), .A(n9587), .ZN(n9595) );
  INV_X1 U7628 ( .A(n9076), .ZN(n7170) );
  AND2_X1 U7629 ( .A1(n6603), .A2(n9237), .ZN(n7166) );
  NOR2_X1 U7630 ( .A1(n7056), .A2(n7055), .ZN(n7054) );
  INV_X1 U7631 ( .A(n14737), .ZN(n7055) );
  INV_X1 U7632 ( .A(n12467), .ZN(n7056) );
  NAND2_X1 U7633 ( .A1(n7150), .A2(n7149), .ZN(n7148) );
  INV_X1 U7634 ( .A(n9326), .ZN(n7149) );
  NAND2_X1 U7635 ( .A1(n7151), .A2(n9327), .ZN(n7150) );
  NAND2_X1 U7636 ( .A1(n7065), .A2(n7069), .ZN(n7064) );
  NAND2_X1 U7637 ( .A1(n12526), .A2(n12938), .ZN(n7069) );
  INV_X1 U7638 ( .A(n12917), .ZN(n7068) );
  INV_X1 U7639 ( .A(n9399), .ZN(n7159) );
  OAI21_X1 U7640 ( .B1(n6758), .B2(n6757), .A(n7080), .ZN(n7079) );
  NAND2_X1 U7641 ( .A1(n12380), .A2(n12546), .ZN(n7080) );
  NAND2_X1 U7642 ( .A1(n8691), .A2(n8690), .ZN(n8710) );
  AOI21_X1 U7643 ( .B1(n8689), .B2(n8688), .A(n8687), .ZN(n8690) );
  NAND2_X1 U7644 ( .A1(n8247), .A2(n10456), .ZN(n6896) );
  NAND2_X1 U7645 ( .A1(n12531), .A2(n12529), .ZN(n12536) );
  INV_X1 U7646 ( .A(n13372), .ZN(n8150) );
  OR2_X1 U7647 ( .A1(n13357), .A2(n13283), .ZN(n12495) );
  NAND2_X1 U7648 ( .A1(n7601), .A2(n13296), .ZN(n7600) );
  OR2_X1 U7649 ( .A1(n13365), .A2(n12712), .ZN(n12484) );
  NOR2_X1 U7650 ( .A1(n7426), .A2(n7421), .ZN(n7420) );
  INV_X1 U7651 ( .A(n7681), .ZN(n7426) );
  INV_X1 U7652 ( .A(n7679), .ZN(n7421) );
  NAND2_X1 U7653 ( .A1(n7397), .A2(n13596), .ZN(n7396) );
  AND2_X1 U7654 ( .A1(n13693), .A2(n9880), .ZN(n7377) );
  NAND2_X1 U7655 ( .A1(n6974), .A2(n8245), .ZN(n6973) );
  NAND2_X1 U7656 ( .A1(n6977), .A2(n6975), .ZN(n6974) );
  NAND2_X1 U7657 ( .A1(n6976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6975) );
  INV_X1 U7658 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8225) );
  OR2_X1 U7659 ( .A1(n14502), .A2(n14010), .ZN(n10052) );
  OR2_X1 U7660 ( .A1(n14104), .A2(n12161), .ZN(n10049) );
  INV_X1 U7661 ( .A(n10047), .ZN(n7553) );
  OR2_X1 U7662 ( .A1(n14136), .A2(n14973), .ZN(n10030) );
  NAND2_X1 U7663 ( .A1(n9428), .A2(n9427), .ZN(n14441) );
  NAND2_X1 U7664 ( .A1(n6792), .A2(n6614), .ZN(n14290) );
  AND2_X1 U7665 ( .A1(n7579), .A2(n7578), .ZN(n7577) );
  INV_X1 U7666 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7578) );
  NAND2_X1 U7667 ( .A1(n7106), .A2(n8789), .ZN(n8807) );
  INV_X1 U7668 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9514) );
  AOI21_X1 U7669 ( .B1(n7515), .B2(n7517), .A(n7513), .ZN(n7512) );
  NOR2_X1 U7670 ( .A1(n7516), .A2(n8597), .ZN(n7515) );
  XNOR2_X1 U7671 ( .A(n8624), .B(SI_16_), .ZN(n8622) );
  INV_X1 U7672 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6832) );
  INV_X1 U7673 ( .A(n8405), .ZN(n7505) );
  INV_X1 U7674 ( .A(n7347), .ZN(n7346) );
  OAI21_X1 U7675 ( .B1(n6591), .B2(n7348), .A(n11552), .ZN(n7347) );
  OAI22_X1 U7676 ( .A1(n10428), .A2(n10122), .B1(n14729), .B2(n10121), .ZN(
        n10437) );
  OR2_X1 U7677 ( .A1(n11191), .A2(n11190), .ZN(n7248) );
  NOR2_X1 U7678 ( .A1(n7299), .A2(n7805), .ZN(n7293) );
  AOI21_X1 U7679 ( .B1(n6498), .B2(n15333), .A(n11828), .ZN(n7231) );
  XNOR2_X1 U7680 ( .A(n12843), .B(n12860), .ZN(n12829) );
  AND2_X1 U7681 ( .A1(n11060), .A2(n11058), .ZN(n11038) );
  NOR2_X1 U7682 ( .A1(n12829), .A2(n12828), .ZN(n12844) );
  OR2_X1 U7683 ( .A1(n12848), .A2(n12847), .ZN(n12871) );
  OR2_X1 U7684 ( .A1(n12900), .A2(n6543), .ZN(n7637) );
  INV_X1 U7685 ( .A(n6714), .ZN(n6713) );
  OAI21_X1 U7686 ( .B1(n12516), .B2(n12507), .A(n12514), .ZN(n6714) );
  NAND2_X1 U7687 ( .A1(n13286), .A2(n7227), .ZN(n6715) );
  NOR2_X1 U7688 ( .A1(n7229), .A2(n7228), .ZN(n7227) );
  INV_X1 U7689 ( .A(n12491), .ZN(n7228) );
  NOR2_X1 U7690 ( .A1(n8129), .A2(n7592), .ZN(n7591) );
  INV_X1 U7691 ( .A(n8128), .ZN(n7592) );
  NAND2_X1 U7692 ( .A1(n11105), .A2(n8117), .ZN(n11229) );
  AND2_X1 U7693 ( .A1(n12530), .A2(n10170), .ZN(n15324) );
  INV_X1 U7694 ( .A(n12555), .ZN(n8210) );
  INV_X1 U7695 ( .A(n10455), .ZN(n6843) );
  AND2_X1 U7696 ( .A1(n13408), .A2(n10414), .ZN(n11219) );
  NAND2_X1 U7697 ( .A1(n7661), .A2(n6720), .ZN(n6719) );
  OAI21_X1 U7698 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(n12259), .A(n8097), .ZN(
        n9530) );
  NAND2_X1 U7699 ( .A1(n7441), .A2(n6692), .ZN(n8055) );
  INV_X1 U7700 ( .A(n8039), .ZN(n8038) );
  OAI21_X1 U7701 ( .B1(n8173), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U7702 ( .A1(n8004), .A2(n8003), .ZN(n8007) );
  NOR2_X1 U7703 ( .A1(n6576), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n7927) );
  OAI21_X1 U7704 ( .B1(n7777), .B2(n7776), .A(n7778), .ZN(n7794) );
  XNOR2_X1 U7705 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7744) );
  XNOR2_X1 U7706 ( .A(n11926), .B(n8834), .ZN(n8574) );
  NAND2_X1 U7707 ( .A1(n6821), .A2(n7396), .ZN(n7395) );
  OR2_X1 U7708 ( .A1(n7397), .A2(n13596), .ZN(n6821) );
  AND2_X1 U7709 ( .A1(n9939), .A2(n9812), .ZN(n13629) );
  AOI21_X1 U7710 ( .B1(n7380), .B2(n7382), .A(n6636), .ZN(n7379) );
  OAI21_X1 U7711 ( .B1(n12191), .B2(n7280), .A(n7278), .ZN(n13755) );
  INV_X1 U7712 ( .A(n7279), .ZN(n7278) );
  OAI21_X1 U7713 ( .B1(n6589), .B2(n7280), .A(n9929), .ZN(n7279) );
  INV_X1 U7714 ( .A(n7285), .ZN(n7284) );
  OAI21_X1 U7715 ( .B1(n9923), .B2(n7286), .A(n9926), .ZN(n7285) );
  NAND2_X1 U7716 ( .A1(n11784), .A2(n6618), .ZN(n11850) );
  XNOR2_X1 U7717 ( .A(n15232), .B(n11477), .ZN(n11491) );
  INV_X2 U7718 ( .A(n10533), .ZN(n8669) );
  OR2_X1 U7719 ( .A1(n6660), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8335) );
  INV_X1 U7720 ( .A(n7474), .ZN(n7473) );
  OAI21_X1 U7721 ( .B1(n12576), .B2(n12577), .A(n13932), .ZN(n7474) );
  XNOR2_X1 U7722 ( .A(n10185), .B(n12589), .ZN(n10193) );
  NAND2_X1 U7723 ( .A1(n12588), .A2(n8985), .ZN(n10183) );
  NAND2_X1 U7724 ( .A1(n14096), .A2(n14095), .ZN(n10298) );
  OR2_X1 U7725 ( .A1(n10224), .A2(n10218), .ZN(n6865) );
  NAND2_X1 U7726 ( .A1(n6864), .A2(n6863), .ZN(n11311) );
  INV_X1 U7727 ( .A(n11314), .ZN(n6863) );
  AND3_X1 U7728 ( .A1(n9296), .A2(n9295), .A3(n9294), .ZN(n13984) );
  AND4_X1 U7729 ( .A1(n9106), .A2(n9105), .A3(n9104), .A4(n9103), .ZN(n11769)
         );
  CLKBUF_X3 U7730 ( .A(n9017), .Z(n9442) );
  NOR2_X1 U7731 ( .A1(n14899), .A2(n14202), .ZN(n14203) );
  XNOR2_X1 U7732 ( .A(n14441), .B(n14109), .ZN(n10062) );
  NAND2_X1 U7733 ( .A1(n9998), .A2(n6619), .ZN(n14330) );
  NAND2_X1 U7734 ( .A1(n14386), .A2(n7583), .ZN(n14369) );
  AND2_X1 U7735 ( .A1(n7208), .A2(n9991), .ZN(n7207) );
  NAND2_X1 U7736 ( .A1(n6789), .A2(n9967), .ZN(n14947) );
  NAND2_X1 U7737 ( .A1(n9522), .A2(n9521), .ZN(n14937) );
  NAND2_X1 U7738 ( .A1(n9396), .A2(n9395), .ZN(n14450) );
  AND2_X1 U7739 ( .A1(n7614), .A2(n9517), .ZN(n7579) );
  NAND2_X1 U7740 ( .A1(n7487), .A2(n7486), .ZN(n9513) );
  NOR2_X1 U7741 ( .A1(n7488), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n7486) );
  INV_X1 U7742 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9263) );
  NAND2_X1 U7743 ( .A1(n14665), .A2(n14664), .ZN(n7364) );
  AOI21_X1 U7744 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14577), .A(n14576), .ZN(
        n14630) );
  NOR2_X1 U7745 ( .A1(n14626), .A2(n14627), .ZN(n14576) );
  AND2_X1 U7746 ( .A1(n7132), .A2(n7134), .ZN(n6733) );
  AND2_X1 U7747 ( .A1(n8092), .A2(n8091), .ZN(n12934) );
  NOR2_X1 U7748 ( .A1(n12376), .A2(n12548), .ZN(n12377) );
  INV_X1 U7749 ( .A(n6904), .ZN(n6903) );
  NAND2_X1 U7750 ( .A1(n9336), .A2(n9335), .ZN(n14472) );
  NOR2_X2 U7751 ( .A1(n6728), .A2(n14668), .ZN(n14672) );
  OAI21_X1 U7752 ( .B1(n9602), .B2(n9601), .A(n9600), .ZN(n9604) );
  NAND2_X1 U7753 ( .A1(n6769), .A2(n6767), .ZN(n9631) );
  INV_X1 U7754 ( .A(n9629), .ZN(n6810) );
  MUX2_X1 U7755 ( .A(n11658), .B(n14131), .S(n9413), .Z(n9055) );
  NAND2_X1 U7756 ( .A1(n9057), .A2(n9058), .ZN(n9056) );
  MUX2_X1 U7757 ( .A(n14129), .B(n11878), .S(n9468), .Z(n9091) );
  NOR2_X1 U7758 ( .A1(n9151), .A2(n9148), .ZN(n7172) );
  INV_X1 U7759 ( .A(n9148), .ZN(n7171) );
  NOR2_X1 U7760 ( .A1(n9681), .A2(n6612), .ZN(n7446) );
  INV_X1 U7761 ( .A(n9300), .ZN(n7162) );
  INV_X1 U7762 ( .A(n9290), .ZN(n7167) );
  NAND2_X1 U7763 ( .A1(n9242), .A2(n7165), .ZN(n7163) );
  AND2_X1 U7764 ( .A1(n6603), .A2(n9241), .ZN(n7165) );
  INV_X1 U7765 ( .A(n7054), .ZN(n7051) );
  INV_X1 U7766 ( .A(n7038), .ZN(n7037) );
  NAND2_X1 U7767 ( .A1(n12440), .A2(n7033), .ZN(n7032) );
  OAI21_X1 U7768 ( .B1(n7039), .B2(n15336), .A(n6675), .ZN(n7038) );
  INV_X1 U7769 ( .A(n6674), .ZN(n7050) );
  AOI21_X1 U7770 ( .B1(n7054), .B2(n8127), .A(n7053), .ZN(n7052) );
  INV_X1 U7771 ( .A(n12471), .ZN(n7053) );
  OAI22_X1 U7772 ( .A1(n9701), .A2(n6759), .B1(n9700), .B2(n9702), .ZN(n9709)
         );
  NOR2_X1 U7773 ( .A1(n9703), .A2(n9699), .ZN(n6759) );
  NAND2_X1 U7774 ( .A1(n9709), .A2(n9708), .ZN(n6860) );
  INV_X1 U7775 ( .A(n9709), .ZN(n6828) );
  MUX2_X1 U7776 ( .A(n14113), .B(n14460), .S(n9468), .Z(n9367) );
  NOR2_X1 U7777 ( .A1(n7061), .A2(n12533), .ZN(n7059) );
  NAND2_X1 U7778 ( .A1(n7063), .A2(n7062), .ZN(n7061) );
  INV_X1 U7779 ( .A(n12532), .ZN(n7062) );
  NAND2_X1 U7780 ( .A1(n9719), .A2(n6678), .ZN(n7455) );
  NAND2_X1 U7781 ( .A1(n12836), .A2(n12834), .ZN(n6999) );
  AND2_X1 U7782 ( .A1(n7657), .A2(n7251), .ZN(n6895) );
  OR2_X1 U7783 ( .A1(n13449), .A2(n7540), .ZN(n7539) );
  INV_X1 U7784 ( .A(n8706), .ZN(n7540) );
  INV_X1 U7785 ( .A(n9871), .ZN(n7384) );
  AND2_X1 U7786 ( .A1(n8362), .A2(n8219), .ZN(n8220) );
  AND2_X1 U7787 ( .A1(n9398), .A2(n9399), .ZN(n7518) );
  NAND2_X1 U7788 ( .A1(n7157), .A2(n9415), .ZN(n7156) );
  INV_X1 U7789 ( .A(n7518), .ZN(n7157) );
  INV_X1 U7790 ( .A(n7155), .ZN(n7154) );
  OAI21_X1 U7791 ( .B1(n7158), .B2(n9416), .A(n9414), .ZN(n7155) );
  NAND2_X1 U7792 ( .A1(n7100), .A2(n6694), .ZN(n7099) );
  NAND2_X1 U7793 ( .A1(n9433), .A2(n7101), .ZN(n7100) );
  NOR2_X1 U7794 ( .A1(n7099), .A2(n8886), .ZN(n7096) );
  NOR2_X1 U7795 ( .A1(n7111), .A2(n8647), .ZN(n7110) );
  INV_X1 U7796 ( .A(n8625), .ZN(n7111) );
  OAI21_X1 U7797 ( .B1(n8247), .B2(n10478), .A(n6825), .ZN(n8284) );
  NAND2_X1 U7798 ( .A1(n8247), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6825) );
  INV_X1 U7799 ( .A(n14557), .ZN(n6724) );
  INV_X1 U7800 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14558) );
  INV_X1 U7801 ( .A(n7328), .ZN(n7327) );
  INV_X1 U7802 ( .A(n12648), .ZN(n7331) );
  AND2_X1 U7803 ( .A1(n6757), .A2(n6549), .ZN(n7449) );
  NOR2_X1 U7804 ( .A1(n12917), .A2(n7451), .ZN(n7450) );
  INV_X1 U7805 ( .A(n12544), .ZN(n6872) );
  INV_X1 U7806 ( .A(n7078), .ZN(n7077) );
  OAI21_X1 U7807 ( .B1(n7079), .B2(n7083), .A(n12547), .ZN(n7078) );
  AND2_X1 U7808 ( .A1(n7079), .A2(n7075), .ZN(n7074) );
  AOI21_X1 U7809 ( .B1(n6758), .B2(n7082), .A(n7081), .ZN(n7076) );
  INV_X1 U7810 ( .A(n12549), .ZN(n7081) );
  INV_X1 U7811 ( .A(n7305), .ZN(n7304) );
  AND3_X1 U7812 ( .A1(n7310), .A2(n7309), .A3(n12808), .ZN(n12810) );
  NOR2_X1 U7813 ( .A1(n12798), .A2(n14701), .ZN(n12799) );
  NAND2_X1 U7814 ( .A1(n12918), .A2(n8149), .ZN(n7613) );
  OR2_X1 U7815 ( .A1(n13375), .A2(n12949), .ZN(n12527) );
  NAND2_X1 U7816 ( .A1(n13375), .A2(n12949), .ZN(n12913) );
  AND2_X1 U7817 ( .A1(n12989), .A2(n8141), .ZN(n7609) );
  NAND2_X1 U7818 ( .A1(n12997), .A2(n12996), .ZN(n12995) );
  INV_X1 U7819 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n13244) );
  OR2_X1 U7820 ( .A1(n12247), .A2(n12713), .ZN(n12412) );
  INV_X1 U7821 ( .A(n7593), .ZN(n7589) );
  NAND2_X1 U7822 ( .A1(n15337), .A2(n8123), .ZN(n7602) );
  NAND2_X1 U7823 ( .A1(n11103), .A2(n15391), .ZN(n12427) );
  NAND2_X1 U7824 ( .A1(n12720), .A2(n10877), .ZN(n12428) );
  OR2_X1 U7825 ( .A1(n8208), .A2(n8210), .ZN(n8206) );
  OR2_X1 U7826 ( .A1(n13350), .A2(n13295), .ZN(n12491) );
  AND2_X1 U7827 ( .A1(n7413), .A2(n7412), .ZN(n7411) );
  INV_X1 U7828 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7661) );
  AND2_X1 U7829 ( .A1(n7418), .A2(n6702), .ZN(n7416) );
  AND2_X1 U7830 ( .A1(n6564), .A2(n7251), .ZN(n7250) );
  NAND2_X1 U7831 ( .A1(n8055), .A2(n8054), .ZN(n8068) );
  NAND2_X1 U7832 ( .A1(n7871), .A2(n7870), .ZN(n6756) );
  NOR2_X1 U7833 ( .A1(n8795), .A2(n13459), .ZN(n8812) );
  AND2_X1 U7834 ( .A1(n8403), .A2(n8381), .ZN(n6943) );
  INV_X1 U7835 ( .A(n13478), .ZN(n7541) );
  INV_X1 U7836 ( .A(n8663), .ZN(n6962) );
  OAI21_X1 U7837 ( .B1(n7539), .B2(n6587), .A(n8726), .ZN(n7538) );
  OR2_X1 U7838 ( .A1(n8725), .A2(n8724), .ZN(n8726) );
  NOR2_X1 U7839 ( .A1(n6961), .A2(n7539), .ZN(n6958) );
  NAND2_X1 U7840 ( .A1(n6958), .A2(n6962), .ZN(n6956) );
  AND2_X1 U7841 ( .A1(n13576), .A2(n15101), .ZN(n13578) );
  NAND2_X1 U7842 ( .A1(n15140), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7398) );
  INV_X1 U7843 ( .A(n9938), .ZN(n7275) );
  INV_X1 U7844 ( .A(n7630), .ZN(n7272) );
  OR2_X1 U7845 ( .A1(n7276), .A2(n7275), .ZN(n7274) );
  INV_X1 U7846 ( .A(n7261), .ZN(n7256) );
  NOR2_X1 U7847 ( .A1(n13697), .A2(n13682), .ZN(n13663) );
  NAND2_X1 U7848 ( .A1(n9934), .A2(n7263), .ZN(n7260) );
  INV_X1 U7849 ( .A(n13792), .ZN(n7281) );
  OR2_X1 U7850 ( .A1(n11855), .A2(n9813), .ZN(n9857) );
  XNOR2_X1 U7851 ( .A(n10897), .B(n11574), .ZN(n11569) );
  NAND2_X1 U7852 ( .A1(n13756), .A2(n6979), .ZN(n13697) );
  NOR2_X1 U7853 ( .A1(n6980), .A2(n6984), .ZN(n6979) );
  INV_X1 U7854 ( .A(n6981), .ZN(n6980) );
  INV_X1 U7855 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8261) );
  OR2_X1 U7856 ( .A1(n8519), .A2(n8261), .ZN(n6978) );
  OAI21_X1 U7857 ( .B1(n8855), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8863) );
  INV_X1 U7858 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6966) );
  INV_X1 U7859 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8224) );
  AND2_X1 U7860 ( .A1(n14027), .A2(n10383), .ZN(n12567) );
  AND2_X1 U7861 ( .A1(n10182), .A2(n10181), .ZN(n10299) );
  NAND2_X1 U7862 ( .A1(n14285), .A2(n7569), .ZN(n7568) );
  INV_X1 U7863 ( .A(n10061), .ZN(n7569) );
  NAND2_X1 U7864 ( .A1(n14355), .A2(n7582), .ZN(n7581) );
  INV_X1 U7865 ( .A(n10057), .ZN(n7582) );
  NOR2_X1 U7866 ( .A1(n14373), .A2(n7584), .ZN(n7583) );
  INV_X1 U7867 ( .A(n10056), .ZN(n7584) );
  NOR2_X1 U7868 ( .A1(n14510), .A2(n14804), .ZN(n7194) );
  NOR2_X1 U7869 ( .A1(n6501), .A2(n7552), .ZN(n7551) );
  NOR2_X1 U7870 ( .A1(n11972), .A2(n7553), .ZN(n7552) );
  INV_X1 U7871 ( .A(n14915), .ZN(n7559) );
  INV_X1 U7872 ( .A(n10032), .ZN(n7560) );
  AND2_X1 U7873 ( .A1(n9477), .A2(n10035), .ZN(n10034) );
  NAND2_X1 U7874 ( .A1(n14322), .A2(n14327), .ZN(n14321) );
  AND2_X1 U7875 ( .A1(n10024), .A2(n11824), .ZN(n10069) );
  AND2_X1 U7876 ( .A1(n8765), .A2(n8764), .ZN(n8768) );
  NAND2_X1 U7877 ( .A1(n8732), .A2(n8731), .ZN(n8748) );
  NAND2_X1 U7878 ( .A1(n8666), .A2(SI_19_), .ZN(n8688) );
  NAND2_X1 U7879 ( .A1(n7109), .A2(n8646), .ZN(n8683) );
  XNOR2_X1 U7880 ( .A(n8598), .B(SI_14_), .ZN(n8576) );
  XNOR2_X1 U7881 ( .A(n8558), .B(SI_13_), .ZN(n8556) );
  OR2_X1 U7882 ( .A1(n9160), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9161) );
  XNOR2_X1 U7883 ( .A(n8540), .B(SI_12_), .ZN(n8538) );
  NAND2_X1 U7884 ( .A1(n8476), .A2(SI_10_), .ZN(n8494) );
  INV_X1 U7885 ( .A(n7504), .ZN(n7503) );
  OAI21_X1 U7886 ( .B1(n8386), .B2(n7505), .A(n8424), .ZN(n7504) );
  OAI21_X1 U7887 ( .B1(n8407), .B2(SI_7_), .A(n8426), .ZN(n8423) );
  NOR2_X1 U7888 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n8914) );
  NAND2_X1 U7889 ( .A1(n8284), .A2(SI_2_), .ZN(n8302) );
  NAND2_X1 U7890 ( .A1(n8246), .A2(SI_1_), .ZN(n8282) );
  NAND2_X1 U7891 ( .A1(n8248), .A2(n8247), .ZN(n6913) );
  INV_X1 U7892 ( .A(n7126), .ZN(n7125) );
  NAND2_X1 U7893 ( .A1(n6850), .A2(n14565), .ZN(n14566) );
  XNOR2_X1 U7894 ( .A(n14566), .B(n13244), .ZN(n14609) );
  NAND2_X1 U7895 ( .A1(n14570), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7142) );
  NAND2_X1 U7896 ( .A1(n7140), .A2(n14575), .ZN(n14627) );
  NAND2_X1 U7897 ( .A1(n14622), .A2(n14623), .ZN(n7140) );
  NOR2_X1 U7898 ( .A1(n6585), .A2(n7325), .ZN(n7321) );
  INV_X1 U7899 ( .A(n7326), .ZN(n7325) );
  OAI21_X1 U7900 ( .B1(n7330), .B2(n7327), .A(n12682), .ZN(n7326) );
  INV_X1 U7901 ( .A(n12921), .ZN(n12529) );
  INV_X1 U7902 ( .A(n10105), .ZN(n7348) );
  OR2_X1 U7903 ( .A1(n7355), .A2(n6651), .ZN(n7354) );
  NAND2_X1 U7904 ( .A1(n10977), .A2(n7335), .ZN(n11148) );
  NOR2_X1 U7905 ( .A1(n7336), .A2(n11150), .ZN(n7335) );
  INV_X1 U7906 ( .A(n10096), .ZN(n7336) );
  INV_X1 U7907 ( .A(n6586), .ZN(n7318) );
  AND2_X1 U7908 ( .A1(n10118), .A2(n7356), .ZN(n7355) );
  INV_X1 U7909 ( .A(n10119), .ZN(n7356) );
  INV_X1 U7910 ( .A(n11447), .ZN(n7349) );
  AND2_X1 U7911 ( .A1(n12352), .A2(n12539), .ZN(n7638) );
  NOR2_X1 U7912 ( .A1(n11175), .A2(n15263), .ZN(n11174) );
  INV_X1 U7913 ( .A(n6800), .ZN(n11026) );
  OR2_X1 U7914 ( .A1(n11193), .A2(n11194), .ZN(n11014) );
  NOR2_X1 U7915 ( .A1(n11174), .A2(n11012), .ZN(n11193) );
  NAND2_X1 U7916 ( .A1(n7248), .A2(n7247), .ZN(n7246) );
  AND2_X1 U7917 ( .A1(n11132), .A2(n11133), .ZN(n11134) );
  NOR2_X1 U7918 ( .A1(n11299), .A2(n11033), .ZN(n11301) );
  AND2_X1 U7919 ( .A1(n11586), .A2(n11585), .ZN(n11587) );
  OAI21_X1 U7920 ( .B1(n11811), .B2(n7305), .A(n7302), .ZN(n6787) );
  NAND2_X1 U7921 ( .A1(n6841), .A2(n6840), .ZN(n12030) );
  XNOR2_X1 U7922 ( .A(n12031), .B(n12045), .ZN(n15292) );
  OR2_X1 U7923 ( .A1(n13420), .A2(n15255), .ZN(n11036) );
  NOR2_X1 U7924 ( .A1(n12861), .A2(n12862), .ZN(n12865) );
  AND2_X1 U7925 ( .A1(n8162), .A2(n8161), .ZN(n14719) );
  NAND2_X1 U7926 ( .A1(n6839), .A2(n7609), .ZN(n12985) );
  AOI21_X1 U7927 ( .B1(n7224), .B2(n7226), .A(n7223), .ZN(n7222) );
  INV_X1 U7928 ( .A(n12495), .ZN(n7223) );
  NAND2_X1 U7929 ( .A1(n6594), .A2(n8138), .ZN(n7595) );
  NAND2_X1 U7930 ( .A1(n7597), .A2(n8138), .ZN(n7594) );
  AND2_X1 U7931 ( .A1(n12495), .A2(n12492), .ZN(n13300) );
  NAND2_X1 U7932 ( .A1(n7599), .A2(n6594), .ZN(n7598) );
  INV_X1 U7933 ( .A(n13010), .ZN(n13295) );
  NAND2_X1 U7934 ( .A1(n12281), .A2(n12392), .ZN(n12280) );
  INV_X1 U7935 ( .A(n12714), .ZN(n14739) );
  AND2_X1 U7936 ( .A1(n12469), .A2(n12472), .ZN(n14737) );
  AND2_X1 U7937 ( .A1(n7852), .A2(n7851), .ZN(n14741) );
  NAND2_X1 U7938 ( .A1(n12530), .A2(n10172), .ZN(n15381) );
  AND2_X1 U7939 ( .A1(n9552), .A2(n12552), .ZN(n15388) );
  INV_X1 U7940 ( .A(n12350), .ZN(n12414) );
  INV_X1 U7941 ( .A(n15388), .ZN(n15341) );
  AND2_X1 U7942 ( .A1(n14718), .A2(n14717), .ZN(n14749) );
  NAND2_X1 U7943 ( .A1(n6848), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7699) );
  INV_X1 U7944 ( .A(n15324), .ZN(n15382) );
  AND2_X1 U7945 ( .A1(n8190), .A2(n8191), .ZN(n10716) );
  NAND2_X1 U7946 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7419), .ZN(n7418) );
  NAND2_X1 U7947 ( .A1(n6737), .A2(n6735), .ZN(n8095) );
  NAND2_X1 U7948 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n6736), .ZN(n6735) );
  NAND2_X1 U7949 ( .A1(n8081), .A2(n8082), .ZN(n6737) );
  INV_X1 U7950 ( .A(n6740), .ZN(n6739) );
  OAI21_X1 U7951 ( .B1(n8006), .B2(n6741), .A(n8032), .ZN(n6740) );
  NAND2_X1 U7952 ( .A1(n8007), .A2(n8006), .ZN(n8019) );
  OR2_X1 U7953 ( .A1(n8154), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8173) );
  AND2_X1 U7954 ( .A1(n7927), .A2(n7027), .ZN(n7644) );
  AND2_X1 U7955 ( .A1(n7029), .A2(n7028), .ZN(n7027) );
  NAND2_X1 U7956 ( .A1(n7992), .A2(n7993), .ZN(n8004) );
  AND2_X1 U7957 ( .A1(n6552), .A2(n7358), .ZN(n7029) );
  NAND2_X1 U7958 ( .A1(n6753), .A2(n7438), .ZN(n7943) );
  AOI21_X1 U7959 ( .B1(n6672), .B2(n7921), .A(n7439), .ZN(n7438) );
  NAND2_X1 U7960 ( .A1(n7922), .A2(n6672), .ZN(n6753) );
  INV_X1 U7961 ( .A(n7939), .ZN(n7439) );
  NAND2_X1 U7962 ( .A1(n7943), .A2(n7942), .ZN(n7958) );
  NAND2_X1 U7963 ( .A1(n7927), .A2(n7654), .ZN(n7944) );
  NAND2_X1 U7964 ( .A1(n7906), .A2(n7905), .ZN(n7922) );
  AND2_X1 U7965 ( .A1(n7641), .A2(n7024), .ZN(n7023) );
  INV_X1 U7966 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7024) );
  OR2_X1 U7967 ( .A1(n7873), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7889) );
  XNOR2_X1 U7968 ( .A(n7779), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n7793) );
  INV_X1 U7969 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U7970 ( .A1(n6751), .A2(n7764), .ZN(n7777) );
  NAND2_X1 U7971 ( .A1(n7762), .A2(n7761), .ZN(n6751) );
  NAND2_X1 U7972 ( .A1(n10483), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U7973 ( .A1(n6645), .A2(n7680), .ZN(n7425) );
  NAND2_X1 U7974 ( .A1(n7678), .A2(n7677), .ZN(n7714) );
  NAND2_X1 U7975 ( .A1(n7702), .A2(n7701), .ZN(n7678) );
  NOR2_X1 U7976 ( .A1(n13643), .A2(n13520), .ZN(n8890) );
  INV_X1 U7977 ( .A(n7529), .ZN(n6954) );
  AND2_X1 U7978 ( .A1(n13643), .A2(n7530), .ZN(n7529) );
  NAND2_X1 U7979 ( .A1(n8883), .A2(n13520), .ZN(n7530) );
  NAND2_X1 U7980 ( .A1(n6943), .A2(n10923), .ZN(n10937) );
  AND2_X1 U7981 ( .A1(n13464), .A2(n13431), .ZN(n7523) );
  NAND2_X1 U7982 ( .A1(n8682), .A2(n6587), .ZN(n13475) );
  NAND2_X1 U7983 ( .A1(n11641), .A2(n8537), .ZN(n11861) );
  NAND2_X1 U7984 ( .A1(n8805), .A2(n6581), .ZN(n13505) );
  NAND2_X1 U7985 ( .A1(n12317), .A2(n8575), .ZN(n8593) );
  AND2_X1 U7986 ( .A1(n9811), .A2(n8271), .ZN(n10532) );
  NOR2_X1 U7987 ( .A1(n9794), .A2(n9764), .ZN(n9795) );
  OAI21_X1 U7988 ( .B1(n6761), .B2(n9741), .A(n9740), .ZN(n6760) );
  NAND2_X1 U7989 ( .A1(n9793), .A2(n9792), .ZN(n7086) );
  OR2_X1 U7990 ( .A1(n10586), .A2(n10585), .ZN(n7178) );
  NOR2_X1 U7991 ( .A1(n10965), .A2(n7392), .ZN(n10969) );
  AND2_X1 U7992 ( .A1(n10966), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7392) );
  OR2_X1 U7993 ( .A1(n11955), .A2(n11956), .ZN(n13575) );
  AND2_X1 U7994 ( .A1(n15101), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7403) );
  INV_X1 U7995 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7394) );
  INV_X1 U7996 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13610) );
  NOR2_X1 U7997 ( .A1(n13693), .A2(n7262), .ZN(n7261) );
  INV_X1 U7998 ( .A(n7263), .ZN(n7262) );
  AND2_X1 U7999 ( .A1(n7375), .A2(n13677), .ZN(n7374) );
  OR2_X1 U8000 ( .A1(n7377), .A2(n7376), .ZN(n7375) );
  INV_X1 U8001 ( .A(n9882), .ZN(n7376) );
  NAND2_X1 U8002 ( .A1(n7264), .A2(n13470), .ZN(n7263) );
  NAND2_X1 U8003 ( .A1(n7377), .A2(n9881), .ZN(n13692) );
  AND2_X1 U8004 ( .A1(n13737), .A2(n9931), .ZN(n7267) );
  NAND2_X1 U8005 ( .A1(n7266), .A2(n7265), .ZN(n13729) );
  AND2_X1 U8006 ( .A1(n13730), .A2(n6606), .ZN(n7265) );
  NAND2_X1 U8007 ( .A1(n12191), .A2(n6589), .ZN(n13789) );
  NAND2_X1 U8008 ( .A1(n9924), .A2(n9923), .ZN(n7289) );
  NAND2_X1 U8009 ( .A1(n12020), .A2(n9858), .ZN(n11918) );
  OR2_X1 U8010 ( .A1(n12014), .A2(n14782), .ZN(n12015) );
  OAI21_X1 U8011 ( .B1(n11791), .B2(n9916), .A(n9917), .ZN(n11846) );
  NAND2_X1 U8012 ( .A1(n9853), .A2(n11790), .ZN(n11784) );
  INV_X1 U8013 ( .A(n9852), .ZN(n7370) );
  CLKBUF_X1 U8014 ( .A(n7618), .Z(n6849) );
  NAND2_X1 U8015 ( .A1(n6849), .A2(n9850), .ZN(n11348) );
  NAND2_X1 U8016 ( .A1(n15146), .A2(n11067), .ZN(n7389) );
  OAI22_X1 U8017 ( .A1(n10925), .A2(n10924), .B1(n13545), .B2(n11689), .ZN(
        n11085) );
  NAND2_X1 U8018 ( .A1(n6971), .A2(n6970), .ZN(n15166) );
  NAND2_X1 U8019 ( .A1(n10533), .A2(n13929), .ZN(n6971) );
  NAND2_X1 U8020 ( .A1(n9754), .A2(n9753), .ZN(n9954) );
  AOI21_X1 U8021 ( .B1(n13622), .B2(n15212), .A(n13627), .ZN(n9946) );
  NAND2_X1 U8022 ( .A1(n8734), .A2(n8733), .ZN(n13836) );
  NAND2_X1 U8023 ( .A1(n8652), .A2(n8651), .ZN(n13857) );
  NAND2_X1 U8024 ( .A1(n8438), .A2(n8437), .ZN(n11712) );
  XNOR2_X1 U8025 ( .A(n8265), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U8026 ( .A1(n8264), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8265) );
  OR2_X1 U8027 ( .A1(n8459), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8496) );
  AND3_X1 U8028 ( .A1(n8364), .A2(n8363), .A3(n8362), .ZN(n8607) );
  AND2_X1 U8029 ( .A1(n8311), .A2(n8335), .ZN(n10572) );
  OR2_X1 U8030 ( .A1(n12180), .A2(n9519), .ZN(n10182) );
  OR2_X1 U8031 ( .A1(n10005), .A2(n12257), .ZN(n9519) );
  NAND2_X1 U8032 ( .A1(n11652), .A2(n7483), .ZN(n7480) );
  INV_X1 U8033 ( .A(n7462), .ZN(n7461) );
  OAI21_X1 U8034 ( .B1(n10261), .B2(n7463), .A(n12204), .ZN(n7462) );
  AND2_X1 U8035 ( .A1(n10297), .A2(n10306), .ZN(n7470) );
  INV_X1 U8036 ( .A(n14003), .ZN(n10306) );
  NAND2_X1 U8037 ( .A1(n10382), .A2(n14027), .ZN(n14032) );
  INV_X1 U8038 ( .A(n14132), .ZN(n11316) );
  NAND2_X1 U8039 ( .A1(n7464), .A2(n10261), .ZN(n12146) );
  NAND2_X1 U8040 ( .A1(n11311), .A2(n10230), .ZN(n10232) );
  AND2_X1 U8041 ( .A1(n14547), .A2(n9520), .ZN(n10513) );
  AOI21_X1 U8042 ( .B1(n6824), .B2(n7493), .A(n6823), .ZN(n7492) );
  NAND2_X1 U8043 ( .A1(n6561), .A2(n6622), .ZN(n6823) );
  AND2_X1 U8044 ( .A1(n7494), .A2(n6661), .ZN(n7493) );
  AND4_X1 U8045 ( .A1(n9322), .A2(n9321), .A3(n9320), .A4(n9319), .ZN(n13983)
         );
  AND4_X1 U8046 ( .A1(n9255), .A2(n9254), .A3(n9253), .A4(n9252), .ZN(n14072)
         );
  INV_X1 U8047 ( .A(n9017), .ZN(n8923) );
  OR2_X1 U8048 ( .A1(n9032), .A2(n11376), .ZN(n8926) );
  OR2_X1 U8049 ( .A1(n10658), .A2(n10657), .ZN(n6929) );
  XNOR2_X1 U8050 ( .A(n14201), .B(n14906), .ZN(n14901) );
  AND2_X1 U8051 ( .A1(n10078), .A2(n14239), .ZN(n14228) );
  AND3_X1 U8052 ( .A1(n7184), .A2(n14259), .A3(n14311), .ZN(n14239) );
  NOR2_X1 U8053 ( .A1(n14446), .A2(n7185), .ZN(n7184) );
  INV_X1 U8054 ( .A(n7186), .ZN(n7185) );
  OAI211_X1 U8055 ( .C1(n14276), .C2(n6797), .A(n6796), .B(n6642), .ZN(n14245)
         );
  OR2_X1 U8056 ( .A1(n7187), .A2(n14450), .ZN(n14255) );
  INV_X1 U8057 ( .A(n7568), .ZN(n7566) );
  INV_X1 U8058 ( .A(n14303), .ZN(n7567) );
  NOR2_X1 U8059 ( .A1(n14314), .A2(n13949), .ZN(n10061) );
  XNOR2_X1 U8060 ( .A(n14460), .B(n14113), .ZN(n14285) );
  NOR2_X1 U8061 ( .A1(n14314), .A2(n14331), .ZN(n14311) );
  NOR2_X1 U8062 ( .A1(n14300), .A2(n14299), .ZN(n14303) );
  INV_X1 U8063 ( .A(n6794), .ZN(n6793) );
  INV_X1 U8064 ( .A(n7217), .ZN(n6795) );
  NOR2_X1 U8065 ( .A1(n7218), .A2(n14355), .ZN(n7217) );
  INV_X1 U8066 ( .A(n9995), .ZN(n7218) );
  NAND2_X1 U8067 ( .A1(n9993), .A2(n9992), .ZN(n14371) );
  OR2_X1 U8068 ( .A1(n14371), .A2(n9994), .ZN(n14372) );
  NAND2_X1 U8069 ( .A1(n10055), .A2(n10054), .ZN(n14386) );
  NAND2_X1 U8070 ( .A1(n12117), .A2(n9986), .ZN(n12167) );
  NAND2_X1 U8071 ( .A1(n10050), .A2(n10049), .ZN(n12159) );
  AND4_X1 U8072 ( .A1(n9233), .A2(n9232), .A3(n9231), .A4(n9230), .ZN(n14011)
         );
  NOR2_X1 U8073 ( .A1(n11773), .A2(n7555), .ZN(n7554) );
  INV_X1 U8074 ( .A(n10039), .ZN(n7555) );
  INV_X1 U8075 ( .A(n7576), .ZN(n11527) );
  AOI21_X1 U8076 ( .B1(n7574), .B2(n7572), .A(n7571), .ZN(n7570) );
  INV_X1 U8077 ( .A(n7574), .ZN(n7573) );
  NAND2_X1 U8078 ( .A1(n11527), .A2(n11526), .ZN(n11525) );
  NOR2_X1 U8079 ( .A1(n11399), .A2(n7575), .ZN(n7574) );
  INV_X1 U8080 ( .A(n10036), .ZN(n7575) );
  NAND2_X1 U8081 ( .A1(n11509), .A2(n11508), .ZN(n11507) );
  NAND2_X1 U8082 ( .A1(n9965), .A2(n9964), .ZN(n11364) );
  NAND2_X1 U8083 ( .A1(n8951), .A2(n6628), .ZN(n8985) );
  OAI22_X1 U8084 ( .A1(n10477), .A2(n10476), .B1(n7212), .B2(n6799), .ZN(n6798) );
  INV_X1 U8085 ( .A(n14231), .ZN(n14438) );
  INV_X1 U8086 ( .A(n7196), .ZN(n6885) );
  AOI21_X1 U8087 ( .B1(n14441), .B2(n14979), .A(n14440), .ZN(n7196) );
  NAND2_X1 U8088 ( .A1(n9258), .A2(n9257), .ZN(n14498) );
  OR2_X1 U8089 ( .A1(n10680), .A2(n14415), .ZN(n14966) );
  NAND2_X1 U8090 ( .A1(n7546), .A2(n7219), .ZN(n8925) );
  NAND2_X1 U8091 ( .A1(n8920), .A2(n6558), .ZN(n7546) );
  XNOR2_X1 U8092 ( .A(n9435), .B(n9456), .ZN(n13912) );
  INV_X1 U8093 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8936) );
  AND4_X1 U8094 ( .A1(n8916), .A2(n8917), .A3(n8915), .A4(n9514), .ZN(n7614)
         );
  XNOR2_X1 U8095 ( .A(n8748), .B(SI_22_), .ZN(n9324) );
  NAND2_X1 U8096 ( .A1(n8964), .A2(n7491), .ZN(n7490) );
  INV_X1 U8097 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7491) );
  INV_X1 U8098 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8963) );
  XNOR2_X1 U8099 ( .A(n8968), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9520) );
  OAI21_X1 U8100 ( .B1(n8969), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8968) );
  NOR2_X1 U8101 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n8910) );
  XNOR2_X1 U8102 ( .A(n8576), .B(n8596), .ZN(n9168) );
  NAND2_X1 U8103 ( .A1(n8452), .A2(n8451), .ZN(n8456) );
  AND3_X1 U8104 ( .A1(n8913), .A2(n8948), .A3(n8914), .ZN(n9072) );
  NAND2_X1 U8105 ( .A1(n8303), .A2(n8302), .ZN(n8308) );
  INV_X1 U8106 ( .A(n8307), .ZN(n7201) );
  INV_X1 U8107 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14560) );
  INV_X1 U8108 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14603) );
  XOR2_X1 U8109 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14609), .Z(n14611) );
  NAND2_X1 U8110 ( .A1(n14620), .A2(n14621), .ZN(n14625) );
  XNOR2_X1 U8111 ( .A(n14627), .B(n7139), .ZN(n14628) );
  INV_X1 U8112 ( .A(n14626), .ZN(n7139) );
  OR2_X1 U8113 ( .A1(n14666), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6729) );
  OAI21_X1 U8114 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n14579), .A(n14578), .ZN(
        n14633) );
  INV_X1 U8115 ( .A(n6814), .ZN(n14638) );
  NOR2_X1 U8116 ( .A1(n7340), .A2(n7343), .ZN(n7339) );
  NAND2_X1 U8117 ( .A1(n7344), .A2(n7345), .ZN(n7341) );
  INV_X1 U8118 ( .A(n12960), .ZN(n12933) );
  NAND2_X1 U8119 ( .A1(n11935), .A2(n10115), .ZN(n11936) );
  NAND2_X1 U8120 ( .A1(n9535), .A2(n9534), .ZN(n12301) );
  NAND2_X1 U8121 ( .A1(n8110), .A2(n10839), .ZN(n11209) );
  NAND2_X1 U8122 ( .A1(n7337), .A2(n10873), .ZN(n10977) );
  AND2_X1 U8123 ( .A1(n10978), .A2(n10976), .ZN(n7337) );
  AND2_X1 U8124 ( .A1(n8051), .A2(n8050), .ZN(n12976) );
  NAND2_X1 U8125 ( .A1(n8024), .A2(n8023), .ZN(n12979) );
  NAND2_X1 U8126 ( .A1(n11336), .A2(n6591), .ZN(n11449) );
  NAND2_X1 U8127 ( .A1(n10156), .A2(n10155), .ZN(n12696) );
  INV_X1 U8128 ( .A(n12696), .ZN(n12691) );
  NAND2_X1 U8129 ( .A1(n11219), .A2(n10158), .ZN(n12706) );
  OR2_X1 U8130 ( .A1(n12557), .A2(n12556), .ZN(n7022) );
  OAI211_X1 U8131 ( .C1(n12363), .C2(n13099), .A(n8002), .B(n8001), .ZN(n13011) );
  NAND2_X1 U8132 ( .A1(n12360), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7741) );
  INV_X1 U8133 ( .A(n15290), .ZN(n15281) );
  NOR2_X1 U8134 ( .A1(n12844), .A2(n12830), .ZN(n12833) );
  AND2_X1 U8135 ( .A1(n12829), .A2(n12828), .ZN(n12830) );
  INV_X1 U8136 ( .A(n12890), .ZN(n7017) );
  NOR2_X1 U8137 ( .A1(n12865), .A2(n12864), .ZN(n12877) );
  NAND2_X1 U8138 ( .A1(n12877), .A2(n12882), .ZN(n6780) );
  NOR2_X1 U8139 ( .A1(n15298), .A2(n6782), .ZN(n6781) );
  AND2_X1 U8140 ( .A1(n12882), .A2(n12876), .ZN(n6782) );
  XNOR2_X1 U8141 ( .A(n12886), .B(n7021), .ZN(n7020) );
  INV_X1 U8142 ( .A(n12885), .ZN(n7021) );
  AOI21_X1 U8143 ( .B1(n13411), .B2(n12370), .A(n12359), .ZN(n14745) );
  NAND2_X1 U8144 ( .A1(n12915), .A2(n7241), .ZN(n9546) );
  AND3_X1 U8145 ( .A1(n7752), .A2(n7751), .A3(n7750), .ZN(n15365) );
  AND2_X1 U8146 ( .A1(n8099), .A2(n8098), .ZN(n13368) );
  NAND2_X1 U8147 ( .A1(n8043), .A2(n8042), .ZN(n13383) );
  NAND2_X1 U8148 ( .A1(n7978), .A2(n7977), .ZN(n13400) );
  OR2_X1 U8149 ( .A1(n8008), .A2(n6843), .ZN(n7734) );
  NAND2_X2 U8150 ( .A1(n8483), .A2(n8482), .ZN(n15232) );
  OR2_X1 U8151 ( .A1(n10525), .A2(n8359), .ZN(n8483) );
  NAND2_X1 U8152 ( .A1(n8671), .A2(n8670), .ZN(n13853) );
  OAI21_X1 U8153 ( .B1(n8805), .B2(n7534), .A(n7531), .ZN(n8854) );
  OR2_X1 U8154 ( .A1(n13424), .A2(n7535), .ZN(n7534) );
  AOI21_X1 U8155 ( .B1(n7533), .B2(n7532), .A(n6633), .ZN(n7531) );
  NAND2_X1 U8156 ( .A1(n8714), .A2(n8713), .ZN(n13744) );
  NAND2_X1 U8157 ( .A1(n8613), .A2(n8612), .ZN(n13869) );
  NAND2_X1 U8158 ( .A1(n8693), .A2(n8692), .ZN(n13757) );
  NOR2_X1 U8159 ( .A1(n15057), .A2(n7400), .ZN(n10557) );
  NAND2_X1 U8160 ( .A1(n6817), .A2(n6815), .ZN(n7182) );
  INV_X1 U8161 ( .A(n6816), .ZN(n6815) );
  NAND2_X1 U8162 ( .A1(n7183), .A2(n13605), .ZN(n6817) );
  OAI21_X1 U8163 ( .B1(n13606), .B2(n15120), .A(n11968), .ZN(n6816) );
  XNOR2_X1 U8164 ( .A(n13617), .B(n13612), .ZN(n13613) );
  NAND2_X1 U8165 ( .A1(n13807), .A2(n9938), .ZN(n13630) );
  AOI22_X1 U8166 ( .A1(n8333), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n8669), .B2(
        n15065), .ZN(n8291) );
  INV_X1 U8167 ( .A(n9946), .ZN(n9947) );
  AND2_X1 U8168 ( .A1(n13797), .A2(n13800), .ZN(n13875) );
  NAND2_X1 U8169 ( .A1(n9946), .A2(n15242), .ZN(n7269) );
  OAI211_X1 U8170 ( .C1(n13806), .C2(n13861), .A(n13805), .B(n13804), .ZN(
        n13881) );
  AOI21_X1 U8171 ( .B1(n11652), .B2(n11653), .A(n10238), .ZN(n11665) );
  OAI21_X1 U8172 ( .B1(n14078), .B2(n12577), .A(n7473), .ZN(n13930) );
  NAND2_X1 U8173 ( .A1(n10336), .A2(n10335), .ZN(n13982) );
  OAI21_X1 U8174 ( .B1(n10488), .B2(n9118), .A(n9031), .ZN(n11287) );
  NAND2_X1 U8175 ( .A1(n9298), .A2(n9297), .ZN(n14492) );
  OR2_X1 U8176 ( .A1(n9118), .A2(n8958), .ZN(n8962) );
  AND2_X1 U8177 ( .A1(n10782), .A2(n10394), .ZN(n14103) );
  INV_X1 U8178 ( .A(n14214), .ZN(n6877) );
  AOI21_X1 U8179 ( .B1(n14215), .B2(n14903), .A(n14218), .ZN(n6876) );
  NAND2_X1 U8180 ( .A1(n14219), .A2(n14218), .ZN(n6878) );
  AND2_X1 U8181 ( .A1(n14110), .A2(n14052), .ZN(n10064) );
  INV_X1 U8182 ( .A(n14443), .ZN(n10027) );
  NAND2_X1 U8183 ( .A1(n14274), .A2(n10002), .ZN(n14260) );
  NAND2_X1 U8184 ( .A1(n14330), .A2(n10000), .ZN(n14307) );
  NAND2_X1 U8185 ( .A1(n14546), .A2(n8983), .ZN(n14348) );
  NAND2_X1 U8186 ( .A1(n9312), .A2(n9311), .ZN(n14486) );
  NAND2_X1 U8187 ( .A1(n9268), .A2(n9267), .ZN(n14502) );
  INV_X1 U8188 ( .A(n14334), .ZN(n14953) );
  OR2_X1 U8189 ( .A1(n14942), .A2(n10680), .ZN(n14432) );
  NAND2_X1 U8190 ( .A1(n15452), .A2(n15453), .ZN(n14599) );
  NAND2_X1 U8191 ( .A1(n7117), .A2(n14557), .ZN(n14595) );
  XNOR2_X1 U8192 ( .A(n14625), .B(n14624), .ZN(n14666) );
  NAND2_X1 U8193 ( .A1(n6870), .A2(n6869), .ZN(n7116) );
  INV_X1 U8194 ( .A(n14671), .ZN(n6869) );
  OR2_X1 U8195 ( .A1(n14854), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7136) );
  INV_X1 U8196 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14694) );
  NAND2_X1 U8197 ( .A1(n7360), .A2(n6673), .ZN(n6915) );
  OAI22_X1 U8198 ( .A1(n9041), .A2(n7168), .B1(n7169), .B2(n9042), .ZN(n9057)
         );
  AND2_X1 U8199 ( .A1(n9042), .A2(n7169), .ZN(n7168) );
  INV_X1 U8200 ( .A(n9040), .ZN(n7169) );
  NAND2_X1 U8201 ( .A1(n6830), .A2(n7436), .ZN(n6766) );
  NAND2_X1 U8202 ( .A1(n9635), .A2(n6562), .ZN(n7436) );
  NAND2_X1 U8203 ( .A1(n6811), .A2(n6810), .ZN(n6809) );
  OAI22_X1 U8204 ( .A1(n9077), .A2(n6557), .B1(n9078), .B2(n7170), .ZN(n9093)
         );
  NAND2_X1 U8205 ( .A1(n7443), .A2(n6565), .ZN(n6920) );
  OAI22_X1 U8206 ( .A1(n9110), .A2(n7174), .B1(n9111), .B2(n7173), .ZN(n9126)
         );
  NOR2_X1 U8207 ( .A1(n9112), .A2(n9109), .ZN(n7174) );
  INV_X1 U8208 ( .A(n9109), .ZN(n7173) );
  NAND2_X1 U8209 ( .A1(n7437), .A2(n6567), .ZN(n6922) );
  OR2_X1 U8210 ( .A1(n9166), .A2(n9167), .ZN(n9197) );
  NAND2_X1 U8211 ( .A1(n9681), .A2(n6612), .ZN(n7444) );
  NAND2_X1 U8212 ( .A1(n6776), .A2(n9686), .ZN(n6775) );
  OAI21_X1 U8213 ( .B1(n12447), .B2(n11700), .A(n7043), .ZN(n7035) );
  INV_X1 U8214 ( .A(n12453), .ZN(n7043) );
  INV_X1 U8215 ( .A(n7040), .ZN(n7039) );
  OAI21_X1 U8216 ( .B1(n12448), .B2(n7036), .A(n7034), .ZN(n7040) );
  INV_X1 U8217 ( .A(n7035), .ZN(n7034) );
  NAND2_X1 U8218 ( .A1(n12454), .A2(n8119), .ZN(n7036) );
  AND2_X1 U8219 ( .A1(n7041), .A2(n7042), .ZN(n7033) );
  NAND2_X1 U8220 ( .A1(n12439), .A2(n12454), .ZN(n7031) );
  MUX2_X1 U8221 ( .A(n14117), .B(n14486), .S(n9468), .Z(n9313) );
  AND2_X1 U8222 ( .A1(n7162), .A2(n7167), .ZN(n7161) );
  AND2_X1 U8223 ( .A1(n7049), .A2(n6569), .ZN(n7046) );
  NOR2_X1 U8224 ( .A1(n7051), .A2(n7050), .ZN(n7049) );
  AOI21_X1 U8225 ( .B1(n7047), .B2(n6569), .A(n6683), .ZN(n7045) );
  OAI21_X1 U8226 ( .B1(n7052), .B2(n7050), .A(n7048), .ZN(n7047) );
  INV_X1 U8227 ( .A(n12474), .ZN(n7048) );
  NAND2_X1 U8228 ( .A1(n6829), .A2(n6826), .ZN(n6772) );
  INV_X1 U8229 ( .A(n9708), .ZN(n6827) );
  NAND2_X1 U8230 ( .A1(n9337), .A2(n9339), .ZN(n7145) );
  MUX2_X1 U8231 ( .A(n14114), .B(n14314), .S(n9468), .Z(n9352) );
  NAND2_X1 U8232 ( .A1(n12526), .A2(n6556), .ZN(n7060) );
  NOR2_X1 U8233 ( .A1(n9719), .A2(n6678), .ZN(n7456) );
  INV_X1 U8234 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7650) );
  NAND2_X1 U8235 ( .A1(n9448), .A2(n11764), .ZN(n9450) );
  AND2_X1 U8236 ( .A1(n9369), .A2(n7508), .ZN(n7507) );
  INV_X1 U8237 ( .A(n9367), .ZN(n7508) );
  INV_X1 U8238 ( .A(n9424), .ZN(n7101) );
  NOR2_X1 U8239 ( .A1(n7112), .A2(n7108), .ZN(n7107) );
  INV_X1 U8240 ( .A(n8646), .ZN(n7108) );
  INV_X1 U8241 ( .A(n8644), .ZN(n8645) );
  INV_X1 U8242 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7094) );
  AOI21_X1 U8243 ( .B1(n7059), .B2(n6626), .A(n6559), .ZN(n7058) );
  NOR2_X1 U8244 ( .A1(n12529), .A2(n12530), .ZN(n7067) );
  AND2_X1 U8245 ( .A1(n12545), .A2(n12530), .ZN(n7082) );
  OR2_X1 U8246 ( .A1(n13383), .A2(n12976), .ZN(n12522) );
  INV_X1 U8247 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7611) );
  INV_X1 U8248 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U8249 ( .A1(n9729), .A2(n6640), .ZN(n7435) );
  NAND2_X1 U8250 ( .A1(n7089), .A2(n7088), .ZN(n7087) );
  INV_X1 U8251 ( .A(n9783), .ZN(n7088) );
  NAND2_X1 U8252 ( .A1(n11672), .A2(n6578), .ZN(n9815) );
  NOR2_X1 U8253 ( .A1(n13713), .A2(n6982), .ZN(n6981) );
  INV_X1 U8254 ( .A(n6983), .ZN(n6982) );
  INV_X1 U8255 ( .A(n9430), .ZN(n7496) );
  NOR2_X1 U8256 ( .A1(n7191), .A2(n12168), .ZN(n14375) );
  OR2_X1 U8257 ( .A1(n7193), .A2(n14498), .ZN(n7191) );
  INV_X1 U8258 ( .A(n9980), .ZN(n7204) );
  INV_X1 U8259 ( .A(n8559), .ZN(n7517) );
  NOR2_X1 U8260 ( .A1(n8556), .A2(n7517), .ZN(n7516) );
  INV_X1 U8261 ( .A(n8603), .ZN(n7513) );
  NOR2_X1 U8262 ( .A1(n8513), .A2(n7510), .ZN(n7509) );
  INV_X1 U8263 ( .A(n8494), .ZN(n7510) );
  OAI21_X1 U8264 ( .B1(n9323), .B2(n10481), .A(n6858), .ZN(n8328) );
  NAND2_X1 U8265 ( .A1(n9323), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6858) );
  AND2_X1 U8266 ( .A1(n7122), .A2(n14593), .ZN(n6851) );
  NAND2_X1 U8267 ( .A1(n7126), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n7122) );
  NAND2_X1 U8268 ( .A1(n14573), .A2(n14572), .ZN(n14574) );
  NAND2_X1 U8269 ( .A1(n14618), .A2(n14619), .ZN(n14572) );
  OR2_X1 U8270 ( .A1(n12301), .A2(n6543), .ZN(n12534) );
  INV_X1 U8271 ( .A(n12237), .ZN(n7353) );
  OR2_X1 U8272 ( .A1(n11197), .A2(n11045), .ZN(n11048) );
  XNOR2_X1 U8273 ( .A(n11303), .B(n11033), .ZN(n11055) );
  AND2_X1 U8274 ( .A1(n12729), .A2(n11053), .ZN(n11303) );
  NOR2_X1 U8275 ( .A1(n11055), .A2(n7668), .ZN(n11304) );
  AND2_X1 U8276 ( .A1(n11605), .A2(n11604), .ZN(n11606) );
  NAND2_X1 U8277 ( .A1(n7305), .A2(n7302), .ZN(n7301) );
  INV_X1 U8278 ( .A(n11609), .ZN(n7300) );
  NOR2_X1 U8279 ( .A1(n11614), .A2(n7788), .ZN(n7305) );
  OR2_X1 U8280 ( .A1(n12036), .A2(n12037), .ZN(n7010) );
  NAND2_X1 U8281 ( .A1(n12757), .A2(n12756), .ZN(n6900) );
  NAND2_X1 U8282 ( .A1(n12797), .A2(n12796), .ZN(n12798) );
  NAND2_X1 U8283 ( .A1(n7000), .A2(n6997), .ZN(n12878) );
  INV_X1 U8284 ( .A(n6998), .ZN(n6997) );
  OAI21_X1 U8285 ( .B1(n12837), .B2(n6999), .A(n12851), .ZN(n6998) );
  AND2_X1 U8286 ( .A1(n12533), .A2(n8151), .ZN(n7612) );
  INV_X1 U8287 ( .A(n12522), .ZN(n8053) );
  INV_X1 U8288 ( .A(n12498), .ZN(n7229) );
  OR2_X1 U8289 ( .A1(n13400), .A2(n12686), .ZN(n12498) );
  INV_X1 U8290 ( .A(n7225), .ZN(n7224) );
  OAI21_X1 U8291 ( .B1(n12392), .B2(n7226), .A(n13300), .ZN(n7225) );
  NAND2_X1 U8292 ( .A1(n11342), .A2(n15365), .ZN(n12437) );
  NAND2_X1 U8293 ( .A1(n15380), .A2(n15379), .ZN(n15378) );
  INV_X1 U8294 ( .A(n8018), .ZN(n6741) );
  INV_X1 U8295 ( .A(n7684), .ZN(n7026) );
  NAND2_X1 U8296 ( .A1(n10491), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7778) );
  INV_X1 U8297 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7605) );
  INV_X1 U8298 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8248) );
  INV_X1 U8299 ( .A(n13507), .ZN(n7536) );
  INV_X1 U8300 ( .A(n9787), .ZN(n9791) );
  NOR2_X1 U8301 ( .A1(n13643), .A2(n6995), .ZN(n6994) );
  INV_X1 U8302 ( .A(n6996), .ZN(n6995) );
  NOR2_X1 U8303 ( .A1(n13809), .A2(n13815), .ZN(n6996) );
  INV_X1 U8304 ( .A(n13891), .ZN(n6984) );
  NOR2_X1 U8305 ( .A1(n13836), .A2(n13744), .ZN(n6983) );
  INV_X1 U8306 ( .A(n7381), .ZN(n7380) );
  OAI21_X1 U8307 ( .B1(n7383), .B2(n7382), .A(n9875), .ZN(n7381) );
  NOR2_X1 U8308 ( .A1(n13736), .A2(n7384), .ZN(n7383) );
  INV_X1 U8309 ( .A(n9874), .ZN(n7382) );
  NAND2_X1 U8310 ( .A1(n6599), .A2(n9928), .ZN(n7280) );
  NOR2_X1 U8311 ( .A1(n6990), .A2(n12340), .ZN(n6989) );
  INV_X1 U8312 ( .A(n6991), .ZN(n6990) );
  INV_X1 U8313 ( .A(n7287), .ZN(n7286) );
  NOR2_X1 U8314 ( .A1(n12109), .A2(n13869), .ZN(n6991) );
  NOR2_X1 U8315 ( .A1(n12015), .A2(n11926), .ZN(n11923) );
  INV_X1 U8316 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8462) );
  AND2_X1 U8317 ( .A1(n9585), .A2(n13700), .ZN(n11250) );
  INV_X1 U8318 ( .A(n11871), .ZN(n7479) );
  INV_X1 U8319 ( .A(n11664), .ZN(n7485) );
  AND2_X1 U8320 ( .A1(n10344), .A2(n10343), .ZN(n10346) );
  NAND2_X1 U8321 ( .A1(n9454), .A2(n7495), .ZN(n7494) );
  NOR2_X1 U8322 ( .A1(n6588), .A2(n7154), .ZN(n7153) );
  AOI22_X1 U8323 ( .A1(n6588), .A2(n7518), .B1(n7154), .B2(n7156), .ZN(n7152)
         );
  AOI21_X1 U8324 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14211), .A(n14879), .ZN(
        n14212) );
  NOR2_X1 U8325 ( .A1(n14883), .A2(n6930), .ZN(n14201) );
  AND2_X1 U8326 ( .A1(n14211), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6930) );
  INV_X1 U8327 ( .A(n7634), .ZN(n7213) );
  NOR2_X1 U8328 ( .A1(n14261), .A2(n7215), .ZN(n7214) );
  INV_X1 U8329 ( .A(n10002), .ZN(n7215) );
  NOR2_X1 U8330 ( .A1(n14455), .A2(n14460), .ZN(n7186) );
  AOI21_X1 U8331 ( .B1(n7217), .B2(n9994), .A(n6630), .ZN(n7216) );
  NOR2_X1 U8332 ( .A1(n6550), .A2(n9276), .ZN(n7211) );
  OR2_X1 U8333 ( .A1(n6550), .A2(n7209), .ZN(n7208) );
  NAND2_X1 U8334 ( .A1(n9990), .A2(n9989), .ZN(n7209) );
  OR2_X1 U8335 ( .A1(n14498), .A2(n14038), .ZN(n9472) );
  NAND2_X1 U8336 ( .A1(n14409), .A2(n7194), .ZN(n7193) );
  NAND2_X1 U8337 ( .A1(n11980), .A2(n10067), .ZN(n12078) );
  NOR2_X1 U8338 ( .A1(n11990), .A2(n14827), .ZN(n11980) );
  AND2_X1 U8339 ( .A1(n7189), .A2(n7190), .ZN(n7188) );
  NOR2_X1 U8340 ( .A1(n12010), .A2(n15022), .ZN(n7190) );
  INV_X1 U8341 ( .A(n10037), .ZN(n7571) );
  INV_X1 U8342 ( .A(n14131), .ZN(n10234) );
  NOR2_X1 U8343 ( .A1(n11721), .A2(n11333), .ZN(n11329) );
  INV_X1 U8344 ( .A(n10476), .ZN(n6799) );
  NAND2_X1 U8345 ( .A1(n14137), .A2(n14964), .ZN(n9479) );
  AND2_X1 U8346 ( .A1(n10066), .A2(n11329), .ZN(n14949) );
  INV_X1 U8347 ( .A(n7543), .ZN(n7220) );
  OAI21_X1 U8348 ( .B1(n7545), .B2(P1_IR_REG_30__SCAN_IN), .A(n7544), .ZN(
        n7543) );
  NAND2_X1 U8349 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n7544) );
  NOR2_X1 U8350 ( .A1(n8921), .A2(n8935), .ZN(n7545) );
  OAI22_X1 U8351 ( .A1(n7097), .A2(n7095), .B1(n7099), .B2(n6688), .ZN(n9457)
         );
  NAND2_X1 U8352 ( .A1(n8828), .A2(n7096), .ZN(n7095) );
  NOR2_X1 U8353 ( .A1(n9425), .A2(n7103), .ZN(n7102) );
  INV_X1 U8354 ( .A(n8885), .ZN(n7103) );
  NAND2_X1 U8355 ( .A1(n7489), .A2(n9504), .ZN(n7488) );
  INV_X1 U8356 ( .A(n7490), .ZN(n7489) );
  NAND2_X1 U8357 ( .A1(n8712), .A2(n8711), .ZN(n8729) );
  OR2_X1 U8358 ( .A1(n8710), .A2(n13024), .ZN(n8711) );
  XNOR2_X1 U8359 ( .A(n8710), .B(SI_20_), .ZN(n8709) );
  OAI21_X1 U8360 ( .B1(n8247), .B2(n10483), .A(n6897), .ZN(n8304) );
  NAND2_X1 U8361 ( .A1(n8247), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6897) );
  INV_X1 U8362 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14556) );
  NAND2_X1 U8363 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n14558), .ZN(n14559) );
  INV_X1 U8364 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14570) );
  XOR2_X1 U8365 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n14574), .Z(n14622) );
  OAI21_X1 U8366 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n14585), .A(n14584), .ZN(
        n14642) );
  NAND2_X1 U8367 ( .A1(n7138), .A2(n7133), .ZN(n7132) );
  NOR2_X1 U8368 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n7133) );
  OR2_X1 U8369 ( .A1(n8025), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8044) );
  NOR2_X1 U8370 ( .A1(n7979), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U8371 ( .A1(n12534), .A2(n9578), .ZN(n12399) );
  AND2_X1 U8372 ( .A1(n10149), .A2(n10148), .ZN(n12630) );
  OR2_X1 U8373 ( .A1(n8044), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U8374 ( .A1(n7333), .A2(n12625), .ZN(n12673) );
  NAND2_X1 U8375 ( .A1(n7357), .A2(n10119), .ZN(n10416) );
  NAND2_X1 U8376 ( .A1(n11936), .A2(n10118), .ZN(n7357) );
  AOI21_X1 U8377 ( .B1(n7331), .B2(n6582), .A(n7329), .ZN(n7328) );
  NOR2_X1 U8378 ( .A1(n10130), .A2(n12644), .ZN(n7329) );
  AND2_X1 U8379 ( .A1(n7331), .A2(n12638), .ZN(n7330) );
  AND4_X1 U8380 ( .A1(n12397), .A2(n12541), .A3(n7636), .A4(n12396), .ZN(
        n12398) );
  AND2_X1 U8381 ( .A1(n12549), .A2(n7449), .ZN(n7448) );
  NAND3_X1 U8382 ( .A1(n7072), .A2(n6871), .A3(n7071), .ZN(n6750) );
  AOI21_X1 U8383 ( .B1(n7077), .B2(n7074), .A(n7073), .ZN(n7072) );
  NAND2_X1 U8384 ( .A1(n6872), .A2(n6624), .ZN(n6871) );
  NAND2_X1 U8385 ( .A1(n6750), .A2(n12550), .ZN(n6749) );
  OR2_X1 U8386 ( .A1(n7755), .A2(n11005), .ZN(n7709) );
  NAND2_X1 U8387 ( .A1(n11039), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11040) );
  AOI21_X1 U8388 ( .B1(n11041), .B2(n11040), .A(n7306), .ZN(n11180) );
  NOR2_X1 U8389 ( .A1(n11040), .A2(n7307), .ZN(n7306) );
  NOR2_X1 U8390 ( .A1(n11198), .A2(n11199), .ZN(n11197) );
  XNOR2_X1 U8391 ( .A(n11048), .B(n11047), .ZN(n11141) );
  NOR2_X1 U8392 ( .A1(n11141), .A2(n11000), .ZN(n11140) );
  NOR2_X1 U8393 ( .A1(n11130), .A2(n11029), .ZN(n12724) );
  NAND2_X1 U8394 ( .A1(n7315), .A2(n6705), .ZN(n11605) );
  INV_X1 U8395 ( .A(n6704), .ZN(n7234) );
  OR2_X1 U8396 ( .A1(n11034), .A2(n11035), .ZN(n7237) );
  OR2_X1 U8397 ( .A1(n7796), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7817) );
  NOR2_X1 U8398 ( .A1(n11610), .A2(n11609), .ZN(n11811) );
  AND2_X1 U8399 ( .A1(n7010), .A2(n12039), .ZN(n15293) );
  OR2_X1 U8400 ( .A1(n15292), .A2(n7841), .ZN(n7291) );
  AND2_X1 U8401 ( .A1(n12030), .A2(n12029), .ZN(n12031) );
  NOR2_X1 U8402 ( .A1(n15284), .A2(n12047), .ZN(n12741) );
  NAND2_X1 U8403 ( .A1(n7221), .A2(n12742), .ZN(n12766) );
  OR2_X1 U8404 ( .A1(n12741), .A2(n12740), .ZN(n7221) );
  NOR2_X1 U8405 ( .A1(n7008), .A2(n12746), .ZN(n7006) );
  AND2_X1 U8406 ( .A1(n6900), .A2(n12772), .ZN(n12765) );
  NOR2_X1 U8407 ( .A1(n12750), .A2(n12751), .ZN(n12776) );
  OR2_X1 U8408 ( .A1(n12776), .A2(n7011), .ZN(n12797) );
  OR2_X1 U8409 ( .A1(n12777), .A2(n12775), .ZN(n7011) );
  OR2_X1 U8410 ( .A1(n12758), .A2(n7311), .ZN(n7310) );
  NAND2_X1 U8411 ( .A1(n7312), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U8412 ( .A1(n12765), .A2(n7312), .ZN(n7309) );
  OAI21_X1 U8413 ( .B1(n14702), .B2(n6785), .A(n6784), .ZN(n12859) );
  NAND2_X1 U8414 ( .A1(n12813), .A2(n12821), .ZN(n6784) );
  NAND2_X1 U8415 ( .A1(n6786), .A2(n12821), .ZN(n6785) );
  INV_X1 U8416 ( .A(n12812), .ZN(n6786) );
  NOR2_X1 U8417 ( .A1(n12837), .A2(n7002), .ZN(n7001) );
  INV_X1 U8418 ( .A(n12834), .ZN(n7002) );
  NAND2_X1 U8419 ( .A1(n7005), .A2(n7004), .ZN(n7003) );
  INV_X1 U8420 ( .A(n12835), .ZN(n7005) );
  AOI21_X1 U8421 ( .B1(n7241), .B2(n7240), .A(n7239), .ZN(n7238) );
  INV_X1 U8422 ( .A(n12536), .ZN(n7239) );
  INV_X1 U8423 ( .A(n8094), .ZN(n7240) );
  NAND2_X1 U8424 ( .A1(n9547), .A2(n9537), .ZN(n9579) );
  INV_X1 U8425 ( .A(n8171), .ZN(n6905) );
  OR2_X1 U8426 ( .A1(n8150), .A2(n12934), .ZN(n12402) );
  NAND2_X1 U8427 ( .A1(n12402), .A2(n12401), .ZN(n12917) );
  INV_X1 U8428 ( .A(n7607), .ZN(n7606) );
  OAI21_X1 U8429 ( .B1(n7609), .B2(n6593), .A(n8143), .ZN(n7607) );
  AND2_X1 U8430 ( .A1(n7998), .A2(n13221), .ZN(n8012) );
  INV_X1 U8431 ( .A(n13001), .ZN(n12996) );
  OR2_X1 U8432 ( .A1(n7965), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7979) );
  AND2_X1 U8433 ( .A1(n7933), .A2(n12640), .ZN(n7951) );
  NOR2_X1 U8434 ( .A1(n7913), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7933) );
  OR2_X1 U8435 ( .A1(n7898), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7913) );
  INV_X1 U8436 ( .A(n12390), .ZN(n12482) );
  NOR2_X1 U8437 ( .A1(n6677), .A2(n7589), .ZN(n7588) );
  OR2_X1 U8438 ( .A1(n7839), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7864) );
  OR2_X1 U8439 ( .A1(n7822), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7839) );
  INV_X1 U8440 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U8441 ( .A1(n7602), .A2(n8125), .ZN(n15321) );
  AND3_X1 U8442 ( .A1(n7821), .A2(n7820), .A3(n7819), .ZN(n15330) );
  INV_X1 U8443 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11600) );
  AND2_X1 U8444 ( .A1(n7786), .A2(n11600), .ZN(n7803) );
  AND3_X1 U8445 ( .A1(n7800), .A2(n7799), .A3(n7798), .ZN(n15347) );
  OR2_X1 U8446 ( .A1(n7753), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U8447 ( .A1(n11224), .A2(n12437), .ZN(n11411) );
  NAND2_X1 U8448 ( .A1(n11411), .A2(n12382), .ZN(n11410) );
  NAND2_X1 U8449 ( .A1(n11097), .A2(n7735), .ZN(n11225) );
  INV_X1 U8450 ( .A(n11228), .ZN(n12435) );
  NAND2_X1 U8451 ( .A1(n11225), .A2(n12435), .ZN(n11224) );
  INV_X1 U8452 ( .A(n12718), .ZN(n11342) );
  NAND2_X1 U8453 ( .A1(n8160), .A2(n8206), .ZN(n15385) );
  OR2_X1 U8454 ( .A1(n8008), .A2(n10469), .ZN(n7703) );
  OR2_X1 U8455 ( .A1(n7729), .A2(n7498), .ZN(n6807) );
  OR2_X1 U8456 ( .A1(n7683), .A2(n11041), .ZN(n7704) );
  NAND2_X1 U8457 ( .A1(n8058), .A2(n8057), .ZN(n12655) );
  NAND2_X1 U8458 ( .A1(n13286), .A2(n12491), .ZN(n13015) );
  NAND2_X1 U8459 ( .A1(n7964), .A2(n7963), .ZN(n13350) );
  OR2_X1 U8460 ( .A1(n15385), .A2(n15426), .ZN(n15411) );
  INV_X1 U8461 ( .A(n15346), .ZN(n15410) );
  INV_X1 U8462 ( .A(n7673), .ZN(n6718) );
  NAND2_X1 U8463 ( .A1(n7410), .A2(n7409), .ZN(n12367) );
  AOI21_X1 U8464 ( .B1(n7411), .B2(n7415), .A(n6573), .ZN(n7409) );
  AOI21_X1 U8465 ( .B1(n7416), .B2(n7414), .A(n6701), .ZN(n7413) );
  INV_X1 U8466 ( .A(n7416), .ZN(n7415) );
  OR2_X1 U8467 ( .A1(n8068), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U8468 ( .A1(n8067), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6738) );
  XNOR2_X1 U8469 ( .A(n8068), .B(n12602), .ZN(n8067) );
  NAND2_X1 U8470 ( .A1(n6755), .A2(n7973), .ZN(n7989) );
  NAND2_X1 U8471 ( .A1(n7972), .A2(n7971), .ZN(n6755) );
  NAND2_X1 U8472 ( .A1(n7958), .A2(n7957), .ZN(n7972) );
  AND2_X1 U8473 ( .A1(n7905), .A2(n7891), .ZN(n7892) );
  INV_X1 U8474 ( .A(n7434), .ZN(n7433) );
  AOI21_X1 U8475 ( .B1(n7434), .B2(n7432), .A(n6641), .ZN(n7431) );
  INV_X1 U8476 ( .A(n7828), .ZN(n7432) );
  INV_X1 U8477 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7812) );
  XNOR2_X1 U8478 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7810) );
  NAND2_X1 U8479 ( .A1(n6752), .A2(n7682), .ZN(n7762) );
  NAND2_X1 U8480 ( .A1(n7425), .A2(n7681), .ZN(n7424) );
  XNOR2_X1 U8481 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7761) );
  CLKBUF_X1 U8482 ( .A(n7684), .Z(n7685) );
  NAND2_X1 U8483 ( .A1(n11039), .A2(n6788), .ZN(n6800) );
  XNOR2_X1 U8484 ( .A(n15209), .B(n8341), .ZN(n8322) );
  INV_X1 U8485 ( .A(n8825), .ZN(n7535) );
  INV_X1 U8486 ( .A(n13424), .ZN(n7533) );
  NOR2_X1 U8487 ( .A1(n6581), .A2(n7535), .ZN(n7532) );
  OR2_X1 U8488 ( .A1(n8440), .A2(n8439), .ZN(n8463) );
  XNOR2_X1 U8489 ( .A(n11712), .B(n8341), .ZN(n11239) );
  NAND2_X1 U8490 ( .A1(n6959), .A2(n6960), .ZN(n8682) );
  OR2_X1 U8491 ( .A1(n12349), .A2(n6962), .ZN(n6959) );
  OR2_X1 U8492 ( .A1(n8527), .A2(n13133), .ZN(n8565) );
  INV_X1 U8493 ( .A(n7538), .ZN(n7537) );
  AND2_X1 U8494 ( .A1(n8493), .A2(n8473), .ZN(n6946) );
  NOR2_X1 U8495 ( .A1(n8463), .A2(n8462), .ZN(n8502) );
  NOR2_X1 U8496 ( .A1(n8371), .A2(n8370), .ZN(n8393) );
  AND2_X1 U8497 ( .A1(n8585), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8614) );
  INV_X1 U8498 ( .A(n9585), .ZN(n9804) );
  NAND4_X1 U8499 ( .A1(n8319), .A2(n8318), .A3(n8317), .A4(n8316), .ZN(n13548)
         );
  NAND2_X1 U8500 ( .A1(n8314), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8275) );
  NOR2_X1 U8501 ( .A1(n15049), .A2(n15050), .ZN(n15048) );
  NOR2_X1 U8502 ( .A1(n15071), .A2(n7176), .ZN(n15085) );
  AND2_X1 U8503 ( .A1(n15076), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7176) );
  NAND2_X1 U8504 ( .A1(n15085), .A2(n15084), .ZN(n15083) );
  NOR2_X1 U8505 ( .A1(n15068), .A2(n7391), .ZN(n15082) );
  AND2_X1 U8506 ( .A1(n15076), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7391) );
  NOR2_X1 U8507 ( .A1(n15080), .A2(n7390), .ZN(n13554) );
  AND2_X1 U8508 ( .A1(n15089), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7390) );
  NAND2_X1 U8509 ( .A1(n15083), .A2(n7175), .ZN(n13557) );
  OR2_X1 U8510 ( .A1(n15089), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7175) );
  NAND2_X1 U8511 ( .A1(n13557), .A2(n13556), .ZN(n13555) );
  OR2_X1 U8512 ( .A1(n13578), .A2(n13577), .ZN(n15097) );
  NOR2_X1 U8513 ( .A1(n15097), .A2(n15098), .ZN(n15096) );
  NOR2_X1 U8514 ( .A1(n15096), .A2(n13578), .ZN(n13579) );
  OR2_X1 U8515 ( .A1(n15122), .A2(n15121), .ZN(n15118) );
  AOI21_X1 U8516 ( .B1(n15125), .B2(P2_REG1_REG_16__SCAN_IN), .A(n15115), .ZN(
        n15137) );
  INV_X1 U8517 ( .A(n7396), .ZN(n13601) );
  AND2_X1 U8518 ( .A1(n6992), .A2(n13663), .ZN(n13618) );
  AND2_X1 U8519 ( .A1(n6994), .A2(n6993), .ZN(n6992) );
  NAND2_X1 U8520 ( .A1(n13618), .A2(n13880), .ZN(n13617) );
  NAND2_X1 U8521 ( .A1(n7270), .A2(n7273), .ZN(n13632) );
  AND2_X1 U8522 ( .A1(n7274), .A2(n13629), .ZN(n7273) );
  NOR2_X1 U8523 ( .A1(n7275), .A2(n7272), .ZN(n7271) );
  NAND2_X1 U8524 ( .A1(n13663), .A2(n6994), .ZN(n13638) );
  AND2_X1 U8525 ( .A1(n13656), .A2(n6604), .ZN(n7276) );
  NAND2_X1 U8526 ( .A1(n7253), .A2(n7252), .ZN(n13671) );
  AOI21_X1 U8527 ( .B1(n7255), .B2(n7259), .A(n6613), .ZN(n7252) );
  AOI21_X1 U8528 ( .B1(n7258), .B2(n7256), .A(n6631), .ZN(n7255) );
  NAND2_X1 U8529 ( .A1(n13663), .A2(n13668), .ZN(n13664) );
  AND2_X1 U8530 ( .A1(n9885), .A2(n9886), .ZN(n13669) );
  AND2_X1 U8531 ( .A1(n8630), .A2(n8224), .ZN(n8233) );
  NAND2_X1 U8532 ( .A1(n13756), .A2(n6983), .ZN(n13724) );
  NAND2_X1 U8533 ( .A1(n13756), .A2(n13899), .ZN(n13741) );
  NAND2_X1 U8534 ( .A1(n9872), .A2(n9871), .ZN(n13751) );
  AND2_X1 U8535 ( .A1(n9874), .A2(n9873), .ZN(n13754) );
  AND2_X1 U8536 ( .A1(n8672), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8694) );
  NOR2_X1 U8537 ( .A1(n8654), .A2(n8653), .ZN(n8672) );
  OR2_X1 U8538 ( .A1(n13857), .A2(n9867), .ZN(n6845) );
  NAND2_X1 U8539 ( .A1(n13771), .A2(n9945), .ZN(n13772) );
  NAND2_X1 U8540 ( .A1(n6989), .A2(n11923), .ZN(n13785) );
  NAND2_X1 U8541 ( .A1(n8614), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8635) );
  AND2_X1 U8542 ( .A1(n9925), .A2(n7288), .ZN(n7287) );
  INV_X1 U8543 ( .A(n12142), .ZN(n7288) );
  NAND2_X1 U8544 ( .A1(n11923), .A2(n9944), .ZN(n12135) );
  AOI21_X1 U8545 ( .B1(n11846), .B2(n11847), .A(n9918), .ZN(n12013) );
  NAND2_X1 U8546 ( .A1(n9915), .A2(n9914), .ZN(n11791) );
  NOR2_X1 U8547 ( .A1(n11887), .A2(n11781), .ZN(n11853) );
  NAND2_X1 U8548 ( .A1(n6968), .A2(n6967), .ZN(n11781) );
  INV_X1 U8549 ( .A(n11496), .ZN(n6968) );
  XNOR2_X1 U8550 ( .A(n11443), .B(n9851), .ZN(n11347) );
  NAND2_X1 U8551 ( .A1(n11083), .A2(n7282), .ZN(n11158) );
  NOR2_X1 U8552 ( .A1(n11160), .A2(n7283), .ZN(n7282) );
  INV_X1 U8553 ( .A(n9910), .ZN(n7283) );
  NOR2_X1 U8554 ( .A1(n11086), .A2(n15146), .ZN(n11164) );
  NAND2_X1 U8555 ( .A1(n11164), .A2(n11168), .ZN(n11351) );
  NAND2_X1 U8556 ( .A1(n11085), .A2(n11084), .ZN(n11083) );
  OAI21_X1 U8557 ( .B1(n11266), .B2(n9909), .A(n9908), .ZN(n10925) );
  CLKBUF_X1 U8558 ( .A(n11569), .Z(n6879) );
  NAND2_X1 U8559 ( .A1(n9899), .A2(n9898), .ZN(n11677) );
  NAND2_X1 U8560 ( .A1(n10953), .A2(n7386), .ZN(n9899) );
  XNOR2_X1 U8561 ( .A(n13549), .B(n11684), .ZN(n11676) );
  INV_X1 U8562 ( .A(n11676), .ZN(n11672) );
  NOR2_X1 U8563 ( .A1(n9589), .A2(n9588), .ZN(n15158) );
  AND3_X1 U8564 ( .A1(n13684), .A2(n13742), .A3(n13683), .ZN(n13820) );
  INV_X1 U8565 ( .A(n15212), .ZN(n13861) );
  AND2_X1 U8566 ( .A1(n10766), .A2(n9773), .ZN(n15200) );
  XNOR2_X1 U8567 ( .A(n9585), .B(n9586), .ZN(n8236) );
  AND2_X1 U8568 ( .A1(n12258), .A2(n8867), .ZN(n15175) );
  AND2_X1 U8569 ( .A1(n10530), .A2(n10531), .ZN(n8903) );
  AOI21_X1 U8570 ( .B1(n8262), .B2(n8261), .A(n6644), .ZN(n6938) );
  NAND2_X1 U8571 ( .A1(n6880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8244) );
  AND2_X1 U8572 ( .A1(n6608), .A2(n6965), .ZN(n6964) );
  NOR2_X1 U8573 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6965) );
  AND2_X1 U8574 ( .A1(n8460), .A2(n8496), .ZN(n11960) );
  AND2_X1 U8575 ( .A1(n8436), .A2(n8459), .ZN(n10966) );
  INV_X1 U8576 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n13134) );
  NOR2_X1 U8577 ( .A1(n13941), .A2(n7469), .ZN(n7468) );
  INV_X1 U8578 ( .A(n10282), .ZN(n7469) );
  AND2_X1 U8579 ( .A1(n14029), .A2(n10359), .ZN(n13954) );
  AOI21_X1 U8580 ( .B1(n7485), .B2(n10238), .A(n7482), .ZN(n7481) );
  NOR2_X1 U8581 ( .A1(n10244), .A2(n10245), .ZN(n7482) );
  CLKBUF_X1 U8582 ( .A(n14000), .Z(n14019) );
  AND2_X1 U8583 ( .A1(n10384), .A2(n10369), .ZN(n14027) );
  NAND2_X1 U8584 ( .A1(n7465), .A2(n6616), .ZN(n13953) );
  NAND2_X1 U8585 ( .A1(n13981), .A2(n14058), .ZN(n7466) );
  NAND2_X1 U8586 ( .A1(n7467), .A2(n10340), .ZN(n14059) );
  INV_X1 U8587 ( .A(n9316), .ZN(n9317) );
  NAND2_X1 U8588 ( .A1(n13938), .A2(n10291), .ZN(n10294) );
  AND4_X1 U8589 ( .A1(n9117), .A2(n9116), .A3(n9115), .A4(n9114), .ZN(n11737)
         );
  AND4_X1 U8590 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(n11528)
         );
  OR2_X1 U8591 ( .A1(n9017), .A2(n8939), .ZN(n8942) );
  OR2_X1 U8592 ( .A1(n9015), .A2(n8940), .ZN(n8941) );
  OR2_X1 U8593 ( .A1(n10623), .A2(n10622), .ZN(n6927) );
  OR2_X1 U8594 ( .A1(n10645), .A2(n10644), .ZN(n6925) );
  AND2_X1 U8595 ( .A1(n6925), .A2(n6924), .ZN(n10711) );
  NAND2_X1 U8596 ( .A1(n10709), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U8597 ( .A1(n11115), .A2(n6931), .ZN(n11120) );
  AND2_X1 U8598 ( .A1(n11116), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6931) );
  NOR2_X1 U8599 ( .A1(n11120), .A2(n11119), .ZN(n11426) );
  NOR2_X1 U8600 ( .A1(n11895), .A2(n6934), .ZN(n11900) );
  AND2_X1 U8601 ( .A1(n11896), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6934) );
  NOR2_X1 U8602 ( .A1(n11900), .A2(n11899), .ZN(n12055) );
  XNOR2_X1 U8603 ( .A(n14198), .B(n14208), .ZN(n12056) );
  NOR2_X1 U8604 ( .A1(n12055), .A2(n6933), .ZN(n14198) );
  AND2_X1 U8605 ( .A1(n12062), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6933) );
  AOI21_X1 U8606 ( .B1(n14874), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14865), .ZN(
        n14880) );
  NOR2_X1 U8607 ( .A1(n14901), .A2(n14900), .ZN(n14899) );
  OR2_X1 U8608 ( .A1(n14243), .A2(n14110), .ZN(n7626) );
  OR2_X1 U8609 ( .A1(n14094), .A2(n14112), .ZN(n7620) );
  OAI21_X1 U8610 ( .B1(n7568), .B2(n7565), .A(n7621), .ZN(n7564) );
  NAND2_X1 U8611 ( .A1(n14311), .A2(n14293), .ZN(n14292) );
  OR2_X1 U8612 ( .A1(n14472), .A2(n14342), .ZN(n14331) );
  INV_X1 U8613 ( .A(n9329), .ZN(n9330) );
  AOI21_X1 U8614 ( .B1(n14386), .B2(n6595), .A(n7580), .ZN(n14338) );
  NAND2_X1 U8615 ( .A1(n7581), .A2(n6611), .ZN(n7580) );
  INV_X1 U8616 ( .A(n9305), .ZN(n9306) );
  AOI21_X1 U8617 ( .B1(n6548), .B2(n12166), .A(n6634), .ZN(n7585) );
  NAND2_X1 U8618 ( .A1(n9250), .A2(n9249), .ZN(n9269) );
  AND4_X1 U8619 ( .A1(n9275), .A2(n9274), .A3(n9273), .A4(n9272), .ZN(n14010)
         );
  NOR2_X1 U8620 ( .A1(n12168), .A2(n7192), .ZN(n14423) );
  INV_X1 U8621 ( .A(n7194), .ZN(n7192) );
  OR2_X1 U8622 ( .A1(n14104), .A2(n12078), .ZN(n12168) );
  NOR2_X1 U8623 ( .A1(n9185), .A2(n9177), .ZN(n9210) );
  INV_X1 U8624 ( .A(n10048), .ZN(n7549) );
  NAND2_X1 U8625 ( .A1(n11974), .A2(n11972), .ZN(n7550) );
  NAND3_X1 U8626 ( .A1(n7188), .A2(n11530), .A3(n13999), .ZN(n11990) );
  AND2_X1 U8627 ( .A1(n7188), .A2(n11530), .ZN(n11991) );
  NAND2_X1 U8628 ( .A1(n11530), .A2(n7190), .ZN(n11775) );
  AND2_X1 U8629 ( .A1(n11516), .A2(n11548), .ZN(n11530) );
  NAND2_X1 U8630 ( .A1(n11530), .A2(n15017), .ZN(n11774) );
  NOR2_X1 U8631 ( .A1(n14928), .A2(n15006), .ZN(n11516) );
  AOI21_X1 U8632 ( .B1(n11387), .B2(n7560), .A(n7559), .ZN(n7558) );
  OR2_X1 U8633 ( .A1(n14927), .A2(n11658), .ZN(n14928) );
  INV_X1 U8634 ( .A(n10034), .ZN(n14916) );
  NAND2_X1 U8635 ( .A1(n10033), .A2(n10032), .ZN(n11386) );
  NAND2_X1 U8636 ( .A1(n11386), .A2(n11387), .ZN(n11385) );
  AND2_X1 U8637 ( .A1(n14949), .A2(n14988), .ZN(n14951) );
  NAND2_X1 U8638 ( .A1(n11720), .A2(n14964), .ZN(n11721) );
  OR2_X1 U8639 ( .A1(n10070), .A2(n14151), .ZN(n14268) );
  AND2_X1 U8640 ( .A1(n6792), .A2(n6600), .ZN(n14289) );
  NAND2_X1 U8641 ( .A1(n7587), .A2(n6548), .ZN(n14421) );
  OR2_X1 U8642 ( .A1(n12159), .A2(n12166), .ZN(n7587) );
  AND2_X1 U8643 ( .A1(n9046), .A2(n9045), .ZN(n14999) );
  NAND2_X1 U8644 ( .A1(n10685), .A2(n14677), .ZN(n14979) );
  INV_X1 U8645 ( .A(n8920), .ZN(n8919) );
  INV_X1 U8646 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8921) );
  XNOR2_X1 U8647 ( .A(n9434), .B(n9433), .ZN(n12332) );
  NAND2_X1 U8648 ( .A1(n7098), .A2(n9424), .ZN(n9434) );
  NAND2_X1 U8649 ( .A1(n7104), .A2(n7102), .ZN(n7098) );
  XNOR2_X1 U8650 ( .A(n8887), .B(n8831), .ZN(n13925) );
  XNOR2_X1 U8651 ( .A(n8827), .B(n8809), .ZN(n12255) );
  NAND2_X1 U8652 ( .A1(n9513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U8653 ( .A1(n8748), .A2(SI_22_), .ZN(n8765) );
  INV_X1 U8654 ( .A(n8747), .ZN(n6868) );
  XNOR2_X1 U8655 ( .A(n7506), .B(n8668), .ZN(n9256) );
  OAI21_X1 U8656 ( .B1(n8664), .B2(n8684), .A(n8665), .ZN(n7506) );
  NAND2_X1 U8657 ( .A1(n8626), .A2(n8625), .ZN(n8648) );
  INV_X1 U8658 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9169) );
  NAND2_X1 U8659 ( .A1(n8495), .A2(n8494), .ZN(n8512) );
  OAI21_X1 U8660 ( .B1(n9202), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9144) );
  AOI21_X1 U8661 ( .B1(n7503), .B2(n7505), .A(n7501), .ZN(n7500) );
  INV_X1 U8662 ( .A(n8426), .ZN(n7501) );
  OR2_X1 U8663 ( .A1(n9087), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U8664 ( .A1(n8406), .A2(n8405), .ZN(n8425) );
  NAND2_X1 U8665 ( .A1(n8387), .A2(n8386), .ZN(n8406) );
  OR2_X1 U8666 ( .A1(n8979), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9008) );
  INV_X1 U8667 ( .A(n8288), .ZN(n8285) );
  NAND2_X1 U8668 ( .A1(n8282), .A2(n7499), .ZN(n8253) );
  AND2_X1 U8669 ( .A1(n7118), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14597) );
  INV_X1 U8670 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7118) );
  INV_X1 U8671 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15258) );
  XNOR2_X1 U8672 ( .A(n14592), .B(n14593), .ZN(n14606) );
  NAND2_X1 U8673 ( .A1(n7127), .A2(n7124), .ZN(n14592) );
  AND2_X1 U8674 ( .A1(n6730), .A2(n6647), .ZN(n14614) );
  OR2_X1 U8675 ( .A1(n15443), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U8676 ( .A1(n14569), .A2(n14568), .ZN(n14612) );
  NAND2_X1 U8677 ( .A1(n14609), .A2(n14567), .ZN(n14568) );
  XNOR2_X1 U8678 ( .A(n14571), .B(n7141), .ZN(n14618) );
  INV_X1 U8679 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n7141) );
  AND2_X1 U8680 ( .A1(n14846), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U8681 ( .A1(n7322), .A2(n7319), .ZN(n12613) );
  INV_X1 U8682 ( .A(n7321), .ZN(n7319) );
  NAND2_X1 U8683 ( .A1(n7323), .A2(n6586), .ZN(n7322) );
  INV_X1 U8684 ( .A(n12639), .ZN(n7323) );
  NAND2_X1 U8685 ( .A1(n7342), .A2(n10153), .ZN(n12304) );
  OAI21_X1 U8686 ( .B1(n11336), .B2(n7348), .A(n7346), .ZN(n10108) );
  INV_X1 U8687 ( .A(n15310), .ZN(n15339) );
  NAND2_X1 U8688 ( .A1(n10869), .A2(n10090), .ZN(n10868) );
  AOI21_X1 U8689 ( .B1(n11936), .B2(n7354), .A(n6551), .ZN(n12236) );
  AOI21_X1 U8690 ( .B1(n12639), .B2(n12638), .A(n6582), .ZN(n12649) );
  AND2_X1 U8691 ( .A1(n8080), .A2(n8079), .ZN(n12949) );
  OAI22_X1 U8692 ( .A1(n6560), .A2(n10144), .B1(n12675), .B2(n7332), .ZN(
        n12660) );
  NAND2_X1 U8693 ( .A1(n7334), .A2(n12625), .ZN(n7332) );
  OR2_X1 U8694 ( .A1(n11910), .A2(n11911), .ZN(n11935) );
  NAND2_X1 U8695 ( .A1(n7316), .A2(n7317), .ZN(n12666) );
  AOI21_X1 U8696 ( .B1(n7320), .B2(n7318), .A(n6635), .ZN(n7317) );
  OR2_X1 U8697 ( .A1(n10173), .A2(n10172), .ZN(n12685) );
  NAND2_X1 U8698 ( .A1(n7324), .A2(n7328), .ZN(n12683) );
  NAND2_X1 U8699 ( .A1(n12639), .A2(n7330), .ZN(n7324) );
  OR2_X1 U8700 ( .A1(n10173), .A2(n10170), .ZN(n12296) );
  NAND2_X1 U8701 ( .A1(n11336), .A2(n10103), .ZN(n11448) );
  INV_X1 U8702 ( .A(n12552), .ZN(n6711) );
  INV_X1 U8703 ( .A(n12934), .ZN(n12708) );
  INV_X1 U8704 ( .A(n12949), .ZN(n12920) );
  INV_X1 U8705 ( .A(n12976), .ZN(n12709) );
  NAND2_X1 U8706 ( .A1(n13408), .A2(n10415), .ZN(n12710) );
  CLKBUF_X1 U8707 ( .A(n12720), .Z(n6803) );
  NAND2_X1 U8708 ( .A1(n6547), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7706) );
  NAND2_X1 U8709 ( .A1(n6547), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7694) );
  OR2_X1 U8710 ( .A1(n7755), .A2(n11009), .ZN(n7693) );
  INV_X1 U8711 ( .A(n11040), .ZN(n15251) );
  INV_X1 U8712 ( .A(n11014), .ZN(n11192) );
  NAND2_X1 U8713 ( .A1(n12732), .A2(n7014), .ZN(n7013) );
  OR2_X1 U8714 ( .A1(n11134), .A2(n7014), .ZN(n12733) );
  NOR2_X1 U8715 ( .A1(n15266), .A2(n15267), .ZN(n15265) );
  NAND2_X1 U8716 ( .A1(n7245), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7244) );
  INV_X1 U8717 ( .A(n11589), .ZN(n7245) );
  NAND2_X1 U8718 ( .A1(n6695), .A2(n7296), .ZN(n11813) );
  OR2_X1 U8719 ( .A1(n11799), .A2(n15333), .ZN(n7232) );
  NAND2_X1 U8720 ( .A1(n7290), .A2(n12034), .ZN(n12757) );
  AND2_X1 U8721 ( .A1(n7007), .A2(n7009), .ZN(n12747) );
  XNOR2_X1 U8722 ( .A(n12766), .B(n12772), .ZN(n12743) );
  NOR2_X1 U8723 ( .A1(n12744), .A2(n12743), .ZN(n12769) );
  OR2_X1 U8724 ( .A1(n12758), .A2(n7883), .ZN(n7314) );
  INV_X1 U8725 ( .A(n12765), .ZN(n7313) );
  NAND2_X1 U8726 ( .A1(n7309), .A2(n7310), .ZN(n12809) );
  OR2_X1 U8727 ( .A1(n12814), .A2(n12813), .ZN(n12822) );
  NOR2_X1 U8728 ( .A1(n14702), .A2(n12812), .ZN(n12814) );
  NOR2_X1 U8729 ( .A1(n12791), .A2(n14697), .ZN(n12793) );
  XNOR2_X1 U8730 ( .A(n12859), .B(n12860), .ZN(n12823) );
  NOR2_X1 U8731 ( .A1(n12823), .A2(n12824), .ZN(n12861) );
  NAND2_X1 U8732 ( .A1(n7003), .A2(n12834), .ZN(n12838) );
  NOR2_X1 U8733 ( .A1(n12867), .A2(n6689), .ZN(n6902) );
  NAND2_X1 U8734 ( .A1(n11038), .A2(n11037), .ZN(n15304) );
  NOR2_X1 U8735 ( .A1(n12845), .A2(n12844), .ZN(n12848) );
  NAND2_X1 U8736 ( .A1(n12875), .A2(n12884), .ZN(n6783) );
  OR2_X1 U8737 ( .A1(n14719), .A2(n8163), .ZN(n12898) );
  AND2_X1 U8738 ( .A1(n12937), .A2(n12936), .ZN(n13314) );
  NAND2_X1 U8739 ( .A1(n12985), .A2(n8142), .ZN(n12973) );
  NAND2_X1 U8740 ( .A1(n8017), .A2(n12507), .ZN(n12977) );
  AND2_X1 U8741 ( .A1(n6839), .A2(n8141), .ZN(n12986) );
  NAND2_X1 U8742 ( .A1(n7949), .A2(n7948), .ZN(n13357) );
  NAND2_X1 U8743 ( .A1(n12280), .A2(n12485), .ZN(n13301) );
  NAND2_X1 U8744 ( .A1(n7598), .A2(n7596), .ZN(n13298) );
  NAND2_X1 U8745 ( .A1(n7912), .A2(n7911), .ZN(n13365) );
  OR2_X1 U8746 ( .A1(n11704), .A2(n15392), .ZN(n12250) );
  NAND2_X1 U8747 ( .A1(n7590), .A2(n7593), .ZN(n14726) );
  NAND2_X1 U8748 ( .A1(n15307), .A2(n8128), .ZN(n14736) );
  INV_X1 U8749 ( .A(n12250), .ZN(n15349) );
  AND3_X1 U8750 ( .A1(n7785), .A2(n7784), .A3(n7783), .ZN(n15409) );
  AND2_X1 U8751 ( .A1(n11227), .A2(n8118), .ZN(n11414) );
  AND2_X1 U8752 ( .A1(n11081), .A2(n12872), .ZN(n15392) );
  INV_X2 U8753 ( .A(n15396), .ZN(n15398) );
  AND2_X1 U8754 ( .A1(n15396), .A2(n15353), .ZN(n13306) );
  NAND2_X1 U8755 ( .A1(n15349), .A2(n15410), .ZN(n13304) );
  AND2_X1 U8756 ( .A1(n14747), .A2(n14746), .ZN(n14764) );
  AOI21_X1 U8757 ( .B1(n12285), .B2(n12370), .A(n9566), .ZN(n12894) );
  INV_X1 U8758 ( .A(n12301), .ZN(n12900) );
  AND2_X1 U8759 ( .A1(n8085), .A2(n8084), .ZN(n13372) );
  AND2_X1 U8760 ( .A1(n8010), .A2(n8009), .ZN(n13393) );
  NAND2_X1 U8761 ( .A1(n7997), .A2(n7996), .ZN(n13396) );
  AND2_X1 U8762 ( .A1(n8193), .A2(n8192), .ZN(n13407) );
  AND2_X1 U8763 ( .A1(n11023), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13408) );
  INV_X1 U8764 ( .A(n7667), .ZN(n12288) );
  XNOR2_X1 U8765 ( .A(n6746), .B(n7412), .ZN(n12285) );
  NAND2_X1 U8766 ( .A1(n6747), .A2(n7413), .ZN(n6746) );
  OR2_X1 U8767 ( .A1(n9530), .A2(n7415), .ZN(n6747) );
  CLKBUF_X1 U8768 ( .A(n8169), .Z(n13420) );
  NAND2_X1 U8769 ( .A1(n7417), .A2(n7418), .ZN(n9565) );
  NAND2_X1 U8770 ( .A1(n7441), .A2(n8035), .ZN(n8040) );
  XNOR2_X1 U8771 ( .A(n7643), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12555) );
  NAND2_X1 U8772 ( .A1(n8019), .A2(n8018), .ZN(n8033) );
  NAND2_X1 U8773 ( .A1(n8156), .A2(n8173), .ZN(n12350) );
  NAND2_X1 U8774 ( .A1(n7927), .A2(n7029), .ZN(n7648) );
  OR2_X1 U8775 ( .A1(n7930), .A2(n7929), .ZN(n12825) );
  AND2_X1 U8776 ( .A1(n7440), .A2(n7923), .ZN(n7926) );
  NAND2_X1 U8777 ( .A1(n7440), .A2(n6672), .ZN(n7940) );
  OR2_X1 U8778 ( .A1(n7922), .A2(n7921), .ZN(n7440) );
  NAND2_X1 U8779 ( .A1(n7889), .A2(n7874), .ZN(n7442) );
  NAND2_X1 U8780 ( .A1(n7423), .A2(n7681), .ZN(n7745) );
  NAND2_X1 U8781 ( .A1(n7428), .A2(n7427), .ZN(n7423) );
  INV_X1 U8782 ( .A(n7425), .ZN(n7427) );
  NAND2_X1 U8783 ( .A1(n7428), .A2(n7680), .ZN(n7728) );
  NAND2_X1 U8784 ( .A1(n13505), .A2(n8825), .ZN(n13425) );
  AND2_X1 U8785 ( .A1(n8844), .A2(n8836), .ZN(n13652) );
  NOR2_X1 U8786 ( .A1(n12314), .A2(n8572), .ZN(n6939) );
  INV_X1 U8787 ( .A(n11926), .ZN(n14776) );
  NAND2_X1 U8788 ( .A1(n11246), .A2(n8473), .ZN(n11647) );
  INV_X1 U8789 ( .A(n6952), .ZN(n6951) );
  OAI21_X1 U8790 ( .B1(n6954), .B2(n8853), .A(n6953), .ZN(n6952) );
  NAND2_X1 U8791 ( .A1(n8890), .A2(n8853), .ZN(n6953) );
  OAI21_X1 U8792 ( .B1(n6954), .B2(n6955), .A(n6950), .ZN(n6949) );
  NAND2_X1 U8793 ( .A1(n8890), .A2(n6955), .ZN(n6950) );
  NAND2_X1 U8794 ( .A1(n7529), .A2(n13518), .ZN(n7528) );
  NAND2_X1 U8795 ( .A1(n10937), .A2(n8404), .ZN(n6944) );
  NAND2_X1 U8796 ( .A1(n13475), .A2(n8706), .ZN(n13448) );
  INV_X1 U8797 ( .A(n7525), .ZN(n7524) );
  NAND2_X1 U8798 ( .A1(n7526), .A2(n8763), .ZN(n13465) );
  NAND2_X1 U8799 ( .A1(n13432), .A2(n13431), .ZN(n7526) );
  INV_X1 U8800 ( .A(n10789), .ZN(n8324) );
  CLKBUF_X1 U8801 ( .A(n10826), .Z(n10915) );
  NAND2_X1 U8802 ( .A1(n8682), .A2(n13439), .ZN(n13477) );
  NAND2_X1 U8803 ( .A1(n8546), .A2(n8545), .ZN(n14782) );
  INV_X1 U8804 ( .A(n13513), .ZN(n13491) );
  NAND2_X1 U8805 ( .A1(n12349), .A2(n6590), .ZN(n13498) );
  NAND2_X1 U8806 ( .A1(n12349), .A2(n8643), .ZN(n13497) );
  NAND2_X1 U8807 ( .A1(n10923), .A2(n8381), .ZN(n10938) );
  NAND2_X1 U8808 ( .A1(n8805), .A2(n8804), .ZN(n13508) );
  XNOR2_X1 U8809 ( .A(n8593), .B(n8592), .ZN(n12108) );
  AND2_X1 U8810 ( .A1(n9802), .A2(n9801), .ZN(n9803) );
  INV_X1 U8811 ( .A(n9586), .ZN(n9811) );
  CLKBUF_X1 U8812 ( .A(n13548), .Z(n6898) );
  NAND2_X1 U8813 ( .A1(n8315), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8267) );
  OR2_X1 U8814 ( .A1(n10553), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8815 ( .A1(n10553), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6890) );
  NOR2_X1 U8816 ( .A1(n15046), .A2(n7401), .ZN(n15059) );
  NOR2_X1 U8817 ( .A1(n10553), .A2(n15243), .ZN(n7401) );
  NOR2_X1 U8818 ( .A1(n10564), .A2(n6625), .ZN(n10586) );
  INV_X1 U8819 ( .A(n7178), .ZN(n10584) );
  NOR2_X1 U8820 ( .A1(n10570), .A2(n10569), .ZN(n10664) );
  AND2_X1 U8821 ( .A1(n7178), .A2(n7177), .ZN(n10570) );
  NAND2_X1 U8822 ( .A1(n10574), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7177) );
  AOI21_X1 U8823 ( .B1(n10574), .B2(P2_REG1_REG_4__SCAN_IN), .A(n10587), .ZN(
        n10577) );
  NOR2_X1 U8824 ( .A1(n10849), .A2(n7393), .ZN(n10853) );
  AND2_X1 U8825 ( .A1(n10850), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7393) );
  NOR2_X1 U8826 ( .A1(n10844), .A2(n7180), .ZN(n10848) );
  AND2_X1 U8827 ( .A1(n10850), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7180) );
  NOR2_X1 U8828 ( .A1(n10848), .A2(n10847), .ZN(n10959) );
  NOR2_X1 U8829 ( .A1(n10959), .A2(n7179), .ZN(n10963) );
  AND2_X1 U8830 ( .A1(n10966), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8831 ( .A1(n10963), .A2(n10962), .ZN(n11948) );
  XNOR2_X1 U8832 ( .A(n13579), .B(n13580), .ZN(n15106) );
  NOR2_X1 U8833 ( .A1(n15106), .A2(n15105), .ZN(n15104) );
  NOR2_X1 U8834 ( .A1(n15107), .A2(n13568), .ZN(n15117) );
  INV_X1 U8835 ( .A(n7395), .ZN(n13571) );
  OAI21_X1 U8836 ( .B1(n15144), .B2(n13610), .A(n13609), .ZN(n7404) );
  AND2_X1 U8837 ( .A1(n7277), .A2(n6604), .ZN(n13657) );
  NAND2_X1 U8838 ( .A1(n7254), .A2(n7258), .ZN(n13675) );
  NAND2_X1 U8839 ( .A1(n13711), .A2(n7261), .ZN(n7254) );
  NAND2_X1 U8840 ( .A1(n13692), .A2(n9882), .ZN(n13678) );
  NAND2_X1 U8841 ( .A1(n7257), .A2(n7263), .ZN(n13691) );
  OR2_X1 U8842 ( .A1(n13711), .A2(n9934), .ZN(n7257) );
  INV_X1 U8843 ( .A(n13891), .ZN(n13703) );
  AND2_X1 U8844 ( .A1(n7266), .A2(n6606), .ZN(n13731) );
  NAND2_X1 U8845 ( .A1(n9932), .A2(n9931), .ZN(n13735) );
  NAND2_X1 U8846 ( .A1(n13789), .A2(n9928), .ZN(n13765) );
  NAND2_X1 U8847 ( .A1(n12191), .A2(n9927), .ZN(n13791) );
  NAND2_X1 U8848 ( .A1(n7289), .A2(n9925), .ZN(n12143) );
  NAND2_X1 U8849 ( .A1(n7289), .A2(n7287), .ZN(n13871) );
  NAND2_X1 U8850 ( .A1(n11784), .A2(n9855), .ZN(n11848) );
  OAI21_X1 U8851 ( .B1(n6849), .B2(n7370), .A(n7368), .ZN(n11494) );
  AND2_X1 U8852 ( .A1(n7388), .A2(n6601), .ZN(n11161) );
  NAND2_X1 U8853 ( .A1(n10927), .A2(n9848), .ZN(n11088) );
  OR2_X1 U8854 ( .A1(n15174), .A2(n11253), .ZN(n15152) );
  INV_X1 U8855 ( .A(n15163), .ZN(n13774) );
  INV_X1 U8856 ( .A(n15152), .ZN(n15170) );
  INV_X1 U8857 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6912) );
  AND2_X1 U8858 ( .A1(n8903), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15187) );
  INV_X1 U8859 ( .A(n8266), .ZN(n13917) );
  OAI211_X1 U8860 ( .C1(P2_IR_REG_27__SCAN_IN), .C2(P2_IR_REG_31__SCAN_IN), 
        .A(n8245), .B(n6972), .ZN(n13926) );
  OR2_X1 U8861 ( .A1(n8244), .A2(n6976), .ZN(n6972) );
  INV_X1 U8862 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n13109) );
  INV_X1 U8863 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10908) );
  INV_X1 U8864 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10517) );
  INV_X1 U8865 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10500) );
  INV_X1 U8866 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10491) );
  AND2_X1 U8867 ( .A1(n8366), .A2(n8365), .ZN(n10670) );
  INV_X1 U8868 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10459) );
  NAND2_X1 U8869 ( .A1(n8519), .A2(n6819), .ZN(n6818) );
  NAND2_X1 U8870 ( .A1(n8290), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n6820) );
  NAND2_X1 U8872 ( .A1(n10283), .A2(n10282), .ZN(n13940) );
  CLKBUF_X1 U8873 ( .A(n12148), .Z(n6919) );
  AOI21_X1 U8874 ( .B1(n7473), .B2(n12577), .A(n12586), .ZN(n7472) );
  NAND2_X1 U8875 ( .A1(n7480), .A2(n7481), .ZN(n11872) );
  XNOR2_X1 U8876 ( .A(n10186), .B(n10193), .ZN(n10885) );
  NAND2_X1 U8877 ( .A1(n10298), .A2(n10297), .ZN(n14002) );
  NAND2_X1 U8878 ( .A1(n9236), .A2(n9235), .ZN(n14804) );
  INV_X1 U8879 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n11284) );
  INV_X1 U8880 ( .A(n10232), .ZN(n11283) );
  NAND2_X1 U8881 ( .A1(n10314), .A2(n14016), .ZN(n14015) );
  INV_X1 U8882 ( .A(n6864), .ZN(n11313) );
  CLKBUF_X1 U8883 ( .A(n12002), .Z(n12004) );
  NAND2_X1 U8884 ( .A1(n13972), .A2(n10329), .ZN(n14035) );
  CLKBUF_X1 U8885 ( .A(n13953), .Z(n14061) );
  NAND2_X1 U8886 ( .A1(n12146), .A2(n10262), .ZN(n12203) );
  CLKBUF_X1 U8887 ( .A(n10777), .Z(n10778) );
  INV_X1 U8888 ( .A(n14073), .ZN(n14097) );
  NAND2_X1 U8889 ( .A1(n10232), .A2(n11280), .ZN(n6842) );
  OAI21_X1 U8890 ( .B1(n10232), .B2(n11280), .A(n11281), .ZN(n10233) );
  AND2_X1 U8891 ( .A1(n10513), .A2(n14151), .ZN(n14052) );
  INV_X1 U8892 ( .A(n9499), .ZN(n9500) );
  NOR3_X1 U8893 ( .A1(n9503), .A2(n9502), .A3(n9501), .ZN(n9509) );
  AND4_X1 U8894 ( .A1(n9216), .A2(n9215), .A3(n9214), .A4(n9213), .ZN(n12161)
         );
  INV_X1 U8895 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11127) );
  NAND4_X1 U8896 ( .A1(n8977), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n14135)
         );
  OR2_X1 U8897 ( .A1(n9032), .A2(n11331), .ZN(n8956) );
  OR2_X1 U8898 ( .A1(n9417), .A2(n10192), .ZN(n8928) );
  NOR2_X1 U8899 ( .A1(n14188), .A2(n6620), .ZN(n10658) );
  INV_X1 U8900 ( .A(n6929), .ZN(n10656) );
  AOI21_X1 U8901 ( .B1(n10613), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14184), .ZN(
        n10651) );
  NOR2_X1 U8902 ( .A1(n10606), .A2(n10605), .ZN(n10621) );
  AND2_X1 U8903 ( .A1(n6929), .A2(n6928), .ZN(n10606) );
  NAND2_X1 U8904 ( .A1(n10653), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6928) );
  INV_X1 U8905 ( .A(n6927), .ZN(n10640) );
  AOI21_X1 U8906 ( .B1(n10625), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10624), .ZN(
        n10627) );
  AND2_X1 U8907 ( .A1(n6927), .A2(n6926), .ZN(n10645) );
  NAND2_X1 U8908 ( .A1(n10641), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6926) );
  INV_X1 U8909 ( .A(n6925), .ZN(n10708) );
  AOI21_X1 U8910 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10641), .A(n10635), .ZN(
        n10638) );
  NOR2_X1 U8911 ( .A1(n10806), .A2(n6932), .ZN(n10810) );
  AND2_X1 U8912 ( .A1(n10813), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6932) );
  NOR2_X1 U8913 ( .A1(n10810), .A2(n10809), .ZN(n11115) );
  AOI21_X1 U8914 ( .B1(n11116), .B2(P1_REG1_REG_10__SCAN_IN), .A(n11109), .ZN(
        n11112) );
  NAND2_X1 U8915 ( .A1(n11424), .A2(n11425), .ZN(n11621) );
  NAND2_X1 U8916 ( .A1(n11621), .A2(n6873), .ZN(n11623) );
  OR2_X1 U8917 ( .A1(n11622), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6873) );
  AOI21_X1 U8918 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n11896), .A(n11890), .ZN(
        n11893) );
  INV_X1 U8919 ( .A(n14868), .ZN(n14903) );
  AOI22_X1 U8920 ( .A1(n14537), .A2(n9466), .B1(P2_DATAO_REG_31__SCAN_IN), 
        .B2(n9465), .ZN(n14435) );
  NAND2_X1 U8921 ( .A1(n9438), .A2(n9437), .ZN(n14231) );
  NOR2_X1 U8922 ( .A1(n14303), .A2(n10061), .ZN(n14283) );
  NAND2_X1 U8923 ( .A1(n7567), .A2(n7566), .ZN(n14284) );
  NAND2_X1 U8924 ( .A1(n9998), .A2(n9997), .ZN(n14328) );
  NAND2_X1 U8925 ( .A1(n14369), .A2(n10057), .ZN(n14356) );
  NAND2_X1 U8926 ( .A1(n14372), .A2(n9995), .ZN(n14354) );
  NAND2_X1 U8927 ( .A1(n14386), .A2(n10056), .ZN(n14367) );
  MUX2_X1 U8928 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8966), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n8967) );
  NAND2_X1 U8929 ( .A1(n7206), .A2(n9989), .ZN(n14403) );
  OR2_X1 U8930 ( .A1(n14420), .A2(n9990), .ZN(n7206) );
  NAND2_X1 U8931 ( .A1(n12085), .A2(n9985), .ZN(n12119) );
  NAND2_X1 U8932 ( .A1(n9168), .A2(n9466), .ZN(n9175) );
  NAND2_X1 U8933 ( .A1(n9163), .A2(n9162), .ZN(n14679) );
  NAND2_X1 U8934 ( .A1(n7205), .A2(n9980), .ZN(n11744) );
  NAND2_X1 U8935 ( .A1(n11525), .A2(n10039), .ZN(n11768) );
  NAND2_X1 U8936 ( .A1(n11507), .A2(n7574), .ZN(n11403) );
  NAND2_X1 U8937 ( .A1(n11507), .A2(n10036), .ZN(n11400) );
  OR2_X1 U8938 ( .A1(n10075), .A2(n14415), .ZN(n14334) );
  INV_X1 U8939 ( .A(n14432), .ZN(n14954) );
  INV_X1 U8940 ( .A(n14944), .ZN(n14417) );
  INV_X1 U8941 ( .A(n14942), .ZN(n14427) );
  INV_X1 U8942 ( .A(n15045), .ZN(n15043) );
  AND2_X1 U8943 ( .A1(n14444), .A2(n6884), .ZN(n6883) );
  NOR2_X1 U8944 ( .A1(n6885), .A2(n14439), .ZN(n6884) );
  OR2_X1 U8945 ( .A1(n14471), .A2(n14470), .ZN(n14521) );
  NAND2_X1 U8946 ( .A1(n8919), .A2(n8921), .ZN(n14534) );
  INV_X1 U8947 ( .A(n8925), .ZN(n14541) );
  NAND2_X1 U8948 ( .A1(n8933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U8949 ( .A1(n8918), .A2(n7579), .ZN(n8931) );
  XNOR2_X1 U8950 ( .A(n9518), .B(n9517), .ZN(n12257) );
  NAND2_X1 U8951 ( .A1(n8918), .A2(n7614), .ZN(n9516) );
  CLKBUF_X1 U8952 ( .A(n10005), .Z(n12604) );
  XNOR2_X1 U8953 ( .A(n9325), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14546) );
  NOR2_X1 U8954 ( .A1(n8969), .A2(n7490), .ZN(n9505) );
  INV_X1 U8955 ( .A(n9520), .ZN(n11824) );
  NOR2_X1 U8956 ( .A1(n8912), .A2(n8911), .ZN(n7542) );
  INV_X1 U8957 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10997) );
  INV_X1 U8958 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10893) );
  INV_X1 U8959 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11128) );
  INV_X1 U8960 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10909) );
  INV_X1 U8961 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n13062) );
  INV_X1 U8962 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10522) );
  INV_X1 U8963 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10518) );
  OR2_X1 U8964 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  INV_X1 U8965 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U8966 ( .A1(n8383), .A2(n8358), .ZN(n10488) );
  NAND2_X1 U8967 ( .A1(n8307), .A2(n8308), .ZN(n8327) );
  NAND2_X1 U8968 ( .A1(n6937), .A2(n6935), .ZN(n8959) );
  NAND2_X1 U8969 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6936), .ZN(n6935) );
  OAI21_X1 U8970 ( .B1(n8948), .B2(n8935), .A(P1_IR_REG_2__SCAN_IN), .ZN(n6937) );
  NAND2_X1 U8971 ( .A1(n8950), .A2(n8949), .ZN(n10608) );
  XNOR2_X1 U8972 ( .A(n14598), .B(n6914), .ZN(n15452) );
  INV_X1 U8973 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6914) );
  XNOR2_X1 U8974 ( .A(n14606), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15441) );
  XNOR2_X1 U8975 ( .A(n14614), .B(n7365), .ZN(n14665) );
  INV_X1 U8976 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7365) );
  XNOR2_X1 U8977 ( .A(n14617), .B(n14616), .ZN(n15447) );
  AND2_X1 U8978 ( .A1(n6729), .A2(n6655), .ZN(n14667) );
  INV_X1 U8979 ( .A(n14634), .ZN(n7114) );
  INV_X1 U8980 ( .A(n14645), .ZN(n7361) );
  NAND2_X1 U8981 ( .A1(n11449), .A2(n10105), .ZN(n11553) );
  OAI21_X1 U8982 ( .B1(n13368), .B2(n12706), .A(n10176), .ZN(n10177) );
  NAND2_X1 U8983 ( .A1(n10977), .A2(n10096), .ZN(n11151) );
  OAI21_X1 U8984 ( .B1(n6710), .B2(n12558), .A(n6708), .ZN(P3_U3296) );
  INV_X1 U8985 ( .A(n6709), .ZN(n6708) );
  OAI21_X1 U8986 ( .B1(n6892), .B2(n12558), .A(n7022), .ZN(n6709) );
  NAND2_X1 U8987 ( .A1(n7020), .A2(n15279), .ZN(n7019) );
  OAI211_X1 U8988 ( .C1(n12877), .C2(n6783), .A(n6781), .B(n6780), .ZN(n7018)
         );
  OAI22_X1 U8989 ( .A1(n13368), .A2(n13339), .B1(n15438), .B2(n8215), .ZN(
        n8216) );
  INV_X1 U8990 ( .A(n6887), .ZN(n6886) );
  OAI22_X1 U8991 ( .A1(n13368), .A2(n13392), .B1(n15430), .B2(n13367), .ZN(
        n6887) );
  INV_X1 U8992 ( .A(n7404), .ZN(n6888) );
  AOI21_X1 U8993 ( .B1(n13622), .B2(n15168), .A(n6805), .ZN(n6804) );
  NAND2_X1 U8994 ( .A1(n13623), .A2(n11353), .ZN(n6806) );
  INV_X1 U8995 ( .A(n13628), .ZN(n6805) );
  MUX2_X1 U8996 ( .A(n13798), .B(n13875), .S(n15250), .Z(n13799) );
  OAI21_X1 U8997 ( .B1(n6993), .B2(n13850), .A(n9956), .ZN(n9957) );
  AOI21_X1 U8998 ( .B1(n13643), .B2(n11886), .A(n6908), .ZN(n6907) );
  NAND2_X1 U8999 ( .A1(n13881), .A2(n15250), .ZN(n6909) );
  NOR2_X1 U9000 ( .A1(n15250), .A2(n13199), .ZN(n6908) );
  OAI21_X1 U9001 ( .B1(n13875), .B2(n15240), .A(n6986), .ZN(P2_U3498) );
  AOI21_X1 U9002 ( .B1(n13611), .B2(n11884), .A(n6987), .ZN(n6986) );
  NOR2_X1 U9003 ( .A1(n15242), .A2(n13876), .ZN(n6987) );
  NAND2_X1 U9004 ( .A1(n7269), .A2(n10406), .ZN(n7268) );
  AOI21_X1 U9005 ( .B1(n13623), .B2(n10406), .A(n6632), .ZN(n7387) );
  NAND2_X1 U9006 ( .A1(n13643), .A2(n11884), .ZN(n6893) );
  INV_X1 U9007 ( .A(n6835), .ZN(n6834) );
  OAI21_X1 U9008 ( .B1(n14259), .B2(n14093), .A(n13937), .ZN(n6835) );
  NAND2_X1 U9009 ( .A1(n6838), .A2(n6837), .ZN(P1_U3229) );
  AOI21_X1 U9010 ( .B1(n14314), .B2(n14103), .A(n14034), .ZN(n6837) );
  INV_X1 U9011 ( .A(n14033), .ZN(n6838) );
  NAND2_X1 U9012 ( .A1(n6878), .A2(n6875), .ZN(n14222) );
  NAND2_X1 U9013 ( .A1(n6877), .A2(n6876), .ZN(n6875) );
  OR2_X1 U9014 ( .A1(n10027), .A2(n14432), .ZN(n7624) );
  INV_X1 U9015 ( .A(n6856), .ZN(n14248) );
  OAI21_X1 U9016 ( .B1(n14449), .B2(n14432), .A(n6857), .ZN(n6856) );
  AOI21_X1 U9017 ( .B1(n14445), .B2(n14953), .A(n14247), .ZN(n6857) );
  AND2_X1 U9018 ( .A1(n6854), .A2(n6853), .ZN(n14264) );
  AOI21_X1 U9019 ( .B1(n14451), .B2(n14263), .A(n14262), .ZN(n6853) );
  OR2_X1 U9020 ( .A1(n14454), .A2(n14432), .ZN(n6854) );
  INV_X1 U9021 ( .A(n7116), .ZN(n14670) );
  NOR2_X1 U9022 ( .A1(n14847), .A2(n14846), .ZN(n14845) );
  OAI21_X1 U9023 ( .B1(n14689), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6915), .ZN(
        n6899) );
  CLKBUF_X3 U9024 ( .A(n8992), .Z(n9468) );
  AND2_X1 U9025 ( .A1(n6553), .A2(n10051), .ZN(n6548) );
  AND2_X1 U9026 ( .A1(n8182), .A2(n7659), .ZN(n8176) );
  AND3_X1 U9027 ( .A1(n9537), .A2(n8152), .A3(n7450), .ZN(n6549) );
  INV_X2 U9028 ( .A(n8247), .ZN(n8945) );
  AND2_X1 U9029 ( .A1(n14502), .A2(n14120), .ZN(n6550) );
  INV_X1 U9030 ( .A(n11508), .ZN(n7572) );
  INV_X1 U9031 ( .A(n12548), .ZN(n7075) );
  INV_X2 U9032 ( .A(n8547), .ZN(n8587) );
  INV_X1 U9033 ( .A(n12382), .ZN(n8119) );
  NOR2_X1 U9034 ( .A1(n10119), .A2(n15309), .ZN(n6551) );
  AND2_X1 U9035 ( .A1(n7654), .A2(n7030), .ZN(n6552) );
  XOR2_X1 U9036 ( .A(n14510), .B(n14072), .Z(n6553) );
  INV_X1 U9037 ( .A(n10042), .ZN(n11743) );
  AND2_X1 U9038 ( .A1(n11160), .A2(n6601), .ZN(n6554) );
  OR3_X1 U9039 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6555) );
  INV_X1 U9040 ( .A(n7259), .ZN(n7258) );
  OAI21_X1 U9041 ( .B1(n13693), .B2(n7260), .A(n9935), .ZN(n7259) );
  AND2_X1 U9042 ( .A1(n12945), .A2(n12938), .ZN(n6556) );
  AND2_X1 U9043 ( .A1(n9078), .A2(n7170), .ZN(n6557) );
  AND2_X1 U9044 ( .A1(n14531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6558) );
  INV_X1 U9045 ( .A(n7299), .ZN(n7298) );
  OAI21_X1 U9046 ( .B1(n7303), .B2(n7300), .A(n7301), .ZN(n7299) );
  AND2_X1 U9047 ( .A1(n13368), .A2(n7067), .ZN(n6559) );
  AND2_X1 U9048 ( .A1(n10141), .A2(n6680), .ZN(n6560) );
  NAND2_X1 U9049 ( .A1(n7494), .A2(n6662), .ZN(n6561) );
  AND2_X1 U9050 ( .A1(n9633), .A2(n9632), .ZN(n6562) );
  INV_X1 U9051 ( .A(n13464), .ZN(n7527) );
  OR2_X1 U9052 ( .A1(n9797), .A2(n9796), .ZN(n6563) );
  AND3_X1 U9053 ( .A1(n7610), .A2(n7659), .A3(n7676), .ZN(n6564) );
  AND2_X1 U9054 ( .A1(n9643), .A2(n9642), .ZN(n6565) );
  AND2_X1 U9055 ( .A1(n6505), .A2(n8125), .ZN(n6566) );
  AND2_X1 U9056 ( .A1(n9658), .A2(n9657), .ZN(n6567) );
  NAND2_X1 U9057 ( .A1(n9397), .A2(n7159), .ZN(n7158) );
  INV_X1 U9058 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13231) );
  INV_X1 U9059 ( .A(n11353), .ZN(n15174) );
  NAND2_X1 U9060 ( .A1(n8752), .A2(n8751), .ZN(n13713) );
  AND2_X1 U9061 ( .A1(n11923), .A2(n6991), .ZN(n6568) );
  OR2_X1 U9062 ( .A1(n12473), .A2(n12547), .ZN(n6569) );
  NAND2_X1 U9063 ( .A1(n7927), .A2(n6552), .ZN(n6570) );
  OR2_X1 U9064 ( .A1(n12107), .A2(n13742), .ZN(n6571) );
  NOR2_X1 U9065 ( .A1(n11609), .A2(n11829), .ZN(n6572) );
  INV_X1 U9066 ( .A(n12774), .ZN(n7312) );
  INV_X1 U9067 ( .A(n9531), .ZN(n7414) );
  AND2_X1 U9068 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n12333), .ZN(n6573) );
  OR2_X1 U9069 ( .A1(n11140), .A2(n11049), .ZN(n6574) );
  NAND2_X2 U9070 ( .A1(n7683), .A2(n10476), .ZN(n7729) );
  AND2_X2 U9071 ( .A1(n8945), .A2(n10533), .ZN(n8333) );
  NAND2_X1 U9072 ( .A1(n7714), .A2(n7679), .ZN(n7428) );
  AND2_X1 U9073 ( .A1(n8258), .A2(n8259), .ZN(n6575) );
  INV_X1 U9074 ( .A(n14299), .ZN(n7565) );
  NAND2_X1 U9075 ( .A1(n9744), .A2(n9743), .ZN(n13611) );
  INV_X1 U9076 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7359) );
  NAND3_X1 U9077 ( .A1(n7025), .A2(n7026), .A3(n7023), .ZN(n6576) );
  OR2_X1 U9078 ( .A1(n9471), .A2(n9470), .ZN(n6577) );
  AND3_X1 U9079 ( .A1(n11471), .A2(n9832), .A3(n7385), .ZN(n6578) );
  NAND2_X1 U9080 ( .A1(n8176), .A2(n7660), .ZN(n8178) );
  AND2_X1 U9081 ( .A1(n12673), .A2(n10141), .ZN(n6579) );
  OR2_X1 U9082 ( .A1(n14625), .A2(n14624), .ZN(n6580) );
  AND2_X1 U9083 ( .A1(n7536), .A2(n8804), .ZN(n6581) );
  AND2_X1 U9084 ( .A1(n10128), .A2(n12711), .ZN(n6582) );
  AND2_X1 U9085 ( .A1(n8941), .A2(n8942), .ZN(n6583) );
  XOR2_X1 U9086 ( .A(n7447), .B(n12889), .Z(n6584) );
  AND2_X1 U9087 ( .A1(n10132), .A2(n13010), .ZN(n6585) );
  NOR2_X1 U9088 ( .A1(n7327), .A2(n6585), .ZN(n6586) );
  AND2_X1 U9089 ( .A1(n7541), .A2(n13439), .ZN(n6587) );
  AND2_X1 U9090 ( .A1(n9416), .A2(n7158), .ZN(n6588) );
  AND2_X1 U9091 ( .A1(n7281), .A2(n9927), .ZN(n6589) );
  AND2_X1 U9092 ( .A1(n8658), .A2(n8643), .ZN(n6590) );
  AND2_X1 U9093 ( .A1(n7349), .A2(n10103), .ZN(n6591) );
  XOR2_X1 U9094 ( .A(n14653), .B(n14652), .Z(n6592) );
  OR2_X1 U9095 ( .A1(n8144), .A2(n7608), .ZN(n6593) );
  NAND2_X1 U9096 ( .A1(n13358), .A2(n12711), .ZN(n6594) );
  AND2_X1 U9097 ( .A1(n14355), .A2(n7583), .ZN(n6595) );
  XNOR2_X1 U9098 ( .A(n14642), .B(n14641), .ZN(n6596) );
  OR2_X1 U9099 ( .A1(n14638), .A2(n14637), .ZN(n6597) );
  INV_X1 U9100 ( .A(n6758), .ZN(n7083) );
  NAND2_X1 U9101 ( .A1(n12542), .A2(n12541), .ZN(n6758) );
  INV_X1 U9102 ( .A(n9453), .ZN(n7495) );
  AND3_X1 U9103 ( .A1(n7742), .A2(n7743), .A3(n7740), .ZN(n6598) );
  OR2_X1 U9104 ( .A1(n13853), .A2(n13532), .ZN(n6599) );
  NAND4_X1 U9105 ( .A1(n7709), .A2(n7712), .A3(n7710), .A4(n7711), .ZN(n12720)
         );
  OR2_X1 U9106 ( .A1(n14314), .A2(n14114), .ZN(n6600) );
  OR2_X1 U9107 ( .A1(n15146), .A2(n11067), .ZN(n6601) );
  AND4_X1 U9108 ( .A1(n8948), .A2(n9263), .A3(n8914), .A4(n8913), .ZN(n6602)
         );
  INV_X1 U9109 ( .A(n12543), .ZN(n6757) );
  INV_X1 U9110 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U9111 ( .A1(n9108), .A2(n9107), .ZN(n12010) );
  NOR2_X1 U9112 ( .A1(n9277), .A2(n9283), .ZN(n6603) );
  NAND2_X1 U9113 ( .A1(n13668), .A2(n9936), .ZN(n6604) );
  AND2_X1 U9114 ( .A1(n14274), .A2(n7214), .ZN(n6605) );
  OR2_X1 U9115 ( .A1(n13744), .A2(n13530), .ZN(n6606) );
  OR2_X1 U9116 ( .A1(n6562), .A2(n9635), .ZN(n6607) );
  AND2_X1 U9117 ( .A1(n8225), .A2(n6966), .ZN(n6608) );
  OR2_X1 U9118 ( .A1(n12045), .A2(n12031), .ZN(n6609) );
  INV_X1 U9119 ( .A(n12109), .ZN(n9944) );
  INV_X1 U9120 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6976) );
  NAND2_X1 U9121 ( .A1(n13663), .A2(n6996), .ZN(n6610) );
  NAND2_X1 U9122 ( .A1(n7603), .A2(n7604), .ZN(n7747) );
  OR2_X1 U9123 ( .A1(n14486), .A2(n14037), .ZN(n6611) );
  AND2_X1 U9124 ( .A1(n9679), .A2(n9678), .ZN(n6612) );
  NAND2_X1 U9125 ( .A1(n8634), .A2(n8633), .ZN(n12340) );
  AND2_X1 U9126 ( .A1(n13682), .A2(n13526), .ZN(n6613) );
  NAND2_X1 U9127 ( .A1(n13756), .A2(n6981), .ZN(n6985) );
  NAND2_X1 U9128 ( .A1(n14311), .A2(n7186), .ZN(n7187) );
  AND2_X1 U9129 ( .A1(n14291), .A2(n6600), .ZN(n6614) );
  INV_X1 U9130 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6936) );
  AND2_X1 U9131 ( .A1(n9389), .A2(n9388), .ZN(n6615) );
  INV_X1 U9132 ( .A(n9314), .ZN(n7521) );
  AND2_X1 U9133 ( .A1(n14056), .A2(n7466), .ZN(n6616) );
  AND2_X1 U9134 ( .A1(n14372), .A2(n7217), .ZN(n6617) );
  AND2_X1 U9135 ( .A1(n9856), .A2(n9855), .ZN(n6618) );
  AND2_X1 U9136 ( .A1(n9999), .A2(n9997), .ZN(n6619) );
  AND2_X1 U9137 ( .A1(n10613), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6620) );
  INV_X1 U9138 ( .A(n6961), .ZN(n6960) );
  OAI21_X1 U9139 ( .B1(n6590), .B2(n6962), .A(n13440), .ZN(n6961) );
  OR2_X1 U9140 ( .A1(n7408), .A2(n9609), .ZN(n6621) );
  OR2_X1 U9141 ( .A1(n9454), .A2(n7495), .ZN(n6622) );
  AND2_X1 U9142 ( .A1(n7082), .A2(n6757), .ZN(n6623) );
  AND2_X1 U9143 ( .A1(n7075), .A2(n6623), .ZN(n6624) );
  AND2_X1 U9144 ( .A1(n10572), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U9145 ( .A1(n7064), .A2(n7068), .ZN(n6626) );
  AND2_X1 U9146 ( .A1(n6956), .A2(n7537), .ZN(n6627) );
  NAND2_X1 U9147 ( .A1(n6798), .A2(n8983), .ZN(n6628) );
  INV_X1 U9148 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10456) );
  OR2_X1 U9149 ( .A1(n9794), .A2(n7086), .ZN(n6629) );
  NOR2_X1 U9150 ( .A1(n14486), .A2(n14117), .ZN(n6630) );
  NOR2_X1 U9151 ( .A1(n13682), .A2(n13526), .ZN(n6631) );
  NOR2_X1 U9152 ( .A1(n6993), .A2(n13903), .ZN(n6632) );
  NOR2_X1 U9153 ( .A1(n8842), .A2(n8841), .ZN(n6633) );
  NOR2_X1 U9154 ( .A1(n14510), .A2(n14072), .ZN(n6634) );
  NOR2_X1 U9155 ( .A1(n10133), .A2(n12686), .ZN(n6635) );
  NOR2_X1 U9156 ( .A1(n13744), .A2(n9876), .ZN(n6636) );
  AND2_X1 U9157 ( .A1(n10522), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6637) );
  XOR2_X1 U9158 ( .A(n14696), .B(n14695), .Z(n6638) );
  INV_X1 U9159 ( .A(n6754), .ZN(n7992) );
  OAI21_X1 U9160 ( .B1(n7989), .B2(n7988), .A(n7990), .ZN(n6754) );
  INV_X1 U9161 ( .A(n10144), .ZN(n7334) );
  NAND2_X1 U9162 ( .A1(n14330), .A2(n6790), .ZN(n6792) );
  AND2_X1 U9163 ( .A1(n6584), .A2(n10084), .ZN(n6639) );
  AND2_X1 U9164 ( .A1(n9727), .A2(n9726), .ZN(n6640) );
  AND2_X1 U9165 ( .A1(n10526), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n6641) );
  AND2_X1 U9166 ( .A1(n14246), .A2(n7213), .ZN(n6642) );
  INV_X1 U9167 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7641) );
  INV_X1 U9168 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10478) );
  INV_X1 U9169 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10481) );
  AND2_X1 U9170 ( .A1(n7613), .A2(n8151), .ZN(n6643) );
  INV_X1 U9171 ( .A(n7478), .ZN(n7477) );
  NAND2_X1 U9172 ( .A1(n7481), .A2(n7479), .ZN(n7478) );
  INV_X1 U9173 ( .A(n7242), .ZN(n7241) );
  NAND2_X1 U9174 ( .A1(n8152), .A2(n12402), .ZN(n7242) );
  INV_X1 U9175 ( .A(n7484), .ZN(n7483) );
  NAND2_X1 U9176 ( .A1(n7485), .A2(n11653), .ZN(n7484) );
  AND2_X1 U9177 ( .A1(n8519), .A2(n8261), .ZN(n6644) );
  INV_X1 U9178 ( .A(n12945), .ZN(n7070) );
  INV_X1 U9179 ( .A(n13368), .ZN(n12531) );
  NAND2_X1 U9180 ( .A1(n10460), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6645) );
  INV_X1 U9181 ( .A(n7597), .ZN(n7596) );
  NAND2_X1 U9182 ( .A1(n12488), .A2(n7600), .ZN(n7597) );
  AND2_X1 U9183 ( .A1(n9478), .A2(n14915), .ZN(n11387) );
  INV_X1 U9184 ( .A(n11387), .ZN(n7561) );
  AND2_X1 U9185 ( .A1(n14448), .A2(n14447), .ZN(n6646) );
  INV_X1 U9186 ( .A(n9954), .ZN(n6993) );
  OR2_X1 U9187 ( .A1(n14610), .A2(n14611), .ZN(n6647) );
  AND2_X1 U9188 ( .A1(n11712), .A2(n9849), .ZN(n6648) );
  OR2_X1 U9189 ( .A1(n13634), .A2(n13633), .ZN(n6649) );
  AND2_X1 U9190 ( .A1(n11133), .A2(n12732), .ZN(n6650) );
  XNOR2_X1 U9191 ( .A(n13611), .B(n9800), .ZN(n9780) );
  AND2_X1 U9192 ( .A1(n10118), .A2(n14728), .ZN(n6651) );
  NOR2_X1 U9193 ( .A1(n11740), .A2(n14126), .ZN(n6652) );
  NOR2_X1 U9194 ( .A1(n15232), .A2(n11477), .ZN(n6653) );
  AND2_X1 U9195 ( .A1(n9881), .A2(n9880), .ZN(n6654) );
  AND2_X1 U9196 ( .A1(n6580), .A2(n14628), .ZN(n6655) );
  AND2_X1 U9197 ( .A1(n7138), .A2(n7137), .ZN(n6656) );
  INV_X1 U9198 ( .A(n10262), .ZN(n7463) );
  INV_X1 U9199 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6819) );
  AND2_X1 U9200 ( .A1(n9848), .A2(n7389), .ZN(n6657) );
  AND2_X1 U9201 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(n8921), .ZN(n6658) );
  AND2_X1 U9202 ( .A1(n6760), .A2(n9795), .ZN(n6659) );
  XNOR2_X1 U9203 ( .A(n8514), .B(SI_11_), .ZN(n8513) );
  AND2_X1 U9204 ( .A1(n8108), .A2(n12536), .ZN(n8152) );
  NAND2_X1 U9205 ( .A1(n8364), .A2(n6819), .ZN(n6660) );
  NOR2_X1 U9206 ( .A1(n7321), .A2(n12612), .ZN(n7320) );
  OR2_X1 U9207 ( .A1(n7496), .A2(n9429), .ZN(n6661) );
  AND2_X1 U9208 ( .A1(n9429), .A2(n7496), .ZN(n6662) );
  OR2_X1 U9209 ( .A1(n9339), .A2(n9337), .ZN(n6663) );
  OR2_X1 U9210 ( .A1(n6640), .A2(n9729), .ZN(n6664) );
  AND2_X1 U9211 ( .A1(n7003), .A2(n7001), .ZN(n6665) );
  OR2_X1 U9212 ( .A1(n7437), .A2(n6567), .ZN(n6666) );
  OR2_X1 U9213 ( .A1(n6565), .A2(n7443), .ZN(n6667) );
  AND2_X1 U9214 ( .A1(n7610), .A2(n7659), .ZN(n6668) );
  AND2_X1 U9215 ( .A1(n7528), .A2(n8907), .ZN(n6669) );
  OR2_X1 U9216 ( .A1(n7521), .A2(n9313), .ZN(n6670) );
  OR2_X1 U9217 ( .A1(n7459), .A2(n7458), .ZN(n6671) );
  INV_X1 U9218 ( .A(n7629), .ZN(n7459) );
  INV_X1 U9219 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11039) );
  INV_X1 U9220 ( .A(n7066), .ZN(n7065) );
  NAND2_X1 U9221 ( .A1(n7060), .A2(n12528), .ZN(n7066) );
  AND2_X1 U9222 ( .A1(n10049), .A2(n9474), .ZN(n12121) );
  INV_X1 U9223 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7676) );
  INV_X1 U9224 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7181) );
  AND2_X1 U9225 ( .A1(n7925), .A2(n7923), .ZN(n6672) );
  INV_X1 U9226 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7212) );
  OAI21_X1 U9227 ( .B1(n10696), .B2(n8008), .A(n7932), .ZN(n13358) );
  INV_X1 U9228 ( .A(n13358), .ZN(n7601) );
  INV_X1 U9229 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7028) );
  INV_X1 U9230 ( .A(n13523), .ZN(n7373) );
  NAND2_X1 U9231 ( .A1(n12223), .A2(n12222), .ZN(n12221) );
  INV_X1 U9232 ( .A(SI_1_), .ZN(n7498) );
  INV_X1 U9233 ( .A(n12485), .ZN(n7226) );
  XOR2_X1 U9234 ( .A(n14691), .B(n14690), .Z(n6673) );
  NAND2_X1 U9235 ( .A1(n8031), .A2(n8030), .ZN(n12987) );
  INV_X1 U9236 ( .A(n12987), .ZN(n12625) );
  NOR2_X2 U9237 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9142) );
  NAND2_X1 U9238 ( .A1(n13498), .A2(n8663), .ZN(n13441) );
  NAND2_X1 U9239 ( .A1(n7586), .A2(n7585), .ZN(n14404) );
  NAND2_X1 U9240 ( .A1(n7550), .A2(n10047), .ZN(n12080) );
  NAND2_X1 U9241 ( .A1(n11770), .A2(n10041), .ZN(n11736) );
  AND2_X1 U9242 ( .A1(n7025), .A2(n7026), .ZN(n7859) );
  OR2_X1 U9243 ( .A1(n14739), .A2(n14730), .ZN(n6674) );
  AND2_X1 U9244 ( .A1(n12457), .A2(n15322), .ZN(n6675) );
  OR2_X1 U9245 ( .A1(n12168), .A2(n14804), .ZN(n6676) );
  NOR2_X1 U9246 ( .A1(n14730), .A2(n12714), .ZN(n6677) );
  AND2_X1 U9247 ( .A1(n9717), .A2(n9716), .ZN(n6678) );
  OR2_X1 U9248 ( .A1(n12168), .A2(n7193), .ZN(n6679) );
  AND3_X1 U9249 ( .A1(n6989), .A2(n6988), .A3(n11923), .ZN(n13771) );
  NAND2_X1 U9250 ( .A1(n7291), .A2(n6609), .ZN(n7290) );
  AND2_X1 U9251 ( .A1(n12491), .A2(n12494), .ZN(n12395) );
  NAND2_X1 U9252 ( .A1(n10143), .A2(n12976), .ZN(n6680) );
  AND2_X1 U9253 ( .A1(n7587), .A2(n10051), .ZN(n6681) );
  NAND2_X1 U9254 ( .A1(n11936), .A2(n7355), .ZN(n6682) );
  NAND2_X1 U9255 ( .A1(n12476), .A2(n12475), .ZN(n6683) );
  INV_X1 U9256 ( .A(n15309), .ZN(n14728) );
  INV_X1 U9257 ( .A(n15336), .ZN(n7042) );
  AND2_X1 U9258 ( .A1(n7314), .A2(n7313), .ZN(n6684) );
  INV_X1 U9259 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10775) );
  INV_X1 U9260 ( .A(n15149), .ZN(n11353) );
  NAND2_X1 U9261 ( .A1(n9147), .A2(n9146), .ZN(n11740) );
  INV_X1 U9262 ( .A(n11740), .ZN(n7189) );
  NAND3_X1 U9263 ( .A1(n11217), .A2(n8214), .A3(n8213), .ZN(n15439) );
  INV_X1 U9264 ( .A(n13857), .ZN(n6988) );
  AND2_X1 U9265 ( .A1(n6944), .A2(n10985), .ZN(n6685) );
  NAND2_X1 U9266 ( .A1(n10874), .A2(n10875), .ZN(n10873) );
  OR2_X1 U9267 ( .A1(n15174), .A2(n11251), .ZN(n13793) );
  INV_X1 U9268 ( .A(n13793), .ZN(n15168) );
  XOR2_X1 U9269 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .Z(n6686) );
  AND2_X1 U9270 ( .A1(n12498), .A2(n12499), .ZN(n13014) );
  INV_X1 U9271 ( .A(n13014), .ZN(n6861) );
  AND2_X1 U9272 ( .A1(n10120), .A2(n14739), .ZN(n6687) );
  AND2_X1 U9273 ( .A1(n7102), .A2(n9433), .ZN(n6688) );
  AND2_X2 U9274 ( .A1(n10404), .A2(n15182), .ZN(n15242) );
  NAND2_X1 U9275 ( .A1(n7542), .A2(n9072), .ZN(n9262) );
  AND2_X1 U9276 ( .A1(n15281), .A2(n12880), .ZN(n6689) );
  AND2_X1 U9277 ( .A1(n9852), .A2(n11348), .ZN(n6690) );
  AND2_X1 U9278 ( .A1(n11083), .A2(n9910), .ZN(n6691) );
  AND2_X1 U9279 ( .A1(n8038), .A2(n8035), .ZN(n6692) );
  INV_X1 U9280 ( .A(n6940), .ZN(n12306) );
  OR2_X1 U9281 ( .A1(n11861), .A2(n11862), .ZN(n6940) );
  NAND2_X1 U9282 ( .A1(n7292), .A2(n6787), .ZN(n6841) );
  AND2_X1 U9283 ( .A1(n7405), .A2(n7406), .ZN(n8604) );
  AND2_X1 U9284 ( .A1(n7480), .A2(n7477), .ZN(n6693) );
  OR2_X1 U9285 ( .A1(n9432), .A2(SI_29_), .ZN(n6694) );
  AND2_X1 U9286 ( .A1(n7294), .A2(n7298), .ZN(n6695) );
  AND2_X1 U9287 ( .A1(n13573), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6696) );
  OR2_X1 U9288 ( .A1(n8969), .A2(n7488), .ZN(n6697) );
  AND2_X1 U9289 ( .A1(n7232), .A2(n6498), .ZN(n6698) );
  INV_X1 U9290 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7419) );
  INV_X1 U9291 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n6736) );
  NOR2_X1 U9292 ( .A1(n9891), .A2(n9890), .ZN(n13769) );
  INV_X1 U9293 ( .A(n13769), .ZN(n15161) );
  INV_X1 U9294 ( .A(n12353), .ZN(n7412) );
  XNOR2_X1 U9295 ( .A(n8937), .B(n8936), .ZN(n9524) );
  INV_X1 U9296 ( .A(n15232), .ZN(n6967) );
  INV_X1 U9297 ( .A(n6507), .ZN(n6848) );
  INV_X1 U9298 ( .A(n11831), .ZN(n6840) );
  INV_X1 U9299 ( .A(n12836), .ZN(n7004) );
  NOR2_X1 U9300 ( .A1(n15265), .A2(n11588), .ZN(n6699) );
  AND2_X1 U9301 ( .A1(n10539), .A2(n10538), .ZN(n15129) );
  NAND2_X1 U9302 ( .A1(n7237), .A2(n7236), .ZN(n6700) );
  OR2_X1 U9303 ( .A1(n11304), .A2(n11305), .ZN(n7315) );
  AND2_X1 U9304 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n9564), .ZN(n6701) );
  OR2_X1 U9305 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n9564), .ZN(n6702) );
  INV_X1 U9306 ( .A(n7009), .ZN(n7008) );
  AOI21_X1 U9307 ( .B1(n12039), .B2(n12037), .A(n12040), .ZN(n7009) );
  INV_X1 U9308 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n6720) );
  INV_X1 U9309 ( .A(n8170), .ZN(n12553) );
  XNOR2_X1 U9310 ( .A(n7649), .B(n7028), .ZN(n12889) );
  OR2_X1 U9311 ( .A1(n8264), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n6777) );
  AND2_X1 U9312 ( .A1(n6891), .A2(n6890), .ZN(n6703) );
  AND2_X1 U9313 ( .A1(n11585), .A2(n11302), .ZN(n6704) );
  AND2_X1 U9314 ( .A1(n11604), .A2(n11306), .ZN(n6705) );
  AND2_X1 U9315 ( .A1(n11053), .A2(n11052), .ZN(n6706) );
  NOR2_X1 U9316 ( .A1(n13412), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n6707) );
  XNOR2_X1 U9317 ( .A(n14135), .B(n14980), .ZN(n11369) );
  INV_X1 U9318 ( .A(n11829), .ZN(n7302) );
  NAND2_X1 U9319 ( .A1(n7304), .A2(n11829), .ZN(n7303) );
  OR2_X1 U9320 ( .A1(n15428), .A2(n15346), .ZN(n13392) );
  MUX2_X1 U9321 ( .A(n9560), .B(P3_REG0_REG_28__SCAN_IN), .S(n15428), .Z(n9558) );
  NAND2_X1 U9322 ( .A1(n6712), .A2(n6711), .ZN(n6710) );
  XNOR2_X1 U9323 ( .A(n12379), .B(n12872), .ZN(n6712) );
  NAND2_X1 U9324 ( .A1(n15378), .A2(n12427), .ZN(n11098) );
  NAND2_X1 U9325 ( .A1(n12214), .A2(n12475), .ZN(n6716) );
  OAI21_X1 U9326 ( .B1(n11458), .B2(n12385), .A(n6717), .ZN(n11752) );
  NOR2_X1 U9327 ( .A1(n6722), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n7025) );
  NOR2_X2 U9328 ( .A1(n7684), .A2(n6722), .ZN(n7857) );
  NAND2_X1 U9329 ( .A1(n6724), .A2(n14594), .ZN(n6723) );
  INV_X1 U9330 ( .A(n14594), .ZN(n6725) );
  NAND2_X1 U9331 ( .A1(n6729), .A2(n6580), .ZN(n6727) );
  NOR2_X2 U9332 ( .A1(n14667), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6728) );
  OAI21_X2 U9333 ( .B1(n14688), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n6731), .ZN(
        n7360) );
  NAND2_X1 U9334 ( .A1(n6732), .A2(n6592), .ZN(n6731) );
  INV_X1 U9335 ( .A(n14852), .ZN(n6734) );
  INV_X1 U9336 ( .A(n6744), .ZN(n6743) );
  XNOR2_X1 U9337 ( .A(n6745), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U9338 ( .B1(n6750), .B2(n12551), .A(n6749), .ZN(n6748) );
  NAND3_X1 U9339 ( .A1(n7422), .A2(n7424), .A3(n7744), .ZN(n6752) );
  NAND2_X1 U9340 ( .A1(n6756), .A2(n7872), .ZN(n7873) );
  NAND2_X1 U9341 ( .A1(n7856), .A2(n7855), .ZN(n7871) );
  AOI21_X1 U9342 ( .B1(n9734), .B2(n9733), .A(n9730), .ZN(n6761) );
  NAND3_X1 U9343 ( .A1(n6764), .A2(n6667), .A3(n6762), .ZN(n6921) );
  NAND2_X1 U9344 ( .A1(n6763), .A2(n9641), .ZN(n6762) );
  INV_X1 U9345 ( .A(n6766), .ZN(n6763) );
  NAND2_X1 U9346 ( .A1(n6765), .A2(n9639), .ZN(n6764) );
  NAND2_X1 U9347 ( .A1(n6766), .A2(n9640), .ZN(n6765) );
  NAND2_X1 U9348 ( .A1(n6768), .A2(n9626), .ZN(n6767) );
  INV_X1 U9349 ( .A(n6771), .ZN(n6768) );
  NAND2_X1 U9350 ( .A1(n6770), .A2(n9624), .ZN(n6769) );
  NAND2_X1 U9351 ( .A1(n6771), .A2(n9625), .ZN(n6770) );
  NAND2_X1 U9352 ( .A1(n9620), .A2(n9619), .ZN(n6771) );
  NOR2_X1 U9353 ( .A1(n6772), .A2(n9713), .ZN(n9714) );
  AOI21_X1 U9354 ( .B1(n6772), .B2(n9713), .A(n9712), .ZN(n9715) );
  NAND2_X1 U9355 ( .A1(n6774), .A2(n6773), .ZN(n9691) );
  NAND2_X1 U9356 ( .A1(n6775), .A2(n9685), .ZN(n6774) );
  OAI21_X1 U9357 ( .B1(n7445), .B2(n9677), .A(n7444), .ZN(n6776) );
  NAND4_X1 U9358 ( .A1(n8243), .A2(n7631), .A3(n6976), .A4(n8261), .ZN(n8264)
         );
  OAI211_X1 U9359 ( .C1(n9833), .C2(n6779), .A(n6778), .B(n9808), .ZN(n6808)
         );
  NAND2_X1 U9360 ( .A1(n9833), .A2(n9807), .ZN(n6778) );
  INV_X1 U9361 ( .A(n9806), .ZN(n6779) );
  NAND2_X1 U9362 ( .A1(n6574), .A2(n6706), .ZN(n12729) );
  NAND2_X1 U9363 ( .A1(n14947), .A2(n14946), .ZN(n9969) );
  NAND2_X1 U9364 ( .A1(n11364), .A2(n9966), .ZN(n6789) );
  NAND3_X1 U9365 ( .A1(n9485), .A2(n9985), .A3(n12085), .ZN(n12117) );
  OAI21_X1 U9366 ( .B1(n6795), .B2(n9992), .A(n7216), .ZN(n6794) );
  NAND2_X1 U9367 ( .A1(n7577), .A2(n8918), .ZN(n8933) );
  NAND2_X1 U9368 ( .A1(n7214), .A2(n14266), .ZN(n6796) );
  INV_X1 U9369 ( .A(n7214), .ZN(n6797) );
  NAND2_X1 U9370 ( .A1(n14245), .A2(n10003), .ZN(n10004) );
  NAND2_X2 U9371 ( .A1(n8983), .A2(n10476), .ZN(n9436) );
  NAND2_X1 U9372 ( .A1(n9988), .A2(n9987), .ZN(n14420) );
  NOR2_X1 U9373 ( .A1(n7771), .A2(n15269), .ZN(n15268) );
  NAND2_X1 U9374 ( .A1(n9982), .A2(n9981), .ZN(n11973) );
  NAND2_X1 U9375 ( .A1(n9962), .A2(n9961), .ZN(n11321) );
  OAI21_X1 U9376 ( .B1(n12866), .B2(n15298), .A(n6902), .ZN(n6901) );
  INV_X1 U9377 ( .A(n6901), .ZN(n12868) );
  XNOR2_X2 U9378 ( .A(n14820), .B(n14123), .ZN(n12086) );
  NAND2_X1 U9379 ( .A1(n8479), .A2(n8478), .ZN(n8495) );
  NAND2_X1 U9380 ( .A1(n8357), .A2(n8356), .ZN(n8383) );
  NAND2_X1 U9381 ( .A1(n8623), .A2(n8622), .ZN(n8626) );
  NAND3_X1 U9382 ( .A1(n6889), .A2(n6888), .A3(n6801), .ZN(P2_U3233) );
  NAND2_X1 U9383 ( .A1(n6802), .A2(n13607), .ZN(n6801) );
  INV_X1 U9384 ( .A(n13608), .ZN(n6802) );
  NOR2_X2 U9385 ( .A1(n13635), .A2(n7372), .ZN(n7371) );
  MUX2_X1 U9386 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8255), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8257) );
  NOR2_X1 U9387 ( .A1(n13623), .A2(n9947), .ZN(n10405) );
  NOR2_X1 U9388 ( .A1(n11963), .A2(n11964), .ZN(n13565) );
  NOR2_X1 U9389 ( .A1(n15094), .A2(n15095), .ZN(n15093) );
  NOR2_X1 U9390 ( .A1(n10673), .A2(n10672), .ZN(n10751) );
  AOI21_X1 U9391 ( .B1(n13647), .B2(n13646), .A(n9889), .ZN(n13634) );
  OAI21_X1 U9392 ( .B1(n7638), .B2(n12378), .A(n12377), .ZN(n12379) );
  NAND2_X1 U9393 ( .A1(n11410), .A2(n12442), .ZN(n11458) );
  NOR2_X1 U9394 ( .A1(n12769), .A2(n12770), .ZN(n12789) );
  NAND4_X1 U9395 ( .A1(n14694), .A2(n7091), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7090) );
  OAI21_X2 U9396 ( .B1(n13781), .B2(n9868), .A(n6845), .ZN(n13767) );
  NAND2_X1 U9397 ( .A1(n8283), .A2(n8282), .ZN(n8288) );
  NAND2_X1 U9398 ( .A1(n7502), .A2(n7500), .ZN(n8430) );
  AOI21_X1 U9399 ( .B1(n7368), .B2(n7370), .A(n6653), .ZN(n7366) );
  NAND2_X1 U9400 ( .A1(n7233), .A2(n7235), .ZN(n11586) );
  NAND2_X1 U9401 ( .A1(n6806), .A2(n6804), .ZN(P2_U3236) );
  NAND2_X1 U9402 ( .A1(n7230), .A2(n7231), .ZN(n12044) );
  NAND2_X1 U9403 ( .A1(n11588), .A2(n7245), .ZN(n7243) );
  NOR2_X2 U9404 ( .A1(n15286), .A2(n15285), .ZN(n15284) );
  OAI21_X1 U9405 ( .B1(n12789), .B2(n12788), .A(n12795), .ZN(n12790) );
  NAND2_X1 U9406 ( .A1(n7249), .A2(n12787), .ZN(n12827) );
  OAI21_X1 U9407 ( .B1(n12891), .B2(n15304), .A(n7017), .ZN(n7016) );
  NAND2_X1 U9408 ( .A1(n8475), .A2(n8474), .ZN(n8479) );
  NAND2_X1 U9409 ( .A1(n8353), .A2(n8352), .ZN(n8357) );
  NAND3_X1 U9410 ( .A1(n9828), .A2(n7087), .A3(n9782), .ZN(n9790) );
  NAND3_X1 U9411 ( .A1(n8282), .A2(n7499), .A3(n8251), .ZN(n8283) );
  NAND2_X1 U9412 ( .A1(n9960), .A2(n11728), .ZN(n9962) );
  INV_X1 U9413 ( .A(n14137), .ZN(n8986) );
  NAND3_X2 U9414 ( .A1(n8943), .A2(n8944), .A3(n6583), .ZN(n14137) );
  NAND3_X2 U9415 ( .A1(n7577), .A2(n8918), .A3(n8936), .ZN(n8920) );
  NAND2_X1 U9416 ( .A1(n8288), .A2(n8287), .ZN(n8303) );
  NAND3_X1 U9417 ( .A1(n7704), .A2(n7703), .A3(n6807), .ZN(n11208) );
  OAI21_X1 U9418 ( .B1(n6615), .B2(n7153), .A(n7152), .ZN(n6824) );
  NOR2_X1 U9419 ( .A1(n9714), .A2(n7456), .ZN(n7453) );
  OAI21_X1 U9420 ( .B1(n6882), .B2(n9723), .A(n7435), .ZN(n9734) );
  NAND2_X1 U9421 ( .A1(n9631), .A2(n9630), .ZN(n6811) );
  NAND2_X1 U9422 ( .A1(n6812), .A2(n6809), .ZN(n6830) );
  INV_X1 U9423 ( .A(n6881), .ZN(n6812) );
  NAND3_X1 U9424 ( .A1(n6808), .A2(n9834), .A3(n9835), .ZN(P2_U3328) );
  AOI21_X1 U9425 ( .B1(n9691), .B2(n9690), .A(n9689), .ZN(n6813) );
  OAI22_X1 U9426 ( .A1(n7457), .A2(n6813), .B1(n9696), .B2(n7629), .ZN(n9701)
         );
  NOR2_X1 U9427 ( .A1(n13602), .A2(n13601), .ZN(n13603) );
  NOR2_X1 U9428 ( .A1(n6703), .A2(n7402), .ZN(n15046) );
  NOR2_X1 U9429 ( .A1(n7395), .A2(n7394), .ZN(n13602) );
  NAND2_X1 U9430 ( .A1(n15307), .A2(n7591), .ZN(n7590) );
  INV_X1 U9431 ( .A(n7663), .ZN(n12562) );
  NAND2_X1 U9432 ( .A1(n13009), .A2(n8140), .ZN(n12997) );
  NAND2_X1 U9433 ( .A1(n11461), .A2(n11460), .ZN(n11459) );
  NAND2_X1 U9434 ( .A1(n11229), .A2(n11228), .ZN(n11227) );
  NAND2_X1 U9435 ( .A1(n7838), .A2(n12465), .ZN(n14735) );
  NAND2_X1 U9436 ( .A1(n6822), .A2(n9500), .ZN(n9510) );
  NAND3_X1 U9437 ( .A1(n9503), .A2(n6577), .A3(n7616), .ZN(n6822) );
  NAND2_X1 U9438 ( .A1(n9238), .A2(n7166), .ZN(n7164) );
  NAND2_X1 U9439 ( .A1(n7104), .A2(n8885), .ZN(n9426) );
  NAND2_X1 U9440 ( .A1(n7519), .A2(n7520), .ZN(n7151) );
  NAND2_X1 U9441 ( .A1(n7146), .A2(n7145), .ZN(n9351) );
  NAND2_X1 U9442 ( .A1(n11824), .A2(n8971), .ZN(n9448) );
  OAI22_X1 U9443 ( .A1(n9368), .A2(n7507), .B1(n9369), .B2(n7508), .ZN(n9384)
         );
  NAND2_X1 U9444 ( .A1(n6828), .A2(n6827), .ZN(n6826) );
  NAND2_X1 U9445 ( .A1(n6860), .A2(n9707), .ZN(n6829) );
  NAND2_X1 U9446 ( .A1(n6921), .A2(n6920), .ZN(n9650) );
  NAND2_X1 U9447 ( .A1(n9650), .A2(n9651), .ZN(n9649) );
  NAND2_X1 U9448 ( .A1(n6923), .A2(n6922), .ZN(n9665) );
  OAI21_X1 U9449 ( .B1(n6659), .B2(n6859), .A(n6563), .ZN(n7113) );
  NAND2_X1 U9450 ( .A1(n7399), .A2(n7398), .ZN(n7397) );
  NOR2_X1 U9451 ( .A1(n15109), .A2(n15108), .ZN(n15107) );
  NAND2_X1 U9452 ( .A1(n10969), .A2(n10968), .ZN(n11959) );
  NAND2_X1 U9453 ( .A1(n7182), .A2(n13700), .ZN(n6889) );
  NAND2_X1 U9454 ( .A1(n10927), .A2(n6657), .ZN(n7388) );
  INV_X1 U9455 ( .A(n13635), .ZN(n6867) );
  NAND2_X1 U9456 ( .A1(n9842), .A2(n9841), .ZN(n11261) );
  NAND2_X1 U9457 ( .A1(n9839), .A2(n9838), .ZN(n11565) );
  NAND2_X1 U9458 ( .A1(n6836), .A2(n6834), .ZN(P1_U3214) );
  NAND2_X1 U9459 ( .A1(n13933), .A2(n14082), .ZN(n6836) );
  NAND2_X1 U9460 ( .A1(n13991), .A2(n10277), .ZN(n14045) );
  NAND2_X1 U9461 ( .A1(n9595), .A2(n9594), .ZN(n9602) );
  NAND2_X1 U9462 ( .A1(n14079), .A2(n12578), .ZN(n13931) );
  NAND2_X1 U9463 ( .A1(n6862), .A2(n6861), .ZN(n13009) );
  NAND2_X1 U9464 ( .A1(n13281), .A2(n8139), .ZN(n13007) );
  NAND2_X1 U9465 ( .A1(n10863), .A2(n12721), .ZN(n12421) );
  NAND2_X1 U9466 ( .A1(n14250), .A2(n14261), .ZN(n14249) );
  NAND2_X1 U9467 ( .A1(n14267), .A2(n14266), .ZN(n14265) );
  NAND2_X1 U9468 ( .A1(n14236), .A2(n14235), .ZN(n14234) );
  INV_X1 U9469 ( .A(n7564), .ZN(n7563) );
  INV_X1 U9470 ( .A(n13007), .ZN(n6862) );
  NAND2_X1 U9471 ( .A1(n12424), .A2(n15377), .ZN(n11100) );
  NAND2_X1 U9472 ( .A1(n13282), .A2(n6502), .ZN(n13281) );
  NAND2_X1 U9473 ( .A1(n11850), .A2(n9857), .ZN(n12022) );
  AOI21_X1 U9474 ( .B1(n7388), .B2(n6554), .A(n6648), .ZN(n7618) );
  NAND2_X1 U9475 ( .A1(n7378), .A2(n7379), .ZN(n13720) );
  NOR2_X1 U9476 ( .A1(n10224), .A2(n10223), .ZN(n13963) );
  NAND2_X1 U9477 ( .A1(n12131), .A2(n12142), .ZN(n6844) );
  NAND2_X1 U9478 ( .A1(n6847), .A2(n15161), .ZN(n6846) );
  XNOR2_X1 U9479 ( .A(n7371), .B(n9940), .ZN(n6847) );
  INV_X1 U9480 ( .A(n14562), .ZN(n7119) );
  NAND3_X1 U9481 ( .A1(n7121), .A2(n7123), .A3(n6851), .ZN(n6850) );
  OAI21_X1 U9482 ( .B1(n14449), .B2(n14825), .A(n6646), .ZN(n14517) );
  OAI21_X1 U9483 ( .B1(n14244), .B2(n14246), .A(n14245), .ZN(n14449) );
  NAND2_X1 U9484 ( .A1(n6852), .A2(n7202), .ZN(n11988) );
  NAND2_X1 U9485 ( .A1(n11772), .A2(n7203), .ZN(n6852) );
  NAND2_X1 U9486 ( .A1(n6855), .A2(n6621), .ZN(n9615) );
  NAND3_X1 U9487 ( .A1(n9604), .A2(n7407), .A3(n9603), .ZN(n6855) );
  INV_X1 U9488 ( .A(n9608), .ZN(n7408) );
  NAND2_X1 U9489 ( .A1(n7084), .A2(n8541), .ZN(n8557) );
  NAND2_X1 U9490 ( .A1(n7514), .A2(n8559), .ZN(n8598) );
  INV_X1 U9491 ( .A(n7497), .ZN(n8246) );
  NAND2_X1 U9492 ( .A1(n7195), .A2(n6883), .ZN(n14516) );
  AOI21_X1 U9493 ( .B1(n7551), .B2(n7553), .A(n7549), .ZN(n7548) );
  NAND2_X1 U9494 ( .A1(n7623), .A2(n6629), .ZN(n6859) );
  NAND2_X1 U9495 ( .A1(n8787), .A2(n8786), .ZN(n7106) );
  OR2_X1 U9496 ( .A1(n9676), .A2(n7446), .ZN(n7445) );
  OAI21_X1 U9497 ( .B1(n9725), .B2(n9724), .A(n6664), .ZN(n6882) );
  NOR2_X2 U9498 ( .A1(n8912), .A2(n8911), .ZN(n6916) );
  NAND3_X1 U9499 ( .A1(n6865), .A2(n6917), .A3(n6918), .ZN(n6864) );
  NAND2_X2 U9500 ( .A1(n10360), .A2(n13954), .ZN(n14030) );
  NOR2_X1 U9501 ( .A1(n10883), .A2(n7617), .ZN(n10777) );
  INV_X1 U9502 ( .A(n8985), .ZN(n14964) );
  INV_X1 U9503 ( .A(n11786), .ZN(n9853) );
  NAND2_X2 U9504 ( .A1(n10540), .A2(n6973), .ZN(n10533) );
  AND2_X2 U9505 ( .A1(n8291), .A2(n8292), .ZN(n11684) );
  NAND2_X1 U9506 ( .A1(n9837), .A2(n9836), .ZN(n11673) );
  XNOR2_X1 U9507 ( .A(n14610), .B(n14611), .ZN(n15443) );
  INV_X1 U9508 ( .A(n14672), .ZN(n6870) );
  NAND4_X1 U9509 ( .A1(n8272), .A2(n8274), .A3(n8275), .A4(n8273), .ZN(n9589)
         );
  AND2_X2 U9510 ( .A1(n6866), .A2(n13637), .ZN(n13805) );
  NAND3_X1 U9511 ( .A1(n6867), .A2(n6649), .A3(n15161), .ZN(n6866) );
  INV_X1 U9512 ( .A(n9781), .ZN(n7089) );
  NAND2_X1 U9513 ( .A1(n8626), .A2(n7110), .ZN(n7109) );
  NAND2_X1 U9514 ( .A1(n7511), .A2(n7512), .ZN(n8623) );
  NAND2_X1 U9515 ( .A1(n7085), .A2(n8516), .ZN(n8539) );
  NAND2_X1 U9516 ( .A1(n8709), .A2(n8708), .ZN(n8712) );
  NAND3_X1 U9517 ( .A1(n8829), .A2(n7105), .A3(n8828), .ZN(n7104) );
  NAND2_X2 U9518 ( .A1(n14948), .A2(n14218), .ZN(n14682) );
  INV_X1 U9519 ( .A(n10219), .ZN(n6917) );
  XNOR2_X1 U9520 ( .A(n10203), .B(n12589), .ZN(n10225) );
  NAND2_X1 U9521 ( .A1(n7893), .A2(n7892), .ZN(n7906) );
  INV_X1 U9522 ( .A(n8918), .ZN(n8965) );
  NOR2_X1 U9523 ( .A1(n7076), .A2(n12548), .ZN(n7073) );
  NAND2_X1 U9524 ( .A1(n7430), .A2(n7429), .ZN(n7856) );
  XNOR2_X1 U9525 ( .A(n6874), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14216) );
  NOR2_X1 U9526 ( .A1(n14894), .A2(n14213), .ZN(n6874) );
  OAI21_X2 U9527 ( .B1(n11268), .B2(n9847), .A(n9846), .ZN(n10929) );
  NAND2_X1 U9528 ( .A1(n7268), .A2(n7387), .ZN(P2_U3496) );
  NAND2_X1 U9529 ( .A1(n6909), .A2(n6907), .ZN(P2_U3527) );
  NAND2_X1 U9530 ( .A1(n8243), .A2(n7631), .ZN(n6880) );
  OAI21_X1 U9531 ( .B1(n9631), .B2(n9630), .A(n6607), .ZN(n6881) );
  INV_X1 U9532 ( .A(n9623), .ZN(n9624) );
  INV_X1 U9533 ( .A(n12793), .ZN(n7249) );
  INV_X1 U9534 ( .A(n7016), .ZN(n7015) );
  XNOR2_X1 U9535 ( .A(n12810), .B(n12811), .ZN(n14703) );
  NAND2_X1 U9536 ( .A1(n7197), .A2(n6501), .ZN(n12085) );
  NAND2_X1 U9537 ( .A1(n7210), .A2(n7207), .ZN(n14385) );
  NAND2_X1 U9538 ( .A1(n9984), .A2(n9983), .ZN(n12087) );
  XNOR2_X1 U9539 ( .A(n10004), .B(n10062), .ZN(n14443) );
  NAND2_X1 U9540 ( .A1(n14443), .A2(n14442), .ZN(n7195) );
  NAND2_X1 U9541 ( .A1(n13554), .A2(n13553), .ZN(n13552) );
  NOR2_X1 U9542 ( .A1(n15082), .A2(n15081), .ZN(n15080) );
  NOR2_X1 U9543 ( .A1(n15117), .A2(n15116), .ZN(n15115) );
  NOR2_X1 U9544 ( .A1(n10853), .A2(n10852), .ZN(n10965) );
  INV_X1 U9545 ( .A(n13604), .ZN(n7183) );
  NOR2_X1 U9546 ( .A1(n13565), .A2(n6696), .ZN(n15094) );
  INV_X1 U9547 ( .A(n15134), .ZN(n7399) );
  NOR2_X1 U9548 ( .A1(n15093), .A2(n7403), .ZN(n13567) );
  XNOR2_X1 U9549 ( .A(n13567), .B(n13580), .ZN(n15109) );
  NAND2_X1 U9550 ( .A1(n8457), .A2(n8475), .ZN(n10519) );
  OAI21_X1 U9551 ( .B1(n11918), .B2(n14776), .A(n13537), .ZN(n9860) );
  NAND2_X1 U9552 ( .A1(n8331), .A2(n8330), .ZN(n8353) );
  NOR2_X1 U9553 ( .A1(n9850), .A2(n7370), .ZN(n7369) );
  NAND2_X1 U9554 ( .A1(n9590), .A2(n9591), .ZN(n9593) );
  NAND2_X1 U9555 ( .A1(n7920), .A2(n12484), .ZN(n12281) );
  NAND2_X1 U9556 ( .A1(n6894), .A2(n6893), .ZN(P2_U3495) );
  NAND2_X1 U9557 ( .A1(n8480), .A2(n8495), .ZN(n10525) );
  NOR2_X1 U9558 ( .A1(n11491), .A2(n7369), .ZN(n7368) );
  OAI21_X1 U9559 ( .B1(n8247), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6913), .ZN(
        n8250) );
  INV_X1 U9560 ( .A(n15171), .ZN(n15192) );
  AND2_X4 U9561 ( .A1(n12588), .A2(n14682), .ZN(n10196) );
  NAND2_X1 U9562 ( .A1(n15158), .A2(n7385), .ZN(n9837) );
  NAND2_X1 U9563 ( .A1(n12909), .A2(n15385), .ZN(n6906) );
  INV_X1 U9564 ( .A(n12720), .ZN(n11103) );
  NAND2_X1 U9565 ( .A1(n8430), .A2(n8429), .ZN(n8452) );
  NAND2_X1 U9566 ( .A1(n8729), .A2(n8728), .ZN(n8732) );
  NAND2_X1 U9567 ( .A1(n14596), .A2(n14597), .ZN(n7117) );
  XNOR2_X1 U9568 ( .A(n6899), .B(n6638), .ZN(SUB_1596_U4) );
  NAND2_X1 U9569 ( .A1(n7120), .A2(n7359), .ZN(n7127) );
  NAND2_X4 U9570 ( .A1(n8924), .A2(n8925), .ZN(n9032) );
  NAND2_X1 U9571 ( .A1(n10224), .A2(n10220), .ZN(n6918) );
  MUX2_X1 U9572 ( .A(n10372), .B(n10822), .S(n10821), .Z(n10884) );
  XNOR2_X1 U9573 ( .A(n6900), .B(n12772), .ZN(n12758) );
  NOR2_X1 U9574 ( .A1(n11180), .A2(n15431), .ZN(n11179) );
  NAND2_X1 U9575 ( .A1(n8233), .A2(n8225), .ZN(n8227) );
  NAND2_X2 U9576 ( .A1(n8229), .A2(n8230), .ZN(n11766) );
  NAND4_X2 U9577 ( .A1(n8346), .A2(n8345), .A3(n8344), .A4(n8343), .ZN(n13547)
         );
  NAND2_X1 U9578 ( .A1(n15240), .A2(n6912), .ZN(n6911) );
  OR2_X2 U9579 ( .A1(n13767), .A2(n9869), .ZN(n9872) );
  NAND2_X1 U9580 ( .A1(n7367), .A2(n7366), .ZN(n11786) );
  INV_X1 U9581 ( .A(n7362), .ZN(n14646) );
  NAND2_X1 U9582 ( .A1(n10298), .A2(n7470), .ZN(n14000) );
  AND2_X4 U9583 ( .A1(n6916), .A2(n6602), .ZN(n8918) );
  OAI21_X2 U9584 ( .B1(n11652), .B2(n7478), .A(n7475), .ZN(n10256) );
  NAND3_X1 U9585 ( .A1(n9655), .A2(n9654), .A3(n6666), .ZN(n6923) );
  NAND2_X1 U9586 ( .A1(n8244), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6977) );
  NAND3_X1 U9587 ( .A1(n6973), .A2(P2_IR_REG_0__SCAN_IN), .A3(n10540), .ZN(
        n6970) );
  NAND2_X2 U9588 ( .A1(n6938), .A2(n6969), .ZN(n10540) );
  AND2_X2 U9589 ( .A1(n12114), .A2(n8594), .ZN(n12223) );
  OR2_X2 U9590 ( .A1(n12108), .A2(n6571), .ZN(n12114) );
  NAND3_X1 U9591 ( .A1(n8447), .A2(n6942), .A3(n6941), .ZN(n11070) );
  NAND2_X1 U9592 ( .A1(n10985), .A2(n6945), .ZN(n6941) );
  NAND3_X1 U9593 ( .A1(n6943), .A2(n10923), .A3(n10985), .ZN(n6942) );
  INV_X1 U9594 ( .A(n8404), .ZN(n6945) );
  NAND2_X1 U9595 ( .A1(n11246), .A2(n6946), .ZN(n11476) );
  NAND2_X2 U9596 ( .A1(n8469), .A2(n11240), .ZN(n11246) );
  NAND3_X1 U9597 ( .A1(n6948), .A2(n6947), .A3(n6669), .ZN(P2_U3192) );
  NAND2_X1 U9598 ( .A1(n8854), .A2(n6949), .ZN(n6947) );
  OR2_X1 U9599 ( .A1(n8854), .A2(n6951), .ZN(n6948) );
  INV_X1 U9600 ( .A(n8853), .ZN(n6955) );
  NAND2_X1 U9601 ( .A1(n12349), .A2(n6958), .ZN(n6957) );
  AND2_X1 U9602 ( .A1(n8630), .A2(n6963), .ZN(n8231) );
  NAND2_X1 U9603 ( .A1(n8631), .A2(n6964), .ZN(n8855) );
  AND2_X1 U9604 ( .A1(n6608), .A2(n8224), .ZN(n6963) );
  INV_X1 U9605 ( .A(n6985), .ZN(n13712) );
  NAND2_X1 U9606 ( .A1(n13613), .A2(n13742), .ZN(n13797) );
  NAND2_X1 U9607 ( .A1(n12835), .A2(n7001), .ZN(n7000) );
  NAND2_X1 U9608 ( .A1(n7007), .A2(n7006), .ZN(n12748) );
  NAND2_X1 U9609 ( .A1(n12036), .A2(n12039), .ZN(n7007) );
  INV_X1 U9610 ( .A(n7010), .ZN(n15294) );
  NAND3_X1 U9611 ( .A1(n7603), .A2(n7640), .A3(n7604), .ZN(n7684) );
  MUX2_X1 U9612 ( .A(n15431), .B(n11221), .S(n12553), .Z(n11008) );
  MUX2_X1 U9613 ( .A(n11009), .B(n11010), .S(n12553), .Z(n11011) );
  MUX2_X1 U9614 ( .A(n11005), .B(n11006), .S(n12553), .Z(n11013) );
  NAND2_X1 U9615 ( .A1(n11132), .A2(n6650), .ZN(n7012) );
  NAND2_X1 U9616 ( .A1(n7012), .A2(n7013), .ZN(n12735) );
  INV_X1 U9617 ( .A(n11016), .ZN(n7014) );
  NAND3_X1 U9618 ( .A1(n7019), .A2(n7018), .A3(n7015), .ZN(P3_U3201) );
  NAND3_X1 U9619 ( .A1(n7025), .A2(n7026), .A3(n7641), .ZN(n7658) );
  NOR2_X1 U9620 ( .A1(n7031), .A2(n12448), .ZN(n7041) );
  NAND2_X1 U9621 ( .A1(n7032), .A2(n7037), .ZN(n12462) );
  NAND2_X1 U9622 ( .A1(n12468), .A2(n7046), .ZN(n7044) );
  NAND2_X1 U9623 ( .A1(n7044), .A2(n7045), .ZN(n12477) );
  NAND2_X1 U9624 ( .A1(n7058), .A2(n7057), .ZN(n12538) );
  NAND2_X1 U9625 ( .A1(n12520), .A2(n7059), .ZN(n7057) );
  NAND3_X1 U9626 ( .A1(n7064), .A2(n7068), .A3(n7066), .ZN(n7063) );
  NAND3_X1 U9627 ( .A1(n12544), .A2(n7077), .A3(n7075), .ZN(n7071) );
  NAND2_X1 U9628 ( .A1(n8539), .A2(n8538), .ZN(n7084) );
  NAND2_X1 U9629 ( .A1(n8495), .A2(n7509), .ZN(n7085) );
  INV_X1 U9630 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7093) );
  INV_X1 U9631 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7091) );
  NAND4_X1 U9632 ( .A1(n13610), .A2(n7094), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n7093), .ZN(n7092) );
  INV_X1 U9633 ( .A(n8829), .ZN(n7097) );
  NAND2_X1 U9634 ( .A1(n8829), .A2(n8828), .ZN(n8887) );
  INV_X1 U9635 ( .A(n8886), .ZN(n7105) );
  OAI21_X2 U9636 ( .B1(n8807), .B2(n8806), .A(n8808), .ZN(n8827) );
  NAND2_X1 U9637 ( .A1(n7109), .A2(n7107), .ZN(n8691) );
  NAND2_X1 U9638 ( .A1(n7628), .A2(n8688), .ZN(n7112) );
  NAND2_X1 U9639 ( .A1(n14631), .A2(n15079), .ZN(n7115) );
  NAND3_X1 U9640 ( .A1(n14562), .A2(n14563), .A3(n7126), .ZN(n7123) );
  NAND2_X1 U9641 ( .A1(n7119), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n7121) );
  NAND2_X1 U9642 ( .A1(n14562), .A2(n14563), .ZN(n7120) );
  NAND2_X1 U9643 ( .A1(n14562), .A2(n7125), .ZN(n7124) );
  NAND2_X1 U9644 ( .A1(n14562), .A2(n14563), .ZN(n14564) );
  OAI21_X2 U9645 ( .B1(n14850), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7128), .ZN(
        n7362) );
  NAND2_X1 U9646 ( .A1(n7129), .A2(n6596), .ZN(n7128) );
  INV_X1 U9647 ( .A(n14851), .ZN(n7138) );
  NAND2_X1 U9648 ( .A1(n14647), .A2(n7135), .ZN(n7130) );
  NOR2_X1 U9649 ( .A1(n6656), .A2(n14647), .ZN(n14853) );
  OAI21_X1 U9650 ( .B1(n14647), .B2(n7135), .A(n15128), .ZN(n7134) );
  INV_X1 U9651 ( .A(n14854), .ZN(n7135) );
  INV_X1 U9652 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7137) );
  NAND2_X2 U9653 ( .A1(n14218), .A2(n14547), .ZN(n10026) );
  XNOR2_X2 U9654 ( .A(n7144), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14547) );
  NAND3_X1 U9655 ( .A1(n7148), .A2(n7147), .A3(n6663), .ZN(n7146) );
  OR2_X1 U9656 ( .A1(n7151), .A2(n9327), .ZN(n7147) );
  NAND2_X1 U9657 ( .A1(n7160), .A2(n9299), .ZN(n9303) );
  NAND3_X1 U9658 ( .A1(n7164), .A2(n7163), .A3(n7161), .ZN(n7160) );
  NAND3_X1 U9659 ( .A1(n7164), .A2(n7163), .A3(n7167), .ZN(n9301) );
  INV_X2 U9660 ( .A(n8992), .ZN(n9413) );
  NAND2_X2 U9661 ( .A1(n9450), .A2(n8972), .ZN(n8992) );
  NAND2_X2 U9662 ( .A1(n8918), .A2(n8963), .ZN(n8969) );
  NAND2_X1 U9663 ( .A1(n9093), .A2(n9094), .ZN(n9092) );
  OAI22_X1 U9664 ( .A1(n9149), .A2(n7172), .B1(n9150), .B2(n7171), .ZN(n9166)
         );
  NAND2_X1 U9665 ( .A1(n9126), .A2(n9127), .ZN(n9125) );
  MUX2_X1 U9666 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7181), .S(n10553), .Z(n15049) );
  INV_X1 U9667 ( .A(n7187), .ZN(n14254) );
  INV_X1 U9668 ( .A(n12087), .ZN(n7197) );
  INV_X1 U9669 ( .A(n8326), .ZN(n7199) );
  INV_X1 U9670 ( .A(n8302), .ZN(n7200) );
  NAND2_X1 U9671 ( .A1(n11772), .A2(n11773), .ZN(n7205) );
  AOI21_X1 U9672 ( .B1(n11743), .B2(n7204), .A(n6652), .ZN(n7202) );
  NOR2_X1 U9673 ( .A1(n10042), .A2(n10040), .ZN(n7203) );
  NAND2_X1 U9674 ( .A1(n14420), .A2(n7211), .ZN(n7210) );
  NOR2_X1 U9675 ( .A1(n6605), .A2(n7634), .ZN(n14244) );
  AOI21_X1 U9676 ( .B1(n8919), .B2(n6658), .A(n7220), .ZN(n7219) );
  XNOR2_X1 U9677 ( .A(n12790), .B(n14701), .ZN(n14698) );
  NAND2_X1 U9678 ( .A1(n6498), .A2(n11799), .ZN(n7230) );
  INV_X1 U9679 ( .A(n7232), .ZN(n11826) );
  NAND2_X1 U9680 ( .A1(n7236), .A2(n11034), .ZN(n7235) );
  INV_X1 U9681 ( .A(n11301), .ZN(n7236) );
  INV_X1 U9682 ( .A(n7237), .ZN(n11300) );
  XNOR2_X2 U9683 ( .A(n11587), .B(n15280), .ZN(n15266) );
  INV_X1 U9684 ( .A(n7248), .ZN(n11189) );
  INV_X1 U9685 ( .A(n7246), .ZN(n11028) );
  NOR2_X2 U9686 ( .A1(n11131), .A2(n11001), .ZN(n11130) );
  NAND2_X1 U9687 ( .A1(n11043), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7247) );
  AND2_X2 U9688 ( .A1(n12827), .A2(n12826), .ZN(n12843) );
  NAND3_X1 U9689 ( .A1(n7250), .A2(n7657), .A3(n7857), .ZN(n7673) );
  NAND2_X1 U9690 ( .A1(n13711), .A2(n7255), .ZN(n7253) );
  INV_X1 U9691 ( .A(n13713), .ZN(n7264) );
  NAND2_X1 U9692 ( .A1(n9932), .A2(n7267), .ZN(n7266) );
  NAND2_X1 U9693 ( .A1(n9937), .A2(n7630), .ZN(n7277) );
  NAND2_X1 U9694 ( .A1(n9937), .A2(n7271), .ZN(n7270) );
  NAND2_X1 U9695 ( .A1(n7277), .A2(n7276), .ZN(n13807) );
  OAI21_X1 U9696 ( .B1(n9924), .B2(n7286), .A(n7284), .ZN(n12189) );
  XNOR2_X2 U9697 ( .A(n15171), .B(n13551), .ZN(n7385) );
  NAND2_X1 U9698 ( .A1(n9014), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U9699 ( .A1(n8314), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8268) );
  INV_X1 U9700 ( .A(n7291), .ZN(n15291) );
  INV_X1 U9701 ( .A(n7292), .ZN(n11830) );
  NAND3_X1 U9702 ( .A1(n7294), .A2(n7293), .A3(n7296), .ZN(n7292) );
  NAND2_X1 U9703 ( .A1(n11610), .A2(n7297), .ZN(n7296) );
  INV_X1 U9704 ( .A(n11610), .ZN(n7295) );
  XNOR2_X2 U9705 ( .A(n7308), .B(P3_IR_REG_1__SCAN_IN), .ZN(n11041) );
  INV_X1 U9706 ( .A(n7314), .ZN(n12764) );
  NAND2_X1 U9707 ( .A1(n12639), .A2(n7320), .ZN(n7316) );
  INV_X1 U9708 ( .A(n12675), .ZN(n7333) );
  NAND2_X1 U9709 ( .A1(n12693), .A2(n10152), .ZN(n7342) );
  OAI211_X1 U9710 ( .C1(n12693), .C2(n7341), .A(n12696), .B(n7338), .ZN(n10179) );
  NAND2_X1 U9711 ( .A1(n12693), .A2(n7339), .ZN(n7338) );
  INV_X1 U9712 ( .A(n7344), .ZN(n7340) );
  NOR2_X1 U9713 ( .A1(n10153), .A2(n10151), .ZN(n7343) );
  NAND2_X1 U9714 ( .A1(n10153), .A2(n10151), .ZN(n7344) );
  INV_X1 U9715 ( .A(n10153), .ZN(n7345) );
  NAND2_X1 U9716 ( .A1(n11936), .A2(n7352), .ZN(n7351) );
  INV_X1 U9717 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U9718 ( .A1(n7618), .A2(n7368), .ZN(n7367) );
  AND2_X2 U9719 ( .A1(n13634), .A2(n13633), .ZN(n13635) );
  NAND2_X1 U9720 ( .A1(n9872), .A2(n7380), .ZN(n7378) );
  INV_X1 U9721 ( .A(n7385), .ZN(n7386) );
  XNOR2_X1 U9722 ( .A(n15158), .B(n7385), .ZN(n15162) );
  XNOR2_X1 U9723 ( .A(n15167), .B(n7385), .ZN(n15196) );
  AND2_X4 U9724 ( .A1(n10533), .A2(n10476), .ZN(n9767) );
  AND2_X1 U9725 ( .A1(n15065), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7400) );
  NOR2_X1 U9726 ( .A1(n15058), .A2(n15059), .ZN(n15057) );
  NAND2_X1 U9727 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n7402) );
  NAND2_X1 U9728 ( .A1(n9609), .A2(n7408), .ZN(n7407) );
  NAND2_X1 U9729 ( .A1(n9530), .A2(n7411), .ZN(n7410) );
  NAND2_X1 U9730 ( .A1(n9530), .A2(n9531), .ZN(n7417) );
  NAND2_X1 U9731 ( .A1(n7714), .A2(n7420), .ZN(n7422) );
  NAND2_X1 U9732 ( .A1(n7830), .A2(n7431), .ZN(n7430) );
  OAI21_X1 U9733 ( .B1(n7830), .B2(n7433), .A(n7431), .ZN(n7853) );
  AOI21_X1 U9734 ( .B1(n7431), .B2(n7433), .A(n6686), .ZN(n7429) );
  OAI21_X1 U9735 ( .B1(n7830), .B2(n7829), .A(n7828), .ZN(n7850) );
  AOI21_X1 U9736 ( .B1(n7829), .B2(n7828), .A(n6637), .ZN(n7434) );
  NAND2_X1 U9737 ( .A1(n9665), .A2(n9666), .ZN(n9664) );
  INV_X1 U9738 ( .A(n9659), .ZN(n7437) );
  NAND3_X1 U9739 ( .A1(n7889), .A2(n7874), .A3(P1_DATAO_REG_13__SCAN_IN), .ZN(
        n7890) );
  NAND2_X1 U9740 ( .A1(n7442), .A2(n10775), .ZN(n7875) );
  INV_X1 U9741 ( .A(n9644), .ZN(n7443) );
  NAND3_X1 U9742 ( .A1(n7075), .A2(n12398), .A3(n7448), .ZN(n7447) );
  NAND3_X1 U9743 ( .A1(n12938), .A2(n12972), .A3(n7070), .ZN(n7451) );
  NAND2_X1 U9744 ( .A1(n7452), .A2(n7455), .ZN(n9725) );
  NAND2_X1 U9745 ( .A1(n7454), .A2(n7453), .ZN(n7452) );
  INV_X1 U9746 ( .A(n9715), .ZN(n7454) );
  OAI21_X1 U9747 ( .B1(n9691), .B2(n9690), .A(n6671), .ZN(n7457) );
  INV_X1 U9748 ( .A(n9696), .ZN(n7458) );
  INV_X1 U9749 ( .A(n6919), .ZN(n7464) );
  NAND2_X1 U9750 ( .A1(n7460), .A2(n7461), .ZN(n12202) );
  NAND2_X1 U9751 ( .A1(n12148), .A2(n10262), .ZN(n7460) );
  INV_X1 U9752 ( .A(n13982), .ZN(n7467) );
  NAND2_X1 U9753 ( .A1(n13982), .A2(n14058), .ZN(n7465) );
  NAND2_X1 U9754 ( .A1(n10283), .A2(n7468), .ZN(n13938) );
  NAND2_X1 U9755 ( .A1(n14000), .A2(n14018), .ZN(n10314) );
  NAND2_X1 U9756 ( .A1(n14078), .A2(n7473), .ZN(n7471) );
  NAND2_X1 U9757 ( .A1(n7471), .A2(n7472), .ZN(n12595) );
  NAND2_X1 U9758 ( .A1(n14078), .A2(n12576), .ZN(n14079) );
  INV_X1 U9759 ( .A(n10252), .ZN(n7476) );
  INV_X1 U9760 ( .A(n8969), .ZN(n7487) );
  INV_X1 U9761 ( .A(n7492), .ZN(n9503) );
  NAND2_X1 U9762 ( .A1(n7497), .A2(n7498), .ZN(n7499) );
  NAND2_X1 U9763 ( .A1(n8387), .A2(n7503), .ZN(n7502) );
  NAND2_X1 U9764 ( .A1(n9351), .A2(n9352), .ZN(n9350) );
  INV_X1 U9765 ( .A(n9384), .ZN(n9387) );
  NAND2_X1 U9766 ( .A1(n8557), .A2(n7515), .ZN(n7511) );
  NAND2_X1 U9767 ( .A1(n8557), .A2(n8556), .ZN(n7514) );
  NAND3_X1 U9768 ( .A1(n9303), .A2(n9302), .A3(n6670), .ZN(n7519) );
  NAND2_X1 U9769 ( .A1(n13432), .A2(n7523), .ZN(n7522) );
  NAND2_X1 U9770 ( .A1(n7524), .A2(n7522), .ZN(n13457) );
  NAND2_X2 U9771 ( .A1(n8639), .A2(n12341), .ZN(n12349) );
  NAND2_X1 U9772 ( .A1(n11974), .A2(n7551), .ZN(n7547) );
  NAND2_X1 U9773 ( .A1(n7547), .A2(n7548), .ZN(n12120) );
  NAND2_X1 U9774 ( .A1(n11525), .A2(n7554), .ZN(n11770) );
  NAND3_X1 U9775 ( .A1(n7557), .A2(n7556), .A3(n10034), .ZN(n14919) );
  NAND2_X1 U9776 ( .A1(n7558), .A2(n7561), .ZN(n7556) );
  NAND2_X1 U9777 ( .A1(n10033), .A2(n7558), .ZN(n7557) );
  NAND2_X1 U9778 ( .A1(n14300), .A2(n7566), .ZN(n7562) );
  NAND2_X1 U9779 ( .A1(n7562), .A2(n7563), .ZN(n14267) );
  OAI21_X1 U9780 ( .B1(n11509), .B2(n7573), .A(n7570), .ZN(n7576) );
  NAND2_X1 U9781 ( .A1(n12159), .A2(n6548), .ZN(n7586) );
  NAND2_X1 U9782 ( .A1(n7590), .A2(n7588), .ZN(n8131) );
  OR2_X1 U9783 ( .A1(n15309), .A2(n14741), .ZN(n7593) );
  OAI21_X1 U9784 ( .B1(n12277), .B2(n7595), .A(n7594), .ZN(n13282) );
  NAND2_X1 U9785 ( .A1(n7598), .A2(n7600), .ZN(n13294) );
  INV_X1 U9786 ( .A(n12278), .ZN(n7599) );
  OAI21_X2 U9787 ( .B1(n12995), .B2(n6593), .A(n7606), .ZN(n12958) );
  NAND2_X1 U9788 ( .A1(n7613), .A2(n7612), .ZN(n9529) );
  NAND3_X1 U9789 ( .A1(n11227), .A2(n8118), .A3(n8119), .ZN(n11413) );
  AND2_X1 U9790 ( .A1(n11413), .A2(n8120), .ZN(n11461) );
  INV_X1 U9791 ( .A(n8616), .ZN(n8720) );
  NAND2_X1 U9792 ( .A1(n7644), .A2(n7642), .ZN(n8154) );
  INV_X1 U9793 ( .A(n10393), .ZN(n10403) );
  NAND2_X1 U9794 ( .A1(n7811), .A2(n7810), .ZN(n7814) );
  INV_X1 U9795 ( .A(n9650), .ZN(n9653) );
  NAND2_X1 U9796 ( .A1(n8210), .A2(n12350), .ZN(n15346) );
  OAI21_X1 U9797 ( .B1(n12533), .B2(n6643), .A(n9529), .ZN(n8153) );
  NAND2_X2 U9798 ( .A1(n8340), .A2(n8339), .ZN(n11259) );
  CLKBUF_X1 U9799 ( .A(n12202), .Z(n13990) );
  CLKBUF_X1 U9800 ( .A(n12277), .Z(n12278) );
  NAND2_X1 U9801 ( .A1(n14265), .A2(n7620), .ZN(n14250) );
  NAND2_X1 U9802 ( .A1(n8925), .A2(n12334), .ZN(n9015) );
  INV_X1 U9803 ( .A(n10081), .ZN(n10082) );
  OAI21_X1 U9804 ( .B1(n14444), .B2(n14942), .A(n10080), .ZN(n10081) );
  NAND2_X2 U9805 ( .A1(n8924), .A2(n14541), .ZN(n9417) );
  INV_X1 U9806 ( .A(n8152), .ZN(n12533) );
  OR2_X1 U9807 ( .A1(n12900), .A2(n13392), .ZN(n7615) );
  INV_X1 U9808 ( .A(n8369), .ZN(n8698) );
  AND2_X1 U9809 ( .A1(n9501), .A2(n9497), .ZN(n7616) );
  AND2_X1 U9810 ( .A1(n10195), .A2(n10194), .ZN(n7617) );
  AND2_X1 U9811 ( .A1(n12605), .A2(n12709), .ZN(n7619) );
  OR2_X1 U9812 ( .A1(n14293), .A2(n14113), .ZN(n7621) );
  AND2_X1 U9813 ( .A1(n8767), .A2(n11539), .ZN(n7622) );
  AND2_X1 U9814 ( .A1(n9791), .A2(n7633), .ZN(n7623) );
  OR2_X1 U9815 ( .A1(n12900), .A2(n13339), .ZN(n7625) );
  OR2_X1 U9816 ( .A1(n14259), .A2(n14111), .ZN(n7627) );
  INV_X1 U9817 ( .A(n13510), .ZN(n13468) );
  INV_X1 U9818 ( .A(n13853), .ZN(n9945) );
  OR2_X1 U9819 ( .A1(n8684), .A2(n10804), .ZN(n7628) );
  AND2_X1 U9820 ( .A1(n9695), .A2(n9694), .ZN(n7629) );
  INV_X1 U9821 ( .A(n11347), .ZN(n9850) );
  OR2_X1 U9822 ( .A1(n13668), .A2(n9936), .ZN(n7630) );
  INV_X1 U9823 ( .A(n15381), .ZN(n15326) );
  INV_X1 U9824 ( .A(n12889), .ZN(n12872) );
  AND2_X1 U9825 ( .A1(n13510), .A2(n9892), .ZN(n7632) );
  NAND2_X1 U9826 ( .A1(n15438), .A2(n15410), .ZN(n13339) );
  OR3_X1 U9827 ( .A1(n9790), .A2(n9789), .A3(n9788), .ZN(n7633) );
  NOR2_X1 U9828 ( .A1(n14450), .A2(n14111), .ZN(n7634) );
  INV_X1 U9829 ( .A(n14820), .ZN(n10067) );
  AND2_X1 U9830 ( .A1(n9165), .A2(n9164), .ZN(n7635) );
  AND4_X1 U9831 ( .A1(n13014), .A2(n12395), .A3(n13001), .A4(n12394), .ZN(
        n7636) );
  OR2_X1 U9832 ( .A1(n8882), .A2(n15163), .ZN(n13518) );
  INV_X1 U9833 ( .A(n13518), .ZN(n8883) );
  INV_X1 U9834 ( .A(n13520), .ZN(n12224) );
  INV_X1 U9835 ( .A(n15166), .ZN(n9588) );
  INV_X1 U9836 ( .A(n9625), .ZN(n9626) );
  MUX2_X1 U9837 ( .A(n14128), .B(n12010), .S(n9468), .Z(n9111) );
  INV_X1 U9838 ( .A(n9640), .ZN(n9641) );
  MUX2_X1 U9839 ( .A(n14127), .B(n15022), .S(n9468), .Z(n9124) );
  INV_X1 U9840 ( .A(n9651), .ZN(n9652) );
  AND2_X1 U9841 ( .A1(n12086), .A2(n9195), .ZN(n9196) );
  AND2_X1 U9842 ( .A1(n9224), .A2(n9223), .ZN(n9225) );
  MUX2_X1 U9843 ( .A(n14115), .B(n14472), .S(n9468), .Z(n9337) );
  INV_X1 U9844 ( .A(n9702), .ZN(n9703) );
  INV_X1 U9845 ( .A(n9397), .ZN(n9398) );
  NAND2_X1 U9846 ( .A1(n13611), .A2(n6542), .ZN(n9765) );
  OAI21_X1 U9847 ( .B1(n13611), .B2(n13614), .A(n9765), .ZN(n9766) );
  INV_X1 U9848 ( .A(n9728), .ZN(n9729) );
  INV_X1 U9849 ( .A(n11048), .ZN(n11046) );
  INV_X1 U9850 ( .A(n12463), .ZN(n8127) );
  INV_X1 U9851 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7640) );
  INV_X1 U9852 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9198) );
  INV_X1 U9853 ( .A(n11054), .ZN(n11033) );
  INV_X1 U9854 ( .A(n12766), .ZN(n12767) );
  NOR2_X1 U9855 ( .A1(n8114), .A2(n8113), .ZN(n8115) );
  INV_X1 U9856 ( .A(n10939), .ZN(n8403) );
  INV_X1 U9857 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8412) );
  INV_X1 U9858 ( .A(n12092), .ZN(n9923) );
  INV_X1 U9859 ( .A(n9893), .ZN(n9894) );
  INV_X1 U9860 ( .A(n11847), .ZN(n9856) );
  NAND2_X1 U9861 ( .A1(n11677), .A2(n11676), .ZN(n9902) );
  AND2_X1 U9862 ( .A1(n13956), .A2(n10349), .ZN(n14056) );
  INV_X1 U9863 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10705) );
  INV_X1 U9864 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U9865 ( .A1(n14375), .A2(n14381), .ZN(n14376) );
  NOR2_X1 U9866 ( .A1(n8645), .A2(SI_17_), .ZN(n8647) );
  NOR2_X1 U9867 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8913) );
  INV_X1 U9868 ( .A(n12363), .ZN(n8164) );
  AOI21_X1 U9869 ( .B1(n9575), .B2(n15326), .A(n9574), .ZN(n9576) );
  INV_X1 U9870 ( .A(n8341), .ZN(n8834) );
  INV_X1 U9871 ( .A(n11648), .ZN(n8493) );
  NAND2_X1 U9872 ( .A1(n13551), .A2(n11852), .ZN(n8279) );
  NOR2_X1 U9873 ( .A1(n8565), .A2(n8564), .ZN(n8585) );
  OR2_X1 U9874 ( .A1(n8413), .A2(n8412), .ZN(n8440) );
  NOR2_X1 U9875 ( .A1(n15164), .A2(n15199), .ZN(n11680) );
  OR2_X1 U9876 ( .A1(n12176), .A2(n8866), .ZN(n8867) );
  INV_X1 U9877 ( .A(n13981), .ZN(n10340) );
  INV_X1 U9878 ( .A(n14999), .ZN(n11658) );
  OR2_X1 U9879 ( .A1(n9269), .A2(n14070), .ZN(n9271) );
  OR2_X1 U9880 ( .A1(n9064), .A2(n13134), .ZN(n9080) );
  INV_X1 U9881 ( .A(n14327), .ZN(n9999) );
  AND2_X1 U9882 ( .A1(n9210), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9250) );
  NOR2_X1 U9883 ( .A1(n9099), .A2(n10705), .ZN(n9135) );
  OR2_X1 U9884 ( .A1(n9080), .A2(n9079), .ZN(n9099) );
  AND2_X1 U9885 ( .A1(n10413), .A2(n9523), .ZN(n10395) );
  NAND2_X1 U9886 ( .A1(n8453), .A2(SI_9_), .ZN(n8474) );
  NAND2_X1 U9887 ( .A1(n8012), .A2(n8011), .ZN(n8025) );
  NAND2_X1 U9888 ( .A1(n7951), .A2(n7950), .ZN(n7965) );
  OR2_X1 U9889 ( .A1(n12658), .A2(n7619), .ZN(n10144) );
  NAND2_X1 U9890 ( .A1(n7881), .A2(n7880), .ZN(n7898) );
  AND2_X1 U9891 ( .A1(n10123), .A2(n12713), .ZN(n10124) );
  INV_X1 U9892 ( .A(n11047), .ZN(n11027) );
  INV_X1 U9893 ( .A(n15274), .ZN(n15287) );
  AND3_X1 U9894 ( .A1(n7987), .A2(n7986), .A3(n7985), .ZN(n12686) );
  NAND2_X1 U9895 ( .A1(n7803), .A2(n7802), .ZN(n7822) );
  INV_X1 U9896 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7664) );
  INV_X1 U9897 ( .A(n15392), .ZN(n12551) );
  NAND2_X1 U9898 ( .A1(n12372), .A2(n12371), .ZN(n12380) );
  AND3_X1 U9899 ( .A1(n7837), .A2(n7836), .A3(n7835), .ZN(n15314) );
  AND3_X1 U9900 ( .A1(n13409), .A2(n13407), .A3(n9554), .ZN(n10157) );
  OR2_X1 U9901 ( .A1(n8835), .A2(n13426), .ZN(n8844) );
  INV_X1 U9902 ( .A(n13496), .ZN(n8658) );
  AND2_X1 U9903 ( .A1(n10532), .A2(n8897), .ZN(n13509) );
  AND2_X1 U9904 ( .A1(n8694), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8715) );
  OR2_X1 U9905 ( .A1(n8635), .A2(n12336), .ZN(n8654) );
  INV_X1 U9906 ( .A(n13611), .ZN(n13612) );
  INV_X1 U9907 ( .A(n9883), .ZN(n13677) );
  INV_X1 U9908 ( .A(n11923), .ZN(n12098) );
  NOR2_X1 U9909 ( .A1(n11852), .A2(n13607), .ZN(n9950) );
  NAND2_X1 U9910 ( .A1(n8855), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8232) );
  AND2_X1 U9911 ( .A1(n13992), .A2(n13989), .ZN(n10273) );
  XNOR2_X1 U9912 ( .A(n10256), .B(n10257), .ZN(n12002) );
  NAND2_X1 U9913 ( .A1(n10274), .A2(n10276), .ZN(n10277) );
  NOR2_X1 U9914 ( .A1(n9271), .A2(n13976), .ZN(n9291) );
  OR2_X1 U9915 ( .A1(n14862), .A2(n14151), .ZN(n14907) );
  AND2_X1 U9916 ( .A1(n10052), .A2(n9473), .ZN(n14402) );
  INV_X1 U9917 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n13041) );
  INV_X1 U9918 ( .A(n14052), .ZN(n14085) );
  INV_X1 U9919 ( .A(n11980), .ZN(n12079) );
  NAND2_X1 U9920 ( .A1(n14948), .A2(n14415), .ZN(n10685) );
  NAND2_X1 U9921 ( .A1(n8931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8932) );
  INV_X1 U9922 ( .A(n8308), .ZN(n8305) );
  OAI21_X1 U9923 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n14700), .A(n14587), .ZN(
        n14650) );
  INV_X1 U9924 ( .A(n12296), .ZN(n12698) );
  NAND2_X1 U9925 ( .A1(n7863), .A2(n7862), .ZN(n14730) );
  INV_X1 U9926 ( .A(n12706), .ZN(n12679) );
  NAND2_X1 U9927 ( .A1(n10168), .A2(n10167), .ZN(n12689) );
  INV_X1 U9928 ( .A(n15296), .ZN(n15279) );
  AND2_X1 U9929 ( .A1(n11038), .A2(n15255), .ZN(n15252) );
  OR2_X1 U9930 ( .A1(n15385), .A2(n15390), .ZN(n15353) );
  INV_X1 U9931 ( .A(n13339), .ZN(n10409) );
  AND3_X1 U9932 ( .A1(n11219), .A2(n8205), .A3(n9554), .ZN(n11217) );
  AND2_X1 U9933 ( .A1(n8210), .A2(n15392), .ZN(n15426) );
  XNOR2_X1 U9934 ( .A(n8175), .B(n8174), .ZN(n11023) );
  NAND2_X1 U9935 ( .A1(n7890), .A2(n7889), .ZN(n7893) );
  NAND2_X1 U9936 ( .A1(n8904), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13515) );
  AND2_X1 U9937 ( .A1(n8814), .A2(n8796), .ZN(n13685) );
  AND2_X1 U9938 ( .A1(n8892), .A2(n9809), .ZN(n13513) );
  AND4_X1 U9939 ( .A1(n8819), .A2(n8818), .A3(n8817), .A4(n8816), .ZN(n9936)
         );
  AND4_X1 U9940 ( .A1(n8780), .A2(n8779), .A3(n8778), .A4(n8777), .ZN(n9732)
         );
  OR2_X1 U9941 ( .A1(n10537), .A2(n10538), .ZN(n15135) );
  INV_X1 U9942 ( .A(n15129), .ZN(n15120) );
  AND2_X1 U9943 ( .A1(n10546), .A2(n10541), .ZN(n15141) );
  AOI21_X1 U9944 ( .B1(n11921), .B2(n9922), .A(n9921), .ZN(n12091) );
  OR3_X1 U9945 ( .A1(n11249), .A2(n11248), .A3(n11247), .ZN(n11254) );
  INV_X1 U9946 ( .A(n15182), .ZN(n11247) );
  AND2_X1 U9947 ( .A1(n9953), .A2(n9952), .ZN(n10404) );
  XNOR2_X1 U9948 ( .A(n8856), .B(P2_IR_REG_24__SCAN_IN), .ZN(n12105) );
  AND2_X1 U9949 ( .A1(n8544), .A2(n8581), .ZN(n13573) );
  INV_X1 U9950 ( .A(n14106), .ZN(n14082) );
  INV_X1 U9951 ( .A(n12071), .ZN(n9508) );
  AND4_X1 U9952 ( .A1(n9346), .A2(n9345), .A3(n9344), .A4(n9343), .ZN(n13949)
         );
  OR2_X1 U9953 ( .A1(n14862), .A2(n14857), .ZN(n14864) );
  INV_X1 U9954 ( .A(n14864), .ZN(n14898) );
  INV_X2 U9955 ( .A(n9436), .ZN(n9465) );
  OR2_X1 U9956 ( .A1(n9152), .A2(n13041), .ZN(n9185) );
  INV_X1 U9957 ( .A(n14268), .ZN(n14071) );
  INV_X1 U9958 ( .A(n14979), .ZN(n15025) );
  AND2_X1 U9959 ( .A1(n14966), .A2(n15013), .ZN(n14825) );
  AND2_X1 U9960 ( .A1(n10021), .A2(n10020), .ZN(n10687) );
  NAND2_X1 U9961 ( .A1(n10008), .A2(n10007), .ZN(n10504) );
  AND2_X1 U9962 ( .A1(n11060), .A2(n11059), .ZN(n15274) );
  INV_X1 U9963 ( .A(n12689), .ZN(n12700) );
  AOI21_X1 U9964 ( .B1(n12898), .B2(n7981), .A(n8168), .ZN(n11489) );
  INV_X1 U9965 ( .A(n15252), .ZN(n15298) );
  NAND2_X1 U9966 ( .A1(n11219), .A2(n11218), .ZN(n15376) );
  NAND2_X1 U9967 ( .A1(n11704), .A2(n15376), .ZN(n15396) );
  AND2_X1 U9968 ( .A1(n9557), .A2(n9556), .ZN(n15428) );
  INV_X2 U9969 ( .A(n15428), .ZN(n15430) );
  INV_X1 U9970 ( .A(SI_12_), .ZN(n10494) );
  INV_X1 U9971 ( .A(n11614), .ZN(n11812) );
  INV_X1 U9972 ( .A(n12722), .ZN(n11050) );
  NAND2_X1 U9973 ( .A1(n8377), .A2(n10917), .ZN(n10923) );
  INV_X1 U9974 ( .A(n9732), .ZN(n13527) );
  OR2_X1 U9975 ( .A1(n10546), .A2(P2_U3088), .ZN(n15144) );
  AND2_X1 U9976 ( .A1(n13774), .A2(n11254), .ZN(n15149) );
  INV_X1 U9977 ( .A(n15250), .ZN(n9959) );
  AND2_X2 U9978 ( .A1(n10404), .A2(n11247), .ZN(n15250) );
  OR3_X1 U9979 ( .A1(n13867), .A2(n13866), .A3(n13865), .ZN(n13907) );
  INV_X1 U9980 ( .A(n15242), .ZN(n15240) );
  NAND2_X1 U9981 ( .A1(n15187), .A2(n15176), .ZN(n15180) );
  NAND2_X1 U9982 ( .A1(n8869), .A2(n8868), .ZN(n15182) );
  INV_X1 U9983 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10998) );
  INV_X1 U9984 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10526) );
  INV_X1 U9985 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10460) );
  AOI21_X1 U9986 ( .B1(n14460), .B2(n14103), .A(n10401), .ZN(n10402) );
  AND2_X1 U9987 ( .A1(n10397), .A2(n12071), .ZN(n14101) );
  NAND2_X1 U9988 ( .A1(n10390), .A2(n10389), .ZN(n14106) );
  CLKBUF_X1 U9989 ( .A(P1_U4016), .Z(n14133) );
  INV_X1 U9990 ( .A(n14860), .ZN(n14912) );
  OR2_X1 U9991 ( .A1(n14942), .A2(n14677), .ZN(n14944) );
  NAND2_X1 U9992 ( .A1(n10505), .A2(n10025), .ZN(n14940) );
  AND2_X2 U9993 ( .A1(n10693), .A2(n10692), .ZN(n15045) );
  AND3_X2 U9994 ( .A1(n10693), .A2(n10781), .A3(n10687), .ZN(n15030) );
  INV_X1 U9995 ( .A(n15030), .ZN(n15029) );
  AND2_X1 U9996 ( .A1(n10514), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10511) );
  INV_X1 U9997 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10773) );
  INV_X2 U9998 ( .A(n12710), .ZN(P3_U3897) );
  NAND2_X1 U9999 ( .A1(n10403), .A2(n10402), .ZN(P1_U3225) );
  NAND2_X1 U10000 ( .A1(n7624), .A2(n10082), .ZN(P1_U3356) );
  INV_X1 U10001 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7642) );
  NAND2_X1 U10002 ( .A1(n8173), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7643) );
  INV_X1 U10003 ( .A(n7644), .ZN(n7645) );
  NAND2_X1 U10004 ( .A1(n7645), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7646) );
  MUX2_X1 U10005 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7646), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n7647) );
  NAND2_X1 U10006 ( .A1(n7647), .A2(n8154), .ZN(n11081) );
  NAND2_X1 U10007 ( .A1(n7648), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7649) );
  NOR2_X1 U10008 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n7653) );
  NAND4_X1 U10009 ( .A1(n7653), .A2(n7652), .A3(n7651), .A4(n7650), .ZN(n7656)
         );
  NAND4_X1 U10010 ( .A1(n7654), .A2(n7030), .A3(n7358), .A4(n7908), .ZN(n7655)
         );
  NAND2_X1 U10011 ( .A1(n7721), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7672) );
  AND2_X2 U10012 ( .A1(n7663), .A2(n7667), .ZN(n7736) );
  NAND2_X1 U10013 ( .A1(n7738), .A2(n7664), .ZN(n7753) );
  OR2_X1 U10014 ( .A1(n7738), .A2(n7664), .ZN(n7665) );
  AND2_X1 U10015 ( .A1(n7753), .A2(n7665), .ZN(n15360) );
  INV_X1 U10016 ( .A(n15360), .ZN(n7666) );
  NAND2_X1 U10017 ( .A1(n7981), .A2(n7666), .ZN(n7671) );
  NAND2_X1 U10018 ( .A1(n12360), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7670) );
  INV_X1 U10019 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n7668) );
  OR2_X1 U10020 ( .A1(n12363), .A2(n7668), .ZN(n7669) );
  NAND2_X1 U10021 ( .A1(n7673), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U10022 ( .A1(n7675), .A2(n13412), .ZN(n8169) );
  NAND2_X1 U10023 ( .A1(n10456), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U10024 ( .A1(n10478), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U10025 ( .A1(n10459), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7680) );
  INV_X1 U10026 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10483) );
  NAND2_X1 U10027 ( .A1(n10481), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7682) );
  XNOR2_X1 U10028 ( .A(n7762), .B(n7761), .ZN(n10470) );
  NAND2_X1 U10029 ( .A1(n7746), .A2(n10470), .ZN(n7692) );
  INV_X4 U10030 ( .A(n8945), .ZN(n10476) );
  OR2_X1 U10031 ( .A1(n12358), .A2(SI_5_), .ZN(n7691) );
  NOR2_X1 U10032 ( .A1(n7685), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7781) );
  INV_X1 U10033 ( .A(n7781), .ZN(n7689) );
  NAND2_X1 U10034 ( .A1(n7685), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7687) );
  MUX2_X1 U10035 ( .A(n7687), .B(P3_IR_REG_31__SCAN_IN), .S(n7686), .Z(n7688)
         );
  NAND2_X1 U10036 ( .A1(n7689), .A2(n7688), .ZN(n11054) );
  OR2_X1 U10037 ( .A1(n6507), .A2(n11033), .ZN(n7690) );
  NAND2_X1 U10038 ( .A1(n11454), .A2(n15358), .ZN(n12442) );
  NAND2_X1 U10039 ( .A1(n7721), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U10040 ( .A1(n7736), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7695) );
  INV_X1 U10041 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11009) );
  INV_X1 U10042 ( .A(SI_0_), .ZN(n10450) );
  INV_X1 U10043 ( .A(n7701), .ZN(n7698) );
  INV_X1 U10044 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U10045 ( .A1(n8249), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U10046 ( .A1(n7698), .A2(n7697), .ZN(n10449) );
  NAND2_X1 U10047 ( .A1(n7746), .A2(n10449), .ZN(n7700) );
  XOR2_X1 U10048 ( .A(n7702), .B(n7701), .Z(n10469) );
  INV_X1 U10049 ( .A(n11208), .ZN(n10863) );
  NAND2_X1 U10050 ( .A1(n7736), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7707) );
  INV_X1 U10051 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15431) );
  OR2_X1 U10052 ( .A1(n7755), .A2(n15431), .ZN(n7705) );
  NAND2_X1 U10053 ( .A1(n6547), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7712) );
  NAND2_X1 U10054 ( .A1(n7736), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7711) );
  NAND2_X1 U10055 ( .A1(n7721), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7710) );
  INV_X1 U10056 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11005) );
  XNOR2_X1 U10057 ( .A(n10459), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n7713) );
  XNOR2_X1 U10058 ( .A(n7714), .B(n7713), .ZN(n10453) );
  NAND2_X1 U10059 ( .A1(n7746), .A2(n10453), .ZN(n7719) );
  OR2_X1 U10060 ( .A1(n7729), .A2(SI_2_), .ZN(n7718) );
  INV_X1 U10061 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7715) );
  XNOR2_X2 U10062 ( .A(n7716), .B(n7715), .ZN(n11043) );
  OR2_X1 U10063 ( .A1(n6507), .A2(n11206), .ZN(n7717) );
  NAND2_X1 U10064 ( .A1(n6547), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7724) );
  INV_X1 U10065 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U10066 ( .A1(n7736), .A2(n7720), .ZN(n7723) );
  NAND2_X1 U10067 ( .A1(n7721), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7722) );
  AND3_X1 U10068 ( .A1(n7724), .A2(n7723), .A3(n7722), .ZN(n7726) );
  INV_X1 U10069 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11000) );
  OR2_X1 U10070 ( .A1(n7755), .A2(n11000), .ZN(n7725) );
  NAND2_X1 U10071 ( .A1(n7726), .A2(n7725), .ZN(n8116) );
  INV_X1 U10072 ( .A(n8116), .ZN(n15383) );
  XNOR2_X1 U10073 ( .A(n10460), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n7727) );
  XNOR2_X1 U10074 ( .A(n7728), .B(n7727), .ZN(n10455) );
  OR2_X1 U10075 ( .A1(n7729), .A2(SI_3_), .ZN(n7733) );
  INV_X1 U10076 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U10077 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6555), .ZN(n7730) );
  XNOR2_X1 U10078 ( .A(n7731), .B(n7730), .ZN(n11047) );
  OR2_X1 U10079 ( .A1(n6507), .A2(n11027), .ZN(n7732) );
  NAND2_X1 U10080 ( .A1(n15383), .A2(n15373), .ZN(n7735) );
  INV_X1 U10081 ( .A(n15373), .ZN(n11561) );
  NAND2_X1 U10082 ( .A1(n8116), .A2(n11561), .ZN(n12431) );
  NAND2_X1 U10083 ( .A1(n11098), .A2(n8114), .ZN(n11097) );
  NAND2_X1 U10084 ( .A1(n7721), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7743) );
  INV_X1 U10085 ( .A(n7736), .ZN(n8000) );
  AND2_X1 U10086 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7737) );
  NOR2_X1 U10087 ( .A1(n7738), .A2(n7737), .ZN(n15367) );
  INV_X1 U10088 ( .A(n15367), .ZN(n11155) );
  NAND2_X1 U10089 ( .A1(n7736), .A2(n11155), .ZN(n7742) );
  INV_X1 U10090 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11051) );
  OR2_X1 U10091 ( .A1(n7755), .A2(n11051), .ZN(n7740) );
  XNOR2_X1 U10092 ( .A(n7745), .B(n7744), .ZN(n10466) );
  NAND2_X1 U10093 ( .A1(n7746), .A2(n10466), .ZN(n7752) );
  OR2_X1 U10094 ( .A1(n7729), .A2(SI_4_), .ZN(n7751) );
  NAND2_X1 U10095 ( .A1(n7747), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7748) );
  MUX2_X1 U10096 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7748), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7749) );
  AND2_X1 U10097 ( .A1(n7749), .A2(n7685), .ZN(n12722) );
  OR2_X1 U10098 ( .A1(n6507), .A2(n12722), .ZN(n7750) );
  INV_X1 U10099 ( .A(n15365), .ZN(n11577) );
  NAND2_X1 U10100 ( .A1(n12718), .A2(n11577), .ZN(n12438) );
  NAND2_X1 U10101 ( .A1(n12437), .A2(n12438), .ZN(n11228) );
  INV_X1 U10102 ( .A(n15358), .ZN(n11581) );
  NAND2_X1 U10103 ( .A1(n12717), .A2(n11581), .ZN(n12441) );
  AND2_X2 U10104 ( .A1(n12442), .A2(n12441), .ZN(n12382) );
  NAND2_X1 U10105 ( .A1(n12360), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7760) );
  NAND2_X1 U10106 ( .A1(n7721), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U10107 ( .A1(n7753), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7754) );
  NAND2_X1 U10108 ( .A1(n7769), .A2(n7754), .ZN(n11446) );
  NAND2_X1 U10109 ( .A1(n7981), .A2(n11446), .ZN(n7758) );
  INV_X1 U10110 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n7756) );
  OR2_X1 U10111 ( .A1(n12363), .A2(n7756), .ZN(n7757) );
  NAND4_X1 U10112 ( .A1(n7760), .A2(n7759), .A3(n7758), .A4(n7757), .ZN(n12716) );
  INV_X1 U10113 ( .A(n12716), .ZN(n11557) );
  INV_X1 U10114 ( .A(SI_6_), .ZN(n10462) );
  INV_X1 U10115 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7763) );
  NAND2_X1 U10116 ( .A1(n7763), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U10117 ( .A1(n10489), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7765) );
  NAND2_X1 U10118 ( .A1(n7778), .A2(n7765), .ZN(n7776) );
  XNOR2_X1 U10119 ( .A(n7777), .B(n7776), .ZN(n10461) );
  NAND2_X1 U10120 ( .A1(n12370), .A2(n10461), .ZN(n7768) );
  OR2_X1 U10121 ( .A1(n7781), .A2(n13231), .ZN(n7766) );
  INV_X1 U10122 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7780) );
  XNOR2_X1 U10123 ( .A(n7766), .B(n7780), .ZN(n11592) );
  OR2_X1 U10124 ( .A1(n6507), .A2(n11592), .ZN(n7767) );
  OAI211_X1 U10125 ( .C1(n12358), .C2(n10462), .A(n7768), .B(n7767), .ZN(
        n11452) );
  NAND2_X1 U10126 ( .A1(n11557), .A2(n11452), .ZN(n12445) );
  INV_X1 U10127 ( .A(n11452), .ZN(n11748) );
  NAND2_X1 U10128 ( .A1(n12716), .A2(n11748), .ZN(n12446) );
  NAND2_X1 U10129 ( .A1(n12445), .A2(n12446), .ZN(n11460) );
  INV_X1 U10130 ( .A(n11460), .ZN(n12385) );
  NAND2_X1 U10131 ( .A1(n7721), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U10132 ( .A1(n12360), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7774) );
  AND2_X1 U10133 ( .A1(n7769), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7770) );
  OR2_X1 U10134 ( .A1(n7770), .A2(n7786), .ZN(n11705) );
  NAND2_X1 U10135 ( .A1(n7981), .A2(n11705), .ZN(n7773) );
  INV_X1 U10136 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n7771) );
  OR2_X1 U10137 ( .A1(n12363), .A2(n7771), .ZN(n7772) );
  NAND4_X1 U10138 ( .A1(n7775), .A2(n7774), .A3(n7773), .A4(n7772), .ZN(n12715) );
  INV_X1 U10139 ( .A(n12715), .ZN(n15338) );
  XNOR2_X1 U10140 ( .A(n7794), .B(n7793), .ZN(n10447) );
  NAND2_X1 U10141 ( .A1(n12370), .A2(n10447), .ZN(n7785) );
  OR2_X1 U10142 ( .A1(n12358), .A2(SI_7_), .ZN(n7784) );
  NAND2_X1 U10143 ( .A1(n7781), .A2(n7780), .ZN(n7796) );
  NAND2_X1 U10144 ( .A1(n7796), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7782) );
  XNOR2_X1 U10145 ( .A(n7782), .B(P3_IR_REG_7__SCAN_IN), .ZN(n15280) );
  OR2_X1 U10146 ( .A1(n6507), .A2(n15280), .ZN(n7783) );
  NAND2_X1 U10147 ( .A1(n15338), .A2(n15409), .ZN(n12450) );
  INV_X1 U10148 ( .A(n15409), .ZN(n11554) );
  NAND2_X1 U10149 ( .A1(n12715), .A2(n11554), .ZN(n12449) );
  NAND2_X1 U10150 ( .A1(n12450), .A2(n12449), .ZN(n11700) );
  INV_X1 U10151 ( .A(n11700), .ZN(n12454) );
  NAND2_X1 U10152 ( .A1(n12360), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U10153 ( .A1(n7721), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7791) );
  NOR2_X1 U10154 ( .A1(n7786), .A2(n11600), .ZN(n7787) );
  OR2_X1 U10155 ( .A1(n7803), .A2(n7787), .ZN(n15348) );
  NAND2_X1 U10156 ( .A1(n7981), .A2(n15348), .ZN(n7790) );
  INV_X1 U10157 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n7788) );
  OR2_X1 U10158 ( .A1(n12363), .A2(n7788), .ZN(n7789) );
  NAND4_X1 U10159 ( .A1(n7792), .A2(n7791), .A3(n7790), .A4(n7789), .ZN(n15325) );
  INV_X1 U10160 ( .A(n7810), .ZN(n7795) );
  XNOR2_X1 U10161 ( .A(n7811), .B(n7795), .ZN(n10467) );
  NAND2_X1 U10162 ( .A1(n12370), .A2(n10467), .ZN(n7800) );
  NAND2_X1 U10163 ( .A1(n7817), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7797) );
  XNOR2_X1 U10164 ( .A(n7797), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11614) );
  OR2_X1 U10165 ( .A1(n6507), .A2(n11812), .ZN(n7799) );
  INV_X1 U10166 ( .A(SI_8_), .ZN(n13233) );
  OR2_X1 U10167 ( .A1(n12358), .A2(n13233), .ZN(n7798) );
  NAND2_X1 U10168 ( .A1(n15325), .A2(n15347), .ZN(n12456) );
  NAND2_X1 U10169 ( .A1(n15335), .A2(n12456), .ZN(n7801) );
  INV_X1 U10170 ( .A(n15325), .ZN(n10110) );
  INV_X1 U10171 ( .A(n15347), .ZN(n8124) );
  NAND2_X1 U10172 ( .A1(n10110), .A2(n8124), .ZN(n12455) );
  NAND2_X1 U10173 ( .A1(n7721), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U10174 ( .A1(n12360), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7808) );
  OR2_X1 U10175 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  NAND2_X1 U10176 ( .A1(n7822), .A2(n7804), .ZN(n15331) );
  NAND2_X1 U10177 ( .A1(n7981), .A2(n15331), .ZN(n7807) );
  INV_X1 U10178 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n7805) );
  OR2_X1 U10179 ( .A1(n12363), .A2(n7805), .ZN(n7806) );
  NAND4_X1 U10180 ( .A1(n7809), .A2(n7808), .A3(n7807), .A4(n7806), .ZN(n15310) );
  NAND2_X1 U10181 ( .A1(n7812), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U10182 ( .A1(n10517), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U10183 ( .A1(n10518), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U10184 ( .A1(n7828), .A2(n7815), .ZN(n7829) );
  INV_X1 U10185 ( .A(n7829), .ZN(n7816) );
  XNOR2_X1 U10186 ( .A(n7830), .B(n7816), .ZN(n10465) );
  NAND2_X1 U10187 ( .A1(n12370), .A2(n10465), .ZN(n7821) );
  OR2_X1 U10188 ( .A1(n12358), .A2(SI_9_), .ZN(n7820) );
  NOR2_X1 U10189 ( .A1(n7817), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7833) );
  OR2_X1 U10190 ( .A1(n7833), .A2(n13231), .ZN(n7818) );
  XNOR2_X1 U10191 ( .A(n7818), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11829) );
  OR2_X1 U10192 ( .A1(n6507), .A2(n11829), .ZN(n7819) );
  XNOR2_X1 U10193 ( .A(n15310), .B(n15330), .ZN(n15322) );
  NAND2_X1 U10194 ( .A1(n15339), .A2(n15330), .ZN(n12459) );
  NAND2_X1 U10195 ( .A1(n7721), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U10196 ( .A1(n12360), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U10197 ( .A1(n7822), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U10198 ( .A1(n7839), .A2(n7823), .ZN(n15315) );
  NAND2_X1 U10199 ( .A1(n7981), .A2(n15315), .ZN(n7825) );
  INV_X1 U10200 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12028) );
  OR2_X1 U10201 ( .A1(n12363), .A2(n12028), .ZN(n7824) );
  NAND4_X1 U10202 ( .A1(n7827), .A2(n7826), .A3(n7825), .A4(n7824), .ZN(n15323) );
  XNOR2_X1 U10203 ( .A(n10526), .B(P2_DATAO_REG_10__SCAN_IN), .ZN(n7831) );
  XNOR2_X1 U10204 ( .A(n7850), .B(n7831), .ZN(n10475) );
  NAND2_X1 U10205 ( .A1(n12370), .A2(n10475), .ZN(n7837) );
  OR2_X1 U10206 ( .A1(n12358), .A2(SI_10_), .ZN(n7836) );
  INV_X1 U10207 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7832) );
  NAND2_X1 U10208 ( .A1(n7833), .A2(n7832), .ZN(n7846) );
  NAND2_X1 U10209 ( .A1(n7846), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7834) );
  XNOR2_X1 U10210 ( .A(n7834), .B(P3_IR_REG_10__SCAN_IN), .ZN(n12042) );
  OR2_X1 U10211 ( .A1(n6507), .A2(n12042), .ZN(n7835) );
  XNOR2_X1 U10212 ( .A(n15323), .B(n15314), .ZN(n12463) );
  INV_X1 U10213 ( .A(n15323), .ZN(n14740) );
  NAND2_X1 U10214 ( .A1(n14740), .A2(n15314), .ZN(n12465) );
  NAND2_X1 U10215 ( .A1(n12360), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10216 ( .A1(n7721), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10217 ( .A1(n7839), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10218 ( .A1(n7864), .A2(n7840), .ZN(n14742) );
  NAND2_X1 U10219 ( .A1(n7981), .A2(n14742), .ZN(n7843) );
  INV_X1 U10220 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n7841) );
  OR2_X1 U10221 ( .A1(n12363), .A2(n7841), .ZN(n7842) );
  NAND4_X1 U10222 ( .A1(n7845), .A2(n7844), .A3(n7843), .A4(n7842), .ZN(n15309) );
  OAI21_X1 U10223 ( .B1(n7846), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7848) );
  INV_X1 U10224 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7847) );
  XNOR2_X1 U10225 ( .A(n7848), .B(n7847), .ZN(n15289) );
  INV_X1 U10226 ( .A(n15289), .ZN(n12045) );
  OAI22_X1 U10227 ( .A1(n12358), .A2(SI_11_), .B1(n12045), .B2(n6507), .ZN(
        n7849) );
  INV_X1 U10228 ( .A(n7849), .ZN(n7852) );
  XNOR2_X1 U10229 ( .A(n7853), .B(n6686), .ZN(n10486) );
  NAND2_X1 U10230 ( .A1(n10486), .A2(n12370), .ZN(n7851) );
  NAND2_X1 U10231 ( .A1(n14728), .A2(n14741), .ZN(n12469) );
  INV_X1 U10232 ( .A(n14741), .ZN(n10419) );
  NAND2_X1 U10233 ( .A1(n15309), .A2(n10419), .ZN(n12472) );
  INV_X1 U10234 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U10235 ( .A1(n7854), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7855) );
  XNOR2_X1 U10236 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n7870) );
  XNOR2_X1 U10237 ( .A(n7871), .B(n7870), .ZN(n10492) );
  NAND2_X1 U10238 ( .A1(n10492), .A2(n12370), .ZN(n7863) );
  NOR2_X1 U10239 ( .A1(n7857), .A2(n13231), .ZN(n7858) );
  MUX2_X1 U10240 ( .A(n13231), .B(n7858), .S(P3_IR_REG_12__SCAN_IN), .Z(n7860)
         );
  OR2_X1 U10241 ( .A1(n7860), .A2(n7859), .ZN(n12755) );
  OAI22_X1 U10242 ( .A1(n7729), .A2(n10494), .B1(n6507), .B2(n12755), .ZN(
        n7861) );
  INV_X1 U10243 ( .A(n7861), .ZN(n7862) );
  NAND2_X1 U10244 ( .A1(n12360), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U10245 ( .A1(n9570), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7868) );
  AND2_X1 U10246 ( .A1(n7864), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7865) );
  OR2_X1 U10247 ( .A1(n7865), .A2(n7881), .ZN(n14731) );
  NAND2_X1 U10248 ( .A1(n7981), .A2(n14731), .ZN(n7867) );
  INV_X1 U10249 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12033) );
  OR2_X1 U10250 ( .A1(n12363), .A2(n12033), .ZN(n7866) );
  NAND4_X1 U10251 ( .A1(n7869), .A2(n7868), .A3(n7867), .A4(n7866), .ZN(n12714) );
  XNOR2_X1 U10252 ( .A(n14730), .B(n12714), .ZN(n14725) );
  NAND2_X1 U10253 ( .A1(n14739), .A2(n14730), .ZN(n12473) );
  NAND2_X1 U10254 ( .A1(n8517), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U10255 ( .A1(n7873), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U10256 ( .A1(n7890), .A2(n7875), .ZN(n10520) );
  NAND2_X1 U10257 ( .A1(n10520), .A2(n12370), .ZN(n7879) );
  OR2_X1 U10258 ( .A1(n7859), .A2(n13231), .ZN(n7876) );
  XNOR2_X1 U10259 ( .A(n7876), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12768) );
  OAI22_X1 U10260 ( .A1(n12358), .A2(SI_13_), .B1(n12768), .B2(n6507), .ZN(
        n7877) );
  INV_X1 U10261 ( .A(n7877), .ZN(n7878) );
  NAND2_X1 U10262 ( .A1(n7879), .A2(n7878), .ZN(n12405) );
  NAND2_X1 U10263 ( .A1(n12360), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U10264 ( .A1(n7721), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7886) );
  INV_X1 U10265 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7880) );
  OR2_X1 U10266 ( .A1(n7881), .A2(n7880), .ZN(n7882) );
  NAND2_X1 U10267 ( .A1(n7898), .A2(n7882), .ZN(n12215) );
  NAND2_X1 U10268 ( .A1(n7981), .A2(n12215), .ZN(n7885) );
  INV_X1 U10269 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n7883) );
  OR2_X1 U10270 ( .A1(n12363), .A2(n7883), .ZN(n7884) );
  NAND4_X1 U10271 ( .A1(n7887), .A2(n7886), .A3(n7885), .A4(n7884), .ZN(n12407) );
  XNOR2_X1 U10272 ( .A(n12405), .B(n12407), .ZN(n12391) );
  INV_X1 U10273 ( .A(n12391), .ZN(n12475) );
  OR2_X1 U10274 ( .A1(n12405), .A2(n12407), .ZN(n7888) );
  NAND2_X1 U10275 ( .A1(n10909), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U10276 ( .A1(n10908), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7891) );
  OAI21_X1 U10277 ( .B1(n7893), .B2(n7892), .A(n7906), .ZN(n10528) );
  NAND2_X1 U10278 ( .A1(n10528), .A2(n12370), .ZN(n7897) );
  NAND2_X1 U10279 ( .A1(n7658), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7894) );
  XNOR2_X1 U10280 ( .A(n7894), .B(P3_IR_REG_14__SCAN_IN), .ZN(n10527) );
  OAI22_X1 U10281 ( .A1(n12358), .A2(SI_14_), .B1(n10527), .B2(n6507), .ZN(
        n7895) );
  INV_X1 U10282 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U10283 ( .A1(n7897), .A2(n7896), .ZN(n12247) );
  NAND2_X1 U10284 ( .A1(n12360), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U10285 ( .A1(n9570), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U10286 ( .A1(n7898), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7899) );
  NAND2_X1 U10287 ( .A1(n7913), .A2(n7899), .ZN(n12248) );
  NAND2_X1 U10288 ( .A1(n7981), .A2(n12248), .ZN(n7902) );
  INV_X1 U10289 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n7900) );
  OR2_X1 U10290 ( .A1(n12363), .A2(n7900), .ZN(n7901) );
  NAND4_X1 U10291 ( .A1(n7904), .A2(n7903), .A3(n7902), .A4(n7901), .ZN(n12713) );
  NAND2_X1 U10292 ( .A1(n12247), .A2(n12713), .ZN(n12411) );
  NAND2_X1 U10293 ( .A1(n12412), .A2(n12411), .ZN(n12408) );
  INV_X1 U10294 ( .A(n12408), .ZN(n12476) );
  XNOR2_X1 U10295 ( .A(n11127), .B(P2_DATAO_REG_15__SCAN_IN), .ZN(n7921) );
  INV_X1 U10296 ( .A(n7921), .ZN(n7907) );
  XNOR2_X1 U10297 ( .A(n7922), .B(n7907), .ZN(n10633) );
  NAND2_X1 U10298 ( .A1(n10633), .A2(n12370), .ZN(n7912) );
  NAND2_X1 U10299 ( .A1(n6576), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7909) );
  XNOR2_X1 U10300 ( .A(n7909), .B(n7908), .ZN(n14701) );
  INV_X1 U10301 ( .A(n14701), .ZN(n12811) );
  OAI22_X1 U10302 ( .A1(n12358), .A2(SI_15_), .B1(n12811), .B2(n6507), .ZN(
        n7910) );
  INV_X1 U10303 ( .A(n7910), .ZN(n7911) );
  NAND2_X1 U10304 ( .A1(n9570), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7919) );
  INV_X1 U10305 ( .A(n7933), .ZN(n7915) );
  NAND2_X1 U10306 ( .A1(n7913), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U10307 ( .A1(n7915), .A2(n7914), .ZN(n12274) );
  NAND2_X1 U10308 ( .A1(n7981), .A2(n12274), .ZN(n7918) );
  NAND2_X1 U10309 ( .A1(n12360), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7917) );
  INV_X1 U10310 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14704) );
  OR2_X1 U10311 ( .A1(n12363), .A2(n14704), .ZN(n7916) );
  NAND4_X1 U10312 ( .A1(n7919), .A2(n7918), .A3(n7917), .A4(n7916), .ZN(n12712) );
  NAND2_X1 U10313 ( .A1(n13365), .A2(n12712), .ZN(n12480) );
  NAND2_X1 U10314 ( .A1(n12484), .A2(n12480), .ZN(n12390) );
  NAND2_X1 U10315 ( .A1(n11127), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U10316 ( .A1(n10893), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10317 ( .A1(n13109), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7924) );
  AND2_X1 U10318 ( .A1(n7939), .A2(n7924), .ZN(n7925) );
  OAI21_X1 U10319 ( .B1(n7926), .B2(n7925), .A(n7940), .ZN(n10696) );
  INV_X1 U10320 ( .A(SI_16_), .ZN(n10697) );
  NOR2_X1 U10321 ( .A1(n7927), .A2(n13231), .ZN(n7928) );
  MUX2_X1 U10322 ( .A(n13231), .B(n7928), .S(P3_IR_REG_16__SCAN_IN), .Z(n7930)
         );
  INV_X1 U10323 ( .A(n7944), .ZN(n7929) );
  OAI22_X1 U10324 ( .A1(n12358), .A2(n10697), .B1(n6507), .B2(n12825), .ZN(
        n7931) );
  INV_X1 U10325 ( .A(n7931), .ZN(n7932) );
  NAND2_X1 U10326 ( .A1(n9570), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U10327 ( .A1(n12360), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7937) );
  INV_X1 U10328 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12640) );
  NOR2_X1 U10329 ( .A1(n7933), .A2(n12640), .ZN(n7934) );
  OR2_X1 U10330 ( .A1(n7951), .A2(n7934), .ZN(n12641) );
  NAND2_X1 U10331 ( .A1(n7981), .A2(n12641), .ZN(n7936) );
  INV_X1 U10332 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12800) );
  OR2_X1 U10333 ( .A1(n12363), .A2(n12800), .ZN(n7935) );
  NAND4_X1 U10334 ( .A1(n7938), .A2(n7937), .A3(n7936), .A4(n7935), .ZN(n12711) );
  XNOR2_X1 U10335 ( .A(n13358), .B(n12711), .ZN(n12392) );
  INV_X1 U10336 ( .A(n12711), .ZN(n13296) );
  NAND2_X1 U10337 ( .A1(n13358), .A2(n13296), .ZN(n12485) );
  NAND2_X1 U10338 ( .A1(n10997), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U10339 ( .A1(n10998), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7941) );
  AND2_X1 U10340 ( .A1(n7957), .A2(n7941), .ZN(n7942) );
  OAI21_X1 U10341 ( .B1(n7943), .B2(n7942), .A(n7958), .ZN(n10762) );
  NAND2_X1 U10342 ( .A1(n10762), .A2(n12370), .ZN(n7949) );
  NAND2_X1 U10343 ( .A1(n7944), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7945) );
  MUX2_X1 U10344 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7945), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n7946) );
  NAND2_X1 U10345 ( .A1(n7946), .A2(n6570), .ZN(n12849) );
  INV_X1 U10346 ( .A(n12849), .ZN(n12860) );
  OAI22_X1 U10347 ( .A1(n12358), .A2(SI_17_), .B1(n12860), .B2(n6507), .ZN(
        n7947) );
  INV_X1 U10348 ( .A(n7947), .ZN(n7948) );
  NAND2_X1 U10349 ( .A1(n12360), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U10350 ( .A1(n9570), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7955) );
  INV_X1 U10351 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7950) );
  OR2_X1 U10352 ( .A1(n7951), .A2(n7950), .ZN(n7952) );
  NAND2_X1 U10353 ( .A1(n7965), .A2(n7952), .ZN(n13302) );
  NAND2_X1 U10354 ( .A1(n7981), .A2(n13302), .ZN(n7954) );
  INV_X1 U10355 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12824) );
  OR2_X1 U10356 ( .A1(n12363), .A2(n12824), .ZN(n7953) );
  NAND4_X1 U10357 ( .A1(n7956), .A2(n7955), .A3(n7954), .A4(n7953), .ZN(n13283) );
  NAND2_X1 U10358 ( .A1(n13357), .A2(n13283), .ZN(n12492) );
  INV_X1 U10359 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n13234) );
  INV_X1 U10360 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U10361 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n13234), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n11420), .ZN(n7959) );
  INV_X1 U10362 ( .A(n7959), .ZN(n7960) );
  XNOR2_X1 U10363 ( .A(n7972), .B(n7960), .ZN(n10803) );
  NAND2_X1 U10364 ( .A1(n10803), .A2(n12370), .ZN(n7964) );
  INV_X1 U10365 ( .A(SI_18_), .ZN(n10804) );
  NAND2_X1 U10366 ( .A1(n6570), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7961) );
  XNOR2_X1 U10367 ( .A(n7961), .B(n7358), .ZN(n12863) );
  OAI22_X1 U10368 ( .A1(n12358), .A2(n10804), .B1(n6507), .B2(n12863), .ZN(
        n7962) );
  INV_X1 U10369 ( .A(n7962), .ZN(n7963) );
  NAND2_X1 U10370 ( .A1(n12360), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10371 ( .A1(n9570), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U10372 ( .A1(n7965), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7966) );
  NAND2_X1 U10373 ( .A1(n7979), .A2(n7966), .ZN(n13289) );
  NAND2_X1 U10374 ( .A1(n7981), .A2(n13289), .ZN(n7968) );
  INV_X1 U10375 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12852) );
  OR2_X1 U10376 ( .A1(n12363), .A2(n12852), .ZN(n7967) );
  NAND4_X1 U10377 ( .A1(n7970), .A2(n7969), .A3(n7968), .A4(n7967), .ZN(n13010) );
  NAND2_X1 U10378 ( .A1(n13350), .A2(n13295), .ZN(n12494) );
  NAND2_X1 U10379 ( .A1(n13234), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U10380 ( .A1(n11420), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7973) );
  INV_X1 U10381 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11505) );
  INV_X1 U10382 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U10383 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11505), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n11503), .ZN(n7974) );
  INV_X1 U10384 ( .A(n7974), .ZN(n7975) );
  XNOR2_X1 U10385 ( .A(n7989), .B(n7975), .ZN(n10860) );
  NAND2_X1 U10386 ( .A1(n10860), .A2(n12370), .ZN(n7978) );
  INV_X1 U10387 ( .A(SI_19_), .ZN(n10861) );
  OAI22_X1 U10388 ( .A1(n7729), .A2(n10861), .B1(n12889), .B2(n6507), .ZN(
        n7976) );
  INV_X1 U10389 ( .A(n7976), .ZN(n7977) );
  AND2_X1 U10390 ( .A1(n7979), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7980) );
  OR2_X1 U10391 ( .A1(n7980), .A2(n7998), .ZN(n13016) );
  NAND2_X1 U10392 ( .A1(n13016), .A2(n7981), .ZN(n7987) );
  NAND2_X1 U10393 ( .A1(n12360), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n7984) );
  INV_X1 U10394 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n7982) );
  OR2_X1 U10395 ( .A1(n12363), .A2(n7982), .ZN(n7983) );
  AND2_X1 U10396 ( .A1(n7984), .A2(n7983), .ZN(n7986) );
  NAND2_X1 U10397 ( .A1(n9570), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U10398 ( .A1(n13400), .A2(n12686), .ZN(n12499) );
  NOR2_X1 U10399 ( .A1(n11505), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U10400 ( .A1(n11505), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7990) );
  INV_X1 U10401 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11763) );
  NAND2_X1 U10402 ( .A1(n11763), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8003) );
  INV_X1 U10403 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U10404 ( .A1(n11767), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7991) );
  AND2_X1 U10405 ( .A1(n8003), .A2(n7991), .ZN(n7993) );
  INV_X1 U10406 ( .A(n7993), .ZN(n7994) );
  NAND2_X1 U10407 ( .A1(n6754), .A2(n7994), .ZN(n7995) );
  AND2_X1 U10408 ( .A1(n8004), .A2(n7995), .ZN(n11080) );
  NAND2_X1 U10409 ( .A1(n11080), .A2(n12370), .ZN(n7997) );
  INV_X1 U10410 ( .A(SI_20_), .ZN(n13024) );
  OR2_X1 U10411 ( .A1(n12358), .A2(n13024), .ZN(n7996) );
  INV_X1 U10412 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13099) );
  INV_X1 U10413 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n13221) );
  NOR2_X1 U10414 ( .A1(n7998), .A2(n13221), .ZN(n7999) );
  OR2_X1 U10415 ( .A1(n8012), .A2(n7999), .ZN(n13003) );
  NAND2_X1 U10416 ( .A1(n13003), .A2(n7736), .ZN(n8002) );
  AOI22_X1 U10417 ( .A1(n12360), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n9570), 
        .B2(P3_REG2_REG_20__SCAN_IN), .ZN(n8001) );
  XNOR2_X1 U10418 ( .A(n13396), .B(n13011), .ZN(n13001) );
  INV_X1 U10419 ( .A(n13011), .ZN(n12615) );
  INV_X1 U10420 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11822) );
  NAND2_X1 U10421 ( .A1(n11822), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8018) );
  INV_X1 U10422 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11821) );
  NAND2_X1 U10423 ( .A1(n11821), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8005) );
  AND2_X1 U10424 ( .A1(n8018), .A2(n8005), .ZN(n8006) );
  OAI21_X1 U10425 ( .B1(n8007), .B2(n8006), .A(n8019), .ZN(n12351) );
  OR2_X1 U10426 ( .A1(n12351), .A2(n8008), .ZN(n8010) );
  INV_X1 U10427 ( .A(SI_21_), .ZN(n13055) );
  OR2_X1 U10428 ( .A1(n12358), .A2(n13055), .ZN(n8009) );
  INV_X1 U10429 ( .A(n13393), .ZN(n8016) );
  INV_X1 U10430 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13337) );
  INV_X1 U10431 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8011) );
  OR2_X1 U10432 ( .A1(n8012), .A2(n8011), .ZN(n8013) );
  NAND2_X1 U10433 ( .A1(n8025), .A2(n8013), .ZN(n12991) );
  NAND2_X1 U10434 ( .A1(n12991), .A2(n7981), .ZN(n8015) );
  AOI22_X1 U10435 ( .A1(n12360), .A2(P3_REG0_REG_21__SCAN_IN), .B1(n9570), 
        .B2(P3_REG2_REG_21__SCAN_IN), .ZN(n8014) );
  OAI211_X1 U10436 ( .C1(n12363), .C2(n13337), .A(n8015), .B(n8014), .ZN(
        n12998) );
  INV_X1 U10437 ( .A(n12998), .ZN(n12975) );
  NAND2_X1 U10438 ( .A1(n8016), .A2(n12975), .ZN(n12506) );
  NAND2_X1 U10439 ( .A1(n13393), .A2(n12998), .ZN(n12507) );
  INV_X1 U10440 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11987) );
  INV_X1 U10441 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8034) );
  AOI22_X1 U10442 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n11987), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n8034), .ZN(n8020) );
  INV_X1 U10443 ( .A(n8020), .ZN(n8021) );
  XNOR2_X1 U10444 ( .A(n8033), .B(n8021), .ZN(n11361) );
  NAND2_X1 U10445 ( .A1(n11361), .A2(n12370), .ZN(n8024) );
  INV_X1 U10446 ( .A(SI_22_), .ZN(n8022) );
  OR2_X1 U10447 ( .A1(n7729), .A2(n8022), .ZN(n8023) );
  NAND2_X1 U10448 ( .A1(n8025), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U10449 ( .A1(n8044), .A2(n8026), .ZN(n12980) );
  NAND2_X1 U10450 ( .A1(n12980), .A2(n7981), .ZN(n8031) );
  INV_X1 U10451 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13386) );
  NAND2_X1 U10452 ( .A1(n8164), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10453 ( .A1(n9570), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8027) );
  OAI211_X1 U10454 ( .C1(n8167), .C2(n13386), .A(n8028), .B(n8027), .ZN(n8029)
         );
  INV_X1 U10455 ( .A(n8029), .ZN(n8030) );
  NAND2_X1 U10456 ( .A1(n12979), .A2(n12625), .ZN(n12513) );
  NAND2_X1 U10457 ( .A1(n11987), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10458 ( .A1(n8034), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8035) );
  INV_X1 U10459 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10460 ( .A1(n8036), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8054) );
  INV_X1 U10461 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12073) );
  NAND2_X1 U10462 ( .A1(n12073), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10463 ( .A1(n8054), .A2(n8037), .ZN(n8039) );
  NAND2_X1 U10464 ( .A1(n8040), .A2(n8039), .ZN(n8041) );
  NAND2_X1 U10465 ( .A1(n8055), .A2(n8041), .ZN(n11537) );
  NAND2_X1 U10466 ( .A1(n11537), .A2(n12370), .ZN(n8043) );
  INV_X1 U10467 ( .A(SI_23_), .ZN(n11539) );
  OR2_X1 U10468 ( .A1(n7729), .A2(n11539), .ZN(n8042) );
  NAND2_X1 U10469 ( .A1(n8044), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U10470 ( .A1(n8059), .A2(n8045), .ZN(n12964) );
  NAND2_X1 U10471 ( .A1(n12964), .A2(n7736), .ZN(n8051) );
  INV_X1 U10472 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10473 ( .A1(n9570), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10474 ( .A1(n8164), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8046) );
  OAI211_X1 U10475 ( .C1(n8048), .C2(n8167), .A(n8047), .B(n8046), .ZN(n8049)
         );
  INV_X1 U10476 ( .A(n8049), .ZN(n8050) );
  NAND2_X1 U10477 ( .A1(n13383), .A2(n12976), .ZN(n8052) );
  INV_X1 U10478 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12602) );
  INV_X1 U10479 ( .A(n8067), .ZN(n8056) );
  XNOR2_X1 U10480 ( .A(n8056), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11905) );
  NAND2_X1 U10481 ( .A1(n11905), .A2(n12370), .ZN(n8058) );
  INV_X1 U10482 ( .A(SI_24_), .ZN(n11906) );
  OR2_X1 U10483 ( .A1(n12358), .A2(n11906), .ZN(n8057) );
  INV_X1 U10484 ( .A(n8074), .ZN(n8061) );
  NAND2_X1 U10485 ( .A1(n8059), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10486 ( .A1(n8061), .A2(n8060), .ZN(n12953) );
  NAND2_X1 U10487 ( .A1(n12953), .A2(n7981), .ZN(n8066) );
  INV_X1 U10488 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13378) );
  NAND2_X1 U10489 ( .A1(n8164), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U10490 ( .A1(n9570), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8062) );
  OAI211_X1 U10491 ( .C1(n8167), .C2(n13378), .A(n8063), .B(n8062), .ZN(n8064)
         );
  INV_X1 U10492 ( .A(n8064), .ZN(n8065) );
  OR2_X1 U10493 ( .A1(n12655), .A2(n12933), .ZN(n12521) );
  NAND2_X1 U10494 ( .A1(n12655), .A2(n12933), .ZN(n12525) );
  NAND2_X1 U10495 ( .A1(n12521), .A2(n12525), .ZN(n12945) );
  INV_X1 U10496 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U10497 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n12178), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n6736), .ZN(n8082) );
  INV_X1 U10498 ( .A(n8082), .ZN(n8070) );
  XNOR2_X1 U10499 ( .A(n8081), .B(n8070), .ZN(n11931) );
  NAND2_X1 U10500 ( .A1(n11931), .A2(n12370), .ZN(n8072) );
  INV_X1 U10501 ( .A(SI_25_), .ZN(n13160) );
  OR2_X1 U10502 ( .A1(n7729), .A2(n13160), .ZN(n8071) );
  INV_X1 U10503 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10504 ( .A1(n8074), .A2(n8073), .ZN(n8086) );
  OR2_X1 U10505 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  NAND2_X1 U10506 ( .A1(n8086), .A2(n8075), .ZN(n12941) );
  NAND2_X1 U10507 ( .A1(n12941), .A2(n7981), .ZN(n8080) );
  INV_X1 U10508 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13315) );
  NAND2_X1 U10509 ( .A1(n12360), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10510 ( .A1(n9570), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8076) );
  OAI211_X1 U10511 ( .C1(n13315), .C2(n12363), .A(n8077), .B(n8076), .ZN(n8078) );
  INV_X1 U10512 ( .A(n8078), .ZN(n8079) );
  INV_X1 U10513 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12259) );
  INV_X1 U10514 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U10515 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n12259), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n12256), .ZN(n8096) );
  INV_X1 U10516 ( .A(n8096), .ZN(n8083) );
  XNOR2_X1 U10517 ( .A(n8095), .B(n8083), .ZN(n12074) );
  NAND2_X1 U10518 ( .A1(n12074), .A2(n12370), .ZN(n8085) );
  INV_X1 U10519 ( .A(SI_26_), .ZN(n12076) );
  OR2_X1 U10520 ( .A1(n12358), .A2(n12076), .ZN(n8084) );
  NAND2_X1 U10521 ( .A1(n8086), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10522 ( .A1(n8100), .A2(n8087), .ZN(n12925) );
  NAND2_X1 U10523 ( .A1(n12925), .A2(n7981), .ZN(n8092) );
  INV_X1 U10524 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13370) );
  NAND2_X1 U10525 ( .A1(n8164), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10526 ( .A1(n9570), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8088) );
  OAI211_X1 U10527 ( .C1(n8167), .C2(n13370), .A(n8089), .B(n8088), .ZN(n8090)
         );
  INV_X1 U10528 ( .A(n8090), .ZN(n8091) );
  NAND2_X1 U10529 ( .A1(n8150), .A2(n12934), .ZN(n12401) );
  INV_X1 U10530 ( .A(n12913), .ZN(n8093) );
  NOR2_X1 U10531 ( .A1(n12917), .A2(n8093), .ZN(n8094) );
  NAND2_X1 U10532 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  INV_X1 U10533 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U10534 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13927), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n7419), .ZN(n9531) );
  XNOR2_X1 U10535 ( .A(n9530), .B(n7414), .ZN(n12329) );
  NAND2_X1 U10536 ( .A1(n12329), .A2(n12370), .ZN(n8099) );
  INV_X1 U10537 ( .A(SI_27_), .ZN(n12330) );
  OR2_X1 U10538 ( .A1(n12358), .A2(n12330), .ZN(n8098) );
  NOR2_X2 U10539 ( .A1(n8100), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8162) );
  INV_X1 U10540 ( .A(n8162), .ZN(n8102) );
  NAND2_X1 U10541 ( .A1(n8100), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U10542 ( .A1(n8102), .A2(n8101), .ZN(n12906) );
  NAND2_X1 U10543 ( .A1(n12906), .A2(n7736), .ZN(n8107) );
  INV_X1 U10544 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13367) );
  NAND2_X1 U10545 ( .A1(n8164), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8104) );
  NAND2_X1 U10546 ( .A1(n9570), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8103) );
  OAI211_X1 U10547 ( .C1(n8167), .C2(n13367), .A(n8104), .B(n8103), .ZN(n8105)
         );
  INV_X1 U10548 ( .A(n8105), .ZN(n8106) );
  NAND2_X1 U10549 ( .A1(n13368), .A2(n12921), .ZN(n8108) );
  NAND2_X1 U10550 ( .A1(n10087), .A2(n11209), .ZN(n8112) );
  NAND2_X1 U10551 ( .A1(n10863), .A2(n8111), .ZN(n10091) );
  NAND2_X1 U10552 ( .A1(n8112), .A2(n10091), .ZN(n15377) );
  NAND2_X1 U10553 ( .A1(n11103), .A2(n10877), .ZN(n11101) );
  INV_X1 U10554 ( .A(n11101), .ZN(n8113) );
  NAND2_X1 U10555 ( .A1(n11100), .A2(n8115), .ZN(n11105) );
  NAND2_X1 U10556 ( .A1(n15373), .A2(n12719), .ZN(n8117) );
  NAND2_X1 U10557 ( .A1(n12718), .A2(n15365), .ZN(n8118) );
  NAND2_X1 U10558 ( .A1(n11454), .A2(n11581), .ZN(n8120) );
  NAND2_X1 U10559 ( .A1(n12716), .A2(n11452), .ZN(n8121) );
  NAND2_X1 U10560 ( .A1(n11459), .A2(n8121), .ZN(n11701) );
  NAND2_X1 U10561 ( .A1(n11701), .A2(n11700), .ZN(n11699) );
  NAND2_X1 U10562 ( .A1(n12715), .A2(n15409), .ZN(n8122) );
  NAND2_X1 U10563 ( .A1(n11699), .A2(n8122), .ZN(n15337) );
  NAND2_X1 U10564 ( .A1(n10110), .A2(n15347), .ZN(n8123) );
  NAND2_X1 U10565 ( .A1(n15325), .A2(n8124), .ZN(n8125) );
  INV_X1 U10566 ( .A(n15330), .ZN(n12458) );
  NAND2_X1 U10567 ( .A1(n15339), .A2(n12458), .ZN(n8126) );
  NAND2_X1 U10568 ( .A1(n15323), .A2(n15314), .ZN(n8128) );
  AND2_X1 U10569 ( .A1(n15309), .A2(n14741), .ZN(n8129) );
  NAND2_X1 U10570 ( .A1(n14730), .A2(n12714), .ZN(n8130) );
  NAND2_X1 U10571 ( .A1(n8131), .A2(n8130), .ZN(n12212) );
  NAND2_X1 U10572 ( .A1(n12212), .A2(n12391), .ZN(n8132) );
  INV_X1 U10573 ( .A(n12407), .ZN(n14729) );
  OR2_X1 U10574 ( .A1(n12405), .A2(n14729), .ZN(n12410) );
  NAND2_X1 U10575 ( .A1(n8132), .A2(n12410), .ZN(n12243) );
  NAND2_X1 U10576 ( .A1(n12243), .A2(n12408), .ZN(n8135) );
  INV_X1 U10577 ( .A(n12247), .ZN(n8133) );
  NAND2_X1 U10578 ( .A1(n8133), .A2(n12713), .ZN(n8134) );
  NAND2_X1 U10579 ( .A1(n8135), .A2(n8134), .ZN(n12262) );
  NAND2_X1 U10580 ( .A1(n12262), .A2(n12390), .ZN(n8137) );
  INV_X1 U10581 ( .A(n12712), .ZN(n12245) );
  OR2_X1 U10582 ( .A1(n13365), .A2(n12245), .ZN(n8136) );
  NAND2_X1 U10583 ( .A1(n8137), .A2(n8136), .ZN(n12277) );
  INV_X1 U10584 ( .A(n13283), .ZN(n12644) );
  OR2_X1 U10585 ( .A1(n13357), .A2(n12644), .ZN(n8138) );
  OR2_X1 U10586 ( .A1(n13350), .A2(n13010), .ZN(n8139) );
  INV_X1 U10587 ( .A(n12686), .ZN(n13284) );
  NAND2_X1 U10588 ( .A1(n13400), .A2(n13284), .ZN(n8140) );
  NAND2_X1 U10589 ( .A1(n13396), .A2(n13011), .ZN(n8141) );
  NAND2_X1 U10590 ( .A1(n12507), .A2(n12506), .ZN(n12989) );
  NAND2_X1 U10591 ( .A1(n13393), .A2(n12975), .ZN(n8142) );
  NOR2_X1 U10592 ( .A1(n12979), .A2(n12987), .ZN(n8144) );
  NAND2_X1 U10593 ( .A1(n12979), .A2(n12987), .ZN(n8143) );
  NAND2_X1 U10594 ( .A1(n12958), .A2(n12519), .ZN(n8146) );
  NAND2_X1 U10595 ( .A1(n13383), .A2(n12709), .ZN(n8145) );
  AND2_X1 U10596 ( .A1(n12655), .A2(n12960), .ZN(n8147) );
  OR2_X2 U10597 ( .A1(n12930), .A2(n12938), .ZN(n12932) );
  NAND2_X1 U10598 ( .A1(n13375), .A2(n12920), .ZN(n8148) );
  NAND2_X1 U10599 ( .A1(n13372), .A2(n12934), .ZN(n8149) );
  NAND2_X1 U10600 ( .A1(n8150), .A2(n12708), .ZN(n8151) );
  INV_X1 U10601 ( .A(n8153), .ZN(n8172) );
  NAND2_X1 U10602 ( .A1(n12555), .A2(n12872), .ZN(n9552) );
  NAND2_X1 U10603 ( .A1(n8154), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8155) );
  MUX2_X1 U10604 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8155), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8156) );
  INV_X1 U10605 ( .A(n11081), .ZN(n9551) );
  NAND2_X1 U10606 ( .A1(n12414), .A2(n9551), .ZN(n12552) );
  NAND2_X1 U10607 ( .A1(n12350), .A2(n11081), .ZN(n8209) );
  XNOR2_X1 U10608 ( .A(n12555), .B(n8209), .ZN(n8158) );
  NAND2_X1 U10609 ( .A1(n12350), .A2(n12889), .ZN(n8157) );
  NAND2_X1 U10610 ( .A1(n8158), .A2(n8157), .ZN(n10162) );
  NAND2_X1 U10611 ( .A1(n11081), .A2(n12889), .ZN(n9550) );
  INV_X1 U10612 ( .A(n9550), .ZN(n12550) );
  AND2_X1 U10613 ( .A1(n15346), .A2(n12550), .ZN(n8159) );
  NAND2_X1 U10614 ( .A1(n10162), .A2(n8159), .ZN(n8160) );
  NAND2_X1 U10615 ( .A1(n9552), .A2(n9550), .ZN(n8208) );
  INV_X1 U10616 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8161) );
  NOR2_X1 U10617 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  INV_X1 U10618 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13162) );
  NAND2_X1 U10619 ( .A1(n9570), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10620 ( .A1(n8164), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8165) );
  OAI211_X1 U10621 ( .C1(n8167), .C2(n13162), .A(n8166), .B(n8165), .ZN(n8168)
         );
  NAND2_X1 U10622 ( .A1(n11036), .A2(n6507), .ZN(n10170) );
  INV_X1 U10623 ( .A(n10170), .ZN(n10172) );
  OAI22_X1 U10624 ( .A1(n6543), .A2(n15382), .B1(n12934), .B2(n15381), .ZN(
        n8171) );
  INV_X1 U10625 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8174) );
  NOR2_X1 U10626 ( .A1(n8176), .A2(n13231), .ZN(n8177) );
  MUX2_X1 U10627 ( .A(n13231), .B(n8177), .S(P3_IR_REG_25__SCAN_IN), .Z(n8180)
         );
  INV_X1 U10628 ( .A(n8178), .ZN(n8179) );
  NOR2_X1 U10629 ( .A1(n8180), .A2(n8179), .ZN(n8187) );
  NAND2_X1 U10630 ( .A1(n8178), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8181) );
  XNOR2_X1 U10631 ( .A(n8181), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8191) );
  INV_X1 U10632 ( .A(n8182), .ZN(n8183) );
  NAND2_X1 U10633 ( .A1(n8183), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8184) );
  MUX2_X1 U10634 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8184), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8185) );
  INV_X1 U10635 ( .A(n8185), .ZN(n8186) );
  NOR2_X1 U10636 ( .A1(n8186), .A2(n8176), .ZN(n8188) );
  NAND3_X1 U10637 ( .A1(n8187), .A2(n8191), .A3(n8188), .ZN(n10414) );
  INV_X1 U10638 ( .A(n8187), .ZN(n11933) );
  INV_X1 U10639 ( .A(n8188), .ZN(n11908) );
  XNOR2_X1 U10640 ( .A(n11908), .B(P3_B_REG_SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10641 ( .A1(n11933), .A2(n8189), .ZN(n8190) );
  INV_X1 U10642 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n13225) );
  NAND2_X1 U10643 ( .A1(n10716), .A2(n13225), .ZN(n8193) );
  INV_X1 U10644 ( .A(n8191), .ZN(n12077) );
  NAND2_X1 U10645 ( .A1(n11933), .A2(n12077), .ZN(n8192) );
  INV_X1 U10646 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n13224) );
  NAND2_X1 U10647 ( .A1(n10716), .A2(n13224), .ZN(n8195) );
  NAND2_X1 U10648 ( .A1(n12077), .A2(n11908), .ZN(n8194) );
  NAND2_X1 U10649 ( .A1(n8195), .A2(n8194), .ZN(n10083) );
  XNOR2_X1 U10650 ( .A(n13407), .B(n10083), .ZN(n8205) );
  NOR2_X1 U10651 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .ZN(
        n13255) );
  NOR4_X1 U10652 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .A3(
        P3_D_REG_26__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n8198) );
  NOR4_X1 U10653 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n8197) );
  NOR4_X1 U10654 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8196) );
  NAND4_X1 U10655 ( .A1(n13255), .A2(n8198), .A3(n8197), .A4(n8196), .ZN(n8204) );
  NOR4_X1 U10656 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8202) );
  NOR4_X1 U10657 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8201) );
  NOR4_X1 U10658 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8200) );
  NOR4_X1 U10659 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8199) );
  NAND4_X1 U10660 ( .A1(n8202), .A2(n8201), .A3(n8200), .A4(n8199), .ZN(n8203)
         );
  OAI21_X1 U10661 ( .B1(n8204), .B2(n8203), .A(n10716), .ZN(n9554) );
  NAND2_X1 U10662 ( .A1(n8206), .A2(n12547), .ZN(n11214) );
  NAND2_X1 U10663 ( .A1(n12530), .A2(n9550), .ZN(n11216) );
  NAND2_X1 U10664 ( .A1(n11214), .A2(n11216), .ZN(n8207) );
  NAND2_X1 U10665 ( .A1(n8207), .A2(n13407), .ZN(n8214) );
  NAND2_X1 U10666 ( .A1(n8208), .A2(n12350), .ZN(n8212) );
  AOI21_X1 U10667 ( .B1(n8210), .B2(n8209), .A(n13407), .ZN(n8211) );
  NAND2_X1 U10668 ( .A1(n8212), .A2(n8211), .ZN(n8213) );
  INV_X2 U10669 ( .A(n15439), .ZN(n15438) );
  INV_X1 U10670 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8215) );
  INV_X1 U10671 ( .A(n8216), .ZN(n8217) );
  NAND2_X1 U10672 ( .A1(n8218), .A2(n8217), .ZN(P3_U3486) );
  NOR2_X1 U10673 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8219) );
  NOR2_X1 U10674 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8223) );
  INV_X1 U10675 ( .A(n8518), .ZN(n8606) );
  NOR2_X2 U10676 ( .A1(n8237), .A2(n8606), .ZN(n8630) );
  XNOR2_X2 U10677 ( .A(n8226), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8271) );
  INV_X1 U10678 ( .A(n8231), .ZN(n8230) );
  NAND2_X1 U10679 ( .A1(n8227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8228) );
  XNOR2_X2 U10680 ( .A(n8232), .B(n8238), .ZN(n9586) );
  INV_X1 U10681 ( .A(n8233), .ZN(n8234) );
  NAND2_X1 U10682 ( .A1(n8234), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8235) );
  XNOR2_X2 U10683 ( .A(n8235), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13700) );
  NAND2_X2 U10684 ( .A1(n8236), .A2(n13607), .ZN(n9942) );
  NAND2_X4 U10685 ( .A1(n9942), .A2(n9804), .ZN(n8341) );
  NOR2_X1 U10686 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n8241) );
  NOR2_X1 U10687 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n8242) );
  INV_X1 U10688 ( .A(n8262), .ZN(n8245) );
  NOR2_X1 U10689 ( .A1(n8250), .A2(n10450), .ZN(n8251) );
  INV_X1 U10690 ( .A(n8251), .ZN(n8252) );
  NAND2_X1 U10691 ( .A1(n8253), .A2(n8252), .ZN(n8254) );
  AND2_X1 U10692 ( .A1(n8283), .A2(n8254), .ZN(n8946) );
  NAND2_X1 U10693 ( .A1(n9767), .A2(n8946), .ZN(n8260) );
  NAND2_X1 U10694 ( .A1(n8333), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10695 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8255) );
  INV_X1 U10696 ( .A(n8364), .ZN(n8256) );
  INV_X1 U10697 ( .A(n10553), .ZN(n15053) );
  NAND2_X1 U10698 ( .A1(n8669), .A2(n15053), .ZN(n8258) );
  XNOR2_X2 U10699 ( .A(n8341), .B(n15171), .ZN(n10899) );
  XNOR2_X2 U10700 ( .A(n8263), .B(P2_IR_REG_30__SCAN_IN), .ZN(n13913) );
  NAND2_X1 U10701 ( .A1(n8616), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8270) );
  AND2_X2 U10702 ( .A1(n13913), .A2(n8266), .ZN(n8392) );
  NAND2_X1 U10703 ( .A1(n8392), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8269) );
  INV_X1 U10704 ( .A(n8271), .ZN(n11820) );
  NAND2_X4 U10705 ( .A1(n10766), .A2(n11766), .ZN(n11852) );
  XNOR2_X1 U10706 ( .A(n10899), .B(n8279), .ZN(n10954) );
  NAND2_X1 U10707 ( .A1(n8616), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U10708 ( .A1(n8315), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U10709 ( .A1(n8392), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U10710 ( .A1(n10476), .A2(SI_0_), .ZN(n8276) );
  XNOR2_X1 U10711 ( .A(n8276), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13929) );
  NAND2_X1 U10712 ( .A1(n9589), .A2(n15166), .ZN(n10953) );
  OR2_X1 U10713 ( .A1(n8341), .A2(n15166), .ZN(n10947) );
  OAI21_X1 U10714 ( .B1(n13742), .B2(n10953), .A(n10947), .ZN(n8277) );
  INV_X1 U10715 ( .A(n8277), .ZN(n8278) );
  NAND2_X1 U10716 ( .A1(n10954), .A2(n8278), .ZN(n10900) );
  INV_X1 U10717 ( .A(n10899), .ZN(n8280) );
  NAND2_X1 U10718 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  NAND2_X1 U10719 ( .A1(n10900), .A2(n8281), .ZN(n8297) );
  OAI21_X1 U10720 ( .B1(n8284), .B2(SI_2_), .A(n8302), .ZN(n8286) );
  NAND2_X1 U10721 ( .A1(n8285), .A2(n8286), .ZN(n8289) );
  INV_X1 U10722 ( .A(n8286), .ZN(n8287) );
  AND2_X1 U10723 ( .A1(n8289), .A2(n8303), .ZN(n10457) );
  NAND2_X1 U10724 ( .A1(n10457), .A2(n9767), .ZN(n8292) );
  NOR2_X1 U10725 ( .A1(n8364), .A2(n8519), .ZN(n8290) );
  XNOR2_X1 U10726 ( .A(n8341), .B(n15199), .ZN(n8298) );
  NAND2_X1 U10727 ( .A1(n8616), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8296) );
  INV_X1 U10728 ( .A(n8392), .ZN(n8547) );
  NAND2_X1 U10729 ( .A1(n8392), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U10730 ( .A1(n8314), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8294) );
  NAND2_X1 U10731 ( .A1(n8315), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U10732 ( .A1(n13549), .A2(n11852), .ZN(n8299) );
  XNOR2_X1 U10733 ( .A(n8298), .B(n8299), .ZN(n10901) );
  NAND2_X1 U10734 ( .A1(n8297), .A2(n10901), .ZN(n10906) );
  INV_X1 U10735 ( .A(n8298), .ZN(n8300) );
  NAND2_X1 U10736 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  NAND2_X1 U10737 ( .A1(n10906), .A2(n8301), .ZN(n10790) );
  INV_X1 U10738 ( .A(n10790), .ZN(n8325) );
  NAND2_X1 U10739 ( .A1(n8304), .A2(SI_3_), .ZN(n8326) );
  OAI21_X1 U10740 ( .B1(n8304), .B2(SI_3_), .A(n8326), .ZN(n8306) );
  NAND2_X1 U10741 ( .A1(n8305), .A2(n7201), .ZN(n8309) );
  INV_X1 U10742 ( .A(n8306), .ZN(n8307) );
  NAND2_X1 U10743 ( .A1(n8309), .A2(n8327), .ZN(n10484) );
  OR2_X1 U10744 ( .A1(n10484), .A2(n8359), .ZN(n8313) );
  NAND2_X1 U10745 ( .A1(n6660), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8310) );
  MUX2_X1 U10746 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8310), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8311) );
  AOI22_X1 U10747 ( .A1(n8333), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8669), .B2(
        n10572), .ZN(n8312) );
  NAND2_X1 U10748 ( .A1(n8313), .A2(n8312), .ZN(n11574) );
  INV_X1 U10749 ( .A(n11574), .ZN(n15209) );
  INV_X1 U10750 ( .A(n8322), .ZN(n10828) );
  INV_X2 U10751 ( .A(n8720), .ZN(n9745) );
  NAND2_X1 U10752 ( .A1(n9745), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8319) );
  INV_X1 U10753 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U10754 ( .A1(n8392), .A2(n11568), .ZN(n8318) );
  NAND2_X1 U10755 ( .A1(n8314), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10756 ( .A1(n8369), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10757 ( .A1(n6898), .A2(n11852), .ZN(n8321) );
  INV_X1 U10758 ( .A(n8321), .ZN(n8320) );
  NAND2_X1 U10759 ( .A1(n10828), .A2(n8320), .ZN(n8347) );
  NAND2_X1 U10760 ( .A1(n8322), .A2(n8321), .ZN(n8323) );
  NAND2_X1 U10761 ( .A1(n8347), .A2(n8323), .ZN(n10789) );
  NAND2_X1 U10762 ( .A1(n8325), .A2(n8324), .ZN(n10787) );
  NAND2_X1 U10763 ( .A1(n8328), .A2(SI_4_), .ZN(n8352) );
  OAI21_X1 U10764 ( .B1(SI_4_), .B2(n8328), .A(n8352), .ZN(n8329) );
  INV_X1 U10765 ( .A(n8329), .ZN(n8330) );
  OR2_X1 U10766 ( .A1(n8331), .A2(n8330), .ZN(n8332) );
  AND2_X1 U10767 ( .A1(n8353), .A2(n8332), .ZN(n10472) );
  NAND2_X1 U10768 ( .A1(n10472), .A2(n9767), .ZN(n8340) );
  NAND2_X1 U10769 ( .A1(n8335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8334) );
  MUX2_X1 U10770 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8334), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8338) );
  INV_X1 U10771 ( .A(n8335), .ZN(n8337) );
  INV_X1 U10772 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U10773 ( .A1(n8337), .A2(n8336), .ZN(n8360) );
  NAND2_X1 U10774 ( .A1(n8338), .A2(n8360), .ZN(n10592) );
  INV_X1 U10775 ( .A(n10592), .ZN(n10574) );
  AOI22_X1 U10776 ( .A1(n8770), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8669), .B2(
        n10574), .ZN(n8339) );
  XNOR2_X1 U10777 ( .A(n11259), .B(n8341), .ZN(n10916) );
  NAND2_X1 U10778 ( .A1(n8369), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U10779 ( .A1(n8616), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8345) );
  NAND2_X1 U10780 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8371) );
  OAI21_X1 U10781 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8371), .ZN(n11257) );
  INV_X1 U10782 ( .A(n11257), .ZN(n8342) );
  NAND2_X1 U10783 ( .A1(n8392), .A2(n8342), .ZN(n8344) );
  NAND2_X1 U10784 ( .A1(n8314), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U10785 ( .A1(n13547), .A2(n11852), .ZN(n8349) );
  XNOR2_X1 U10786 ( .A(n10916), .B(n8349), .ZN(n10827) );
  AND2_X1 U10787 ( .A1(n10827), .A2(n8347), .ZN(n8348) );
  NAND2_X1 U10788 ( .A1(n10787), .A2(n8348), .ZN(n10826) );
  INV_X1 U10789 ( .A(n10916), .ZN(n8350) );
  NAND2_X1 U10790 ( .A1(n8350), .A2(n8349), .ZN(n8351) );
  NAND2_X1 U10791 ( .A1(n10826), .A2(n8351), .ZN(n8377) );
  MUX2_X1 U10792 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9323), .Z(n8354) );
  NAND2_X1 U10793 ( .A1(n8354), .A2(SI_5_), .ZN(n8382) );
  OAI21_X1 U10794 ( .B1(n8354), .B2(SI_5_), .A(n8382), .ZN(n8355) );
  INV_X1 U10795 ( .A(n8355), .ZN(n8356) );
  OR2_X1 U10796 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  OR2_X1 U10797 ( .A1(n10488), .A2(n8359), .ZN(n8368) );
  NAND2_X1 U10798 ( .A1(n8360), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8361) );
  MUX2_X1 U10799 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8361), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8366) );
  INV_X1 U10800 ( .A(n8607), .ZN(n8365) );
  AOI22_X1 U10801 ( .A1(n8770), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8669), .B2(
        n10670), .ZN(n8367) );
  NAND2_X1 U10802 ( .A1(n8368), .A2(n8367), .ZN(n11274) );
  XNOR2_X1 U10803 ( .A(n11274), .B(n8341), .ZN(n8378) );
  INV_X2 U10804 ( .A(n8698), .ZN(n9746) );
  NAND2_X1 U10805 ( .A1(n9746), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U10806 ( .A1(n6910), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8375) );
  INV_X1 U10807 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8370) );
  AND2_X1 U10808 ( .A1(n8371), .A2(n8370), .ZN(n8372) );
  NOR2_X1 U10809 ( .A1(n8393), .A2(n8372), .ZN(n11275) );
  NAND2_X1 U10810 ( .A1(n8587), .A2(n11275), .ZN(n8374) );
  NAND2_X1 U10811 ( .A1(n6545), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8373) );
  NAND4_X1 U10812 ( .A1(n8376), .A2(n8375), .A3(n8374), .A4(n8373), .ZN(n13546) );
  NAND2_X1 U10813 ( .A1(n13546), .A2(n11852), .ZN(n8379) );
  XNOR2_X1 U10814 ( .A(n8378), .B(n8379), .ZN(n10917) );
  INV_X1 U10815 ( .A(n8378), .ZN(n8380) );
  NAND2_X1 U10816 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  MUX2_X1 U10817 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9323), .Z(n8384) );
  NAND2_X1 U10818 ( .A1(n8384), .A2(SI_6_), .ZN(n8405) );
  OAI21_X1 U10819 ( .B1(n8384), .B2(SI_6_), .A(n8405), .ZN(n8385) );
  INV_X1 U10820 ( .A(n8385), .ZN(n8386) );
  OR2_X1 U10821 ( .A1(n8387), .A2(n8386), .ZN(n8388) );
  NAND2_X1 U10822 ( .A1(n8406), .A2(n8388), .ZN(n9043) );
  OR2_X1 U10823 ( .A1(n9043), .A2(n8359), .ZN(n8391) );
  OR2_X1 U10824 ( .A1(n8607), .A2(n8519), .ZN(n8389) );
  XNOR2_X1 U10825 ( .A(n8389), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U10826 ( .A1(n8770), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8669), .B2(
        n10752), .ZN(n8390) );
  XNOR2_X1 U10827 ( .A(n11689), .B(n8341), .ZN(n10984) );
  NAND2_X1 U10828 ( .A1(n8369), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10829 ( .A1(n6910), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10830 ( .A1(n8393), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8413) );
  OR2_X1 U10831 ( .A1(n8393), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8394) );
  AND2_X1 U10832 ( .A1(n8413), .A2(n8394), .ZN(n11688) );
  NAND2_X1 U10833 ( .A1(n8392), .A2(n11688), .ZN(n8396) );
  NAND2_X1 U10834 ( .A1(n6545), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8395) );
  NAND4_X1 U10835 ( .A1(n8398), .A2(n8397), .A3(n8396), .A4(n8395), .ZN(n13545) );
  AND2_X1 U10836 ( .A1(n13545), .A2(n11852), .ZN(n8399) );
  NAND2_X1 U10837 ( .A1(n10984), .A2(n8399), .ZN(n8404) );
  INV_X1 U10838 ( .A(n10984), .ZN(n8401) );
  INV_X1 U10839 ( .A(n8399), .ZN(n8400) );
  NAND2_X1 U10840 ( .A1(n8401), .A2(n8400), .ZN(n8402) );
  NAND2_X1 U10841 ( .A1(n8404), .A2(n8402), .ZN(n10939) );
  MUX2_X1 U10842 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9323), .Z(n8407) );
  NAND2_X1 U10843 ( .A1(n8407), .A2(SI_7_), .ZN(n8426) );
  XNOR2_X1 U10844 ( .A(n8425), .B(n8423), .ZN(n10495) );
  NAND2_X1 U10845 ( .A1(n10495), .A2(n9767), .ZN(n8411) );
  INV_X1 U10846 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10847 ( .A1(n8607), .A2(n8408), .ZN(n8432) );
  NAND2_X1 U10848 ( .A1(n8432), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8409) );
  XNOR2_X1 U10849 ( .A(n8409), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U10850 ( .A1(n8770), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8669), .B2(
        n10850), .ZN(n8410) );
  XNOR2_X1 U10851 ( .A(n15146), .B(n8341), .ZN(n8419) );
  NAND2_X1 U10852 ( .A1(n8369), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U10853 ( .A1(n6910), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8417) );
  NAND2_X1 U10854 ( .A1(n8413), .A2(n8412), .ZN(n8414) );
  AND2_X1 U10855 ( .A1(n8440), .A2(n8414), .ZN(n15148) );
  NAND2_X1 U10856 ( .A1(n8392), .A2(n15148), .ZN(n8416) );
  NAND2_X1 U10857 ( .A1(n6545), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8415) );
  NAND4_X1 U10858 ( .A1(n8418), .A2(n8417), .A3(n8416), .A4(n8415), .ZN(n13544) );
  AND2_X1 U10859 ( .A1(n13544), .A2(n11852), .ZN(n8420) );
  NAND2_X1 U10860 ( .A1(n8419), .A2(n8420), .ZN(n8446) );
  INV_X1 U10861 ( .A(n8419), .ZN(n11068) );
  INV_X1 U10862 ( .A(n8420), .ZN(n8421) );
  NAND2_X1 U10863 ( .A1(n11068), .A2(n8421), .ZN(n8422) );
  AND2_X1 U10864 ( .A1(n8446), .A2(n8422), .ZN(n10985) );
  INV_X1 U10865 ( .A(n8423), .ZN(n8424) );
  MUX2_X1 U10866 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10476), .Z(n8427) );
  NAND2_X1 U10867 ( .A1(n8427), .A2(SI_8_), .ZN(n8451) );
  OAI21_X1 U10868 ( .B1(SI_8_), .B2(n8427), .A(n8451), .ZN(n8428) );
  INV_X1 U10869 ( .A(n8428), .ZN(n8429) );
  OR2_X1 U10870 ( .A1(n8430), .A2(n8429), .ZN(n8431) );
  NAND2_X1 U10871 ( .A1(n8452), .A2(n8431), .ZN(n10502) );
  OR2_X1 U10872 ( .A1(n10502), .A2(n8359), .ZN(n8438) );
  NOR2_X1 U10873 ( .A1(n8432), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8435) );
  OR2_X1 U10874 ( .A1(n8435), .A2(n8519), .ZN(n8433) );
  MUX2_X1 U10875 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8433), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8436) );
  INV_X1 U10876 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U10877 ( .A1(n8435), .A2(n8434), .ZN(n8459) );
  AOI22_X1 U10878 ( .A1(n8770), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8669), .B2(
        n10966), .ZN(n8437) );
  NAND2_X1 U10879 ( .A1(n8369), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10880 ( .A1(n6910), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8444) );
  INV_X1 U10881 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10882 ( .A1(n8440), .A2(n8439), .ZN(n8441) );
  NAND2_X1 U10883 ( .A1(n8463), .A2(n8441), .ZN(n11075) );
  INV_X1 U10884 ( .A(n11075), .ZN(n11711) );
  NAND2_X1 U10885 ( .A1(n8587), .A2(n11711), .ZN(n8443) );
  NAND2_X1 U10886 ( .A1(n6545), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8442) );
  NAND4_X1 U10887 ( .A1(n8445), .A2(n8444), .A3(n8443), .A4(n8442), .ZN(n13543) );
  NAND2_X1 U10888 ( .A1(n13543), .A2(n11852), .ZN(n8448) );
  XNOR2_X1 U10889 ( .A(n11239), .B(n8448), .ZN(n11078) );
  AND2_X1 U10890 ( .A1(n11078), .A2(n8446), .ZN(n8447) );
  INV_X1 U10891 ( .A(n11239), .ZN(n8449) );
  NAND2_X1 U10892 ( .A1(n8449), .A2(n8448), .ZN(n8450) );
  NAND2_X1 U10893 ( .A1(n11070), .A2(n8450), .ZN(n8469) );
  MUX2_X1 U10894 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10476), .Z(n8453) );
  OAI21_X1 U10895 ( .B1(n8453), .B2(SI_9_), .A(n8474), .ZN(n8454) );
  INV_X1 U10896 ( .A(n8454), .ZN(n8455) );
  NAND2_X1 U10897 ( .A1(n8456), .A2(n8455), .ZN(n8475) );
  NAND2_X1 U10898 ( .A1(n8459), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8458) );
  MUX2_X1 U10899 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8458), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8460) );
  AOI22_X1 U10900 ( .A1(n8770), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8669), .B2(
        n11960), .ZN(n8461) );
  XNOR2_X1 U10901 ( .A(n11443), .B(n8341), .ZN(n8470) );
  NAND2_X1 U10902 ( .A1(n8369), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10903 ( .A1(n6910), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8467) );
  AND2_X1 U10904 ( .A1(n8463), .A2(n8462), .ZN(n8464) );
  NOR2_X1 U10905 ( .A1(n8502), .A2(n8464), .ZN(n11354) );
  NAND2_X1 U10906 ( .A1(n8587), .A2(n11354), .ZN(n8466) );
  NAND2_X1 U10907 ( .A1(n6545), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8465) );
  NAND4_X1 U10908 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(n13542) );
  NAND2_X1 U10909 ( .A1(n13542), .A2(n11852), .ZN(n8471) );
  XNOR2_X1 U10910 ( .A(n8470), .B(n8471), .ZN(n11240) );
  INV_X1 U10911 ( .A(n8470), .ZN(n8472) );
  NAND2_X1 U10912 ( .A1(n8472), .A2(n8471), .ZN(n8473) );
  MUX2_X1 U10913 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10476), .Z(n8476) );
  OAI21_X1 U10914 ( .B1(n8476), .B2(SI_10_), .A(n8494), .ZN(n8477) );
  INV_X1 U10915 ( .A(n8477), .ZN(n8478) );
  OR2_X1 U10916 ( .A1(n8479), .A2(n8478), .ZN(n8480) );
  NAND2_X1 U10917 ( .A1(n8496), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8481) );
  XNOR2_X1 U10918 ( .A(n8481), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15076) );
  AOI22_X1 U10919 ( .A1(n8770), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8669), 
        .B2(n15076), .ZN(n8482) );
  XNOR2_X1 U10920 ( .A(n15232), .B(n8341), .ZN(n8489) );
  NAND2_X1 U10921 ( .A1(n8369), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10922 ( .A1(n6910), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8487) );
  INV_X1 U10923 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8484) );
  XNOR2_X1 U10924 ( .A(n8502), .B(n8484), .ZN(n11642) );
  NAND2_X1 U10925 ( .A1(n8392), .A2(n11642), .ZN(n8486) );
  NAND2_X1 U10926 ( .A1(n6545), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8485) );
  NAND4_X1 U10927 ( .A1(n8488), .A2(n8487), .A3(n8486), .A4(n8485), .ZN(n13541) );
  AND2_X1 U10928 ( .A1(n13541), .A2(n11852), .ZN(n8490) );
  NAND2_X1 U10929 ( .A1(n8489), .A2(n8490), .ZN(n8508) );
  INV_X1 U10930 ( .A(n8489), .ZN(n11478) );
  INV_X1 U10931 ( .A(n8490), .ZN(n8491) );
  NAND2_X1 U10932 ( .A1(n11478), .A2(n8491), .ZN(n8492) );
  NAND2_X1 U10933 ( .A1(n8508), .A2(n8492), .ZN(n11648) );
  MUX2_X1 U10934 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10476), .Z(n8514) );
  XNOR2_X1 U10935 ( .A(n8512), .B(n8513), .ZN(n10596) );
  NAND2_X1 U10936 ( .A1(n10596), .A2(n9767), .ZN(n8499) );
  OAI21_X1 U10937 ( .B1(n8496), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8497) );
  XNOR2_X1 U10938 ( .A(n8497), .B(P2_IR_REG_11__SCAN_IN), .ZN(n15089) );
  AOI22_X1 U10939 ( .A1(n8669), .A2(n15089), .B1(n8770), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8498) );
  XNOR2_X1 U10940 ( .A(n11887), .B(n8341), .ZN(n11634) );
  NAND2_X1 U10941 ( .A1(n8369), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U10942 ( .A1(n6910), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8506) );
  NAND2_X1 U10943 ( .A1(n8502), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8500) );
  INV_X1 U10944 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U10945 ( .A1(n8500), .A2(n11481), .ZN(n8503) );
  AND2_X1 U10946 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n8501) );
  NAND2_X1 U10947 ( .A1(n8502), .A2(n8501), .ZN(n8527) );
  AND2_X1 U10948 ( .A1(n8503), .A2(n8527), .ZN(n11792) );
  NAND2_X1 U10949 ( .A1(n8392), .A2(n11792), .ZN(n8505) );
  NAND2_X1 U10950 ( .A1(n6545), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8504) );
  NAND4_X1 U10951 ( .A1(n8507), .A2(n8506), .A3(n8505), .A4(n8504), .ZN(n13540) );
  NAND2_X1 U10952 ( .A1(n13540), .A2(n11852), .ZN(n8509) );
  XNOR2_X1 U10953 ( .A(n11634), .B(n8509), .ZN(n11486) );
  NAND3_X1 U10954 ( .A1(n11476), .A2(n11486), .A3(n8508), .ZN(n11480) );
  INV_X1 U10955 ( .A(n11634), .ZN(n8510) );
  NAND2_X1 U10956 ( .A1(n8510), .A2(n8509), .ZN(n8511) );
  NAND2_X1 U10957 ( .A1(n11480), .A2(n8511), .ZN(n8533) );
  INV_X1 U10958 ( .A(n8514), .ZN(n8515) );
  INV_X1 U10959 ( .A(SI_11_), .ZN(n10485) );
  NAND2_X1 U10960 ( .A1(n8515), .A2(n10485), .ZN(n8516) );
  MUX2_X1 U10961 ( .A(n13062), .B(n8517), .S(n10476), .Z(n8540) );
  XNOR2_X1 U10962 ( .A(n8539), .B(n8538), .ZN(n10698) );
  NAND2_X1 U10963 ( .A1(n10698), .A2(n9767), .ZN(n8526) );
  AND2_X1 U10964 ( .A1(n8518), .A2(n8607), .ZN(n8522) );
  NOR2_X1 U10965 ( .A1(n8522), .A2(n8519), .ZN(n8520) );
  MUX2_X1 U10966 ( .A(n8519), .B(n8520), .S(P2_IR_REG_12__SCAN_IN), .Z(n8524)
         );
  INV_X1 U10967 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U10968 ( .A1(n8522), .A2(n8521), .ZN(n8543) );
  INV_X1 U10969 ( .A(n8543), .ZN(n8523) );
  NOR2_X1 U10970 ( .A1(n8524), .A2(n8523), .ZN(n13560) );
  AOI22_X1 U10971 ( .A1(n8770), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8669), 
        .B2(n13560), .ZN(n8525) );
  XNOR2_X1 U10972 ( .A(n11855), .B(n8341), .ZN(n8534) );
  NAND2_X1 U10973 ( .A1(n8369), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U10974 ( .A1(n6910), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8531) );
  INV_X1 U10975 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n13133) );
  NAND2_X1 U10976 ( .A1(n8527), .A2(n13133), .ZN(n8528) );
  AND2_X1 U10977 ( .A1(n8565), .A2(n8528), .ZN(n11854) );
  NAND2_X1 U10978 ( .A1(n8587), .A2(n11854), .ZN(n8530) );
  NAND2_X1 U10979 ( .A1(n6545), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8529) );
  NAND4_X1 U10980 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n13539) );
  NAND2_X1 U10981 ( .A1(n13539), .A2(n11852), .ZN(n8535) );
  XNOR2_X1 U10982 ( .A(n8534), .B(n8535), .ZN(n11635) );
  INV_X1 U10983 ( .A(n8534), .ZN(n8536) );
  NAND2_X1 U10984 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  NAND2_X1 U10985 ( .A1(n8540), .A2(n10494), .ZN(n8541) );
  MUX2_X1 U10986 ( .A(n10773), .B(n10775), .S(n10476), .Z(n8558) );
  XNOR2_X1 U10987 ( .A(n8557), .B(n8556), .ZN(n10772) );
  NAND2_X1 U10988 ( .A1(n10772), .A2(n9767), .ZN(n8546) );
  NAND2_X1 U10989 ( .A1(n8543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8542) );
  MUX2_X1 U10990 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8542), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8544) );
  OR2_X1 U10991 ( .A1(n8543), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8581) );
  AOI22_X1 U10992 ( .A1(n8770), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8669), 
        .B2(n13573), .ZN(n8545) );
  XNOR2_X1 U10993 ( .A(n14782), .B(n8341), .ZN(n12307) );
  NAND2_X1 U10994 ( .A1(n6910), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8551) );
  XNOR2_X1 U10995 ( .A(n8565), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n12017) );
  NAND2_X1 U10996 ( .A1(n8587), .A2(n12017), .ZN(n8550) );
  NAND2_X1 U10997 ( .A1(n6545), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10998 ( .A1(n8369), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8548) );
  NAND4_X1 U10999 ( .A1(n8551), .A2(n8550), .A3(n8549), .A4(n8548), .ZN(n13538) );
  AND2_X1 U11000 ( .A1(n13538), .A2(n11852), .ZN(n8552) );
  NAND2_X1 U11001 ( .A1(n12307), .A2(n8552), .ZN(n8571) );
  INV_X1 U11002 ( .A(n12307), .ZN(n8554) );
  INV_X1 U11003 ( .A(n8552), .ZN(n8553) );
  NAND2_X1 U11004 ( .A1(n8554), .A2(n8553), .ZN(n8555) );
  NAND2_X1 U11005 ( .A1(n8571), .A2(n8555), .ZN(n11862) );
  INV_X1 U11006 ( .A(SI_13_), .ZN(n10521) );
  NAND2_X1 U11007 ( .A1(n8558), .A2(n10521), .ZN(n8559) );
  MUX2_X1 U11008 ( .A(n10909), .B(n10908), .S(n10476), .Z(n8596) );
  NAND2_X1 U11009 ( .A1(n9168), .A2(n9767), .ZN(n8562) );
  NAND2_X1 U11010 ( .A1(n8581), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8560) );
  XNOR2_X1 U11011 ( .A(n8560), .B(P2_IR_REG_14__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U11012 ( .A1(n8770), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8669), 
        .B2(n15101), .ZN(n8561) );
  INV_X1 U11013 ( .A(n8565), .ZN(n8563) );
  AOI21_X1 U11014 ( .B1(n8563), .B2(P2_REG3_REG_13__SCAN_IN), .A(
        P2_REG3_REG_14__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U11015 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n8564) );
  OR2_X1 U11016 ( .A1(n8566), .A2(n8585), .ZN(n12311) );
  INV_X1 U11017 ( .A(n12311), .ZN(n11925) );
  NAND2_X1 U11018 ( .A1(n11925), .A2(n8587), .ZN(n8570) );
  NAND2_X1 U11019 ( .A1(n9746), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U11020 ( .A1(n9745), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U11021 ( .A1(n6545), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8567) );
  NAND4_X1 U11022 ( .A1(n8570), .A2(n8569), .A3(n8568), .A4(n8567), .ZN(n13537) );
  NAND2_X1 U11023 ( .A1(n13537), .A2(n11852), .ZN(n8573) );
  XNOR2_X1 U11024 ( .A(n8574), .B(n8573), .ZN(n12314) );
  INV_X1 U11025 ( .A(n8571), .ZN(n8572) );
  NAND2_X1 U11026 ( .A1(n8574), .A2(n8573), .ZN(n8575) );
  INV_X1 U11027 ( .A(n8576), .ZN(n8578) );
  INV_X1 U11028 ( .A(n8596), .ZN(n8599) );
  INV_X1 U11029 ( .A(n8598), .ZN(n8577) );
  OAI22_X1 U11030 ( .A1(n8578), .A2(n8599), .B1(n8577), .B2(SI_14_), .ZN(n8580) );
  MUX2_X1 U11031 ( .A(n11128), .B(n11127), .S(n10476), .Z(n8600) );
  XNOR2_X1 U11032 ( .A(n8600), .B(SI_15_), .ZN(n8579) );
  XNOR2_X1 U11033 ( .A(n8580), .B(n8579), .ZN(n11126) );
  NAND2_X1 U11034 ( .A1(n11126), .A2(n9767), .ZN(n8584) );
  OAI21_X1 U11035 ( .B1(n8581), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8582) );
  XNOR2_X1 U11036 ( .A(n8582), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15112) );
  AOI22_X1 U11037 ( .A1(n8770), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8669), 
        .B2(n15112), .ZN(n8583) );
  XNOR2_X1 U11038 ( .A(n12109), .B(n8834), .ZN(n8592) );
  NOR2_X1 U11039 ( .A1(n8585), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8586) );
  OR2_X1 U11040 ( .A1(n8614), .A2(n8586), .ZN(n12112) );
  NAND2_X1 U11041 ( .A1(n8369), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U11042 ( .A1(n9745), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8588) );
  AND2_X1 U11043 ( .A1(n8589), .A2(n8588), .ZN(n8591) );
  NAND2_X1 U11044 ( .A1(n6545), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8590) );
  OAI211_X1 U11045 ( .C1(n12112), .C2(n8547), .A(n8591), .B(n8590), .ZN(n13536) );
  INV_X1 U11046 ( .A(n13536), .ZN(n12107) );
  OR2_X1 U11047 ( .A1(n8593), .A2(n8592), .ZN(n8594) );
  INV_X1 U11048 ( .A(SI_14_), .ZN(n13168) );
  INV_X1 U11049 ( .A(n8600), .ZN(n8595) );
  NAND2_X1 U11050 ( .A1(n8595), .A2(SI_15_), .ZN(n8601) );
  OAI21_X1 U11051 ( .B1(n8596), .B2(n13168), .A(n8601), .ZN(n8597) );
  NOR2_X1 U11052 ( .A1(n8599), .A2(SI_14_), .ZN(n8602) );
  INV_X1 U11053 ( .A(SI_15_), .ZN(n10634) );
  AOI22_X1 U11054 ( .A1(n8602), .A2(n8601), .B1(n8600), .B2(n10634), .ZN(n8603) );
  MUX2_X1 U11055 ( .A(n10893), .B(n13109), .S(n10476), .Z(n8624) );
  XNOR2_X1 U11056 ( .A(n8623), .B(n8622), .ZN(n10891) );
  NAND2_X1 U11057 ( .A1(n10891), .A2(n9767), .ZN(n8613) );
  INV_X1 U11058 ( .A(n8604), .ZN(n8605) );
  NOR2_X1 U11059 ( .A1(n8606), .A2(n8605), .ZN(n8608) );
  NAND2_X1 U11060 ( .A1(n8608), .A2(n8607), .ZN(n8610) );
  NAND2_X1 U11061 ( .A1(n8610), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8609) );
  MUX2_X1 U11062 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8609), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8611) );
  OR2_X1 U11063 ( .A1(n8610), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8628) );
  AND2_X1 U11064 ( .A1(n8611), .A2(n8628), .ZN(n15125) );
  AOI22_X1 U11065 ( .A1(n8770), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8669), 
        .B2(n15125), .ZN(n8612) );
  XNOR2_X1 U11066 ( .A(n13869), .B(n8341), .ZN(n8619) );
  OR2_X1 U11067 ( .A1(n8614), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U11068 ( .A1(n8635), .A2(n8615), .ZN(n12138) );
  AOI22_X1 U11069 ( .A1(n9746), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n9745), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U11070 ( .A1(n6545), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8617) );
  OAI211_X1 U11071 ( .C1(n12138), .C2(n8547), .A(n8618), .B(n8617), .ZN(n13535) );
  NAND2_X1 U11072 ( .A1(n13535), .A2(n11852), .ZN(n8620) );
  XNOR2_X1 U11073 ( .A(n8619), .B(n8620), .ZN(n12222) );
  INV_X1 U11074 ( .A(n8619), .ZN(n12344) );
  NAND2_X1 U11075 ( .A1(n12344), .A2(n8620), .ZN(n8621) );
  NAND2_X1 U11076 ( .A1(n12221), .A2(n8621), .ZN(n8639) );
  NAND2_X1 U11077 ( .A1(n8624), .A2(n10697), .ZN(n8625) );
  MUX2_X1 U11078 ( .A(n10997), .B(n10998), .S(n10476), .Z(n8644) );
  XNOR2_X1 U11079 ( .A(n8644), .B(SI_17_), .ZN(n8627) );
  XNOR2_X1 U11080 ( .A(n8648), .B(n8627), .ZN(n10996) );
  NAND2_X1 U11081 ( .A1(n10996), .A2(n9767), .ZN(n8634) );
  NAND2_X1 U11082 ( .A1(n8628), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8629) );
  MUX2_X1 U11083 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8629), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8632) );
  INV_X1 U11084 ( .A(n8631), .ZN(n8649) );
  NAND2_X1 U11085 ( .A1(n8632), .A2(n8649), .ZN(n13587) );
  INV_X1 U11086 ( .A(n13587), .ZN(n15140) );
  AOI22_X1 U11087 ( .A1(n8770), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8669), 
        .B2(n15140), .ZN(n8633) );
  XNOR2_X1 U11088 ( .A(n12340), .B(n8341), .ZN(n8640) );
  INV_X1 U11089 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U11090 ( .A1(n8635), .A2(n12336), .ZN(n8636) );
  NAND2_X1 U11091 ( .A1(n8654), .A2(n8636), .ZN(n12335) );
  AOI22_X1 U11092 ( .A1(n9746), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n6910), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U11093 ( .A1(n6545), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8637) );
  OAI211_X1 U11094 ( .C1(n12335), .C2(n8547), .A(n8638), .B(n8637), .ZN(n13534) );
  NAND2_X1 U11095 ( .A1(n13534), .A2(n11852), .ZN(n8641) );
  XNOR2_X1 U11096 ( .A(n8640), .B(n8641), .ZN(n12341) );
  INV_X1 U11097 ( .A(n8640), .ZN(n8642) );
  NAND2_X1 U11098 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  NAND2_X1 U11099 ( .A1(n8645), .A2(SI_17_), .ZN(n8646) );
  XNOR2_X1 U11100 ( .A(n8683), .B(SI_18_), .ZN(n8664) );
  MUX2_X1 U11101 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10476), .Z(n8685) );
  XNOR2_X1 U11102 ( .A(n8664), .B(n8685), .ZN(n11419) );
  NAND2_X1 U11103 ( .A1(n11419), .A2(n9767), .ZN(n8652) );
  NAND2_X1 U11104 ( .A1(n8649), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8650) );
  XNOR2_X1 U11105 ( .A(n8650), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U11106 ( .A1(n8770), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8669), 
        .B2(n13596), .ZN(n8651) );
  XNOR2_X1 U11107 ( .A(n13857), .B(n8834), .ZN(n8659) );
  INV_X1 U11108 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8653) );
  AND2_X1 U11109 ( .A1(n8654), .A2(n8653), .ZN(n8655) );
  OR2_X1 U11110 ( .A1(n8655), .A2(n8672), .ZN(n13786) );
  AOI22_X1 U11111 ( .A1(n9746), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n6910), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U11112 ( .A1(n6545), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8656) );
  OAI211_X1 U11113 ( .C1(n13786), .C2(n8547), .A(n8657), .B(n8656), .ZN(n13533) );
  NAND2_X1 U11114 ( .A1(n13533), .A2(n11852), .ZN(n8660) );
  XNOR2_X1 U11115 ( .A(n8659), .B(n8660), .ZN(n13496) );
  INV_X1 U11116 ( .A(n8659), .ZN(n8662) );
  INV_X1 U11117 ( .A(n8660), .ZN(n8661) );
  NAND2_X1 U11118 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  NAND2_X1 U11119 ( .A1(n8683), .A2(SI_18_), .ZN(n8665) );
  MUX2_X1 U11120 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10476), .Z(n8666) );
  INV_X1 U11121 ( .A(n8666), .ZN(n8667) );
  NAND2_X1 U11122 ( .A1(n8667), .A2(n10861), .ZN(n8686) );
  NAND2_X1 U11123 ( .A1(n8688), .A2(n8686), .ZN(n8668) );
  NAND2_X1 U11124 ( .A1(n9256), .A2(n9767), .ZN(n8671) );
  AOI22_X1 U11125 ( .A1(n8770), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8669), 
        .B2(n13700), .ZN(n8670) );
  XNOR2_X1 U11126 ( .A(n13853), .B(n8834), .ZN(n8678) );
  NOR2_X1 U11127 ( .A1(n8672), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8673) );
  OR2_X1 U11128 ( .A1(n8694), .A2(n8673), .ZN(n13775) );
  INV_X1 U11129 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13776) );
  NAND2_X1 U11130 ( .A1(n8369), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11131 ( .A1(n6545), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8674) );
  OAI211_X1 U11132 ( .C1(n8720), .C2(n13776), .A(n8675), .B(n8674), .ZN(n8676)
         );
  INV_X1 U11133 ( .A(n8676), .ZN(n8677) );
  OAI21_X1 U11134 ( .B1(n13775), .B2(n8547), .A(n8677), .ZN(n13532) );
  NAND2_X1 U11135 ( .A1(n13532), .A2(n11852), .ZN(n8679) );
  NAND2_X1 U11136 ( .A1(n8678), .A2(n8679), .ZN(n13440) );
  INV_X1 U11137 ( .A(n8678), .ZN(n8681) );
  INV_X1 U11138 ( .A(n8679), .ZN(n8680) );
  NAND2_X1 U11139 ( .A1(n8681), .A2(n8680), .ZN(n13439) );
  INV_X1 U11140 ( .A(n8685), .ZN(n8684) );
  NOR2_X1 U11141 ( .A1(n8685), .A2(SI_18_), .ZN(n8689) );
  INV_X1 U11142 ( .A(n8686), .ZN(n8687) );
  MUX2_X1 U11143 ( .A(n11763), .B(n11767), .S(n10476), .Z(n8707) );
  XNOR2_X1 U11144 ( .A(n8709), .B(n8707), .ZN(n11762) );
  NAND2_X1 U11145 ( .A1(n11762), .A2(n9767), .ZN(n8693) );
  NAND2_X1 U11146 ( .A1(n8770), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8692) );
  XNOR2_X1 U11147 ( .A(n13757), .B(n8834), .ZN(n8701) );
  NOR2_X1 U11148 ( .A1(n8694), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8695) );
  OR2_X1 U11149 ( .A1(n8715), .A2(n8695), .ZN(n13758) );
  INV_X1 U11150 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n13901) );
  NAND2_X1 U11151 ( .A1(n9745), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U11152 ( .A1(n6545), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8696) );
  OAI211_X1 U11153 ( .C1(n8698), .C2(n13901), .A(n8697), .B(n8696), .ZN(n8699)
         );
  INV_X1 U11154 ( .A(n8699), .ZN(n8700) );
  OAI21_X1 U11155 ( .B1(n13758), .B2(n8547), .A(n8700), .ZN(n13531) );
  NAND2_X1 U11156 ( .A1(n13531), .A2(n11852), .ZN(n8702) );
  NAND2_X1 U11157 ( .A1(n8701), .A2(n8702), .ZN(n8706) );
  INV_X1 U11158 ( .A(n8701), .ZN(n8704) );
  INV_X1 U11159 ( .A(n8702), .ZN(n8703) );
  NAND2_X1 U11160 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  NAND2_X1 U11161 ( .A1(n8706), .A2(n8705), .ZN(n13478) );
  INV_X1 U11162 ( .A(n8707), .ZN(n8708) );
  MUX2_X1 U11163 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10476), .Z(n8730) );
  XNOR2_X1 U11164 ( .A(n8730), .B(SI_21_), .ZN(n8727) );
  XNOR2_X1 U11165 ( .A(n8729), .B(n8727), .ZN(n11819) );
  NAND2_X1 U11166 ( .A1(n11819), .A2(n9767), .ZN(n8714) );
  NAND2_X1 U11167 ( .A1(n8770), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8713) );
  XNOR2_X1 U11168 ( .A(n13744), .B(n8834), .ZN(n8725) );
  OR2_X1 U11169 ( .A1(n8715), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U11170 ( .A1(n8715), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8735) );
  AND2_X1 U11171 ( .A1(n8716), .A2(n8735), .ZN(n13743) );
  NAND2_X1 U11172 ( .A1(n13743), .A2(n8587), .ZN(n8723) );
  INV_X1 U11173 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11174 ( .A1(n8369), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11175 ( .A1(n6545), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8717) );
  OAI211_X1 U11176 ( .C1(n8720), .C2(n8719), .A(n8718), .B(n8717), .ZN(n8721)
         );
  INV_X1 U11177 ( .A(n8721), .ZN(n8722) );
  NAND2_X1 U11178 ( .A1(n8723), .A2(n8722), .ZN(n13530) );
  NAND2_X1 U11179 ( .A1(n13530), .A2(n11852), .ZN(n8724) );
  XNOR2_X1 U11180 ( .A(n8725), .B(n8724), .ZN(n13449) );
  INV_X1 U11181 ( .A(n8727), .ZN(n8728) );
  NAND2_X1 U11182 ( .A1(n8730), .A2(SI_21_), .ZN(n8731) );
  MUX2_X1 U11183 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10476), .Z(n8747) );
  XNOR2_X1 U11184 ( .A(n9324), .B(n8747), .ZN(n11985) );
  NAND2_X1 U11185 ( .A1(n11985), .A2(n9767), .ZN(n8734) );
  NAND2_X1 U11186 ( .A1(n8333), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8733) );
  XNOR2_X1 U11187 ( .A(n13836), .B(n8834), .ZN(n8742) );
  XNOR2_X1 U11188 ( .A(n8744), .B(n8742), .ZN(n13486) );
  NAND2_X1 U11189 ( .A1(n9745), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U11190 ( .A1(n9746), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8740) );
  INV_X1 U11191 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13490) );
  NAND2_X1 U11192 ( .A1(n13490), .A2(n8735), .ZN(n8737) );
  INV_X1 U11193 ( .A(n8735), .ZN(n8736) );
  NAND2_X1 U11194 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(n8736), .ZN(n8754) );
  AND2_X1 U11195 ( .A1(n8737), .A2(n8754), .ZN(n13726) );
  NAND2_X1 U11196 ( .A1(n8587), .A2(n13726), .ZN(n8739) );
  NAND2_X1 U11197 ( .A1(n6545), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8738) );
  NAND4_X1 U11198 ( .A1(n8741), .A2(n8740), .A3(n8739), .A4(n8738), .ZN(n13529) );
  AND2_X1 U11199 ( .A1(n13529), .A2(n11852), .ZN(n13485) );
  NAND2_X1 U11200 ( .A1(n13486), .A2(n13485), .ZN(n8746) );
  INV_X1 U11201 ( .A(n8742), .ZN(n8743) );
  NAND2_X1 U11202 ( .A1(n8744), .A2(n8743), .ZN(n8745) );
  NAND2_X1 U11203 ( .A1(n8769), .A2(n8765), .ZN(n8750) );
  MUX2_X1 U11204 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10476), .Z(n8766) );
  XNOR2_X1 U11205 ( .A(n8766), .B(SI_23_), .ZN(n8749) );
  NAND2_X1 U11206 ( .A1(n12070), .A2(n9767), .ZN(n8752) );
  NAND2_X1 U11207 ( .A1(n8770), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8751) );
  XNOR2_X1 U11208 ( .A(n13713), .B(n8834), .ZN(n8760) );
  NAND2_X1 U11209 ( .A1(n8369), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U11210 ( .A1(n9745), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8758) );
  INV_X1 U11211 ( .A(n8754), .ZN(n8753) );
  NAND2_X1 U11212 ( .A1(n8753), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8775) );
  INV_X1 U11213 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13435) );
  NAND2_X1 U11214 ( .A1(n8754), .A2(n13435), .ZN(n8755) );
  AND2_X1 U11215 ( .A1(n8775), .A2(n8755), .ZN(n13714) );
  NAND2_X1 U11216 ( .A1(n8587), .A2(n13714), .ZN(n8757) );
  NAND2_X1 U11217 ( .A1(n6545), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8756) );
  NAND4_X1 U11218 ( .A1(n8759), .A2(n8758), .A3(n8757), .A4(n8756), .ZN(n13528) );
  AND2_X1 U11219 ( .A1(n13528), .A2(n11852), .ZN(n13431) );
  INV_X1 U11220 ( .A(n8760), .ZN(n8761) );
  NAND2_X1 U11221 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  NAND2_X1 U11222 ( .A1(n8766), .A2(SI_23_), .ZN(n8764) );
  INV_X1 U11223 ( .A(n8766), .ZN(n8767) );
  AOI21_X2 U11224 ( .B1(n8769), .B2(n8768), .A(n7622), .ZN(n8787) );
  MUX2_X1 U11225 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10476), .Z(n8788) );
  XNOR2_X1 U11226 ( .A(n8788), .B(SI_24_), .ZN(n8785) );
  XNOR2_X1 U11227 ( .A(n8787), .B(n8785), .ZN(n12104) );
  NAND2_X1 U11228 ( .A1(n12104), .A2(n9767), .ZN(n8772) );
  NAND2_X1 U11229 ( .A1(n8770), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8771) );
  XNOR2_X1 U11230 ( .A(n13891), .B(n8341), .ZN(n8781) );
  NAND2_X1 U11231 ( .A1(n9745), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U11232 ( .A1(n6545), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8779) );
  INV_X1 U11233 ( .A(n8775), .ZN(n8773) );
  NAND2_X1 U11234 ( .A1(n8773), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8795) );
  INV_X1 U11235 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U11236 ( .A1(n8775), .A2(n8774), .ZN(n8776) );
  AND2_X1 U11237 ( .A1(n8795), .A2(n8776), .ZN(n13466) );
  NAND2_X1 U11238 ( .A1(n8587), .A2(n13466), .ZN(n8778) );
  NAND2_X1 U11239 ( .A1(n9746), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8777) );
  NOR2_X1 U11240 ( .A1(n9732), .A2(n13742), .ZN(n8782) );
  XNOR2_X1 U11241 ( .A(n8781), .B(n8782), .ZN(n13464) );
  INV_X1 U11242 ( .A(n8781), .ZN(n8783) );
  NAND2_X1 U11243 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  INV_X1 U11244 ( .A(n8785), .ZN(n8786) );
  NAND2_X1 U11245 ( .A1(n8788), .A2(SI_24_), .ZN(n8789) );
  MUX2_X1 U11246 ( .A(n6736), .B(n12178), .S(n10476), .Z(n8790) );
  NAND2_X1 U11247 ( .A1(n8790), .A2(n13160), .ZN(n8808) );
  INV_X1 U11248 ( .A(n8790), .ZN(n8791) );
  NAND2_X1 U11249 ( .A1(n8791), .A2(SI_25_), .ZN(n8792) );
  NAND2_X1 U11250 ( .A1(n8808), .A2(n8792), .ZN(n8806) );
  NAND2_X1 U11251 ( .A1(n12175), .A2(n9767), .ZN(n8794) );
  NAND2_X1 U11252 ( .A1(n8333), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8793) );
  XNOR2_X1 U11253 ( .A(n13682), .B(n8341), .ZN(n8803) );
  NAND2_X1 U11254 ( .A1(n9745), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U11255 ( .A1(n6545), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8799) );
  INV_X1 U11256 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13459) );
  INV_X1 U11257 ( .A(n8812), .ZN(n8814) );
  NAND2_X1 U11258 ( .A1(n8795), .A2(n13459), .ZN(n8796) );
  NAND2_X1 U11259 ( .A1(n8587), .A2(n13685), .ZN(n8798) );
  NAND2_X1 U11260 ( .A1(n9746), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8797) );
  NAND4_X1 U11261 ( .A1(n8800), .A2(n8799), .A3(n8798), .A4(n8797), .ZN(n13526) );
  NAND2_X1 U11262 ( .A1(n13526), .A2(n11852), .ZN(n8801) );
  XNOR2_X1 U11263 ( .A(n8803), .B(n8801), .ZN(n13458) );
  NAND2_X1 U11264 ( .A1(n13457), .A2(n13458), .ZN(n8805) );
  INV_X1 U11265 ( .A(n8801), .ZN(n8802) );
  NAND2_X1 U11266 ( .A1(n8803), .A2(n8802), .ZN(n8804) );
  MUX2_X1 U11267 ( .A(n12256), .B(n12259), .S(n10476), .Z(n8826) );
  XNOR2_X1 U11268 ( .A(n8826), .B(SI_26_), .ZN(n8809) );
  NAND2_X1 U11269 ( .A1(n12255), .A2(n9767), .ZN(n8811) );
  NAND2_X1 U11270 ( .A1(n8333), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8810) );
  XNOR2_X1 U11271 ( .A(n13668), .B(n8341), .ZN(n8820) );
  NAND2_X1 U11272 ( .A1(n9745), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U11273 ( .A1(n9746), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U11274 ( .A1(n8812), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8835) );
  INV_X1 U11275 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U11276 ( .A1(n8814), .A2(n8813), .ZN(n8815) );
  AND2_X1 U11277 ( .A1(n8835), .A2(n8815), .ZN(n13666) );
  NAND2_X1 U11278 ( .A1(n8587), .A2(n13666), .ZN(n8817) );
  NAND2_X1 U11279 ( .A1(n6545), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8816) );
  OR2_X1 U11280 ( .A1(n13742), .A2(n9936), .ZN(n8821) );
  NAND2_X1 U11281 ( .A1(n8820), .A2(n8821), .ZN(n8825) );
  INV_X1 U11282 ( .A(n8820), .ZN(n8823) );
  INV_X1 U11283 ( .A(n8821), .ZN(n8822) );
  NAND2_X1 U11284 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  NAND2_X1 U11285 ( .A1(n8825), .A2(n8824), .ZN(n13507) );
  NAND2_X1 U11286 ( .A1(n8827), .A2(n12076), .ZN(n8828) );
  MUX2_X1 U11287 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10476), .Z(n8884) );
  INV_X1 U11288 ( .A(n8884), .ZN(n8830) );
  XNOR2_X1 U11289 ( .A(n8830), .B(SI_27_), .ZN(n8831) );
  NAND2_X1 U11290 ( .A1(n13925), .A2(n9767), .ZN(n8833) );
  NAND2_X1 U11291 ( .A1(n8333), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8832) );
  NAND2_X2 U11292 ( .A1(n8833), .A2(n8832), .ZN(n13809) );
  XNOR2_X1 U11293 ( .A(n13809), .B(n8834), .ZN(n8842) );
  NAND2_X1 U11294 ( .A1(n9746), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8840) );
  NAND2_X1 U11295 ( .A1(n9745), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8839) );
  INV_X1 U11296 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13426) );
  NAND2_X1 U11297 ( .A1(n8835), .A2(n13426), .ZN(n8836) );
  NAND2_X1 U11298 ( .A1(n8587), .A2(n13652), .ZN(n8838) );
  NAND2_X1 U11299 ( .A1(n6545), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8837) );
  NAND4_X1 U11300 ( .A1(n8840), .A2(n8839), .A3(n8838), .A4(n8837), .ZN(n13524) );
  NAND2_X1 U11301 ( .A1(n13524), .A2(n11852), .ZN(n8841) );
  XNOR2_X1 U11302 ( .A(n8842), .B(n8841), .ZN(n13424) );
  NAND2_X1 U11303 ( .A1(n9746), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11304 ( .A1(n9745), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8850) );
  INV_X1 U11305 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8843) );
  NOR2_X1 U11306 ( .A1(n8844), .A2(n8843), .ZN(n13624) );
  INV_X1 U11307 ( .A(n13624), .ZN(n8846) );
  NAND2_X1 U11308 ( .A1(n8844), .A2(n8843), .ZN(n8845) );
  NAND2_X1 U11309 ( .A1(n8846), .A2(n8845), .ZN(n13640) );
  INV_X1 U11310 ( .A(n13640), .ZN(n8847) );
  NAND2_X1 U11311 ( .A1(n8587), .A2(n8847), .ZN(n8849) );
  NAND2_X1 U11312 ( .A1(n6545), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8848) );
  NAND4_X1 U11313 ( .A1(n8851), .A2(n8850), .A3(n8849), .A4(n8848), .ZN(n13523) );
  AND2_X1 U11314 ( .A1(n13523), .A2(n11852), .ZN(n8852) );
  XNOR2_X1 U11315 ( .A(n8341), .B(n8852), .ZN(n8853) );
  INV_X1 U11316 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11317 ( .A1(n8863), .A2(n8862), .ZN(n8865) );
  NAND2_X1 U11318 ( .A1(n8865), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U11319 ( .A1(n8631), .A2(n8857), .ZN(n8859) );
  OAI21_X1 U11320 ( .B1(n8859), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8858) );
  XNOR2_X1 U11321 ( .A(n8858), .B(P2_IR_REG_26__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U11322 ( .A1(n8859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8860) );
  XNOR2_X1 U11323 ( .A(n8860), .B(P2_IR_REG_25__SCAN_IN), .ZN(n12176) );
  AND2_X1 U11324 ( .A1(n12258), .A2(n12176), .ZN(n8861) );
  NAND2_X1 U11325 ( .A1(n12105), .A2(n8861), .ZN(n10530) );
  OR2_X1 U11326 ( .A1(n8863), .A2(n8862), .ZN(n8864) );
  NAND2_X1 U11327 ( .A1(n8865), .A2(n8864), .ZN(n10531) );
  OR2_X1 U11328 ( .A1(n12105), .A2(n12258), .ZN(n8869) );
  XNOR2_X1 U11329 ( .A(P2_B_REG_SCAN_IN), .B(n12105), .ZN(n8866) );
  INV_X1 U11330 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15181) );
  NAND2_X1 U11331 ( .A1(n15175), .A2(n15181), .ZN(n8868) );
  INV_X1 U11332 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15185) );
  NAND2_X1 U11333 ( .A1(n15175), .A2(n15185), .ZN(n8871) );
  OR2_X1 U11334 ( .A1(n12258), .A2(n12176), .ZN(n8870) );
  AND2_X1 U11335 ( .A1(n8871), .A2(n8870), .ZN(n15183) );
  NOR4_X1 U11336 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8875) );
  NOR4_X1 U11337 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n8874) );
  NOR4_X1 U11338 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8873) );
  NOR4_X1 U11339 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8872) );
  NAND4_X1 U11340 ( .A1(n8875), .A2(n8874), .A3(n8873), .A4(n8872), .ZN(n8881)
         );
  NOR2_X1 U11341 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .ZN(
        n8879) );
  NOR4_X1 U11342 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8878) );
  NOR4_X1 U11343 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n8877) );
  NOR4_X1 U11344 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8876) );
  NAND4_X1 U11345 ( .A1(n8879), .A2(n8878), .A3(n8877), .A4(n8876), .ZN(n8880)
         );
  OAI21_X1 U11346 ( .B1(n8881), .B2(n8880), .A(n15175), .ZN(n9953) );
  NAND2_X1 U11347 ( .A1(n15183), .A2(n9953), .ZN(n11248) );
  NOR2_X1 U11348 ( .A1(n15182), .A2(n11248), .ZN(n8900) );
  NAND2_X1 U11349 ( .A1(n15187), .A2(n8900), .ZN(n8891) );
  NAND2_X1 U11350 ( .A1(n11766), .A2(n13607), .ZN(n9773) );
  OR3_X2 U11351 ( .A1(n8891), .A2(n10532), .A3(n15200), .ZN(n13520) );
  INV_X1 U11352 ( .A(n11766), .ZN(n9832) );
  NAND2_X1 U11353 ( .A1(n10766), .A2(n9832), .ZN(n11253) );
  NOR2_X1 U11354 ( .A1(n8891), .A2(n11253), .ZN(n8882) );
  AND2_X2 U11355 ( .A1(n15187), .A2(n9950), .ZN(n15163) );
  NOR2_X1 U11356 ( .A1(n8884), .A2(SI_27_), .ZN(n8886) );
  NAND2_X1 U11357 ( .A1(n8884), .A2(SI_27_), .ZN(n8885) );
  MUX2_X1 U11358 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10476), .Z(n9422) );
  XNOR2_X1 U11359 ( .A(n9422), .B(SI_28_), .ZN(n9425) );
  NAND2_X1 U11360 ( .A1(n12290), .A2(n9767), .ZN(n8889) );
  NAND2_X1 U11361 ( .A1(n8333), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8888) );
  NAND2_X2 U11362 ( .A1(n8889), .A2(n8888), .ZN(n13643) );
  INV_X1 U11363 ( .A(n8891), .ZN(n8892) );
  INV_X1 U11364 ( .A(n9773), .ZN(n9809) );
  AND2_X2 U11365 ( .A1(n10532), .A2(n10540), .ZN(n13510) );
  NAND2_X1 U11366 ( .A1(n9746), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U11367 ( .A1(n9745), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U11368 ( .A1(n8587), .A2(n13624), .ZN(n8894) );
  NAND2_X1 U11369 ( .A1(n6545), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8893) );
  NAND4_X1 U11370 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8893), .ZN(n13522) );
  NAND2_X1 U11371 ( .A1(n13510), .A2(n13522), .ZN(n8899) );
  INV_X1 U11372 ( .A(n10540), .ZN(n8897) );
  NAND2_X1 U11373 ( .A1(n13509), .A2(n13524), .ZN(n8898) );
  NAND2_X1 U11374 ( .A1(n8899), .A2(n8898), .ZN(n13636) );
  AOI22_X1 U11375 ( .A1(n13513), .A2(n13636), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n8906) );
  INV_X1 U11376 ( .A(n8900), .ZN(n8902) );
  INV_X1 U11377 ( .A(n9950), .ZN(n8901) );
  AND2_X1 U11378 ( .A1(n10532), .A2(n9773), .ZN(n9948) );
  AOI21_X1 U11379 ( .B1(n8902), .B2(n8901), .A(n9948), .ZN(n10796) );
  NAND2_X1 U11380 ( .A1(n10796), .A2(n8903), .ZN(n8904) );
  OR2_X1 U11381 ( .A1(n13640), .A2(n13515), .ZN(n8905) );
  AND2_X1 U11382 ( .A1(n8906), .A2(n8905), .ZN(n8907) );
  NAND2_X1 U11383 ( .A1(n8910), .A2(n9142), .ZN(n8911) );
  NOR2_X1 U11384 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8917) );
  NOR2_X1 U11385 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n8916) );
  NOR2_X1 U11386 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n8915) );
  INV_X1 U11387 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14531) );
  NAND2_X1 U11388 ( .A1(n8920), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8922) );
  XNOR2_X2 U11389 ( .A(n8922), .B(n8921), .ZN(n12334) );
  NAND2_X1 U11390 ( .A1(n8923), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8929) );
  INV_X1 U11391 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10192) );
  INV_X1 U11392 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n11377) );
  OR2_X1 U11393 ( .A1(n9015), .A2(n11377), .ZN(n8927) );
  INV_X1 U11394 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11376) );
  INV_X1 U11395 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14858) );
  NOR2_X1 U11396 ( .A1(n10476), .A2(n10450), .ZN(n8930) );
  XNOR2_X1 U11397 ( .A(n8930), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14548) );
  INV_X1 U11398 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8935) );
  MUX2_X1 U11399 ( .A(n14858), .B(n14548), .S(n8983), .Z(n11720) );
  NAND2_X1 U11400 ( .A1(n8938), .A2(n11380), .ZN(n8987) );
  INV_X1 U11401 ( .A(n8987), .ZN(n8952) );
  INV_X1 U11402 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11730) );
  OR2_X1 U11403 ( .A1(n9032), .A2(n11730), .ZN(n8943) );
  INV_X1 U11404 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8939) );
  INV_X1 U11405 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n8940) );
  INV_X1 U11406 ( .A(n8946), .ZN(n10477) );
  NAND2_X1 U11407 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8947) );
  MUX2_X1 U11408 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8947), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8950) );
  INV_X1 U11409 ( .A(n8948), .ZN(n8949) );
  OR2_X1 U11410 ( .A1(n8983), .A2(n10608), .ZN(n8951) );
  NAND2_X1 U11411 ( .A1(n8952), .A2(n9479), .ZN(n10029) );
  NAND2_X1 U11412 ( .A1(n9014), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8957) );
  INV_X1 U11413 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11331) );
  INV_X1 U11414 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8953) );
  OR2_X1 U11415 ( .A1(n9017), .A2(n8953), .ZN(n8955) );
  INV_X1 U11416 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11328) );
  OR2_X1 U11417 ( .A1(n9015), .A2(n11328), .ZN(n8954) );
  NAND4_X2 U11418 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n14136) );
  INV_X1 U11419 ( .A(n10457), .ZN(n8958) );
  OR2_X1 U11420 ( .A1(n9436), .A2(n10478), .ZN(n8961) );
  NAND2_X1 U11421 ( .A1(n8948), .A2(n6936), .ZN(n8979) );
  NAND2_X1 U11422 ( .A1(n8959), .A2(n8979), .ZN(n14157) );
  OR2_X1 U11423 ( .A1(n8983), .A2(n14157), .ZN(n8960) );
  AND3_X2 U11424 ( .A1(n8962), .A2(n8961), .A3(n8960), .ZN(n14973) );
  NAND2_X1 U11425 ( .A1(n14136), .A2(n14973), .ZN(n8994) );
  INV_X1 U11426 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8964) );
  NAND2_X1 U11427 ( .A1(n8965), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8966) );
  INV_X1 U11428 ( .A(n14547), .ZN(n10024) );
  NAND2_X1 U11429 ( .A1(n10024), .A2(n14415), .ZN(n10682) );
  NAND2_X1 U11430 ( .A1(n10026), .A2(n10682), .ZN(n8971) );
  NAND2_X1 U11431 ( .A1(n8969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U11432 ( .A1(n8971), .A2(n10681), .ZN(n8972) );
  INV_X1 U11433 ( .A(n8992), .ZN(n9447) );
  NAND2_X1 U11434 ( .A1(n8994), .A2(n9447), .ZN(n8997) );
  NAND2_X1 U11435 ( .A1(n9014), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8977) );
  OR2_X1 U11436 ( .A1(n9032), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8976) );
  INV_X1 U11437 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8973) );
  OR2_X1 U11438 ( .A1(n9017), .A2(n8973), .ZN(n8975) );
  OR2_X1 U11439 ( .A1(n9015), .A2(n13071), .ZN(n8974) );
  NAND2_X1 U11440 ( .A1(n8979), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8978) );
  MUX2_X1 U11441 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8978), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8980) );
  NAND2_X1 U11442 ( .A1(n8980), .A2(n9008), .ZN(n10611) );
  OR2_X1 U11443 ( .A1(n10484), .A2(n9118), .ZN(n8982) );
  OR2_X1 U11444 ( .A1(n9436), .A2(n10483), .ZN(n8981) );
  OAI211_X1 U11445 ( .C1(n8983), .C2(n10611), .A(n8982), .B(n8981), .ZN(n14980) );
  OAI21_X1 U11446 ( .B1(n10029), .B2(n8997), .A(n11369), .ZN(n8984) );
  INV_X1 U11447 ( .A(n8984), .ZN(n9002) );
  AND4_X1 U11448 ( .A1(n10028), .A2(n10030), .A3(n8987), .A4(n8992), .ZN(n8990) );
  NAND2_X1 U11449 ( .A1(n14138), .A2(n11380), .ZN(n11728) );
  OR2_X1 U11450 ( .A1(n14138), .A2(n11380), .ZN(n8988) );
  NAND2_X1 U11451 ( .A1(n11728), .A2(n8988), .ZN(n11383) );
  INV_X1 U11452 ( .A(n10180), .ZN(n10181) );
  NAND2_X1 U11453 ( .A1(n11383), .A2(n10181), .ZN(n8989) );
  NAND2_X1 U11454 ( .A1(n8990), .A2(n8989), .ZN(n9001) );
  INV_X1 U11455 ( .A(n9479), .ZN(n8991) );
  NAND3_X1 U11456 ( .A1(n11324), .A2(n8991), .A3(n8992), .ZN(n9000) );
  INV_X1 U11457 ( .A(n10030), .ZN(n8993) );
  NAND2_X1 U11458 ( .A1(n8993), .A2(n9413), .ZN(n8996) );
  OR2_X1 U11459 ( .A1(n8994), .A2(n9413), .ZN(n8995) );
  OAI211_X1 U11460 ( .C1(n8997), .C2(n10028), .A(n8996), .B(n8995), .ZN(n8998)
         );
  INV_X1 U11461 ( .A(n8998), .ZN(n8999) );
  NAND4_X1 U11462 ( .A1(n9002), .A2(n9001), .A3(n9000), .A4(n8999), .ZN(n9006)
         );
  NAND2_X1 U11463 ( .A1(n8992), .A2(n14980), .ZN(n9004) );
  INV_X1 U11464 ( .A(n14980), .ZN(n10066) );
  NAND2_X1 U11465 ( .A1(n10066), .A2(n9447), .ZN(n9003) );
  MUX2_X1 U11466 ( .A(n9004), .B(n9003), .S(n14135), .Z(n9005) );
  NAND2_X1 U11467 ( .A1(n9006), .A2(n9005), .ZN(n9026) );
  NAND2_X1 U11468 ( .A1(n10472), .A2(n9466), .ZN(n9013) );
  NAND2_X1 U11469 ( .A1(n9008), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9007) );
  MUX2_X1 U11470 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9007), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9011) );
  INV_X1 U11471 ( .A(n9008), .ZN(n9010) );
  INV_X1 U11472 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U11473 ( .A1(n9010), .A2(n9009), .ZN(n9029) );
  NAND2_X1 U11474 ( .A1(n9011), .A2(n9029), .ZN(n14182) );
  INV_X1 U11475 ( .A(n14182), .ZN(n10613) );
  AOI22_X1 U11476 ( .A1(n9465), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9266), .B2(
        n10613), .ZN(n9012) );
  NAND2_X1 U11477 ( .A1(n9013), .A2(n9012), .ZN(n10206) );
  NAND2_X1 U11478 ( .A1(n9014), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9022) );
  INV_X1 U11479 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9016) );
  OR2_X1 U11480 ( .A1(n9015), .A2(n9016), .ZN(n9021) );
  NAND2_X1 U11481 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9033) );
  OAI21_X1 U11482 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9033), .ZN(n14939) );
  OR2_X1 U11483 ( .A1(n9032), .A2(n14939), .ZN(n9020) );
  INV_X1 U11484 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9018) );
  OR2_X1 U11485 ( .A1(n9442), .A2(n9018), .ZN(n9019) );
  NAND4_X1 U11486 ( .A1(n9022), .A2(n9021), .A3(n9020), .A4(n9019), .ZN(n14134) );
  MUX2_X1 U11487 ( .A(n10206), .B(n14134), .S(n8992), .Z(n9023) );
  INV_X1 U11488 ( .A(n9023), .ZN(n9025) );
  MUX2_X1 U11489 ( .A(n10206), .B(n14134), .S(n9413), .Z(n9024) );
  OAI21_X1 U11490 ( .B1(n9026), .B2(n9025), .A(n9024), .ZN(n9028) );
  NAND2_X1 U11491 ( .A1(n9026), .A2(n9025), .ZN(n9027) );
  NAND2_X1 U11492 ( .A1(n9028), .A2(n9027), .ZN(n9041) );
  NAND2_X1 U11493 ( .A1(n9029), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9030) );
  XNOR2_X1 U11494 ( .A(n9030), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U11495 ( .A1(n9465), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9266), .B2(
        n10653), .ZN(n9031) );
  NAND2_X1 U11496 ( .A1(n9439), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9039) );
  INV_X1 U11497 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10614) );
  OR2_X1 U11498 ( .A1(n9417), .A2(n10614), .ZN(n9038) );
  AND2_X1 U11499 ( .A1(n9033), .A2(n11284), .ZN(n9034) );
  NOR2_X1 U11500 ( .A1(n9033), .A2(n11284), .ZN(n9048) );
  OR2_X1 U11501 ( .A1(n9034), .A2(n9048), .ZN(n11391) );
  OR2_X1 U11502 ( .A1(n9032), .A2(n11391), .ZN(n9037) );
  INV_X1 U11503 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9035) );
  OR2_X1 U11504 ( .A1(n9442), .A2(n9035), .ZN(n9036) );
  NAND4_X1 U11505 ( .A1(n9039), .A2(n9038), .A3(n9037), .A4(n9036), .ZN(n14132) );
  MUX2_X1 U11506 ( .A(n11287), .B(n14132), .S(n9413), .Z(n9042) );
  MUX2_X1 U11507 ( .A(n11287), .B(n14132), .S(n9468), .Z(n9040) );
  OR2_X1 U11508 ( .A1(n9043), .A2(n9118), .ZN(n9046) );
  OR2_X1 U11509 ( .A1(n9072), .A2(n8935), .ZN(n9044) );
  XNOR2_X1 U11510 ( .A(n9044), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U11511 ( .A1(n9465), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9266), .B2(
        n10625), .ZN(n9045) );
  NAND2_X1 U11512 ( .A1(n9014), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9054) );
  INV_X1 U11513 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9047) );
  OR2_X1 U11514 ( .A1(n9015), .A2(n9047), .ZN(n9053) );
  NAND2_X1 U11515 ( .A1(n9048), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9064) );
  OR2_X1 U11516 ( .A1(n9048), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U11517 ( .A1(n9064), .A2(n9049), .ZN(n14922) );
  OR2_X1 U11518 ( .A1(n9032), .A2(n14922), .ZN(n9052) );
  INV_X1 U11519 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9050) );
  OR2_X1 U11520 ( .A1(n9442), .A2(n9050), .ZN(n9051) );
  NAND4_X1 U11521 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n9051), .ZN(n14131) );
  MUX2_X1 U11522 ( .A(n11658), .B(n14131), .S(n9468), .Z(n9058) );
  NAND2_X1 U11523 ( .A1(n9056), .A2(n9055), .ZN(n9062) );
  INV_X1 U11524 ( .A(n9057), .ZN(n9060) );
  INV_X1 U11525 ( .A(n9058), .ZN(n9059) );
  NAND2_X1 U11526 ( .A1(n9060), .A2(n9059), .ZN(n9061) );
  NAND2_X1 U11527 ( .A1(n9062), .A2(n9061), .ZN(n9077) );
  NAND2_X1 U11528 ( .A1(n9439), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9070) );
  INV_X1 U11529 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9063) );
  OR2_X1 U11530 ( .A1(n9443), .A2(n9063), .ZN(n9069) );
  NAND2_X1 U11531 ( .A1(n9064), .A2(n13134), .ZN(n9065) );
  NAND2_X1 U11532 ( .A1(n9080), .A2(n9065), .ZN(n11668) );
  OR2_X1 U11533 ( .A1(n9032), .A2(n11668), .ZN(n9068) );
  INV_X1 U11534 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9066) );
  OR2_X1 U11535 ( .A1(n9442), .A2(n9066), .ZN(n9067) );
  NAND4_X1 U11536 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n14130) );
  NAND2_X1 U11537 ( .A1(n10495), .A2(n9466), .ZN(n9075) );
  INV_X1 U11538 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U11539 ( .A1(n9072), .A2(n9071), .ZN(n9087) );
  NAND2_X1 U11540 ( .A1(n9087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9073) );
  XNOR2_X1 U11541 ( .A(n9073), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U11542 ( .A1(n9465), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9266), .B2(
        n10641), .ZN(n9074) );
  MUX2_X1 U11543 ( .A(n14130), .B(n15006), .S(n9468), .Z(n9078) );
  MUX2_X1 U11544 ( .A(n14130), .B(n15006), .S(n9413), .Z(n9076) );
  NAND2_X1 U11545 ( .A1(n9439), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9086) );
  INV_X1 U11546 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10636) );
  OR2_X1 U11547 ( .A1(n9417), .A2(n10636), .ZN(n9085) );
  NAND2_X1 U11548 ( .A1(n9080), .A2(n9079), .ZN(n9081) );
  NAND2_X1 U11549 ( .A1(n9099), .A2(n9081), .ZN(n11876) );
  OR2_X1 U11550 ( .A1(n9032), .A2(n11876), .ZN(n9084) );
  INV_X1 U11551 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9082) );
  OR2_X1 U11552 ( .A1(n9442), .A2(n9082), .ZN(n9083) );
  INV_X1 U11553 ( .A(n11528), .ZN(n14129) );
  OR2_X1 U11554 ( .A1(n10502), .A2(n9118), .ZN(n9090) );
  NAND2_X1 U11555 ( .A1(n9202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9088) );
  XNOR2_X1 U11556 ( .A(n9088), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U11557 ( .A1(n9465), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9266), .B2(
        n10709), .ZN(n9089) );
  MUX2_X1 U11558 ( .A(n14129), .B(n11878), .S(n9413), .Z(n9094) );
  NAND2_X1 U11559 ( .A1(n9092), .A2(n9091), .ZN(n9098) );
  INV_X1 U11560 ( .A(n9093), .ZN(n9096) );
  INV_X1 U11561 ( .A(n9094), .ZN(n9095) );
  NAND2_X1 U11562 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  NAND2_X1 U11563 ( .A1(n9098), .A2(n9097), .ZN(n9110) );
  NAND2_X1 U11564 ( .A1(n9439), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9106) );
  INV_X1 U11565 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10701) );
  OR2_X1 U11566 ( .A1(n9443), .A2(n10701), .ZN(n9105) );
  INV_X1 U11567 ( .A(n9135), .ZN(n9101) );
  NAND2_X1 U11568 ( .A1(n9099), .A2(n10705), .ZN(n9100) );
  NAND2_X1 U11569 ( .A1(n9101), .A2(n9100), .ZN(n12008) );
  OR2_X1 U11570 ( .A1(n9032), .A2(n12008), .ZN(n9104) );
  INV_X1 U11571 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9102) );
  OR2_X1 U11572 ( .A1(n9442), .A2(n9102), .ZN(n9103) );
  INV_X1 U11573 ( .A(n11769), .ZN(n14128) );
  OR2_X1 U11574 ( .A1(n10519), .A2(n9118), .ZN(n9108) );
  XNOR2_X1 U11575 ( .A(n9144), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U11576 ( .A1(n9465), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9266), .B2(
        n10813), .ZN(n9107) );
  MUX2_X1 U11577 ( .A(n14128), .B(n12010), .S(n9413), .Z(n9109) );
  INV_X1 U11578 ( .A(n9111), .ZN(n9112) );
  NAND2_X1 U11579 ( .A1(n9439), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9117) );
  INV_X1 U11580 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10811) );
  OR2_X1 U11581 ( .A1(n9417), .A2(n10811), .ZN(n9116) );
  XNOR2_X1 U11582 ( .A(n9135), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n12150) );
  OR2_X1 U11583 ( .A1(n9032), .A2(n12150), .ZN(n9115) );
  INV_X1 U11584 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9113) );
  OR2_X1 U11585 ( .A1(n9442), .A2(n9113), .ZN(n9114) );
  INV_X1 U11586 ( .A(n11737), .ZN(n14127) );
  OR2_X1 U11587 ( .A1(n10525), .A2(n9118), .ZN(n9123) );
  INV_X1 U11588 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U11589 ( .A1(n9144), .A2(n9119), .ZN(n9120) );
  NAND2_X1 U11590 ( .A1(n9120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9121) );
  XNOR2_X1 U11591 ( .A(n9121), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U11592 ( .A1(n9465), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9266), 
        .B2(n11116), .ZN(n9122) );
  MUX2_X1 U11593 ( .A(n14127), .B(n15022), .S(n9413), .Z(n9127) );
  NAND2_X1 U11594 ( .A1(n9125), .A2(n9124), .ZN(n9131) );
  INV_X1 U11595 ( .A(n9126), .ZN(n9129) );
  INV_X1 U11596 ( .A(n9127), .ZN(n9128) );
  NAND2_X1 U11597 ( .A1(n9129), .A2(n9128), .ZN(n9130) );
  NAND2_X1 U11598 ( .A1(n9131), .A2(n9130), .ZN(n9149) );
  NAND2_X1 U11599 ( .A1(n9439), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9141) );
  INV_X1 U11600 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11110) );
  OR2_X1 U11601 ( .A1(n9443), .A2(n11110), .ZN(n9140) );
  NAND2_X1 U11602 ( .A1(n9135), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9133) );
  INV_X1 U11603 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U11604 ( .A1(n9133), .A2(n9132), .ZN(n9136) );
  AND2_X1 U11605 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n9134) );
  NAND2_X1 U11606 ( .A1(n9135), .A2(n9134), .ZN(n9152) );
  NAND2_X1 U11607 ( .A1(n9136), .A2(n9152), .ZN(n12206) );
  OR2_X1 U11608 ( .A1(n9032), .A2(n12206), .ZN(n9139) );
  INV_X1 U11609 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9137) );
  OR2_X1 U11610 ( .A1(n9442), .A2(n9137), .ZN(n9138) );
  NAND4_X1 U11611 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n14126) );
  NAND2_X1 U11612 ( .A1(n10596), .A2(n9466), .ZN(n9147) );
  OR2_X1 U11613 ( .A1(n9142), .A2(n8935), .ZN(n9143) );
  NAND2_X1 U11614 ( .A1(n9144), .A2(n9143), .ZN(n9160) );
  INV_X1 U11615 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9145) );
  XNOR2_X1 U11616 ( .A(n9160), .B(n9145), .ZN(n11427) );
  AOI22_X1 U11617 ( .A1(n9465), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9266), 
        .B2(n11427), .ZN(n9146) );
  MUX2_X1 U11618 ( .A(n14126), .B(n11740), .S(n9468), .Z(n9150) );
  MUX2_X1 U11619 ( .A(n14126), .B(n11740), .S(n9413), .Z(n9148) );
  INV_X1 U11620 ( .A(n9150), .ZN(n9151) );
  NAND2_X1 U11621 ( .A1(n8923), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U11622 ( .A1(n9152), .A2(n13041), .ZN(n9153) );
  NAND2_X1 U11623 ( .A1(n9185), .A2(n9153), .ZN(n14687) );
  OR2_X1 U11624 ( .A1(n9032), .A2(n14687), .ZN(n9158) );
  INV_X1 U11625 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9154) );
  OR2_X1 U11626 ( .A1(n9015), .A2(n9154), .ZN(n9157) );
  INV_X1 U11627 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9155) );
  OR2_X1 U11628 ( .A1(n9417), .A2(n9155), .ZN(n9156) );
  NAND4_X1 U11629 ( .A1(n9159), .A2(n9158), .A3(n9157), .A4(n9156), .ZN(n14125) );
  NAND2_X1 U11630 ( .A1(n10698), .A2(n9466), .ZN(n9163) );
  NAND2_X1 U11631 ( .A1(n9161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9170) );
  XNOR2_X1 U11632 ( .A(n9170), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U11633 ( .A1(n9465), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9266), 
        .B2(n11622), .ZN(n9162) );
  MUX2_X1 U11634 ( .A(n14125), .B(n14679), .S(n9413), .Z(n9167) );
  NAND2_X1 U11635 ( .A1(n9166), .A2(n9167), .ZN(n9165) );
  MUX2_X1 U11636 ( .A(n14125), .B(n14679), .S(n9468), .Z(n9164) );
  NAND2_X1 U11637 ( .A1(n9170), .A2(n9169), .ZN(n9171) );
  NAND2_X1 U11638 ( .A1(n9171), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U11639 ( .A1(n9191), .A2(n6833), .ZN(n9172) );
  NAND2_X1 U11640 ( .A1(n9172), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9173) );
  XNOR2_X1 U11641 ( .A(n9173), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U11642 ( .A1(n9266), .A2(n12062), .B1(n9465), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U11643 ( .A1(n9439), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9183) );
  INV_X1 U11644 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11891) );
  OR2_X1 U11645 ( .A1(n9443), .A2(n11891), .ZN(n9182) );
  INV_X1 U11646 ( .A(n9185), .ZN(n9176) );
  AOI21_X1 U11647 ( .B1(n9176), .B2(P1_REG3_REG_13__SCAN_IN), .A(
        P1_REG3_REG_14__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U11648 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n9177) );
  OR2_X1 U11649 ( .A1(n9178), .A2(n9210), .ZN(n13945) );
  OR2_X1 U11650 ( .A1(n9032), .A2(n13945), .ZN(n9181) );
  INV_X1 U11651 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9179) );
  OR2_X1 U11652 ( .A1(n9442), .A2(n9179), .ZN(n9180) );
  NAND4_X1 U11653 ( .A1(n9183), .A2(n9182), .A3(n9181), .A4(n9180), .ZN(n14123) );
  NAND2_X1 U11654 ( .A1(n9439), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9190) );
  INV_X1 U11655 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11620) );
  OR2_X1 U11656 ( .A1(n9443), .A2(n11620), .ZN(n9189) );
  INV_X1 U11657 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9184) );
  XNOR2_X1 U11658 ( .A(n9185), .B(n9184), .ZN(n14046) );
  OR2_X1 U11659 ( .A1(n9032), .A2(n14046), .ZN(n9188) );
  INV_X1 U11660 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9186) );
  OR2_X1 U11661 ( .A1(n9442), .A2(n9186), .ZN(n9187) );
  NAND4_X1 U11662 ( .A1(n9190), .A2(n9189), .A3(n9188), .A4(n9187), .ZN(n14124) );
  INV_X1 U11663 ( .A(n14124), .ZN(n12081) );
  NAND2_X1 U11664 ( .A1(n10772), .A2(n9466), .ZN(n9193) );
  XNOR2_X1 U11665 ( .A(n9191), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U11666 ( .A1(n9465), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9266), 
        .B2(n11896), .ZN(n9192) );
  MUX2_X1 U11667 ( .A(n14124), .B(n14827), .S(n9468), .Z(n9220) );
  NAND2_X1 U11668 ( .A1(n14827), .A2(n9447), .ZN(n9194) );
  OAI211_X1 U11669 ( .C1(n9447), .C2(n12081), .A(n9220), .B(n9194), .ZN(n9195)
         );
  NAND2_X1 U11670 ( .A1(n9197), .A2(n9196), .ZN(n9226) );
  NAND2_X1 U11671 ( .A1(n11126), .A2(n9466), .ZN(n9209) );
  NOR2_X1 U11672 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .ZN(n9199) );
  NAND4_X1 U11673 ( .A1(n9200), .A2(n9142), .A3(n9199), .A4(n9198), .ZN(n9201)
         );
  NOR2_X1 U11674 ( .A1(n9202), .A2(n9201), .ZN(n9205) );
  NOR2_X1 U11675 ( .A1(n9205), .A2(n8935), .ZN(n9203) );
  MUX2_X1 U11676 ( .A(n8935), .B(n9203), .S(P1_IR_REG_15__SCAN_IN), .Z(n9207)
         );
  INV_X1 U11677 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U11678 ( .A1(n9205), .A2(n9204), .ZN(n9243) );
  INV_X1 U11679 ( .A(n9243), .ZN(n9206) );
  OR2_X1 U11680 ( .A1(n9207), .A2(n9206), .ZN(n12058) );
  INV_X1 U11681 ( .A(n12058), .ZN(n14208) );
  AOI22_X1 U11682 ( .A1(n9465), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9266), 
        .B2(n14208), .ZN(n9208) );
  NAND2_X1 U11683 ( .A1(n9014), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9216) );
  INV_X1 U11684 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12125) );
  OR2_X1 U11685 ( .A1(n9015), .A2(n12125), .ZN(n9215) );
  NOR2_X1 U11686 ( .A1(n9210), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9211) );
  OR2_X1 U11687 ( .A1(n9250), .A2(n9211), .ZN(n14100) );
  OR2_X1 U11688 ( .A1(n9032), .A2(n14100), .ZN(n9214) );
  INV_X1 U11689 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9212) );
  OR2_X1 U11690 ( .A1(n9442), .A2(n9212), .ZN(n9213) );
  INV_X1 U11691 ( .A(n14123), .ZN(n10287) );
  OR2_X1 U11692 ( .A1(n14820), .A2(n10287), .ZN(n10048) );
  AOI21_X1 U11693 ( .B1(n10049), .B2(n10048), .A(n9447), .ZN(n9219) );
  NAND2_X1 U11694 ( .A1(n14104), .A2(n12161), .ZN(n9474) );
  NAND2_X1 U11695 ( .A1(n14820), .A2(n10287), .ZN(n9217) );
  AOI21_X1 U11696 ( .B1(n9474), .B2(n9217), .A(n9468), .ZN(n9218) );
  NOR2_X1 U11697 ( .A1(n9219), .A2(n9218), .ZN(n9224) );
  INV_X1 U11698 ( .A(n9220), .ZN(n9222) );
  MUX2_X1 U11699 ( .A(n14124), .B(n14827), .S(n9447), .Z(n9221) );
  NAND3_X1 U11700 ( .A1(n12086), .A2(n9222), .A3(n9221), .ZN(n9223) );
  OAI21_X1 U11701 ( .B1(n7635), .B2(n9226), .A(n9225), .ZN(n9228) );
  MUX2_X1 U11702 ( .A(n9474), .B(n10049), .S(n9413), .Z(n9227) );
  NAND2_X1 U11703 ( .A1(n9228), .A2(n9227), .ZN(n9239) );
  NAND2_X1 U11704 ( .A1(n9439), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9233) );
  INV_X1 U11705 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14204) );
  OR2_X1 U11706 ( .A1(n9443), .A2(n14204), .ZN(n9232) );
  XNOR2_X1 U11707 ( .A(n9250), .B(P1_REG3_REG_16__SCAN_IN), .ZN(n14006) );
  OR2_X1 U11708 ( .A1(n9032), .A2(n14006), .ZN(n9231) );
  INV_X1 U11709 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9229) );
  OR2_X1 U11710 ( .A1(n9442), .A2(n9229), .ZN(n9230) );
  INV_X1 U11711 ( .A(n14011), .ZN(n14122) );
  NAND2_X1 U11712 ( .A1(n10891), .A2(n9466), .ZN(n9236) );
  NAND2_X1 U11713 ( .A1(n9243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9234) );
  XNOR2_X1 U11714 ( .A(n9234), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14874) );
  AOI22_X1 U11715 ( .A1(n9465), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9266), 
        .B2(n14874), .ZN(n9235) );
  MUX2_X1 U11716 ( .A(n14122), .B(n14804), .S(n9468), .Z(n9240) );
  NAND2_X1 U11717 ( .A1(n9239), .A2(n9240), .ZN(n9238) );
  MUX2_X1 U11718 ( .A(n14122), .B(n14804), .S(n9413), .Z(n9237) );
  INV_X1 U11719 ( .A(n9239), .ZN(n9242) );
  INV_X1 U11720 ( .A(n9240), .ZN(n9241) );
  NAND2_X1 U11721 ( .A1(n10996), .A2(n9466), .ZN(n9246) );
  OAI21_X1 U11722 ( .B1(n9243), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9244) );
  XNOR2_X1 U11723 ( .A(n9244), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14211) );
  AOI22_X1 U11724 ( .A1(n9465), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9266), 
        .B2(n14211), .ZN(n9245) );
  NAND2_X1 U11725 ( .A1(n8923), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9255) );
  INV_X1 U11726 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14426) );
  OR2_X1 U11727 ( .A1(n9015), .A2(n14426), .ZN(n9254) );
  INV_X1 U11728 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14210) );
  OR2_X1 U11729 ( .A1(n9443), .A2(n14210), .ZN(n9253) );
  NAND2_X1 U11730 ( .A1(n9250), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9248) );
  INV_X1 U11731 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U11732 ( .A1(n9248), .A2(n9247), .ZN(n9251) );
  AND2_X1 U11733 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n9249) );
  NAND2_X1 U11734 ( .A1(n9251), .A2(n9269), .ZN(n14425) );
  OR2_X1 U11735 ( .A1(n9032), .A2(n14425), .ZN(n9252) );
  INV_X1 U11736 ( .A(n14072), .ZN(n14121) );
  NAND2_X1 U11737 ( .A1(n14510), .A2(n14121), .ZN(n9989) );
  INV_X1 U11738 ( .A(n9989), .ZN(n9276) );
  NOR2_X1 U11739 ( .A1(n14510), .A2(n14121), .ZN(n9990) );
  NAND2_X1 U11740 ( .A1(n9256), .A2(n9466), .ZN(n9258) );
  AOI22_X1 U11741 ( .A1(n9465), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14415), 
        .B2(n9266), .ZN(n9257) );
  INV_X1 U11742 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n14070) );
  INV_X1 U11743 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13976) );
  AND2_X1 U11744 ( .A1(n9271), .A2(n13976), .ZN(n9259) );
  OR2_X1 U11745 ( .A1(n9259), .A2(n9291), .ZN(n14395) );
  AOI22_X1 U11746 ( .A1(n9439), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9014), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U11747 ( .A1(n8923), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9260) );
  OAI211_X1 U11748 ( .C1(n14395), .C2(n9032), .A(n9261), .B(n9260), .ZN(n14119) );
  INV_X1 U11749 ( .A(n14119), .ZN(n14038) );
  NAND2_X1 U11750 ( .A1(n11419), .A2(n9466), .ZN(n9268) );
  NAND2_X1 U11751 ( .A1(n9262), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9264) );
  XNOR2_X1 U11752 ( .A(n9264), .B(n9263), .ZN(n14906) );
  INV_X1 U11753 ( .A(n14906), .ZN(n9265) );
  AOI22_X1 U11754 ( .A1(n9465), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9266), 
        .B2(n9265), .ZN(n9267) );
  NAND2_X1 U11755 ( .A1(n8923), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11756 ( .A1(n9269), .A2(n14070), .ZN(n9270) );
  NAND2_X1 U11757 ( .A1(n9271), .A2(n9270), .ZN(n14069) );
  OR2_X1 U11758 ( .A1(n14069), .A2(n9032), .ZN(n9274) );
  INV_X1 U11759 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14900) );
  OR2_X1 U11760 ( .A1(n9015), .A2(n14900), .ZN(n9273) );
  INV_X1 U11761 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14895) );
  OR2_X1 U11762 ( .A1(n9443), .A2(n14895), .ZN(n9272) );
  OAI211_X1 U11763 ( .C1(n9276), .C2(n9990), .A(n9472), .B(n10052), .ZN(n9277)
         );
  NAND2_X1 U11764 ( .A1(n14498), .A2(n14038), .ZN(n10056) );
  NAND2_X1 U11765 ( .A1(n14502), .A2(n14010), .ZN(n9473) );
  NAND2_X1 U11766 ( .A1(n10056), .A2(n9473), .ZN(n9283) );
  NAND3_X1 U11767 ( .A1(n14510), .A2(n14072), .A3(n9413), .ZN(n9278) );
  NAND2_X1 U11768 ( .A1(n14010), .A2(n9447), .ZN(n9279) );
  NAND2_X1 U11769 ( .A1(n9278), .A2(n9279), .ZN(n9281) );
  NOR2_X1 U11770 ( .A1(n9279), .A2(n14121), .ZN(n9280) );
  AOI22_X1 U11771 ( .A1(n14502), .A2(n9281), .B1(n9280), .B2(n14510), .ZN(
        n9282) );
  MUX2_X1 U11772 ( .A(n9413), .B(n9282), .S(n9472), .Z(n9289) );
  INV_X1 U11773 ( .A(n9283), .ZN(n9287) );
  INV_X1 U11774 ( .A(n14010), .ZN(n14120) );
  NAND2_X1 U11775 ( .A1(n14120), .A2(n9468), .ZN(n9285) );
  OR3_X1 U11776 ( .A1(n14510), .A2(n9447), .A3(n14072), .ZN(n9284) );
  OAI21_X1 U11777 ( .B1(n14502), .B2(n9285), .A(n9284), .ZN(n9286) );
  NAND2_X1 U11778 ( .A1(n9287), .A2(n9286), .ZN(n9288) );
  OAI211_X1 U11779 ( .C1(n10056), .C2(n9468), .A(n9289), .B(n9288), .ZN(n9290)
         );
  OR2_X1 U11780 ( .A1(n9291), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U11781 ( .A1(n9291), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9305) );
  AND2_X1 U11782 ( .A1(n9292), .A2(n9305), .ZN(n14378) );
  INV_X1 U11783 ( .A(n9032), .ZN(n9293) );
  NAND2_X1 U11784 ( .A1(n14378), .A2(n9293), .ZN(n9296) );
  AOI22_X1 U11785 ( .A1(n9014), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n8923), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n9295) );
  NAND2_X1 U11786 ( .A1(n9439), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11787 ( .A1(n11762), .A2(n9466), .ZN(n9298) );
  OR2_X1 U11788 ( .A1(n9436), .A2(n11763), .ZN(n9297) );
  INV_X1 U11789 ( .A(n14492), .ZN(n14381) );
  MUX2_X1 U11790 ( .A(n13984), .B(n14381), .S(n9468), .Z(n9300) );
  INV_X1 U11791 ( .A(n13984), .ZN(n14118) );
  MUX2_X1 U11792 ( .A(n14492), .B(n14118), .S(n9468), .Z(n9299) );
  NAND2_X1 U11793 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  INV_X1 U11794 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n13082) );
  OR2_X1 U11795 ( .A1(n9417), .A2(n13082), .ZN(n9310) );
  INV_X1 U11796 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9304) );
  OR2_X1 U11797 ( .A1(n9015), .A2(n9304), .ZN(n9309) );
  NAND2_X1 U11798 ( .A1(n9306), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9316) );
  OAI21_X1 U11799 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n9306), .A(n9316), .ZN(
        n14363) );
  OR2_X1 U11800 ( .A1(n9032), .A2(n14363), .ZN(n9308) );
  INV_X1 U11801 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n13033) );
  OR2_X1 U11802 ( .A1(n9442), .A2(n13033), .ZN(n9307) );
  NAND4_X1 U11803 ( .A1(n9310), .A2(n9309), .A3(n9308), .A4(n9307), .ZN(n14117) );
  NAND2_X1 U11804 ( .A1(n11819), .A2(n9466), .ZN(n9312) );
  OR2_X1 U11805 ( .A1(n9436), .A2(n11822), .ZN(n9311) );
  MUX2_X1 U11806 ( .A(n14117), .B(n14486), .S(n9413), .Z(n9314) );
  NAND2_X1 U11807 ( .A1(n9439), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9322) );
  INV_X1 U11808 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9315) );
  OR2_X1 U11809 ( .A1(n9443), .A2(n9315), .ZN(n9321) );
  NAND2_X1 U11810 ( .A1(n9317), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9329) );
  OAI21_X1 U11811 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n9317), .A(n9329), .ZN(
        n14345) );
  OR2_X1 U11812 ( .A1(n9032), .A2(n14345), .ZN(n9320) );
  INV_X1 U11813 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9318) );
  OR2_X1 U11814 ( .A1(n9442), .A2(n9318), .ZN(n9319) );
  INV_X1 U11815 ( .A(n13983), .ZN(n14116) );
  OR2_X1 U11816 ( .A1(n9324), .A2(n10476), .ZN(n9325) );
  INV_X1 U11817 ( .A(n14348), .ZN(n14482) );
  MUX2_X1 U11818 ( .A(n14116), .B(n14482), .S(n9468), .Z(n9327) );
  MUX2_X1 U11819 ( .A(n13983), .B(n14348), .S(n9413), .Z(n9326) );
  NAND2_X1 U11820 ( .A1(n9014), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9334) );
  INV_X1 U11821 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9328) );
  OR2_X1 U11822 ( .A1(n9015), .A2(n9328), .ZN(n9333) );
  NAND2_X1 U11823 ( .A1(n9330), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9340) );
  OAI21_X1 U11824 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9330), .A(n9340), .ZN(
        n14320) );
  OR2_X1 U11825 ( .A1(n9032), .A2(n14320), .ZN(n9332) );
  INV_X1 U11826 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n14523) );
  OR2_X1 U11827 ( .A1(n9442), .A2(n14523), .ZN(n9331) );
  NAND4_X1 U11828 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n14115) );
  NAND2_X1 U11829 ( .A1(n12070), .A2(n9466), .ZN(n9336) );
  OR2_X1 U11830 ( .A1(n9436), .A2(n12073), .ZN(n9335) );
  MUX2_X1 U11831 ( .A(n14115), .B(n14472), .S(n9447), .Z(n9338) );
  INV_X1 U11832 ( .A(n9338), .ZN(n9339) );
  NAND2_X1 U11833 ( .A1(n9439), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9346) );
  INV_X1 U11834 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n13211) );
  OR2_X1 U11835 ( .A1(n9417), .A2(n13211), .ZN(n9345) );
  INV_X1 U11836 ( .A(n9340), .ZN(n9341) );
  NAND2_X1 U11837 ( .A1(n9341), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9358) );
  OAI21_X1 U11838 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9341), .A(n9358), .ZN(
        n14312) );
  OR2_X1 U11839 ( .A1(n9032), .A2(n14312), .ZN(n9344) );
  INV_X1 U11840 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9342) );
  OR2_X1 U11841 ( .A1(n9442), .A2(n9342), .ZN(n9343) );
  INV_X1 U11842 ( .A(n13949), .ZN(n14114) );
  NAND2_X1 U11843 ( .A1(n12104), .A2(n9466), .ZN(n9348) );
  OR2_X1 U11844 ( .A1(n9436), .A2(n12602), .ZN(n9347) );
  MUX2_X1 U11845 ( .A(n14114), .B(n14314), .S(n9413), .Z(n9349) );
  NAND2_X1 U11846 ( .A1(n9350), .A2(n9349), .ZN(n9356) );
  INV_X1 U11847 ( .A(n9351), .ZN(n9354) );
  INV_X1 U11848 ( .A(n9352), .ZN(n9353) );
  NAND2_X1 U11849 ( .A1(n9354), .A2(n9353), .ZN(n9355) );
  NAND2_X1 U11850 ( .A1(n9356), .A2(n9355), .ZN(n9368) );
  NAND2_X1 U11851 ( .A1(n9439), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9364) );
  INV_X1 U11852 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9357) );
  OR2_X1 U11853 ( .A1(n9417), .A2(n9357), .ZN(n9363) );
  INV_X1 U11854 ( .A(n9358), .ZN(n9359) );
  NAND2_X1 U11855 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n9359), .ZN(n9373) );
  OAI21_X1 U11856 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9359), .A(n9373), .ZN(
        n14288) );
  OR2_X1 U11857 ( .A1(n9032), .A2(n14288), .ZN(n9362) );
  INV_X1 U11858 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9360) );
  OR2_X1 U11859 ( .A1(n9442), .A2(n9360), .ZN(n9361) );
  NAND4_X1 U11860 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n14113) );
  NAND2_X1 U11861 ( .A1(n12175), .A2(n9466), .ZN(n9366) );
  OR2_X1 U11862 ( .A1(n9436), .A2(n6736), .ZN(n9365) );
  NAND2_X2 U11863 ( .A1(n9366), .A2(n9365), .ZN(n14460) );
  MUX2_X1 U11864 ( .A(n14113), .B(n14460), .S(n9413), .Z(n9369) );
  NAND2_X1 U11865 ( .A1(n9014), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9379) );
  INV_X1 U11866 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9370) );
  OR2_X1 U11867 ( .A1(n9015), .A2(n9370), .ZN(n9378) );
  INV_X1 U11868 ( .A(n9373), .ZN(n9371) );
  NAND2_X1 U11869 ( .A1(n9371), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9402) );
  INV_X1 U11870 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9372) );
  NAND2_X1 U11871 ( .A1(n9373), .A2(n9372), .ZN(n9374) );
  NAND2_X1 U11872 ( .A1(n9402), .A2(n9374), .ZN(n14084) );
  OR2_X1 U11873 ( .A1(n9032), .A2(n14084), .ZN(n9377) );
  INV_X1 U11874 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9375) );
  OR2_X1 U11875 ( .A1(n9442), .A2(n9375), .ZN(n9376) );
  NAND4_X1 U11876 ( .A1(n9379), .A2(n9378), .A3(n9377), .A4(n9376), .ZN(n14112) );
  NAND2_X1 U11877 ( .A1(n12255), .A2(n9466), .ZN(n9381) );
  OR2_X1 U11878 ( .A1(n9436), .A2(n12256), .ZN(n9380) );
  MUX2_X1 U11879 ( .A(n14112), .B(n14455), .S(n9468), .Z(n9385) );
  NAND2_X1 U11880 ( .A1(n9384), .A2(n9385), .ZN(n9383) );
  MUX2_X1 U11881 ( .A(n14112), .B(n14455), .S(n9413), .Z(n9382) );
  NAND2_X1 U11882 ( .A1(n9383), .A2(n9382), .ZN(n9389) );
  INV_X1 U11883 ( .A(n9385), .ZN(n9386) );
  NAND2_X1 U11884 ( .A1(n9387), .A2(n9386), .ZN(n9388) );
  NAND2_X1 U11885 ( .A1(n9014), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9394) );
  INV_X1 U11886 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9390) );
  OR2_X1 U11887 ( .A1(n9015), .A2(n9390), .ZN(n9393) );
  INV_X1 U11888 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13935) );
  XNOR2_X1 U11889 ( .A(n9402), .B(n13935), .ZN(n13934) );
  OR2_X1 U11890 ( .A1(n9032), .A2(n13934), .ZN(n9392) );
  INV_X1 U11891 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n13208) );
  OR2_X1 U11892 ( .A1(n9442), .A2(n13208), .ZN(n9391) );
  NAND4_X1 U11893 ( .A1(n9394), .A2(n9393), .A3(n9392), .A4(n9391), .ZN(n14111) );
  NAND2_X1 U11894 ( .A1(n13925), .A2(n9466), .ZN(n9396) );
  OR2_X1 U11895 ( .A1(n9436), .A2(n7419), .ZN(n9395) );
  MUX2_X1 U11896 ( .A(n14111), .B(n14450), .S(n9413), .Z(n9399) );
  MUX2_X1 U11897 ( .A(n14111), .B(n14450), .S(n9468), .Z(n9397) );
  NAND2_X1 U11898 ( .A1(n9439), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9410) );
  INV_X1 U11899 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9400) );
  OR2_X1 U11900 ( .A1(n9443), .A2(n9400), .ZN(n9409) );
  INV_X1 U11901 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9401) );
  OAI21_X1 U11902 ( .B1(n9402), .B2(n13935), .A(n9401), .ZN(n9405) );
  INV_X1 U11903 ( .A(n9402), .ZN(n9404) );
  AND2_X1 U11904 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9403) );
  NAND2_X1 U11905 ( .A1(n9404), .A2(n9403), .ZN(n10073) );
  NAND2_X1 U11906 ( .A1(n9405), .A2(n10073), .ZN(n14240) );
  OR2_X1 U11907 ( .A1(n9032), .A2(n14240), .ZN(n9408) );
  INV_X1 U11908 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9406) );
  OR2_X1 U11909 ( .A1(n9442), .A2(n9406), .ZN(n9407) );
  NAND4_X1 U11910 ( .A1(n9410), .A2(n9409), .A3(n9408), .A4(n9407), .ZN(n14110) );
  NAND2_X1 U11911 ( .A1(n12290), .A2(n9466), .ZN(n9412) );
  INV_X1 U11912 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13127) );
  OR2_X1 U11913 ( .A1(n9436), .A2(n13127), .ZN(n9411) );
  MUX2_X1 U11914 ( .A(n14110), .B(n14446), .S(n9468), .Z(n9415) );
  MUX2_X1 U11915 ( .A(n14110), .B(n14446), .S(n9413), .Z(n9414) );
  INV_X1 U11916 ( .A(n9415), .ZN(n9416) );
  NAND2_X1 U11917 ( .A1(n9439), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U11918 ( .A1(n8923), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9420) );
  INV_X1 U11919 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n13096) );
  OR2_X1 U11920 ( .A1(n9417), .A2(n13096), .ZN(n9419) );
  OR2_X1 U11921 ( .A1(n9032), .A2(n10073), .ZN(n9418) );
  NAND4_X1 U11922 ( .A1(n9421), .A2(n9420), .A3(n9419), .A4(n9418), .ZN(n14109) );
  INV_X1 U11923 ( .A(n9422), .ZN(n9423) );
  INV_X1 U11924 ( .A(SI_28_), .ZN(n13422) );
  NAND2_X1 U11925 ( .A1(n9423), .A2(n13422), .ZN(n9424) );
  INV_X1 U11926 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12333) );
  INV_X1 U11927 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13916) );
  MUX2_X1 U11928 ( .A(n12333), .B(n13916), .S(n10476), .Z(n9431) );
  XNOR2_X1 U11929 ( .A(n9431), .B(SI_29_), .ZN(n9433) );
  NAND2_X1 U11930 ( .A1(n12332), .A2(n9466), .ZN(n9428) );
  OR2_X1 U11931 ( .A1(n9436), .A2(n12333), .ZN(n9427) );
  MUX2_X1 U11932 ( .A(n14109), .B(n14441), .S(n9447), .Z(n9429) );
  MUX2_X1 U11933 ( .A(n14109), .B(n14441), .S(n9468), .Z(n9430) );
  INV_X1 U11934 ( .A(n9431), .ZN(n9432) );
  INV_X1 U11935 ( .A(n9457), .ZN(n9435) );
  INV_X1 U11936 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14539) );
  INV_X1 U11937 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13914) );
  MUX2_X1 U11938 ( .A(n14539), .B(n13914), .S(n10476), .Z(n9458) );
  XNOR2_X1 U11939 ( .A(n9458), .B(SI_30_), .ZN(n9456) );
  NAND2_X1 U11940 ( .A1(n13912), .A2(n9466), .ZN(n9438) );
  OR2_X1 U11941 ( .A1(n9436), .A2(n14539), .ZN(n9437) );
  INV_X1 U11942 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n13084) );
  NAND2_X1 U11943 ( .A1(n9439), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U11944 ( .A1(n9014), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9440) );
  OAI211_X1 U11945 ( .C1(n9442), .C2(n13084), .A(n9441), .B(n9440), .ZN(n14108) );
  INV_X1 U11946 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U11947 ( .A1(n8923), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9445) );
  INV_X1 U11948 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n13080) );
  OR2_X1 U11949 ( .A1(n9443), .A2(n13080), .ZN(n9444) );
  OAI211_X1 U11950 ( .C1(n9015), .C2(n9446), .A(n9445), .B(n9444), .ZN(n14224)
         );
  NAND2_X1 U11951 ( .A1(n14224), .A2(n9447), .ZN(n9469) );
  NAND2_X1 U11952 ( .A1(n9469), .A2(n9448), .ZN(n9449) );
  AOI22_X1 U11953 ( .A1(n14231), .A2(n9468), .B1(n14108), .B2(n9449), .ZN(
        n9453) );
  INV_X1 U11954 ( .A(n9450), .ZN(n9451) );
  OAI21_X1 U11955 ( .B1(n14224), .B2(n9451), .A(n14108), .ZN(n9452) );
  MUX2_X1 U11956 ( .A(n14438), .B(n9452), .S(n9468), .Z(n9454) );
  NOR2_X1 U11957 ( .A1(n14547), .A2(n10681), .ZN(n9455) );
  OR2_X1 U11958 ( .A1(n10180), .A2(n14218), .ZN(n14674) );
  OAI21_X1 U11959 ( .B1(n9455), .B2(n10513), .A(n14674), .ZN(n9501) );
  OR2_X1 U11960 ( .A1(n9520), .A2(n11764), .ZN(n9497) );
  INV_X1 U11961 ( .A(n14224), .ZN(n9467) );
  NAND2_X1 U11962 ( .A1(n9457), .A2(n9456), .ZN(n9461) );
  INV_X1 U11963 ( .A(n9458), .ZN(n9459) );
  NAND2_X1 U11964 ( .A1(n9459), .A2(SI_30_), .ZN(n9460) );
  NAND2_X1 U11965 ( .A1(n9461), .A2(n9460), .ZN(n9464) );
  MUX2_X1 U11966 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10476), .Z(n9462) );
  XNOR2_X1 U11967 ( .A(n9462), .B(SI_31_), .ZN(n9463) );
  XNOR2_X1 U11968 ( .A(n9464), .B(n9463), .ZN(n9742) );
  MUX2_X1 U11969 ( .A(n9468), .B(n9467), .S(n14435), .Z(n9471) );
  INV_X1 U11970 ( .A(n9469), .ZN(n9470) );
  XNOR2_X1 U11971 ( .A(n14435), .B(n14224), .ZN(n9502) );
  XOR2_X1 U11972 ( .A(n14108), .B(n14231), .Z(n9493) );
  XNOR2_X1 U11973 ( .A(n14455), .B(n14112), .ZN(n14266) );
  INV_X1 U11974 ( .A(n14266), .ZN(n14275) );
  INV_X1 U11975 ( .A(n14285), .ZN(n14291) );
  XNOR2_X1 U11976 ( .A(n14314), .B(n13949), .ZN(n14299) );
  XNOR2_X1 U11977 ( .A(n14472), .B(n14115), .ZN(n14327) );
  XNOR2_X1 U11978 ( .A(n14348), .B(n13983), .ZN(n14350) );
  XNOR2_X1 U11979 ( .A(n14492), .B(n13984), .ZN(n14373) );
  NAND2_X1 U11980 ( .A1(n9472), .A2(n10056), .ZN(n14389) );
  INV_X1 U11981 ( .A(n12121), .ZN(n9485) );
  XNOR2_X1 U11982 ( .A(n14827), .B(n14124), .ZN(n11972) );
  INV_X1 U11983 ( .A(n11972), .ZN(n11975) );
  XNOR2_X1 U11984 ( .A(n14804), .B(n14011), .ZN(n12166) );
  OR2_X1 U11985 ( .A1(n15022), .A2(n11737), .ZN(n10041) );
  NAND2_X1 U11986 ( .A1(n15022), .A2(n11737), .ZN(n9475) );
  NAND2_X1 U11987 ( .A1(n10041), .A2(n9475), .ZN(n11773) );
  XNOR2_X1 U11988 ( .A(n15006), .B(n14130), .ZN(n11508) );
  OR2_X1 U11989 ( .A1(n11878), .A2(n11528), .ZN(n10037) );
  NAND2_X1 U11990 ( .A1(n11878), .A2(n11528), .ZN(n9476) );
  NAND2_X1 U11991 ( .A1(n10037), .A2(n9476), .ZN(n11399) );
  NAND2_X1 U11992 ( .A1(n14999), .A2(n14131), .ZN(n9477) );
  NAND2_X1 U11993 ( .A1(n11658), .A2(n10234), .ZN(n10035) );
  NAND2_X1 U11994 ( .A1(n14994), .A2(n14132), .ZN(n9478) );
  NAND2_X1 U11995 ( .A1(n11287), .A2(n11316), .ZN(n14915) );
  INV_X1 U11996 ( .A(n11324), .ZN(n9963) );
  INV_X1 U11997 ( .A(n11369), .ZN(n9966) );
  INV_X1 U11998 ( .A(n11383), .ZN(n9480) );
  NOR4_X1 U11999 ( .A1(n9963), .A2(n9966), .A3(n9480), .A4(n9960), .ZN(n9481)
         );
  XNOR2_X1 U12000 ( .A(n14134), .B(n10206), .ZN(n14935) );
  NAND4_X1 U12001 ( .A1(n10034), .A2(n11387), .A3(n9481), .A4(n14935), .ZN(
        n9482) );
  NOR4_X1 U12002 ( .A1(n11773), .A2(n7572), .A3(n11399), .A4(n9482), .ZN(n9483) );
  XNOR2_X1 U12003 ( .A(n14679), .B(n14125), .ZN(n11993) );
  XNOR2_X1 U12004 ( .A(n11740), .B(n14126), .ZN(n10042) );
  XNOR2_X1 U12005 ( .A(n12010), .B(n11769), .ZN(n10038) );
  INV_X1 U12006 ( .A(n10038), .ZN(n11526) );
  NAND4_X1 U12007 ( .A1(n9483), .A2(n11993), .A3(n10042), .A4(n11526), .ZN(
        n9484) );
  NOR4_X1 U12008 ( .A1(n9485), .A2(n11975), .A3(n12166), .A4(n9484), .ZN(n9486) );
  NAND4_X1 U12009 ( .A1(n14402), .A2(n9486), .A3(n12086), .A4(n6553), .ZN(
        n9487) );
  NOR3_X1 U12010 ( .A1(n14373), .A2(n14389), .A3(n9487), .ZN(n9488) );
  XNOR2_X1 U12011 ( .A(n14486), .B(n14117), .ZN(n14355) );
  NAND4_X1 U12012 ( .A1(n14327), .A2(n14350), .A3(n9488), .A4(n14355), .ZN(
        n9489) );
  NOR4_X1 U12013 ( .A1(n14275), .A2(n14291), .A3(n14299), .A4(n9489), .ZN(
        n9491) );
  XNOR2_X1 U12014 ( .A(n14450), .B(n14111), .ZN(n14261) );
  NAND2_X1 U12015 ( .A1(n14446), .A2(n14110), .ZN(n10003) );
  OR2_X1 U12016 ( .A1(n14446), .A2(n14110), .ZN(n9490) );
  NAND2_X1 U12017 ( .A1(n10003), .A2(n9490), .ZN(n14235) );
  NAND4_X1 U12018 ( .A1(n10062), .A2(n9491), .A3(n14261), .A4(n14235), .ZN(
        n9492) );
  NOR3_X1 U12019 ( .A1(n9502), .A2(n9493), .A3(n9492), .ZN(n9494) );
  XNOR2_X1 U12020 ( .A(n9494), .B(n14415), .ZN(n9498) );
  NAND2_X1 U12021 ( .A1(n9502), .A2(n7616), .ZN(n9495) );
  MUX2_X1 U12022 ( .A(n9501), .B(n9495), .S(n6577), .Z(n9496) );
  OAI21_X1 U12023 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9499) );
  INV_X1 U12024 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U12025 ( .A1(n6697), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9506) );
  MUX2_X1 U12026 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9506), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9507) );
  NAND2_X1 U12027 ( .A1(n9507), .A2(n9513), .ZN(n10514) );
  OR2_X1 U12028 ( .A1(n10514), .A2(P1_U3086), .ZN(n12071) );
  OAI21_X1 U12029 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9527) );
  INV_X1 U12030 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9511) );
  XNOR2_X1 U12031 ( .A(n9515), .B(n9514), .ZN(n10005) );
  NAND2_X1 U12032 ( .A1(n9516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9518) );
  INV_X1 U12033 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9517) );
  NAND2_X1 U12034 ( .A1(n14547), .A2(n14415), .ZN(n9522) );
  NAND2_X1 U12035 ( .A1(n9520), .A2(n10681), .ZN(n9521) );
  NAND2_X1 U12036 ( .A1(n14937), .A2(n10513), .ZN(n9523) );
  NAND2_X1 U12037 ( .A1(n10395), .A2(n10511), .ZN(n10691) );
  INV_X1 U12038 ( .A(n10691), .ZN(n10781) );
  INV_X1 U12039 ( .A(n9524), .ZN(n14151) );
  INV_X1 U12040 ( .A(n14545), .ZN(n14857) );
  NAND3_X1 U12041 ( .A1(n10781), .A2(n14052), .A3(n14857), .ZN(n9525) );
  OAI211_X1 U12042 ( .C1(n14547), .C2(n12071), .A(n9525), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9526) );
  NAND2_X1 U12043 ( .A1(n9527), .A2(n9526), .ZN(P1_U3242) );
  NAND2_X1 U12044 ( .A1(n13368), .A2(n12529), .ZN(n9528) );
  INV_X1 U12045 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9564) );
  AOI22_X1 U12046 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n9564), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n13127), .ZN(n9532) );
  INV_X1 U12047 ( .A(n9532), .ZN(n9533) );
  XNOR2_X1 U12048 ( .A(n9565), .B(n9533), .ZN(n13417) );
  NAND2_X1 U12049 ( .A1(n13417), .A2(n12370), .ZN(n9535) );
  OR2_X1 U12050 ( .A1(n12358), .A2(n13422), .ZN(n9534) );
  NAND2_X1 U12051 ( .A1(n12301), .A2(n6543), .ZN(n9578) );
  INV_X1 U12052 ( .A(n9536), .ZN(n9538) );
  INV_X1 U12053 ( .A(n12399), .ZN(n9537) );
  NAND2_X1 U12054 ( .A1(n9538), .A2(n9537), .ZN(n9539) );
  NAND3_X1 U12055 ( .A1(n9563), .A2(n15341), .A3(n9539), .ZN(n9545) );
  NAND2_X1 U12056 ( .A1(n14719), .A2(n7736), .ZN(n12366) );
  INV_X1 U12057 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n13187) );
  NAND2_X1 U12058 ( .A1(n12360), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U12059 ( .A1(n9570), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9540) );
  OAI211_X1 U12060 ( .C1(n13187), .C2(n12363), .A(n9541), .B(n9540), .ZN(n9542) );
  INV_X1 U12061 ( .A(n9542), .ZN(n9543) );
  NAND2_X1 U12062 ( .A1(n12366), .A2(n9543), .ZN(n12707) );
  AOI22_X1 U12063 ( .A1(n15326), .A2(n12921), .B1(n12707), .B2(n15324), .ZN(
        n9544) );
  OR2_X1 U12064 ( .A1(n9547), .A2(n9537), .ZN(n9548) );
  NAND2_X1 U12065 ( .A1(n9579), .A2(n9548), .ZN(n12902) );
  NAND2_X1 U12066 ( .A1(n12902), .A2(n15411), .ZN(n9549) );
  NAND2_X1 U12067 ( .A1(n12904), .A2(n9549), .ZN(n9560) );
  NOR2_X1 U12068 ( .A1(n12547), .A2(n9550), .ZN(n12318) );
  NAND2_X1 U12069 ( .A1(n11219), .A2(n12318), .ZN(n12554) );
  NAND2_X1 U12070 ( .A1(n12350), .A2(n9551), .ZN(n12400) );
  NOR2_X1 U12071 ( .A1(n12400), .A2(n9552), .ZN(n10160) );
  NAND2_X1 U12072 ( .A1(n11219), .A2(n10160), .ZN(n10154) );
  NAND2_X1 U12073 ( .A1(n12554), .A2(n10154), .ZN(n9553) );
  INV_X1 U12074 ( .A(n10083), .ZN(n13409) );
  NAND2_X1 U12075 ( .A1(n9553), .A2(n10157), .ZN(n9557) );
  NAND2_X1 U12076 ( .A1(n10083), .A2(n9554), .ZN(n9555) );
  NOR2_X1 U12077 ( .A1(n9555), .A2(n13407), .ZN(n10159) );
  NAND3_X1 U12078 ( .A1(n11219), .A2(n10159), .A3(n10162), .ZN(n9556) );
  INV_X1 U12079 ( .A(n9558), .ZN(n9559) );
  NAND2_X1 U12080 ( .A1(n9559), .A2(n7615), .ZN(P3_U3455) );
  INV_X1 U12081 ( .A(n9561), .ZN(n9562) );
  NAND2_X1 U12082 ( .A1(n9562), .A2(n7625), .ZN(P3_U3487) );
  NAND2_X1 U12083 ( .A1(n9563), .A2(n7637), .ZN(n9569) );
  OAI22_X1 U12084 ( .A1(n12333), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n13916), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12353) );
  INV_X1 U12085 ( .A(SI_29_), .ZN(n12286) );
  NOR2_X1 U12086 ( .A1(n7729), .A2(n12286), .ZN(n9566) );
  NAND2_X1 U12087 ( .A1(n12894), .A2(n12707), .ZN(n12539) );
  INV_X1 U12088 ( .A(n12894), .ZN(n9568) );
  INV_X1 U12089 ( .A(n12707), .ZN(n9567) );
  NAND2_X1 U12090 ( .A1(n9568), .A2(n9567), .ZN(n12540) );
  NAND2_X1 U12091 ( .A1(n12539), .A2(n12540), .ZN(n12543) );
  XNOR2_X1 U12092 ( .A(n9569), .B(n12543), .ZN(n9577) );
  INV_X1 U12093 ( .A(n6543), .ZN(n9575) );
  INV_X1 U12094 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14750) );
  AOI22_X1 U12095 ( .A1(n12360), .A2(P3_REG0_REG_30__SCAN_IN), .B1(n9570), 
        .B2(P3_REG2_REG_30__SCAN_IN), .ZN(n9571) );
  OAI211_X1 U12096 ( .C1(n12363), .C2(n14750), .A(n12366), .B(n9571), .ZN(
        n12381) );
  INV_X1 U12097 ( .A(n12381), .ZN(n12546) );
  INV_X1 U12098 ( .A(P3_B_REG_SCAN_IN), .ZN(n9572) );
  OR2_X1 U12099 ( .A1(n13420), .A2(n9572), .ZN(n9573) );
  NAND2_X1 U12100 ( .A1(n15324), .A2(n9573), .ZN(n14716) );
  NOR2_X1 U12101 ( .A1(n12546), .A2(n14716), .ZN(n9574) );
  INV_X1 U12102 ( .A(n15430), .ZN(n9580) );
  OR2_X1 U12103 ( .A1(n10407), .A2(n9580), .ZN(n9584) );
  INV_X1 U12104 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9581) );
  OAI22_X1 U12105 ( .A1(n12894), .A2(n13392), .B1(n15430), .B2(n9581), .ZN(
        n9582) );
  INV_X1 U12106 ( .A(n9582), .ZN(n9583) );
  NAND2_X1 U12107 ( .A1(n9584), .A2(n9583), .ZN(P3_U3456) );
  NAND2_X1 U12108 ( .A1(n9589), .A2(n9799), .ZN(n9592) );
  AOI21_X1 U12109 ( .B1(n13700), .B2(n9586), .A(n9804), .ZN(n9587) );
  NAND2_X1 U12110 ( .A1(n9799), .A2(n15166), .ZN(n9591) );
  NAND2_X1 U12111 ( .A1(n9589), .A2(n9588), .ZN(n9590) );
  NAND2_X1 U12112 ( .A1(n9593), .A2(n9592), .ZN(n9594) );
  NAND2_X1 U12113 ( .A1(n13551), .A2(n6542), .ZN(n9597) );
  NAND2_X1 U12114 ( .A1(n9798), .A2(n15171), .ZN(n9596) );
  AND2_X1 U12115 ( .A1(n9597), .A2(n9596), .ZN(n9601) );
  NAND2_X1 U12116 ( .A1(n9798), .A2(n13551), .ZN(n9599) );
  NAND2_X1 U12117 ( .A1(n6542), .A2(n15171), .ZN(n9598) );
  NAND2_X1 U12118 ( .A1(n9599), .A2(n9598), .ZN(n9600) );
  NAND2_X1 U12119 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  NAND2_X1 U12120 ( .A1(n9798), .A2(n13549), .ZN(n9606) );
  NAND2_X1 U12121 ( .A1(n6542), .A2(n15199), .ZN(n9605) );
  NAND2_X1 U12122 ( .A1(n9606), .A2(n9605), .ZN(n9609) );
  NAND2_X1 U12123 ( .A1(n13549), .A2(n9799), .ZN(n9607) );
  OAI21_X1 U12124 ( .B1(n6542), .B2(n11684), .A(n9607), .ZN(n9608) );
  NAND2_X1 U12125 ( .A1(n11574), .A2(n9798), .ZN(n9611) );
  NAND2_X1 U12126 ( .A1(n6898), .A2(n9656), .ZN(n9610) );
  NAND2_X1 U12127 ( .A1(n9611), .A2(n9610), .ZN(n9616) );
  NAND2_X1 U12128 ( .A1(n9615), .A2(n9616), .ZN(n9614) );
  INV_X1 U12129 ( .A(n13548), .ZN(n10897) );
  NAND2_X1 U12130 ( .A1(n11574), .A2(n6542), .ZN(n9612) );
  OAI21_X1 U12131 ( .B1(n10897), .B2(n6542), .A(n9612), .ZN(n9613) );
  NAND2_X1 U12132 ( .A1(n9614), .A2(n9613), .ZN(n9620) );
  INV_X1 U12133 ( .A(n9615), .ZN(n9618) );
  INV_X1 U12134 ( .A(n9616), .ZN(n9617) );
  NAND2_X1 U12135 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  NAND2_X1 U12136 ( .A1(n11259), .A2(n9656), .ZN(n9622) );
  NAND2_X1 U12137 ( .A1(n6544), .A2(n13547), .ZN(n9621) );
  NAND2_X1 U12138 ( .A1(n9622), .A2(n9621), .ZN(n9625) );
  AOI22_X1 U12139 ( .A1(n11259), .A2(n6544), .B1(n13547), .B2(n9656), .ZN(
        n9623) );
  NAND2_X1 U12140 ( .A1(n11274), .A2(n6544), .ZN(n9628) );
  NAND2_X1 U12141 ( .A1(n13546), .A2(n9656), .ZN(n9627) );
  NAND2_X1 U12142 ( .A1(n9628), .A2(n9627), .ZN(n9630) );
  AOI22_X1 U12143 ( .A1(n11274), .A2(n6542), .B1(n6544), .B2(n13546), .ZN(
        n9629) );
  NAND2_X1 U12144 ( .A1(n11689), .A2(n9656), .ZN(n9633) );
  NAND2_X1 U12145 ( .A1(n6544), .A2(n13545), .ZN(n9632) );
  INV_X1 U12146 ( .A(n13545), .ZN(n10912) );
  NAND2_X1 U12147 ( .A1(n11689), .A2(n6544), .ZN(n9634) );
  OAI21_X1 U12148 ( .B1(n10912), .B2(n6544), .A(n9634), .ZN(n9635) );
  NAND2_X1 U12149 ( .A1(n15146), .A2(n6544), .ZN(n9637) );
  NAND2_X1 U12150 ( .A1(n13544), .A2(n9656), .ZN(n9636) );
  NAND2_X1 U12151 ( .A1(n9637), .A2(n9636), .ZN(n9640) );
  AOI22_X1 U12152 ( .A1(n15146), .A2(n9656), .B1(n6544), .B2(n13544), .ZN(
        n9638) );
  INV_X1 U12153 ( .A(n9638), .ZN(n9639) );
  NAND2_X1 U12154 ( .A1(n11712), .A2(n9656), .ZN(n9643) );
  NAND2_X1 U12155 ( .A1(n6544), .A2(n13543), .ZN(n9642) );
  AOI22_X1 U12156 ( .A1(n11712), .A2(n6544), .B1(n13543), .B2(n9656), .ZN(
        n9644) );
  NAND2_X1 U12157 ( .A1(n11443), .A2(n6544), .ZN(n9646) );
  NAND2_X1 U12158 ( .A1(n13542), .A2(n9656), .ZN(n9645) );
  NAND2_X1 U12159 ( .A1(n9646), .A2(n9645), .ZN(n9651) );
  INV_X1 U12160 ( .A(n13542), .ZN(n9851) );
  NAND2_X1 U12161 ( .A1(n11443), .A2(n9656), .ZN(n9647) );
  OAI21_X1 U12162 ( .B1(n9851), .B2(n6542), .A(n9647), .ZN(n9648) );
  NAND2_X1 U12163 ( .A1(n9649), .A2(n9648), .ZN(n9655) );
  NAND2_X1 U12164 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  NAND2_X1 U12165 ( .A1(n15232), .A2(n9656), .ZN(n9658) );
  NAND2_X1 U12166 ( .A1(n6544), .A2(n13541), .ZN(n9657) );
  AOI22_X1 U12167 ( .A1(n15232), .A2(n6544), .B1(n13541), .B2(n9656), .ZN(
        n9659) );
  NAND2_X1 U12168 ( .A1(n11887), .A2(n6544), .ZN(n9661) );
  NAND2_X1 U12169 ( .A1(n13540), .A2(n9656), .ZN(n9660) );
  NAND2_X1 U12170 ( .A1(n9661), .A2(n9660), .ZN(n9666) );
  INV_X1 U12171 ( .A(n13540), .ZN(n9854) );
  NAND2_X1 U12172 ( .A1(n11887), .A2(n9656), .ZN(n9662) );
  OAI21_X1 U12173 ( .B1(n9854), .B2(n6542), .A(n9662), .ZN(n9663) );
  NAND2_X1 U12174 ( .A1(n9664), .A2(n9663), .ZN(n9670) );
  INV_X1 U12175 ( .A(n9665), .ZN(n9668) );
  INV_X1 U12176 ( .A(n9666), .ZN(n9667) );
  NAND2_X1 U12177 ( .A1(n9668), .A2(n9667), .ZN(n9669) );
  NAND2_X1 U12178 ( .A1(n9670), .A2(n9669), .ZN(n9675) );
  NAND2_X1 U12179 ( .A1(n11855), .A2(n6542), .ZN(n9672) );
  NAND2_X1 U12180 ( .A1(n6544), .A2(n13539), .ZN(n9671) );
  NAND2_X1 U12181 ( .A1(n9672), .A2(n9671), .ZN(n9674) );
  AOI22_X1 U12182 ( .A1(n11855), .A2(n6544), .B1(n13539), .B2(n6542), .ZN(
        n9673) );
  AOI21_X1 U12183 ( .B1(n9675), .B2(n9674), .A(n9673), .ZN(n9677) );
  NOR2_X1 U12184 ( .A1(n9675), .A2(n9674), .ZN(n9676) );
  NAND2_X1 U12185 ( .A1(n14782), .A2(n6544), .ZN(n9679) );
  NAND2_X1 U12186 ( .A1(n13538), .A2(n6542), .ZN(n9678) );
  INV_X1 U12187 ( .A(n13538), .ZN(n11919) );
  NAND2_X1 U12188 ( .A1(n14782), .A2(n6542), .ZN(n9680) );
  OAI21_X1 U12189 ( .B1(n11919), .B2(n6542), .A(n9680), .ZN(n9681) );
  NAND2_X1 U12190 ( .A1(n11926), .A2(n6542), .ZN(n9683) );
  NAND2_X1 U12191 ( .A1(n6544), .A2(n13537), .ZN(n9682) );
  NAND2_X1 U12192 ( .A1(n9683), .A2(n9682), .ZN(n9686) );
  AOI22_X1 U12193 ( .A1(n11926), .A2(n6544), .B1(n13537), .B2(n6542), .ZN(
        n9684) );
  INV_X1 U12194 ( .A(n9684), .ZN(n9685) );
  NAND2_X1 U12195 ( .A1(n12109), .A2(n6544), .ZN(n9688) );
  NAND2_X1 U12196 ( .A1(n13536), .A2(n6542), .ZN(n9687) );
  NAND2_X1 U12197 ( .A1(n9688), .A2(n9687), .ZN(n9690) );
  AOI22_X1 U12198 ( .A1(n12109), .A2(n6542), .B1(n6544), .B2(n13536), .ZN(
        n9689) );
  NAND2_X1 U12199 ( .A1(n13869), .A2(n6542), .ZN(n9693) );
  NAND2_X1 U12200 ( .A1(n13535), .A2(n6544), .ZN(n9692) );
  NAND2_X1 U12201 ( .A1(n9693), .A2(n9692), .ZN(n9696) );
  NAND2_X1 U12202 ( .A1(n13869), .A2(n6544), .ZN(n9695) );
  NAND2_X1 U12203 ( .A1(n13535), .A2(n6542), .ZN(n9694) );
  NAND2_X1 U12204 ( .A1(n12340), .A2(n6544), .ZN(n9698) );
  NAND2_X1 U12205 ( .A1(n13534), .A2(n6542), .ZN(n9697) );
  NAND2_X1 U12206 ( .A1(n9698), .A2(n9697), .ZN(n9700) );
  INV_X1 U12207 ( .A(n9700), .ZN(n9699) );
  AOI22_X1 U12208 ( .A1(n12340), .A2(n6542), .B1(n6544), .B2(n13534), .ZN(
        n9702) );
  NAND2_X1 U12209 ( .A1(n13857), .A2(n6542), .ZN(n9705) );
  NAND2_X1 U12210 ( .A1(n13533), .A2(n6544), .ZN(n9704) );
  NAND2_X1 U12211 ( .A1(n9705), .A2(n9704), .ZN(n9708) );
  INV_X1 U12212 ( .A(n13533), .ZN(n9867) );
  NAND2_X1 U12213 ( .A1(n13857), .A2(n6544), .ZN(n9706) );
  OAI21_X1 U12214 ( .B1(n9867), .B2(n6544), .A(n9706), .ZN(n9707) );
  NAND2_X1 U12215 ( .A1(n13853), .A2(n6544), .ZN(n9711) );
  NAND2_X1 U12216 ( .A1(n13532), .A2(n9656), .ZN(n9710) );
  NAND2_X1 U12217 ( .A1(n9711), .A2(n9710), .ZN(n9713) );
  AOI22_X1 U12218 ( .A1(n13853), .A2(n6542), .B1(n6544), .B2(n13532), .ZN(
        n9712) );
  NAND2_X1 U12219 ( .A1(n13757), .A2(n6542), .ZN(n9717) );
  NAND2_X1 U12220 ( .A1(n13531), .A2(n6544), .ZN(n9716) );
  INV_X1 U12221 ( .A(n13531), .ZN(n13451) );
  NAND2_X1 U12222 ( .A1(n13757), .A2(n6544), .ZN(n9718) );
  OAI21_X1 U12223 ( .B1(n13451), .B2(n6544), .A(n9718), .ZN(n9719) );
  NAND2_X1 U12224 ( .A1(n13744), .A2(n6544), .ZN(n9721) );
  NAND2_X1 U12225 ( .A1(n13530), .A2(n6542), .ZN(n9720) );
  NAND2_X1 U12226 ( .A1(n9721), .A2(n9720), .ZN(n9724) );
  AOI22_X1 U12227 ( .A1(n13744), .A2(n6542), .B1(n6544), .B2(n13530), .ZN(
        n9722) );
  AOI21_X1 U12228 ( .B1(n9725), .B2(n9724), .A(n9722), .ZN(n9723) );
  NAND2_X1 U12229 ( .A1(n13836), .A2(n9656), .ZN(n9727) );
  NAND2_X1 U12230 ( .A1(n6544), .A2(n13529), .ZN(n9726) );
  AOI22_X1 U12231 ( .A1(n13836), .A2(n6544), .B1(n13529), .B2(n6542), .ZN(
        n9728) );
  AOI22_X1 U12232 ( .A1(n13713), .A2(n6544), .B1(n13528), .B2(n6542), .ZN(
        n9731) );
  AOI22_X1 U12233 ( .A1(n13713), .A2(n6542), .B1(n6544), .B2(n13528), .ZN(
        n9730) );
  INV_X1 U12234 ( .A(n9731), .ZN(n9733) );
  OAI22_X1 U12235 ( .A1(n13891), .A2(n6542), .B1(n9732), .B2(n6544), .ZN(n9738) );
  AOI22_X1 U12236 ( .A1(n13703), .A2(n6542), .B1(n6544), .B2(n13527), .ZN(
        n9739) );
  OAI22_X1 U12237 ( .A1(n9734), .A2(n9733), .B1(n9738), .B2(n9739), .ZN(n9741)
         );
  AND2_X1 U12238 ( .A1(n6544), .A2(n13526), .ZN(n9735) );
  AOI21_X1 U12239 ( .B1(n13682), .B2(n6542), .A(n9735), .ZN(n9763) );
  NAND2_X1 U12240 ( .A1(n13682), .A2(n6544), .ZN(n9737) );
  NAND2_X1 U12241 ( .A1(n13526), .A2(n6542), .ZN(n9736) );
  NAND2_X1 U12242 ( .A1(n9737), .A2(n9736), .ZN(n9762) );
  AOI22_X1 U12243 ( .A1(n9763), .A2(n9762), .B1(n9739), .B2(n9738), .ZN(n9740)
         );
  NAND2_X1 U12244 ( .A1(n9742), .A2(n9767), .ZN(n9744) );
  NAND2_X1 U12245 ( .A1(n8333), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U12246 ( .A1(n6545), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U12247 ( .A1(n9745), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U12248 ( .A1(n9746), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9747) );
  AND3_X1 U12249 ( .A1(n9749), .A2(n9748), .A3(n9747), .ZN(n9800) );
  AND2_X1 U12250 ( .A1(n6544), .A2(n13523), .ZN(n9750) );
  AOI21_X1 U12251 ( .B1(n13643), .B2(n6542), .A(n9750), .ZN(n9783) );
  NAND2_X1 U12252 ( .A1(n13643), .A2(n6544), .ZN(n9752) );
  NAND2_X1 U12253 ( .A1(n13523), .A2(n6542), .ZN(n9751) );
  NAND2_X1 U12254 ( .A1(n9752), .A2(n9751), .ZN(n9781) );
  NAND2_X1 U12255 ( .A1(n12332), .A2(n9767), .ZN(n9754) );
  NAND2_X1 U12256 ( .A1(n8333), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9753) );
  AND2_X1 U12257 ( .A1(n13522), .A2(n6542), .ZN(n9755) );
  AOI21_X1 U12258 ( .B1(n9954), .B2(n6544), .A(n9755), .ZN(n9777) );
  NAND2_X1 U12259 ( .A1(n9954), .A2(n9656), .ZN(n9757) );
  NAND2_X1 U12260 ( .A1(n6544), .A2(n13522), .ZN(n9756) );
  NAND2_X1 U12261 ( .A1(n9757), .A2(n9756), .ZN(n9776) );
  NAND2_X1 U12262 ( .A1(n9777), .A2(n9776), .ZN(n9782) );
  AND2_X1 U12263 ( .A1(n13524), .A2(n9656), .ZN(n9758) );
  AOI21_X1 U12264 ( .B1(n13809), .B2(n6544), .A(n9758), .ZN(n9789) );
  NAND2_X1 U12265 ( .A1(n13809), .A2(n6542), .ZN(n9760) );
  NAND2_X1 U12266 ( .A1(n6544), .A2(n13524), .ZN(n9759) );
  NAND2_X1 U12267 ( .A1(n9760), .A2(n9759), .ZN(n9788) );
  AND2_X1 U12268 ( .A1(n9789), .A2(n9788), .ZN(n9761) );
  OAI22_X1 U12269 ( .A1(n13668), .A2(n6542), .B1(n9936), .B2(n6544), .ZN(n9792) );
  INV_X1 U12270 ( .A(n9936), .ZN(n13525) );
  AOI22_X1 U12271 ( .A1(n13815), .A2(n6542), .B1(n6544), .B2(n13525), .ZN(
        n9793) );
  OAI22_X1 U12272 ( .A1(n9792), .A2(n9793), .B1(n9763), .B2(n9762), .ZN(n9764)
         );
  INV_X1 U12273 ( .A(n9800), .ZN(n13614) );
  AOI21_X1 U12274 ( .B1(n6544), .B2(n13614), .A(n9766), .ZN(n9786) );
  NAND2_X1 U12275 ( .A1(n13912), .A2(n9767), .ZN(n9769) );
  NAND2_X1 U12276 ( .A1(n8333), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9768) );
  NAND2_X1 U12277 ( .A1(n6545), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U12278 ( .A1(n6910), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U12279 ( .A1(n9746), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9770) );
  AND3_X1 U12280 ( .A1(n9772), .A2(n9771), .A3(n9770), .ZN(n9893) );
  OAI211_X1 U12281 ( .C1(n9586), .C2(n9832), .A(n8271), .B(n9773), .ZN(n9774)
         );
  AOI21_X1 U12282 ( .B1(n6542), .B2(n13614), .A(n9774), .ZN(n9775) );
  OAI22_X1 U12283 ( .A1(n13880), .A2(n6542), .B1(n9893), .B2(n9775), .ZN(n9797) );
  INV_X1 U12284 ( .A(n13880), .ZN(n9825) );
  AOI22_X1 U12285 ( .A1(n9825), .A2(n6542), .B1(n6544), .B2(n9894), .ZN(n9796)
         );
  INV_X1 U12286 ( .A(n9776), .ZN(n9779) );
  INV_X1 U12287 ( .A(n9777), .ZN(n9778) );
  AOI22_X1 U12288 ( .A1(n9797), .A2(n9796), .B1(n9779), .B2(n9778), .ZN(n9785)
         );
  INV_X1 U12289 ( .A(n9780), .ZN(n9828) );
  NAND4_X1 U12290 ( .A1(n9828), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(n9784)
         );
  OAI21_X1 U12291 ( .B1(n9786), .B2(n9785), .A(n9784), .ZN(n9787) );
  NAND3_X1 U12292 ( .A1(n13612), .A2(n9798), .A3(n13614), .ZN(n9802) );
  NAND3_X1 U12293 ( .A1(n13611), .A2(n9800), .A3(n6542), .ZN(n9801) );
  NOR2_X1 U12294 ( .A1(n9811), .A2(n9804), .ZN(n9805) );
  AOI211_X1 U12295 ( .C1(n8271), .C2(n13607), .A(n9809), .B(n9805), .ZN(n9806)
         );
  INV_X1 U12296 ( .A(n10531), .ZN(n10529) );
  NAND2_X1 U12297 ( .A1(n10529), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12067) );
  INV_X1 U12298 ( .A(n12067), .ZN(n9808) );
  AND2_X1 U12299 ( .A1(n9811), .A2(n13700), .ZN(n9891) );
  AND2_X1 U12300 ( .A1(n8271), .A2(n9832), .ZN(n9890) );
  AOI22_X1 U12301 ( .A1(n9891), .A2(n11766), .B1(n9890), .B2(n13700), .ZN(
        n9807) );
  INV_X1 U12302 ( .A(n13926), .ZN(n10538) );
  NAND4_X1 U12303 ( .A1(n15187), .A2(n10538), .A3(n9809), .A4(n13509), .ZN(
        n9810) );
  OAI211_X1 U12304 ( .C1(n9811), .C2(n12067), .A(n9810), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9835) );
  NAND2_X1 U12305 ( .A1(n13643), .A2(n13523), .ZN(n9939) );
  OR2_X1 U12306 ( .A1(n13643), .A2(n13523), .ZN(n9812) );
  INV_X1 U12307 ( .A(n13524), .ZN(n9888) );
  XNOR2_X1 U12308 ( .A(n13809), .B(n9888), .ZN(n13656) );
  INV_X1 U12309 ( .A(n13526), .ZN(n13467) );
  XNOR2_X1 U12310 ( .A(n13682), .B(n13467), .ZN(n9883) );
  OR2_X1 U12311 ( .A1(n13815), .A2(n9936), .ZN(n9885) );
  NAND2_X1 U12312 ( .A1(n13815), .A2(n9936), .ZN(n9886) );
  INV_X1 U12313 ( .A(n13529), .ZN(n13450) );
  XNOR2_X1 U12314 ( .A(n13836), .B(n13450), .ZN(n13730) );
  INV_X1 U12315 ( .A(n13530), .ZN(n9876) );
  XNOR2_X1 U12316 ( .A(n13744), .B(n9876), .ZN(n13737) );
  XOR2_X1 U12317 ( .A(n13532), .B(n13853), .Z(n13766) );
  OR2_X1 U12318 ( .A1(n13757), .A2(n13451), .ZN(n9874) );
  NAND2_X1 U12319 ( .A1(n13757), .A2(n13451), .ZN(n9873) );
  XOR2_X1 U12320 ( .A(n13537), .B(n11926), .Z(n11922) );
  INV_X1 U12321 ( .A(n13534), .ZN(n9865) );
  XNOR2_X1 U12322 ( .A(n12340), .B(n9865), .ZN(n12192) );
  XNOR2_X1 U12323 ( .A(n13869), .B(n13535), .ZN(n12142) );
  INV_X1 U12324 ( .A(n13539), .ZN(n9813) );
  NAND2_X1 U12325 ( .A1(n11855), .A2(n9813), .ZN(n9814) );
  NAND2_X1 U12326 ( .A1(n9857), .A2(n9814), .ZN(n11847) );
  INV_X1 U12327 ( .A(n13541), .ZN(n11477) );
  XNOR2_X1 U12328 ( .A(n11712), .B(n13543), .ZN(n11160) );
  INV_X1 U12329 ( .A(n13546), .ZN(n9845) );
  XNOR2_X1 U12330 ( .A(n11274), .B(n9845), .ZN(n11267) );
  OAI21_X1 U12331 ( .B1(n9589), .B2(n15166), .A(n10953), .ZN(n11471) );
  NOR4_X1 U12332 ( .A1(n11267), .A2(n9905), .A3(n6879), .A4(n9815), .ZN(n9816)
         );
  XNOR2_X1 U12333 ( .A(n15146), .B(n13544), .ZN(n11087) );
  XNOR2_X1 U12334 ( .A(n11689), .B(n13545), .ZN(n10924) );
  NAND4_X1 U12335 ( .A1(n11160), .A2(n9816), .A3(n11087), .A4(n10924), .ZN(
        n9817) );
  NOR4_X1 U12336 ( .A1(n11847), .A2(n11347), .A3(n11491), .A4(n9817), .ZN(
        n9818) );
  XNOR2_X1 U12337 ( .A(n14782), .B(n13538), .ZN(n12021) );
  XNOR2_X1 U12338 ( .A(n11887), .B(n13540), .ZN(n11790) );
  NAND4_X1 U12339 ( .A1(n12142), .A2(n9818), .A3(n12021), .A4(n11790), .ZN(
        n9819) );
  NOR3_X1 U12340 ( .A1(n11922), .A2(n12192), .A3(n9819), .ZN(n9820) );
  XNOR2_X1 U12341 ( .A(n13857), .B(n13533), .ZN(n13792) );
  XNOR2_X1 U12342 ( .A(n12109), .B(n13536), .ZN(n12092) );
  NAND4_X1 U12343 ( .A1(n13754), .A2(n9820), .A3(n13792), .A4(n12092), .ZN(
        n9821) );
  NOR4_X1 U12344 ( .A1(n13730), .A2(n13737), .A3(n13766), .A4(n9821), .ZN(
        n9823) );
  NAND2_X1 U12345 ( .A1(n13703), .A2(n13527), .ZN(n9935) );
  OR2_X1 U12346 ( .A1(n6984), .A2(n13527), .ZN(n9822) );
  NAND2_X1 U12347 ( .A1(n9935), .A2(n9822), .ZN(n13693) );
  XNOR2_X1 U12348 ( .A(n13713), .B(n13528), .ZN(n13710) );
  NAND4_X1 U12349 ( .A1(n13669), .A2(n9823), .A3(n13693), .A4(n13710), .ZN(
        n9824) );
  NOR4_X1 U12350 ( .A1(n13629), .A2(n13656), .A3(n9883), .A4(n9824), .ZN(n9827) );
  XNOR2_X1 U12351 ( .A(n9825), .B(n9894), .ZN(n9826) );
  XNOR2_X1 U12352 ( .A(n9954), .B(n13522), .ZN(n9940) );
  NAND4_X1 U12353 ( .A1(n9828), .A2(n9827), .A3(n9826), .A4(n9940), .ZN(n9829)
         );
  XOR2_X1 U12354 ( .A(n13700), .B(n9829), .Z(n9830) );
  NOR3_X1 U12355 ( .A1(n9830), .A2(n8271), .A3(n12067), .ZN(n9831) );
  OAI21_X1 U12356 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n9834) );
  INV_X1 U12357 ( .A(n13551), .ZN(n10896) );
  NAND2_X1 U12358 ( .A1(n10896), .A2(n15171), .ZN(n9836) );
  NAND2_X1 U12359 ( .A1(n11673), .A2(n11672), .ZN(n9839) );
  INV_X1 U12360 ( .A(n13549), .ZN(n9900) );
  NAND2_X1 U12361 ( .A1(n9900), .A2(n15199), .ZN(n9838) );
  INV_X1 U12362 ( .A(n11569), .ZN(n9840) );
  NAND2_X1 U12363 ( .A1(n11565), .A2(n9840), .ZN(n9842) );
  NAND2_X1 U12364 ( .A1(n10897), .A2(n11574), .ZN(n9841) );
  INV_X1 U12365 ( .A(n9905), .ZN(n11260) );
  NAND2_X1 U12366 ( .A1(n11261), .A2(n11260), .ZN(n9844) );
  NAND2_X1 U12367 ( .A1(n11259), .A2(n10913), .ZN(n9843) );
  NAND2_X1 U12368 ( .A1(n9844), .A2(n9843), .ZN(n11268) );
  AND2_X1 U12369 ( .A1(n11274), .A2(n9845), .ZN(n9847) );
  INV_X1 U12370 ( .A(n11274), .ZN(n15227) );
  NAND2_X1 U12371 ( .A1(n15227), .A2(n13546), .ZN(n9846) );
  INV_X1 U12372 ( .A(n10924), .ZN(n10930) );
  OR2_X2 U12373 ( .A1(n10929), .A2(n10930), .ZN(n10927) );
  NAND2_X1 U12374 ( .A1(n11689), .A2(n10912), .ZN(n9848) );
  INV_X1 U12375 ( .A(n13544), .ZN(n11067) );
  INV_X1 U12376 ( .A(n13543), .ZN(n9849) );
  OR2_X1 U12377 ( .A1(n11443), .A2(n9851), .ZN(n9852) );
  INV_X1 U12378 ( .A(n11790), .ZN(n11787) );
  NAND2_X1 U12379 ( .A1(n11887), .A2(n9854), .ZN(n9855) );
  NAND2_X1 U12380 ( .A1(n12022), .A2(n12021), .ZN(n12020) );
  OR2_X1 U12381 ( .A1(n14782), .A2(n11919), .ZN(n9858) );
  NAND2_X1 U12382 ( .A1(n11918), .A2(n14776), .ZN(n9859) );
  NAND2_X1 U12383 ( .A1(n9860), .A2(n9859), .ZN(n12093) );
  NAND2_X1 U12384 ( .A1(n12093), .A2(n12092), .ZN(n9862) );
  OR2_X1 U12385 ( .A1(n12109), .A2(n12107), .ZN(n9861) );
  NAND2_X1 U12386 ( .A1(n9862), .A2(n9861), .ZN(n12131) );
  INV_X1 U12387 ( .A(n13535), .ZN(n12343) );
  OR2_X1 U12388 ( .A1(n13869), .A2(n12343), .ZN(n9863) );
  NOR2_X1 U12389 ( .A1(n12340), .A2(n9865), .ZN(n9864) );
  NAND2_X1 U12390 ( .A1(n12340), .A2(n9865), .ZN(n9866) );
  AND2_X1 U12391 ( .A1(n13857), .A2(n9867), .ZN(n9868) );
  INV_X1 U12392 ( .A(n13532), .ZN(n9870) );
  NOR2_X1 U12393 ( .A1(n13853), .A2(n9870), .ZN(n9869) );
  NAND2_X1 U12394 ( .A1(n13853), .A2(n9870), .ZN(n9871) );
  INV_X1 U12395 ( .A(n9873), .ZN(n13736) );
  NAND2_X1 U12396 ( .A1(n13744), .A2(n9876), .ZN(n9875) );
  INV_X1 U12397 ( .A(n13730), .ZN(n9877) );
  NAND2_X1 U12398 ( .A1(n13720), .A2(n9877), .ZN(n9879) );
  OR2_X1 U12399 ( .A1(n13836), .A2(n13450), .ZN(n9878) );
  NAND2_X1 U12400 ( .A1(n9879), .A2(n9878), .ZN(n13707) );
  INV_X1 U12401 ( .A(n13528), .ZN(n13470) );
  OR2_X1 U12402 ( .A1(n13713), .A2(n13470), .ZN(n9880) );
  OR2_X1 U12403 ( .A1(n13891), .A2(n13527), .ZN(n9882) );
  NAND2_X1 U12404 ( .A1(n13682), .A2(n13467), .ZN(n9884) );
  NAND2_X1 U12405 ( .A1(n13676), .A2(n9884), .ZN(n13660) );
  NAND2_X1 U12406 ( .A1(n13660), .A2(n9885), .ZN(n9887) );
  NAND2_X1 U12407 ( .A1(n9887), .A2(n9886), .ZN(n13647) );
  INV_X1 U12408 ( .A(n13656), .ZN(n13646) );
  AND2_X1 U12409 ( .A1(n13809), .A2(n9888), .ZN(n9889) );
  INV_X1 U12410 ( .A(n13629), .ZN(n13633) );
  INV_X1 U12411 ( .A(n13509), .ZN(n13469) );
  OR2_X1 U12412 ( .A1(n7373), .A2(n13469), .ZN(n9896) );
  NAND2_X1 U12413 ( .A1(n10538), .A2(P2_B_REG_SCAN_IN), .ZN(n9892) );
  NAND2_X1 U12414 ( .A1(n7632), .A2(n9894), .ZN(n9895) );
  AND2_X1 U12415 ( .A1(n9896), .A2(n9895), .ZN(n9897) );
  INV_X1 U12416 ( .A(n10953), .ZN(n15167) );
  NAND2_X1 U12417 ( .A1(n10896), .A2(n15192), .ZN(n9898) );
  NAND2_X1 U12418 ( .A1(n9900), .A2(n11684), .ZN(n9901) );
  NAND2_X1 U12419 ( .A1(n9902), .A2(n9901), .ZN(n11570) );
  NAND2_X1 U12420 ( .A1(n11570), .A2(n6879), .ZN(n9904) );
  NAND2_X1 U12421 ( .A1(n15209), .A2(n10897), .ZN(n9903) );
  NAND2_X1 U12422 ( .A1(n9904), .A2(n9903), .ZN(n11252) );
  NAND2_X1 U12423 ( .A1(n11252), .A2(n9905), .ZN(n9907) );
  INV_X1 U12424 ( .A(n11259), .ZN(n15217) );
  NAND2_X1 U12425 ( .A1(n15217), .A2(n10913), .ZN(n9906) );
  NAND2_X1 U12426 ( .A1(n9907), .A2(n9906), .ZN(n11266) );
  NOR2_X1 U12427 ( .A1(n11274), .A2(n13546), .ZN(n9909) );
  NAND2_X1 U12428 ( .A1(n11274), .A2(n13546), .ZN(n9908) );
  INV_X1 U12429 ( .A(n11087), .ZN(n11084) );
  OR2_X1 U12430 ( .A1(n15146), .A2(n13544), .ZN(n9910) );
  NAND2_X1 U12431 ( .A1(n11712), .A2(n13543), .ZN(n9911) );
  NAND2_X1 U12432 ( .A1(n11158), .A2(n9911), .ZN(n11346) );
  NAND2_X1 U12433 ( .A1(n11346), .A2(n11347), .ZN(n9913) );
  NAND2_X1 U12434 ( .A1(n11443), .A2(n13542), .ZN(n9912) );
  NAND2_X1 U12435 ( .A1(n9913), .A2(n9912), .ZN(n11490) );
  NAND2_X1 U12436 ( .A1(n11490), .A2(n11491), .ZN(n9915) );
  NAND2_X1 U12437 ( .A1(n15232), .A2(n13541), .ZN(n9914) );
  AND2_X1 U12438 ( .A1(n11887), .A2(n13540), .ZN(n9916) );
  OR2_X1 U12439 ( .A1(n11887), .A2(n13540), .ZN(n9917) );
  NOR2_X1 U12440 ( .A1(n11855), .A2(n13539), .ZN(n9918) );
  OR2_X1 U12441 ( .A1(n14782), .A2(n13538), .ZN(n9920) );
  AND2_X1 U12442 ( .A1(n14782), .A2(n13538), .ZN(n9919) );
  AOI21_X1 U12443 ( .B1(n12013), .B2(n9920), .A(n9919), .ZN(n11921) );
  NAND2_X1 U12444 ( .A1(n11926), .A2(n13537), .ZN(n9922) );
  NOR2_X1 U12445 ( .A1(n11926), .A2(n13537), .ZN(n9921) );
  INV_X1 U12446 ( .A(n12091), .ZN(n9924) );
  OR2_X1 U12447 ( .A1(n12109), .A2(n13536), .ZN(n9925) );
  NAND2_X1 U12448 ( .A1(n13869), .A2(n13535), .ZN(n9926) );
  NAND2_X1 U12449 ( .A1(n12189), .A2(n12192), .ZN(n12191) );
  NAND2_X1 U12450 ( .A1(n12340), .A2(n13534), .ZN(n9927) );
  OR2_X1 U12451 ( .A1(n13857), .A2(n13533), .ZN(n9928) );
  NAND2_X1 U12452 ( .A1(n13853), .A2(n13532), .ZN(n9929) );
  OR2_X1 U12453 ( .A1(n13757), .A2(n13531), .ZN(n9930) );
  NAND2_X1 U12454 ( .A1(n13755), .A2(n9930), .ZN(n9932) );
  NAND2_X1 U12455 ( .A1(n13757), .A2(n13531), .ZN(n9931) );
  NAND2_X1 U12456 ( .A1(n13836), .A2(n13529), .ZN(n9933) );
  NAND2_X1 U12457 ( .A1(n13729), .A2(n9933), .ZN(n13711) );
  AND2_X1 U12458 ( .A1(n13713), .A2(n13528), .ZN(n9934) );
  INV_X1 U12459 ( .A(n13671), .ZN(n9937) );
  NAND2_X1 U12460 ( .A1(n13809), .A2(n13524), .ZN(n9938) );
  NAND2_X1 U12461 ( .A1(n13632), .A2(n9939), .ZN(n9941) );
  XNOR2_X1 U12462 ( .A(n9941), .B(n9940), .ZN(n13622) );
  AND2_X1 U12463 ( .A1(n11766), .A2(n13700), .ZN(n9943) );
  AND2_X1 U12464 ( .A1(n9586), .A2(n9943), .ZN(n15239) );
  INV_X1 U12465 ( .A(n15239), .ZN(n15223) );
  NAND2_X1 U12466 ( .A1(n9942), .A2(n15223), .ZN(n15212) );
  INV_X1 U12467 ( .A(n11855), .ZN(n14793) );
  INV_X1 U12468 ( .A(n11712), .ZN(n11168) );
  NAND2_X1 U12469 ( .A1(n15192), .A2(n9588), .ZN(n15164) );
  NAND2_X1 U12470 ( .A1(n11680), .A2(n15209), .ZN(n11571) );
  NOR2_X1 U12471 ( .A1(n11571), .A2(n11259), .ZN(n11255) );
  NAND2_X1 U12472 ( .A1(n15227), .A2(n11255), .ZN(n11271) );
  OR2_X1 U12473 ( .A1(n11689), .A2(n11271), .ZN(n11086) );
  NAND2_X1 U12474 ( .A1(n14793), .A2(n11853), .ZN(n12014) );
  INV_X1 U12475 ( .A(n12340), .ZN(n13864) );
  NOR2_X1 U12476 ( .A1(n13772), .A2(n13757), .ZN(n13756) );
  INV_X1 U12477 ( .A(n13744), .ZN(n13899) );
  AOI211_X1 U12478 ( .C1(n9954), .C2(n13638), .A(n11852), .B(n13618), .ZN(
        n13627) );
  INV_X1 U12479 ( .A(n9948), .ZN(n9949) );
  NAND2_X1 U12480 ( .A1(n15187), .A2(n9949), .ZN(n11249) );
  OR2_X1 U12481 ( .A1(n9950), .A2(n15183), .ZN(n9951) );
  NOR2_X1 U12482 ( .A1(n11249), .A2(n9951), .ZN(n9952) );
  NAND2_X1 U12483 ( .A1(n15250), .A2(n15200), .ZN(n13850) );
  INV_X1 U12484 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9955) );
  OR2_X1 U12485 ( .A1(n15250), .A2(n9955), .ZN(n9956) );
  INV_X1 U12486 ( .A(n9957), .ZN(n9958) );
  OAI21_X1 U12487 ( .B1(n10405), .B2(n9959), .A(n9958), .ZN(P2_U3528) );
  OR2_X1 U12488 ( .A1(n14137), .A2(n8985), .ZN(n9961) );
  NAND2_X1 U12489 ( .A1(n11321), .A2(n9963), .ZN(n9965) );
  INV_X1 U12490 ( .A(n14973), .ZN(n11333) );
  OR2_X1 U12491 ( .A1(n14136), .A2(n11333), .ZN(n9964) );
  OR2_X1 U12492 ( .A1(n14135), .A2(n14980), .ZN(n9967) );
  INV_X1 U12493 ( .A(n14935), .ZN(n14946) );
  OR2_X1 U12494 ( .A1(n10206), .A2(n14134), .ZN(n9968) );
  NAND2_X1 U12495 ( .A1(n9969), .A2(n9968), .ZN(n11384) );
  NAND2_X1 U12496 ( .A1(n11384), .A2(n7561), .ZN(n9971) );
  NAND2_X1 U12497 ( .A1(n14994), .A2(n11316), .ZN(n9970) );
  NAND2_X1 U12498 ( .A1(n9971), .A2(n9970), .ZN(n14914) );
  NAND2_X1 U12499 ( .A1(n14914), .A2(n14916), .ZN(n9973) );
  NAND2_X1 U12500 ( .A1(n14999), .A2(n10234), .ZN(n9972) );
  NAND2_X1 U12501 ( .A1(n9973), .A2(n9972), .ZN(n11506) );
  NAND2_X1 U12502 ( .A1(n11506), .A2(n7572), .ZN(n9975) );
  OR2_X1 U12503 ( .A1(n15006), .A2(n14130), .ZN(n9974) );
  NAND2_X1 U12504 ( .A1(n9975), .A2(n9974), .ZN(n11398) );
  NAND2_X1 U12505 ( .A1(n11398), .A2(n11399), .ZN(n9977) );
  OR2_X1 U12506 ( .A1(n11878), .A2(n14129), .ZN(n9976) );
  NAND2_X1 U12507 ( .A1(n9977), .A2(n9976), .ZN(n11524) );
  NAND2_X1 U12508 ( .A1(n11524), .A2(n10038), .ZN(n9979) );
  OR2_X1 U12509 ( .A1(n12010), .A2(n14128), .ZN(n9978) );
  NAND2_X1 U12510 ( .A1(n9979), .A2(n9978), .ZN(n11772) );
  OR2_X1 U12511 ( .A1(n15022), .A2(n14127), .ZN(n9980) );
  INV_X1 U12512 ( .A(n11993), .ZN(n11989) );
  NAND2_X1 U12513 ( .A1(n11988), .A2(n11989), .ZN(n9982) );
  OR2_X1 U12514 ( .A1(n14679), .A2(n14125), .ZN(n9981) );
  NAND2_X1 U12515 ( .A1(n11973), .A2(n11975), .ZN(n9984) );
  OR2_X1 U12516 ( .A1(n14827), .A2(n14124), .ZN(n9983) );
  NAND2_X1 U12517 ( .A1(n14820), .A2(n14123), .ZN(n9985) );
  INV_X1 U12518 ( .A(n12161), .ZN(n10292) );
  OR2_X1 U12519 ( .A1(n14104), .A2(n10292), .ZN(n9986) );
  NAND2_X1 U12520 ( .A1(n12167), .A2(n12166), .ZN(n9988) );
  OR2_X1 U12521 ( .A1(n14804), .A2(n14122), .ZN(n9987) );
  OR2_X1 U12522 ( .A1(n14502), .A2(n14120), .ZN(n9991) );
  NAND2_X1 U12523 ( .A1(n14385), .A2(n14389), .ZN(n9993) );
  OR2_X1 U12524 ( .A1(n14498), .A2(n14119), .ZN(n9992) );
  INV_X1 U12525 ( .A(n14373), .ZN(n9994) );
  NAND2_X1 U12526 ( .A1(n14492), .A2(n14118), .ZN(n9995) );
  INV_X1 U12527 ( .A(n14350), .ZN(n9996) );
  NAND2_X1 U12528 ( .A1(n14348), .A2(n13983), .ZN(n9997) );
  NAND2_X1 U12529 ( .A1(n14472), .A2(n14115), .ZN(n10000) );
  NAND2_X1 U12530 ( .A1(n14460), .A2(n14113), .ZN(n10001) );
  NAND2_X1 U12531 ( .A1(n14290), .A2(n10001), .ZN(n14276) );
  NAND2_X1 U12532 ( .A1(n14455), .A2(n14112), .ZN(n10002) );
  INV_X1 U12533 ( .A(n14235), .ZN(n14246) );
  NAND3_X1 U12534 ( .A1(n12180), .A2(P1_B_REG_SCAN_IN), .A3(n12604), .ZN(
        n10008) );
  INV_X1 U12535 ( .A(n12604), .ZN(n10006) );
  INV_X1 U12536 ( .A(P1_B_REG_SCAN_IN), .ZN(n10071) );
  AOI21_X1 U12537 ( .B1(n10006), .B2(n10071), .A(n12257), .ZN(n10007) );
  NAND2_X1 U12538 ( .A1(n12604), .A2(n12257), .ZN(n10506) );
  OAI21_X1 U12539 ( .B1(n10504), .B2(P1_D_REG_0__SCAN_IN), .A(n10506), .ZN(
        n10021) );
  NOR4_X1 U12540 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10012) );
  NOR4_X1 U12541 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10011) );
  NOR4_X1 U12542 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10010) );
  NOR4_X1 U12543 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10009) );
  AND4_X1 U12544 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10018) );
  NOR2_X1 U12545 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .ZN(
        n10016) );
  NOR4_X1 U12546 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n10015) );
  NOR4_X1 U12547 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10014) );
  NOR4_X1 U12548 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n10013) );
  AND4_X1 U12549 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n10017) );
  NAND2_X1 U12550 ( .A1(n10018), .A2(n10017), .ZN(n10385) );
  INV_X1 U12551 ( .A(n10385), .ZN(n10019) );
  OR2_X1 U12552 ( .A1(n10504), .A2(n10019), .ZN(n10020) );
  OR2_X1 U12553 ( .A1(n10504), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10022) );
  NAND2_X1 U12554 ( .A1(n12180), .A2(n12257), .ZN(n10509) );
  NAND2_X1 U12555 ( .A1(n10022), .A2(n10509), .ZN(n10686) );
  INV_X1 U12556 ( .A(n10686), .ZN(n10023) );
  NAND3_X1 U12557 ( .A1(n10687), .A2(n10781), .A3(n10023), .ZN(n10075) );
  NAND2_X1 U12558 ( .A1(n10413), .A2(n10511), .ZN(n10512) );
  INV_X1 U12559 ( .A(n10512), .ZN(n10505) );
  AND2_X4 U12560 ( .A1(n10069), .A2(n11764), .ZN(n14948) );
  INV_X1 U12561 ( .A(n10685), .ZN(n10025) );
  AND2_X2 U12562 ( .A1(n10075), .A2(n14940), .ZN(n14942) );
  OAI21_X1 U12563 ( .B1(n10026), .B2(n10180), .A(n12589), .ZN(n10680) );
  NAND2_X1 U12564 ( .A1(n10029), .A2(n10028), .ZN(n11323) );
  NAND2_X1 U12565 ( .A1(n11323), .A2(n11324), .ZN(n11322) );
  NAND2_X1 U12566 ( .A1(n11322), .A2(n10030), .ZN(n11370) );
  NAND2_X1 U12567 ( .A1(n11370), .A2(n11369), .ZN(n11368) );
  OR2_X1 U12568 ( .A1(n14135), .A2(n10066), .ZN(n10031) );
  NAND2_X1 U12569 ( .A1(n11368), .A2(n10031), .ZN(n14934) );
  NAND2_X1 U12570 ( .A1(n14934), .A2(n14935), .ZN(n10033) );
  INV_X1 U12571 ( .A(n14134), .ZN(n11372) );
  NAND2_X1 U12572 ( .A1(n11372), .A2(n10206), .ZN(n10032) );
  NAND2_X1 U12573 ( .A1(n14919), .A2(n10035), .ZN(n11509) );
  INV_X1 U12574 ( .A(n14130), .ZN(n10242) );
  NAND2_X1 U12575 ( .A1(n15006), .A2(n10242), .ZN(n10036) );
  NAND2_X1 U12576 ( .A1(n12010), .A2(n11769), .ZN(n10039) );
  INV_X1 U12577 ( .A(n11773), .ZN(n10040) );
  NAND2_X1 U12578 ( .A1(n11736), .A2(n10042), .ZN(n10044) );
  INV_X1 U12579 ( .A(n14126), .ZN(n12154) );
  OR2_X1 U12580 ( .A1(n11740), .A2(n12154), .ZN(n10043) );
  NAND2_X1 U12581 ( .A1(n10044), .A2(n10043), .ZN(n11992) );
  NAND2_X1 U12582 ( .A1(n11992), .A2(n11993), .ZN(n10046) );
  INV_X1 U12583 ( .A(n14125), .ZN(n11738) );
  OR2_X1 U12584 ( .A1(n14679), .A2(n11738), .ZN(n10045) );
  NAND2_X1 U12585 ( .A1(n10046), .A2(n10045), .ZN(n11974) );
  OR2_X1 U12586 ( .A1(n14827), .A2(n12081), .ZN(n10047) );
  NAND2_X1 U12587 ( .A1(n12120), .A2(n12121), .ZN(n10050) );
  NAND2_X1 U12588 ( .A1(n14804), .A2(n14011), .ZN(n10051) );
  NAND2_X1 U12589 ( .A1(n14404), .A2(n14402), .ZN(n10053) );
  NAND2_X1 U12590 ( .A1(n10053), .A2(n10052), .ZN(n14388) );
  INV_X1 U12591 ( .A(n14388), .ZN(n10055) );
  INV_X1 U12592 ( .A(n14389), .ZN(n10054) );
  OR2_X1 U12593 ( .A1(n14492), .A2(n13984), .ZN(n10057) );
  INV_X1 U12594 ( .A(n14117), .ZN(n14037) );
  NAND2_X1 U12595 ( .A1(n14338), .A2(n14350), .ZN(n10059) );
  OR2_X1 U12596 ( .A1(n14348), .A2(n14116), .ZN(n10058) );
  NAND2_X1 U12597 ( .A1(n10059), .A2(n10058), .ZN(n14322) );
  INV_X1 U12598 ( .A(n14115), .ZN(n10353) );
  NAND2_X1 U12599 ( .A1(n14472), .A2(n10353), .ZN(n10060) );
  NAND2_X1 U12600 ( .A1(n14321), .A2(n10060), .ZN(n14300) );
  INV_X1 U12601 ( .A(n14314), .ZN(n14469) );
  INV_X1 U12602 ( .A(n14460), .ZN(n14293) );
  INV_X1 U12603 ( .A(n14455), .ZN(n14094) );
  INV_X1 U12604 ( .A(n14450), .ZN(n14259) );
  NAND2_X1 U12605 ( .A1(n14249), .A2(n7627), .ZN(n14236) );
  INV_X1 U12606 ( .A(n14446), .ZN(n14243) );
  NAND2_X1 U12607 ( .A1(n14234), .A2(n7626), .ZN(n10063) );
  XNOR2_X1 U12608 ( .A(n10063), .B(n10062), .ZN(n10065) );
  INV_X1 U12609 ( .A(n14679), .ZN(n13999) );
  INV_X1 U12610 ( .A(n10206), .ZN(n14988) );
  NAND2_X1 U12611 ( .A1(n14951), .A2(n14994), .ZN(n14927) );
  INV_X1 U12612 ( .A(n11878), .ZN(n11548) );
  INV_X1 U12613 ( .A(n12010), .ZN(n15017) );
  INV_X1 U12614 ( .A(n14502), .ZN(n14409) );
  NOR2_X1 U12615 ( .A1(n14376), .A2(n14486), .ZN(n14360) );
  NAND2_X1 U12616 ( .A1(n14348), .A2(n14360), .ZN(n14342) );
  INV_X1 U12617 ( .A(n14239), .ZN(n10068) );
  INV_X1 U12618 ( .A(n14948), .ZN(n14829) );
  INV_X1 U12619 ( .A(n14441), .ZN(n10078) );
  AOI211_X1 U12620 ( .C1(n14441), .C2(n10068), .A(n14829), .B(n14228), .ZN(
        n14439) );
  INV_X1 U12621 ( .A(n10069), .ZN(n10683) );
  OR2_X1 U12622 ( .A1(n10683), .A2(n11764), .ZN(n14677) );
  INV_X1 U12623 ( .A(n10513), .ZN(n10070) );
  NOR2_X1 U12624 ( .A1(n14545), .A2(n10071), .ZN(n10072) );
  NOR2_X1 U12625 ( .A1(n14268), .A2(n10072), .ZN(n14223) );
  AND2_X1 U12626 ( .A1(n14108), .A2(n14223), .ZN(n14440) );
  INV_X1 U12627 ( .A(n14440), .ZN(n10074) );
  OAI22_X1 U12628 ( .A1(n10075), .A2(n10074), .B1(n10073), .B2(n14940), .ZN(
        n10076) );
  AOI21_X1 U12629 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14942), .A(n10076), 
        .ZN(n10077) );
  OAI21_X1 U12630 ( .B1(n10078), .B2(n14944), .A(n10077), .ZN(n10079) );
  AOI21_X1 U12631 ( .B1(n14439), .B2(n14953), .A(n10079), .ZN(n10080) );
  INV_X1 U12632 ( .A(n12400), .ZN(n10084) );
  NAND2_X1 U12633 ( .A1(n10084), .A2(n13409), .ZN(n10086) );
  OAI21_X1 U12634 ( .B1(n12414), .B2(n12889), .A(n11081), .ZN(n10085) );
  XNOR2_X1 U12635 ( .A(n13368), .B(n10865), .ZN(n12297) );
  NOR2_X1 U12636 ( .A1(n12297), .A2(n12921), .ZN(n12292) );
  AOI21_X1 U12637 ( .B1(n12297), .B2(n12921), .A(n12292), .ZN(n10153) );
  MUX2_X1 U12638 ( .A(n10087), .B(n8109), .S(n10097), .Z(n10869) );
  NAND2_X1 U12639 ( .A1(n10109), .A2(n11209), .ZN(n10089) );
  NAND2_X1 U12640 ( .A1(n10088), .A2(n10089), .ZN(n10090) );
  MUX2_X1 U12641 ( .A(n10091), .B(n8109), .S(n10097), .Z(n10092) );
  NAND2_X1 U12642 ( .A1(n10868), .A2(n10092), .ZN(n10874) );
  XNOR2_X1 U12643 ( .A(n10097), .B(n15391), .ZN(n10093) );
  XNOR2_X1 U12644 ( .A(n10093), .B(n6803), .ZN(n10875) );
  XNOR2_X1 U12645 ( .A(n10097), .B(n15373), .ZN(n10094) );
  XNOR2_X1 U12646 ( .A(n10094), .B(n12719), .ZN(n10978) );
  NAND2_X1 U12647 ( .A1(n10093), .A2(n11103), .ZN(n10976) );
  INV_X1 U12648 ( .A(n10094), .ZN(n10095) );
  NAND2_X1 U12649 ( .A1(n10095), .A2(n12719), .ZN(n10096) );
  XNOR2_X1 U12650 ( .A(n10097), .B(n15365), .ZN(n10098) );
  NAND2_X1 U12651 ( .A1(n10098), .A2(n11342), .ZN(n10101) );
  INV_X1 U12652 ( .A(n10098), .ZN(n10099) );
  NAND2_X1 U12653 ( .A1(n10099), .A2(n12718), .ZN(n10100) );
  NAND2_X1 U12654 ( .A1(n10101), .A2(n10100), .ZN(n11150) );
  NAND2_X1 U12655 ( .A1(n11148), .A2(n10101), .ZN(n11337) );
  XNOR2_X1 U12656 ( .A(n10097), .B(n15358), .ZN(n10102) );
  XNOR2_X1 U12657 ( .A(n10102), .B(n12717), .ZN(n11338) );
  NAND2_X1 U12658 ( .A1(n11337), .A2(n11338), .ZN(n11336) );
  NAND2_X1 U12659 ( .A1(n10102), .A2(n11454), .ZN(n10103) );
  XNOR2_X1 U12660 ( .A(n10097), .B(n11748), .ZN(n10104) );
  XNOR2_X1 U12661 ( .A(n10104), .B(n12716), .ZN(n11447) );
  NAND2_X1 U12662 ( .A1(n10104), .A2(n12716), .ZN(n10105) );
  XNOR2_X1 U12663 ( .A(n11700), .B(n10109), .ZN(n11552) );
  XNOR2_X1 U12664 ( .A(n10865), .B(n11554), .ZN(n10106) );
  NAND2_X1 U12665 ( .A1(n10106), .A2(n12715), .ZN(n10107) );
  NAND2_X1 U12666 ( .A1(n10108), .A2(n10107), .ZN(n11755) );
  INV_X2 U12667 ( .A(n10109), .ZN(n10865) );
  XNOR2_X1 U12668 ( .A(n10865), .B(n15347), .ZN(n10111) );
  XNOR2_X1 U12669 ( .A(n10111), .B(n10110), .ZN(n11754) );
  NAND2_X1 U12670 ( .A1(n11755), .A2(n11754), .ZN(n10113) );
  NAND2_X1 U12671 ( .A1(n10111), .A2(n15325), .ZN(n10112) );
  NAND2_X1 U12672 ( .A1(n10113), .A2(n10112), .ZN(n11910) );
  XNOR2_X1 U12673 ( .A(n10865), .B(n15330), .ZN(n10114) );
  XNOR2_X1 U12674 ( .A(n10114), .B(n15339), .ZN(n11911) );
  XNOR2_X1 U12675 ( .A(n10865), .B(n15314), .ZN(n10116) );
  XNOR2_X1 U12676 ( .A(n10116), .B(n15323), .ZN(n11937) );
  NAND2_X1 U12677 ( .A1(n10114), .A2(n15339), .ZN(n11934) );
  AND2_X1 U12678 ( .A1(n11937), .A2(n11934), .ZN(n10115) );
  INV_X1 U12679 ( .A(n10116), .ZN(n10117) );
  NAND2_X1 U12680 ( .A1(n10117), .A2(n15323), .ZN(n10118) );
  XNOR2_X1 U12681 ( .A(n10419), .B(n10865), .ZN(n10119) );
  XNOR2_X1 U12682 ( .A(n14730), .B(n10865), .ZN(n10120) );
  NOR2_X1 U12683 ( .A1(n10120), .A2(n14739), .ZN(n12237) );
  XNOR2_X1 U12684 ( .A(n12405), .B(n10865), .ZN(n10426) );
  NOR2_X1 U12685 ( .A1(n10426), .A2(n12407), .ZN(n10122) );
  INV_X1 U12686 ( .A(n10426), .ZN(n10121) );
  XNOR2_X1 U12687 ( .A(n12247), .B(n10865), .ZN(n10123) );
  XOR2_X1 U12688 ( .A(n12713), .B(n10123), .Z(n10436) );
  XNOR2_X1 U12689 ( .A(n13365), .B(n10865), .ZN(n10125) );
  XNOR2_X1 U12690 ( .A(n10125), .B(n12712), .ZN(n12268) );
  INV_X1 U12691 ( .A(n10125), .ZN(n10126) );
  XNOR2_X1 U12692 ( .A(n13358), .B(n10865), .ZN(n10127) );
  XNOR2_X1 U12693 ( .A(n10127), .B(n12711), .ZN(n12638) );
  INV_X1 U12694 ( .A(n10127), .ZN(n10128) );
  XNOR2_X1 U12695 ( .A(n13357), .B(n10865), .ZN(n10129) );
  XNOR2_X1 U12696 ( .A(n10129), .B(n13283), .ZN(n12648) );
  INV_X1 U12697 ( .A(n10129), .ZN(n10130) );
  XNOR2_X1 U12698 ( .A(n13350), .B(n10865), .ZN(n10131) );
  XNOR2_X1 U12699 ( .A(n10131), .B(n13010), .ZN(n12682) );
  INV_X1 U12700 ( .A(n10131), .ZN(n10132) );
  XNOR2_X1 U12701 ( .A(n13400), .B(n10865), .ZN(n10133) );
  XNOR2_X1 U12702 ( .A(n10133), .B(n12686), .ZN(n12612) );
  XNOR2_X1 U12703 ( .A(n13396), .B(n10865), .ZN(n10134) );
  XNOR2_X1 U12704 ( .A(n10134), .B(n13011), .ZN(n12667) );
  INV_X1 U12705 ( .A(n10134), .ZN(n10135) );
  AOI22_X1 U12706 ( .A1(n12666), .A2(n12667), .B1(n10135), .B2(n13011), .ZN(
        n12621) );
  XNOR2_X1 U12707 ( .A(n13393), .B(n10865), .ZN(n10136) );
  NOR2_X1 U12708 ( .A1(n10136), .A2(n12998), .ZN(n10137) );
  AOI21_X1 U12709 ( .B1(n10136), .B2(n12998), .A(n10137), .ZN(n12622) );
  NAND2_X1 U12710 ( .A1(n12621), .A2(n12622), .ZN(n12620) );
  INV_X1 U12711 ( .A(n10137), .ZN(n10138) );
  NAND2_X1 U12712 ( .A1(n12620), .A2(n10138), .ZN(n10140) );
  XNOR2_X1 U12713 ( .A(n12979), .B(n10865), .ZN(n10139) );
  NAND2_X1 U12714 ( .A1(n10140), .A2(n10139), .ZN(n10141) );
  OAI21_X1 U12715 ( .B1(n10140), .B2(n10139), .A(n10141), .ZN(n12675) );
  XNOR2_X1 U12716 ( .A(n13383), .B(n10865), .ZN(n10143) );
  XNOR2_X1 U12717 ( .A(n12655), .B(n10865), .ZN(n10142) );
  NAND2_X1 U12718 ( .A1(n10142), .A2(n12933), .ZN(n10145) );
  OAI21_X1 U12719 ( .B1(n10142), .B2(n12933), .A(n10145), .ZN(n12658) );
  INV_X1 U12720 ( .A(n10143), .ZN(n12605) );
  INV_X1 U12721 ( .A(n10145), .ZN(n12631) );
  XNOR2_X1 U12722 ( .A(n13375), .B(n10865), .ZN(n10146) );
  NAND2_X1 U12723 ( .A1(n10146), .A2(n12949), .ZN(n10149) );
  INV_X1 U12724 ( .A(n10146), .ZN(n10147) );
  NAND2_X1 U12725 ( .A1(n10147), .A2(n12920), .ZN(n10148) );
  OAI21_X1 U12726 ( .B1(n12660), .B2(n12631), .A(n12630), .ZN(n12629) );
  NAND2_X1 U12727 ( .A1(n12629), .A2(n10149), .ZN(n12694) );
  XNOR2_X1 U12728 ( .A(n13372), .B(n10865), .ZN(n10150) );
  NOR2_X1 U12729 ( .A1(n10150), .A2(n12708), .ZN(n10151) );
  AOI21_X1 U12730 ( .B1(n10150), .B2(n12708), .A(n10151), .ZN(n12695) );
  NAND2_X1 U12731 ( .A1(n12694), .A2(n12695), .ZN(n12693) );
  INV_X1 U12732 ( .A(n10151), .ZN(n10152) );
  INV_X1 U12733 ( .A(n10159), .ZN(n10169) );
  OR2_X1 U12734 ( .A1(n10154), .A2(n10169), .ZN(n10156) );
  NAND4_X1 U12735 ( .A1(n11219), .A2(n10157), .A3(n10162), .A4(n15346), .ZN(
        n10155) );
  INV_X1 U12736 ( .A(n10157), .ZN(n10161) );
  AOI21_X1 U12737 ( .B1(n10161), .B2(n12551), .A(n15346), .ZN(n10158) );
  OR2_X1 U12738 ( .A1(n12554), .A2(n10159), .ZN(n10168) );
  NAND2_X1 U12739 ( .A1(n10160), .A2(n10169), .ZN(n10165) );
  AND2_X1 U12740 ( .A1(n11023), .A2(n10414), .ZN(n10164) );
  NAND2_X1 U12741 ( .A1(n10162), .A2(n10161), .ZN(n10163) );
  NAND4_X1 U12742 ( .A1(n10165), .A2(n10164), .A3(n11216), .A4(n10163), .ZN(
        n10166) );
  NAND2_X1 U12743 ( .A1(n10166), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10167) );
  OR2_X1 U12744 ( .A1(n12554), .A2(n10169), .ZN(n10173) );
  INV_X1 U12745 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n10171) );
  OAI22_X1 U12746 ( .A1(n12934), .A2(n12296), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10171), .ZN(n10175) );
  NOR2_X1 U12747 ( .A1(n6543), .A2(n12685), .ZN(n10174) );
  AOI211_X1 U12748 ( .C1(n12906), .C2(n12689), .A(n10175), .B(n10174), .ZN(
        n10176) );
  INV_X1 U12749 ( .A(n10177), .ZN(n10178) );
  NAND2_X1 U12750 ( .A1(n10179), .A2(n10178), .ZN(P3_U3154) );
  AND2_X4 U12751 ( .A1(n10182), .A2(n10180), .ZN(n12588) );
  AOI22_X1 U12752 ( .A1(n10196), .A2(n14137), .B1(n10299), .B2(n8985), .ZN(
        n10195) );
  INV_X1 U12753 ( .A(n10195), .ZN(n10186) );
  NAND2_X1 U12754 ( .A1(n14137), .A2(n10299), .ZN(n10184) );
  NAND2_X1 U12755 ( .A1(n10184), .A2(n10183), .ZN(n10185) );
  NAND2_X1 U12756 ( .A1(n10196), .A2(n14138), .ZN(n10189) );
  INV_X1 U12757 ( .A(n10413), .ZN(n10187) );
  AOI22_X1 U12758 ( .A1(n10299), .A2(n11380), .B1(n10187), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10188) );
  NAND2_X1 U12759 ( .A1(n10189), .A2(n10188), .ZN(n10822) );
  NAND2_X1 U12760 ( .A1(n14138), .A2(n10299), .ZN(n10191) );
  NAND2_X1 U12761 ( .A1(n12588), .A2(n11380), .ZN(n10190) );
  OAI211_X1 U12762 ( .C1(n10192), .C2(n10413), .A(n10191), .B(n10190), .ZN(
        n10821) );
  INV_X1 U12763 ( .A(n10193), .ZN(n10194) );
  NOR2_X1 U12764 ( .A1(n10254), .A2(n14973), .ZN(n10197) );
  AOI21_X1 U12765 ( .B1(n10196), .B2(n14136), .A(n10197), .ZN(n10212) );
  NAND2_X1 U12766 ( .A1(n14136), .A2(n10299), .ZN(n10199) );
  NAND2_X1 U12767 ( .A1(n11333), .A2(n12588), .ZN(n10198) );
  NAND2_X1 U12768 ( .A1(n10199), .A2(n10198), .ZN(n10200) );
  XNOR2_X1 U12769 ( .A(n10200), .B(n12589), .ZN(n10211) );
  XOR2_X1 U12770 ( .A(n10212), .B(n10211), .Z(n10779) );
  NOR2_X1 U12771 ( .A1(n10777), .A2(n10779), .ZN(n10224) );
  NAND2_X1 U12772 ( .A1(n14135), .A2(n10299), .ZN(n10202) );
  NAND2_X1 U12773 ( .A1(n12588), .A2(n14980), .ZN(n10201) );
  NAND2_X1 U12774 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  NAND2_X1 U12775 ( .A1(n10196), .A2(n14135), .ZN(n10205) );
  NAND2_X1 U12776 ( .A1(n10299), .A2(n14980), .ZN(n10204) );
  NAND2_X1 U12777 ( .A1(n10205), .A2(n10204), .ZN(n10226) );
  NAND2_X1 U12778 ( .A1(n10225), .A2(n10226), .ZN(n10227) );
  NAND2_X1 U12779 ( .A1(n10196), .A2(n14134), .ZN(n10208) );
  NAND2_X1 U12780 ( .A1(n10206), .A2(n10299), .ZN(n10207) );
  AND2_X1 U12781 ( .A1(n10208), .A2(n10207), .ZN(n10217) );
  INV_X1 U12782 ( .A(n10217), .ZN(n10228) );
  NAND2_X1 U12783 ( .A1(n10227), .A2(n10228), .ZN(n10214) );
  INV_X1 U12784 ( .A(n10214), .ZN(n10220) );
  INV_X1 U12785 ( .A(n10226), .ZN(n10209) );
  AOI21_X1 U12786 ( .B1(n10209), .B2(n10228), .A(n10225), .ZN(n10216) );
  INV_X1 U12787 ( .A(n10225), .ZN(n10210) );
  AOI21_X1 U12788 ( .B1(n10217), .B2(n10226), .A(n10210), .ZN(n10215) );
  INV_X1 U12789 ( .A(n10211), .ZN(n10213) );
  NAND2_X1 U12790 ( .A1(n10213), .A2(n10212), .ZN(n10222) );
  OAI22_X1 U12791 ( .A1(n10216), .A2(n10215), .B1(n10214), .B2(n10222), .ZN(
        n10219) );
  OAI211_X1 U12792 ( .C1(n10225), .C2(n10226), .A(n10222), .B(n10217), .ZN(
        n10218) );
  INV_X1 U12793 ( .A(n12588), .ZN(n10341) );
  OAI22_X1 U12794 ( .A1(n11372), .A2(n10254), .B1(n14988), .B2(n10341), .ZN(
        n10221) );
  XOR2_X1 U12795 ( .A(n12589), .B(n10221), .Z(n11314) );
  INV_X1 U12796 ( .A(n10222), .ZN(n10223) );
  XOR2_X1 U12797 ( .A(n10226), .B(n10225), .Z(n13962) );
  NAND2_X1 U12798 ( .A1(n13963), .A2(n13962), .ZN(n13961) );
  NAND2_X1 U12799 ( .A1(n13961), .A2(n10227), .ZN(n10229) );
  NAND2_X1 U12800 ( .A1(n10229), .A2(n10228), .ZN(n10230) );
  OAI22_X1 U12801 ( .A1(n14994), .A2(n10254), .B1(n11316), .B2(n10374), .ZN(
        n11280) );
  OAI22_X1 U12802 ( .A1(n14994), .A2(n10341), .B1(n11316), .B2(n10254), .ZN(
        n10231) );
  XNOR2_X1 U12803 ( .A(n10231), .B(n12589), .ZN(n11281) );
  OAI22_X1 U12804 ( .A1(n14999), .A2(n10254), .B1(n10234), .B2(n10374), .ZN(
        n10237) );
  OAI22_X1 U12805 ( .A1(n14999), .A2(n10341), .B1(n10234), .B2(n10254), .ZN(
        n10235) );
  XNOR2_X1 U12806 ( .A(n10235), .B(n12589), .ZN(n10236) );
  XOR2_X1 U12807 ( .A(n10237), .B(n10236), .Z(n11653) );
  AND2_X1 U12808 ( .A1(n10237), .A2(n10236), .ZN(n10238) );
  NAND2_X1 U12809 ( .A1(n15006), .A2(n12588), .ZN(n10240) );
  NAND2_X1 U12810 ( .A1(n14130), .A2(n10299), .ZN(n10239) );
  NAND2_X1 U12811 ( .A1(n10240), .A2(n10239), .ZN(n10241) );
  XNOR2_X1 U12812 ( .A(n10241), .B(n10372), .ZN(n10244) );
  NOR2_X1 U12813 ( .A1(n10242), .A2(n10374), .ZN(n10243) );
  AOI21_X1 U12814 ( .B1(n15006), .B2(n12591), .A(n10243), .ZN(n10245) );
  XNOR2_X1 U12815 ( .A(n10244), .B(n10245), .ZN(n11664) );
  NAND2_X1 U12816 ( .A1(n11878), .A2(n12588), .ZN(n10247) );
  OR2_X1 U12817 ( .A1(n11528), .A2(n10254), .ZN(n10246) );
  NAND2_X1 U12818 ( .A1(n10247), .A2(n10246), .ZN(n10248) );
  XNOR2_X1 U12819 ( .A(n10248), .B(n10372), .ZN(n10251) );
  NOR2_X1 U12820 ( .A1(n11528), .A2(n10374), .ZN(n10249) );
  AOI21_X1 U12821 ( .B1(n11878), .B2(n12591), .A(n10249), .ZN(n10250) );
  NAND2_X1 U12822 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  OAI21_X1 U12823 ( .B1(n10251), .B2(n10250), .A(n10252), .ZN(n11871) );
  NOR2_X1 U12824 ( .A1(n11769), .A2(n10374), .ZN(n10253) );
  AOI21_X1 U12825 ( .B1(n12010), .B2(n12591), .A(n10253), .ZN(n10257) );
  OAI22_X1 U12826 ( .A1(n15017), .A2(n10341), .B1(n11769), .B2(n10254), .ZN(
        n10255) );
  XOR2_X1 U12827 ( .A(n12589), .B(n10255), .Z(n12003) );
  OAI22_X1 U12828 ( .A1(n12002), .A2(n12003), .B1(n10257), .B2(n10256), .ZN(
        n12148) );
  AOI22_X1 U12829 ( .A1(n15022), .A2(n12588), .B1(n12591), .B2(n14127), .ZN(
        n10258) );
  XNOR2_X1 U12830 ( .A(n10258), .B(n12589), .ZN(n10260) );
  AOI22_X1 U12831 ( .A1(n15022), .A2(n12591), .B1(n10196), .B2(n14127), .ZN(
        n10259) );
  NAND2_X1 U12832 ( .A1(n10260), .A2(n10259), .ZN(n10262) );
  OAI21_X1 U12833 ( .B1(n10260), .B2(n10259), .A(n10262), .ZN(n12149) );
  INV_X1 U12834 ( .A(n12149), .ZN(n10261) );
  NAND2_X1 U12835 ( .A1(n11740), .A2(n12588), .ZN(n10264) );
  NAND2_X1 U12836 ( .A1(n14126), .A2(n12591), .ZN(n10263) );
  NAND2_X1 U12837 ( .A1(n10264), .A2(n10263), .ZN(n10265) );
  XNOR2_X1 U12838 ( .A(n10265), .B(n12589), .ZN(n10270) );
  AOI22_X1 U12839 ( .A1(n11740), .A2(n12591), .B1(n10196), .B2(n14126), .ZN(
        n10271) );
  XNOR2_X1 U12840 ( .A(n10270), .B(n10271), .ZN(n12204) );
  NAND2_X1 U12841 ( .A1(n14679), .A2(n12588), .ZN(n10267) );
  NAND2_X1 U12842 ( .A1(n14125), .A2(n12591), .ZN(n10266) );
  NAND2_X1 U12843 ( .A1(n10267), .A2(n10266), .ZN(n10268) );
  XNOR2_X1 U12844 ( .A(n10268), .B(n12589), .ZN(n10274) );
  NOR2_X1 U12845 ( .A1(n11738), .A2(n10374), .ZN(n10269) );
  AOI21_X1 U12846 ( .B1(n14679), .B2(n12591), .A(n10269), .ZN(n10275) );
  XNOR2_X1 U12847 ( .A(n10274), .B(n10275), .ZN(n13992) );
  INV_X1 U12848 ( .A(n10270), .ZN(n10272) );
  NAND2_X1 U12849 ( .A1(n10272), .A2(n10271), .ZN(n13989) );
  NAND2_X1 U12850 ( .A1(n12202), .A2(n10273), .ZN(n13991) );
  INV_X1 U12851 ( .A(n10275), .ZN(n10276) );
  NOR2_X1 U12852 ( .A1(n12081), .A2(n10374), .ZN(n10278) );
  AOI21_X1 U12853 ( .B1(n14827), .B2(n12591), .A(n10278), .ZN(n10280) );
  AOI22_X1 U12854 ( .A1(n14827), .A2(n12588), .B1(n12591), .B2(n14124), .ZN(
        n10279) );
  XNOR2_X1 U12855 ( .A(n10279), .B(n12589), .ZN(n10281) );
  XOR2_X1 U12856 ( .A(n10280), .B(n10281), .Z(n14044) );
  NAND2_X1 U12857 ( .A1(n14045), .A2(n14044), .ZN(n10283) );
  OR2_X1 U12858 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  NAND2_X1 U12859 ( .A1(n14820), .A2(n12588), .ZN(n10285) );
  NAND2_X1 U12860 ( .A1(n14123), .A2(n12591), .ZN(n10284) );
  NAND2_X1 U12861 ( .A1(n10285), .A2(n10284), .ZN(n10286) );
  XNOR2_X1 U12862 ( .A(n10286), .B(n10372), .ZN(n10290) );
  NOR2_X1 U12863 ( .A1(n10287), .A2(n10374), .ZN(n10288) );
  AOI21_X1 U12864 ( .B1(n14820), .B2(n12591), .A(n10288), .ZN(n10289) );
  NAND2_X1 U12865 ( .A1(n10290), .A2(n10289), .ZN(n10291) );
  OAI21_X1 U12866 ( .B1(n10290), .B2(n10289), .A(n10291), .ZN(n13941) );
  AOI22_X1 U12867 ( .A1(n14104), .A2(n12588), .B1(n12591), .B2(n10292), .ZN(
        n10293) );
  XOR2_X1 U12868 ( .A(n12589), .B(n10293), .Z(n10295) );
  XNOR2_X2 U12869 ( .A(n10294), .B(n10295), .ZN(n14096) );
  INV_X1 U12870 ( .A(n14104), .ZN(n14814) );
  OAI22_X1 U12871 ( .A1(n14814), .A2(n10254), .B1(n12161), .B2(n10374), .ZN(
        n14095) );
  INV_X1 U12872 ( .A(n10294), .ZN(n10296) );
  NAND2_X1 U12873 ( .A1(n10296), .A2(n10295), .ZN(n10297) );
  NAND2_X1 U12874 ( .A1(n14804), .A2(n12588), .ZN(n10301) );
  OR2_X1 U12875 ( .A1(n14011), .A2(n10254), .ZN(n10300) );
  NAND2_X1 U12876 ( .A1(n10301), .A2(n10300), .ZN(n10302) );
  XNOR2_X1 U12877 ( .A(n10302), .B(n10372), .ZN(n10305) );
  NOR2_X1 U12878 ( .A1(n14011), .A2(n10374), .ZN(n10303) );
  AOI21_X1 U12879 ( .B1(n14804), .B2(n12591), .A(n10303), .ZN(n10304) );
  NAND2_X1 U12880 ( .A1(n10305), .A2(n10304), .ZN(n14018) );
  OAI21_X1 U12881 ( .B1(n10305), .B2(n10304), .A(n14018), .ZN(n14003) );
  NAND2_X1 U12882 ( .A1(n14510), .A2(n12588), .ZN(n10308) );
  OR2_X1 U12883 ( .A1(n14072), .A2(n10254), .ZN(n10307) );
  NAND2_X1 U12884 ( .A1(n10308), .A2(n10307), .ZN(n10309) );
  XNOR2_X1 U12885 ( .A(n10309), .B(n12589), .ZN(n10313) );
  NAND2_X1 U12886 ( .A1(n14510), .A2(n12591), .ZN(n10311) );
  NAND2_X1 U12887 ( .A1(n14121), .A2(n10196), .ZN(n10310) );
  NAND2_X1 U12888 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  NOR2_X1 U12889 ( .A1(n10313), .A2(n10312), .ZN(n10315) );
  AOI21_X1 U12890 ( .B1(n10313), .B2(n10312), .A(n10315), .ZN(n14016) );
  INV_X1 U12891 ( .A(n10315), .ZN(n10316) );
  NAND2_X1 U12892 ( .A1(n14015), .A2(n10316), .ZN(n14066) );
  OAI22_X1 U12893 ( .A1(n14409), .A2(n10254), .B1(n14010), .B2(n10374), .ZN(
        n10323) );
  NAND2_X1 U12894 ( .A1(n14502), .A2(n12588), .ZN(n10318) );
  NAND2_X1 U12895 ( .A1(n14120), .A2(n12591), .ZN(n10317) );
  NAND2_X1 U12896 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  XNOR2_X1 U12897 ( .A(n10319), .B(n12589), .ZN(n10324) );
  XOR2_X1 U12898 ( .A(n10323), .B(n10324), .Z(n14067) );
  NAND2_X1 U12899 ( .A1(n14066), .A2(n14067), .ZN(n13968) );
  AOI22_X1 U12900 ( .A1(n14498), .A2(n12591), .B1(n10196), .B2(n14119), .ZN(
        n10326) );
  NAND2_X1 U12901 ( .A1(n14498), .A2(n12588), .ZN(n10321) );
  NAND2_X1 U12902 ( .A1(n14119), .A2(n12591), .ZN(n10320) );
  NAND2_X1 U12903 ( .A1(n10321), .A2(n10320), .ZN(n10322) );
  XNOR2_X1 U12904 ( .A(n10322), .B(n12589), .ZN(n10328) );
  XOR2_X1 U12905 ( .A(n10326), .B(n10328), .Z(n13969) );
  NOR2_X1 U12906 ( .A1(n10324), .A2(n10323), .ZN(n13970) );
  NOR2_X1 U12907 ( .A1(n13969), .A2(n13970), .ZN(n10325) );
  NAND2_X1 U12908 ( .A1(n13968), .A2(n10325), .ZN(n13972) );
  INV_X1 U12909 ( .A(n10326), .ZN(n10327) );
  NAND2_X1 U12910 ( .A1(n10328), .A2(n10327), .ZN(n10329) );
  OAI22_X1 U12911 ( .A1(n14381), .A2(n10254), .B1(n13984), .B2(n10374), .ZN(
        n10333) );
  NAND2_X1 U12912 ( .A1(n14492), .A2(n12588), .ZN(n10331) );
  OR2_X1 U12913 ( .A1(n13984), .A2(n10254), .ZN(n10330) );
  NAND2_X1 U12914 ( .A1(n10331), .A2(n10330), .ZN(n10332) );
  XNOR2_X1 U12915 ( .A(n10332), .B(n12589), .ZN(n10334) );
  XOR2_X1 U12916 ( .A(n10333), .B(n10334), .Z(n14036) );
  NAND2_X1 U12917 ( .A1(n14035), .A2(n14036), .ZN(n10336) );
  NAND2_X1 U12918 ( .A1(n10334), .A2(n10333), .ZN(n10335) );
  AOI22_X1 U12919 ( .A1(n14486), .A2(n12588), .B1(n12591), .B2(n14117), .ZN(
        n10337) );
  XNOR2_X1 U12920 ( .A(n10337), .B(n12589), .ZN(n10339) );
  AOI22_X1 U12921 ( .A1(n14486), .A2(n12591), .B1(n10196), .B2(n14117), .ZN(
        n10338) );
  NAND2_X1 U12922 ( .A1(n10339), .A2(n10338), .ZN(n14058) );
  OAI21_X1 U12923 ( .B1(n10339), .B2(n10338), .A(n14058), .ZN(n13981) );
  OAI22_X1 U12924 ( .A1(n14348), .A2(n10341), .B1(n13983), .B2(n10254), .ZN(
        n10342) );
  XNOR2_X1 U12925 ( .A(n10342), .B(n10372), .ZN(n10345) );
  OR2_X1 U12926 ( .A1(n14348), .A2(n10254), .ZN(n10344) );
  NAND2_X1 U12927 ( .A1(n14116), .A2(n10196), .ZN(n10343) );
  NAND2_X1 U12928 ( .A1(n10345), .A2(n10346), .ZN(n13956) );
  INV_X1 U12929 ( .A(n10345), .ZN(n10348) );
  INV_X1 U12930 ( .A(n10346), .ZN(n10347) );
  NAND2_X1 U12931 ( .A1(n10348), .A2(n10347), .ZN(n10349) );
  NAND2_X1 U12932 ( .A1(n13953), .A2(n13956), .ZN(n10360) );
  NAND2_X1 U12933 ( .A1(n14472), .A2(n12588), .ZN(n10351) );
  NAND2_X1 U12934 ( .A1(n14115), .A2(n12591), .ZN(n10350) );
  NAND2_X1 U12935 ( .A1(n10351), .A2(n10350), .ZN(n10352) );
  XNOR2_X1 U12936 ( .A(n10352), .B(n10372), .ZN(n10355) );
  NOR2_X1 U12937 ( .A1(n10353), .A2(n10374), .ZN(n10354) );
  AOI21_X1 U12938 ( .B1(n14472), .B2(n12591), .A(n10354), .ZN(n10356) );
  NAND2_X1 U12939 ( .A1(n10355), .A2(n10356), .ZN(n14029) );
  INV_X1 U12940 ( .A(n10355), .ZN(n10358) );
  INV_X1 U12941 ( .A(n10356), .ZN(n10357) );
  NAND2_X1 U12942 ( .A1(n10358), .A2(n10357), .ZN(n10359) );
  NAND2_X1 U12943 ( .A1(n14030), .A2(n14029), .ZN(n10382) );
  NAND2_X1 U12944 ( .A1(n14314), .A2(n12588), .ZN(n10362) );
  OR2_X1 U12945 ( .A1(n13949), .A2(n10254), .ZN(n10361) );
  NAND2_X1 U12946 ( .A1(n10362), .A2(n10361), .ZN(n10363) );
  XNOR2_X1 U12947 ( .A(n10363), .B(n10372), .ZN(n10365) );
  NOR2_X1 U12948 ( .A1(n13949), .A2(n10374), .ZN(n10364) );
  AOI21_X1 U12949 ( .B1(n14314), .B2(n12591), .A(n10364), .ZN(n10366) );
  NAND2_X1 U12950 ( .A1(n10365), .A2(n10366), .ZN(n10384) );
  INV_X1 U12951 ( .A(n10365), .ZN(n10368) );
  INV_X1 U12952 ( .A(n10366), .ZN(n10367) );
  NAND2_X1 U12953 ( .A1(n10368), .A2(n10367), .ZN(n10369) );
  NAND2_X1 U12954 ( .A1(n14460), .A2(n12588), .ZN(n10371) );
  NAND2_X1 U12955 ( .A1(n14113), .A2(n12591), .ZN(n10370) );
  NAND2_X1 U12956 ( .A1(n10371), .A2(n10370), .ZN(n10373) );
  XNOR2_X1 U12957 ( .A(n10373), .B(n10372), .ZN(n10376) );
  INV_X1 U12958 ( .A(n14113), .ZN(n14086) );
  NOR2_X1 U12959 ( .A1(n14086), .A2(n10374), .ZN(n10375) );
  AOI21_X1 U12960 ( .B1(n14460), .B2(n12591), .A(n10375), .ZN(n10377) );
  NAND2_X1 U12961 ( .A1(n10376), .A2(n10377), .ZN(n12563) );
  INV_X1 U12962 ( .A(n10376), .ZN(n10379) );
  INV_X1 U12963 ( .A(n10377), .ZN(n10378) );
  NAND2_X1 U12964 ( .A1(n10379), .A2(n10378), .ZN(n10380) );
  NAND2_X1 U12965 ( .A1(n10382), .A2(n12567), .ZN(n10381) );
  AND2_X1 U12966 ( .A1(n10381), .A2(n12564), .ZN(n10392) );
  NAND3_X1 U12967 ( .A1(n14032), .A2(n10384), .A3(n6499), .ZN(n10391) );
  INV_X1 U12968 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10508) );
  NOR2_X1 U12969 ( .A1(n10385), .A2(n10508), .ZN(n10386) );
  OR2_X1 U12970 ( .A1(n10504), .A2(n10386), .ZN(n10387) );
  NAND2_X1 U12971 ( .A1(n10387), .A2(n10506), .ZN(n10690) );
  OR2_X1 U12972 ( .A1(n10686), .A2(n10690), .ZN(n10399) );
  INV_X1 U12973 ( .A(n10399), .ZN(n10390) );
  OR2_X1 U12974 ( .A1(n14979), .A2(n10513), .ZN(n10388) );
  NOR2_X1 U12975 ( .A1(n10388), .A2(n10512), .ZN(n10389) );
  AOI21_X1 U12976 ( .B1(n10392), .B2(n10391), .A(n14106), .ZN(n10393) );
  NAND2_X1 U12977 ( .A1(n10399), .A2(n10685), .ZN(n10782) );
  NOR2_X1 U12978 ( .A1(n15025), .A2(n10512), .ZN(n10394) );
  NAND2_X1 U12979 ( .A1(n10782), .A2(n10395), .ZN(n10396) );
  NAND2_X1 U12980 ( .A1(n10396), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10397) );
  INV_X1 U12981 ( .A(n14112), .ZN(n10398) );
  OAI22_X1 U12982 ( .A1(n10398), .A2(n14268), .B1(n13949), .B2(n14085), .ZN(
        n14286) );
  OR2_X1 U12983 ( .A1(n10399), .A2(n10691), .ZN(n14073) );
  AOI22_X1 U12984 ( .A1(n14286), .A2(n14097), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10400) );
  OAI21_X1 U12985 ( .B1(n14101), .B2(n14288), .A(n10400), .ZN(n10401) );
  OR2_X1 U12986 ( .A1(n15242), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n10406) );
  NAND2_X1 U12987 ( .A1(n15242), .A2(n15200), .ZN(n13903) );
  OR2_X1 U12988 ( .A1(n10407), .A2(n15439), .ZN(n10411) );
  NOR2_X1 U12989 ( .A1(n15438), .A2(n13187), .ZN(n10408) );
  AOI21_X1 U12990 ( .B1(n9568), .B2(n10409), .A(n10408), .ZN(n10410) );
  NAND2_X1 U12991 ( .A1(n10411), .A2(n10410), .ZN(P3_U3488) );
  INV_X1 U12992 ( .A(n10511), .ZN(n10412) );
  NOR2_X2 U12993 ( .A1(n10413), .A2(n10412), .ZN(P1_U4016) );
  INV_X1 U12994 ( .A(n10414), .ZN(n10415) );
  NAND2_X1 U12995 ( .A1(n6682), .A2(n10416), .ZN(n10417) );
  XNOR2_X1 U12996 ( .A(n10417), .B(n14728), .ZN(n10418) );
  NOR2_X1 U12997 ( .A1(n10418), .A2(n12691), .ZN(n10425) );
  NOR2_X1 U12998 ( .A1(n12706), .A2(n10419), .ZN(n10424) );
  AND2_X1 U12999 ( .A1(n12689), .A2(n14742), .ZN(n10423) );
  INV_X1 U13000 ( .A(n12685), .ZN(n12703) );
  NAND2_X1 U13001 ( .A1(n12703), .A2(n12714), .ZN(n10421) );
  AND2_X1 U13002 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n15302) );
  INV_X1 U13003 ( .A(n15302), .ZN(n10420) );
  OAI211_X1 U13004 ( .C1(n14740), .C2(n12296), .A(n10421), .B(n10420), .ZN(
        n10422) );
  OR4_X1 U13005 ( .A1(n10425), .A2(n10424), .A3(n10423), .A4(n10422), .ZN(
        P3_U3176) );
  XNOR2_X1 U13006 ( .A(n10426), .B(n12407), .ZN(n10427) );
  XNOR2_X1 U13007 ( .A(n10428), .B(n10427), .ZN(n10429) );
  NOR2_X1 U13008 ( .A1(n10429), .A2(n12691), .ZN(n10435) );
  NOR2_X1 U13009 ( .A1(n12405), .A2(n12706), .ZN(n10434) );
  AND2_X1 U13010 ( .A1(n12689), .A2(n12215), .ZN(n10433) );
  INV_X1 U13011 ( .A(n12713), .ZN(n12271) );
  NAND2_X1 U13012 ( .A1(n12698), .A2(n12714), .ZN(n10431) );
  AND2_X1 U13013 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12752) );
  INV_X1 U13014 ( .A(n12752), .ZN(n10430) );
  OAI211_X1 U13015 ( .C1(n12271), .C2(n12685), .A(n10431), .B(n10430), .ZN(
        n10432) );
  OR4_X1 U13016 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        P3_U3174) );
  XNOR2_X1 U13017 ( .A(n10437), .B(n10436), .ZN(n10438) );
  NOR2_X1 U13018 ( .A1(n10438), .A2(n12691), .ZN(n10444) );
  NOR2_X1 U13019 ( .A1(n12247), .A2(n12706), .ZN(n10443) );
  AND2_X1 U13020 ( .A1(n12689), .A2(n12248), .ZN(n10442) );
  NAND2_X1 U13021 ( .A1(n12698), .A2(n12407), .ZN(n10440) );
  INV_X1 U13022 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n10439) );
  OR2_X1 U13023 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10439), .ZN(n12780) );
  OAI211_X1 U13024 ( .C1(n12245), .C2(n12685), .A(n10440), .B(n12780), .ZN(
        n10441) );
  OR4_X1 U13025 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        P3_U3155) );
  NAND2_X1 U13026 ( .A1(n10531), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10445) );
  OR2_X2 U13027 ( .A1(n10530), .A2(n10445), .ZN(n13550) );
  INV_X1 U13028 ( .A(n13550), .ZN(P2_U3947) );
  INV_X1 U13029 ( .A(n15280), .ZN(n10448) );
  NOR2_X1 U13030 ( .A1(n10476), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13410) );
  INV_X2 U13031 ( .A(n13410), .ZN(n13419) );
  INV_X1 U13032 ( .A(SI_7_), .ZN(n10446) );
  OAI222_X1 U13033 ( .A1(P3_U3151), .A2(n10448), .B1(n13419), .B2(n10447), 
        .C1(n13423), .C2(n10446), .ZN(P3_U3288) );
  INV_X1 U13034 ( .A(n10449), .ZN(n10451) );
  OAI222_X1 U13035 ( .A1(P3_U3151), .A2(n11039), .B1(n13419), .B2(n10451), 
        .C1(n10450), .C2(n13423), .ZN(P3_U3295) );
  INV_X1 U13036 ( .A(SI_2_), .ZN(n10452) );
  OAI222_X1 U13037 ( .A1(n11043), .A2(P3_U3151), .B1(n13419), .B2(n10453), 
        .C1(n10452), .C2(n13423), .ZN(P3_U3293) );
  INV_X1 U13038 ( .A(SI_3_), .ZN(n10454) );
  OAI222_X1 U13039 ( .A1(n11047), .A2(P3_U3151), .B1(n13419), .B2(n10455), 
        .C1(n10454), .C2(n13423), .ZN(P3_U3292) );
  NOR2_X1 U13040 ( .A1(n10476), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13922) );
  INV_X1 U13041 ( .A(n13922), .ZN(n13928) );
  OAI222_X1 U13042 ( .A1(n13928), .A2(n10456), .B1(n13920), .B2(n10477), .C1(
        n10553), .C2(P2_U3088), .ZN(P2_U3326) );
  INV_X1 U13043 ( .A(n15065), .ZN(n10458) );
  OAI222_X1 U13044 ( .A1(n13928), .A2(n10459), .B1(n13920), .B2(n8958), .C1(
        n10458), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U13045 ( .A(n10572), .ZN(n10560) );
  OAI222_X1 U13046 ( .A1(n13928), .A2(n10460), .B1(n13920), .B2(n10484), .C1(
        n10560), .C2(P2_U3088), .ZN(P2_U3324) );
  INV_X1 U13047 ( .A(n10461), .ZN(n10463) );
  OAI222_X1 U13048 ( .A1(P3_U3151), .A2(n11592), .B1(n13419), .B2(n10463), 
        .C1(n10462), .C2(n13423), .ZN(P3_U3289) );
  INV_X1 U13049 ( .A(SI_9_), .ZN(n10464) );
  OAI222_X1 U13050 ( .A1(n7302), .A2(P3_U3151), .B1(n13419), .B2(n10465), .C1(
        n10464), .C2(n13423), .ZN(P3_U3286) );
  INV_X1 U13051 ( .A(SI_4_), .ZN(n13184) );
  OAI222_X1 U13052 ( .A1(P3_U3151), .A2(n11050), .B1(n13423), .B2(n13184), 
        .C1(n13419), .C2(n10466), .ZN(P3_U3291) );
  INV_X1 U13053 ( .A(n10467), .ZN(n10468) );
  OAI222_X1 U13054 ( .A1(P3_U3151), .A2(n11812), .B1(n13423), .B2(n13233), 
        .C1(n13419), .C2(n10468), .ZN(P3_U3287) );
  OAI222_X1 U13055 ( .A1(n13419), .A2(n10469), .B1(n13423), .B2(n7498), .C1(
        P3_U3151), .C2(n11041), .ZN(P3_U3294) );
  INV_X1 U13056 ( .A(SI_5_), .ZN(n10471) );
  OAI222_X1 U13057 ( .A1(P3_U3151), .A2(n11054), .B1(n13423), .B2(n10471), 
        .C1(n13419), .C2(n10470), .ZN(P3_U3290) );
  INV_X1 U13058 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10473) );
  INV_X1 U13059 ( .A(n10472), .ZN(n10482) );
  OAI222_X1 U13060 ( .A1(n13928), .A2(n10473), .B1(n13920), .B2(n10482), .C1(
        n10592), .C2(P2_U3088), .ZN(P2_U3323) );
  INV_X1 U13061 ( .A(n12042), .ZN(n11841) );
  INV_X1 U13062 ( .A(SI_10_), .ZN(n10474) );
  OAI222_X1 U13063 ( .A1(n11841), .A2(P3_U3151), .B1(n13419), .B2(n10475), 
        .C1(n10474), .C2(n13423), .ZN(P3_U3285) );
  NAND2_X2 U13064 ( .A1(n10476), .A2(P1_U3086), .ZN(n14542) );
  NOR2_X1 U13065 ( .A1(n10476), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14536) );
  OAI222_X1 U13066 ( .A1(n14542), .A2(n7212), .B1(n14544), .B2(n10477), .C1(
        P1_U3086), .C2(n10608), .ZN(P1_U3354) );
  OAI222_X1 U13067 ( .A1(n14542), .A2(n10478), .B1(n14544), .B2(n8958), .C1(
        P1_U3086), .C2(n14157), .ZN(P1_U3353) );
  INV_X1 U13068 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10480) );
  INV_X1 U13069 ( .A(n10670), .ZN(n10479) );
  OAI222_X1 U13070 ( .A1(n13928), .A2(n10480), .B1(n13920), .B2(n10488), .C1(
        n10479), .C2(P2_U3088), .ZN(P2_U3322) );
  OAI222_X1 U13071 ( .A1(P1_U3086), .A2(n14182), .B1(n14544), .B2(n10482), 
        .C1(n10481), .C2(n14542), .ZN(P1_U3351) );
  OAI222_X1 U13072 ( .A1(P1_U3086), .A2(n10611), .B1(n14544), .B2(n10484), 
        .C1(n10483), .C2(n14542), .ZN(P1_U3352) );
  OAI222_X1 U13073 ( .A1(n15289), .A2(P3_U3151), .B1(n13419), .B2(n10486), 
        .C1(n10485), .C2(n13423), .ZN(P3_U3284) );
  INV_X1 U13074 ( .A(n14542), .ZN(n10497) );
  AOI22_X1 U13075 ( .A1(n10653), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10497), .ZN(n10487) );
  OAI21_X1 U13076 ( .B1(n10488), .B2(n14544), .A(n10487), .ZN(P1_U3350) );
  INV_X1 U13077 ( .A(n10625), .ZN(n10490) );
  OAI222_X1 U13078 ( .A1(P1_U3086), .A2(n10490), .B1(n14544), .B2(n9043), .C1(
        n10489), .C2(n14542), .ZN(P1_U3349) );
  INV_X1 U13079 ( .A(n10752), .ZN(n10676) );
  OAI222_X1 U13080 ( .A1(n13928), .A2(n10491), .B1(n13920), .B2(n9043), .C1(
        n10676), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U13081 ( .A(n10492), .ZN(n10493) );
  OAI222_X1 U13082 ( .A1(n13423), .A2(n10494), .B1(n13419), .B2(n10493), .C1(
        P3_U3151), .C2(n12755), .ZN(P3_U3283) );
  INV_X1 U13083 ( .A(n10495), .ZN(n10499) );
  AOI22_X1 U13084 ( .A1(n10641), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10497), .ZN(n10496) );
  OAI21_X1 U13085 ( .B1(n10499), .B2(n14544), .A(n10496), .ZN(P1_U3348) );
  AOI22_X1 U13086 ( .A1(n10709), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10497), .ZN(n10498) );
  OAI21_X1 U13087 ( .B1(n10502), .B2(n14544), .A(n10498), .ZN(P1_U3347) );
  INV_X1 U13088 ( .A(n10850), .ZN(n10758) );
  OAI222_X1 U13089 ( .A1(n13928), .A2(n10500), .B1(n13920), .B2(n10499), .C1(
        P2_U3088), .C2(n10758), .ZN(P2_U3320) );
  NAND2_X1 U13090 ( .A1(P2_U3947), .A2(n9589), .ZN(n10501) );
  OAI21_X1 U13091 ( .B1(P2_U3947), .B2(n8249), .A(n10501), .ZN(P2_U3531) );
  INV_X1 U13092 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10503) );
  INV_X1 U13093 ( .A(n10966), .ZN(n10856) );
  OAI222_X1 U13094 ( .A1(n13928), .A2(n10503), .B1(n13920), .B2(n10502), .C1(
        n10856), .C2(P2_U3088), .ZN(P2_U3319) );
  NAND2_X1 U13095 ( .A1(n10505), .A2(n10504), .ZN(n14962) );
  INV_X1 U13096 ( .A(n10506), .ZN(n10507) );
  AOI22_X1 U13097 ( .A1(n14962), .A2(n10508), .B1(n10511), .B2(n10507), .ZN(
        P1_U3445) );
  INV_X1 U13098 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n13197) );
  INV_X1 U13099 ( .A(n10509), .ZN(n10510) );
  AOI22_X1 U13100 ( .A1(n14962), .A2(n13197), .B1(n10511), .B2(n10510), .ZN(
        P1_U3446) );
  NAND2_X1 U13101 ( .A1(n10512), .A2(n12071), .ZN(n10603) );
  NAND2_X1 U13102 ( .A1(n10514), .A2(n10513), .ZN(n10515) );
  AND2_X1 U13103 ( .A1(n10515), .A2(n8983), .ZN(n10602) );
  INV_X1 U13104 ( .A(n10602), .ZN(n10516) );
  AND2_X1 U13105 ( .A1(n10603), .A2(n10516), .ZN(n14860) );
  NOR2_X1 U13106 ( .A1(n14860), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13107 ( .A(n11960), .ZN(n10971) );
  OAI222_X1 U13108 ( .A1(n13928), .A2(n10517), .B1(n13920), .B2(n10519), .C1(
        n10971), .C2(P2_U3088), .ZN(P2_U3318) );
  INV_X1 U13109 ( .A(n10813), .ZN(n10707) );
  OAI222_X1 U13110 ( .A1(P1_U3086), .A2(n10707), .B1(n14544), .B2(n10519), 
        .C1(n10518), .C2(n14542), .ZN(P1_U3346) );
  INV_X1 U13111 ( .A(n12768), .ZN(n12772) );
  OAI222_X1 U13112 ( .A1(P3_U3151), .A2(n12772), .B1(n13423), .B2(n10521), 
        .C1(n13419), .C2(n10520), .ZN(P3_U3282) );
  INV_X1 U13113 ( .A(n11116), .ZN(n10523) );
  OAI222_X1 U13114 ( .A1(P1_U3086), .A2(n10523), .B1(n14544), .B2(n10525), 
        .C1(n10522), .C2(n14542), .ZN(P1_U3345) );
  INV_X1 U13115 ( .A(n15076), .ZN(n10524) );
  OAI222_X1 U13116 ( .A1(n13928), .A2(n10526), .B1(n13920), .B2(n10525), .C1(
        n10524), .C2(P2_U3088), .ZN(P2_U3317) );
  INV_X1 U13117 ( .A(n10527), .ZN(n12771) );
  OAI222_X1 U13118 ( .A1(P3_U3151), .A2(n12771), .B1(n13423), .B2(n13168), 
        .C1(n13419), .C2(n10528), .ZN(P3_U3281) );
  OR2_X1 U13119 ( .A1(n10530), .A2(n10529), .ZN(n10536) );
  NAND2_X1 U13120 ( .A1(n10532), .A2(n10531), .ZN(n10534) );
  NAND2_X1 U13121 ( .A1(n10534), .A2(n10533), .ZN(n10535) );
  NAND2_X1 U13122 ( .A1(n10536), .A2(n10535), .ZN(n10546) );
  NOR2_X1 U13123 ( .A1(n10540), .A2(P2_U3088), .ZN(n13921) );
  NAND2_X1 U13124 ( .A1(n10546), .A2(n13921), .ZN(n10537) );
  INV_X1 U13125 ( .A(n15135), .ZN(n13605) );
  INV_X1 U13126 ( .A(n10537), .ZN(n10539) );
  AOI22_X1 U13127 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n13605), .B1(n15129), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10545) );
  INV_X1 U13128 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11467) );
  NAND2_X1 U13129 ( .A1(n15129), .A2(n11467), .ZN(n10542) );
  AND2_X1 U13130 ( .A1(n10540), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10541) );
  INV_X1 U13131 ( .A(n15141), .ZN(n11968) );
  OAI211_X1 U13132 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15135), .A(n10542), .B(
        n11968), .ZN(n10543) );
  INV_X1 U13133 ( .A(n10543), .ZN(n10544) );
  MUX2_X1 U13134 ( .A(n10545), .B(n10544), .S(P2_IR_REG_0__SCAN_IN), .Z(n10548) );
  INV_X1 U13135 ( .A(n15144), .ZN(n15056) );
  AOI22_X1 U13136 ( .A1(n15056), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10547) );
  NAND2_X1 U13137 ( .A1(n10548), .A2(n10547), .ZN(P2_U3214) );
  NAND2_X1 U13138 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15050) );
  AOI21_X1 U13139 ( .B1(n15053), .B2(P2_REG2_REG_1__SCAN_IN), .A(n15048), .ZN(
        n15062) );
  INV_X1 U13140 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10549) );
  MUX2_X1 U13141 ( .A(n10549), .B(P2_REG2_REG_2__SCAN_IN), .S(n15065), .Z(
        n15061) );
  NOR2_X1 U13142 ( .A1(n15062), .A2(n15061), .ZN(n15060) );
  AOI21_X1 U13143 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n15065), .A(n15060), .ZN(
        n10552) );
  INV_X1 U13144 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10550) );
  MUX2_X1 U13145 ( .A(n10550), .B(P2_REG2_REG_3__SCAN_IN), .S(n10572), .Z(
        n10551) );
  NOR2_X1 U13146 ( .A1(n10552), .A2(n10551), .ZN(n10564) );
  AOI211_X1 U13147 ( .C1(n10552), .C2(n10551), .A(n10564), .B(n15120), .ZN(
        n10563) );
  INV_X1 U13148 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n15243) );
  INV_X1 U13149 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10554) );
  MUX2_X1 U13150 ( .A(n10554), .B(P2_REG1_REG_2__SCAN_IN), .S(n15065), .Z(
        n15058) );
  INV_X1 U13151 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10555) );
  MUX2_X1 U13152 ( .A(n10555), .B(P2_REG1_REG_3__SCAN_IN), .S(n10572), .Z(
        n10556) );
  NOR2_X1 U13153 ( .A1(n10557), .A2(n10556), .ZN(n10571) );
  AOI211_X1 U13154 ( .C1(n10557), .C2(n10556), .A(n10571), .B(n15135), .ZN(
        n10562) );
  NAND2_X1 U13155 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n10559) );
  NAND2_X1 U13156 ( .A1(n15056), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n10558) );
  OAI211_X1 U13157 ( .C1(n11968), .C2(n10560), .A(n10559), .B(n10558), .ZN(
        n10561) );
  OR3_X1 U13158 ( .A1(n10563), .A2(n10562), .A3(n10561), .ZN(P2_U3217) );
  INV_X1 U13159 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10565) );
  MUX2_X1 U13160 ( .A(n10565), .B(P2_REG2_REG_4__SCAN_IN), .S(n10592), .Z(
        n10566) );
  INV_X1 U13161 ( .A(n10566), .ZN(n10585) );
  INV_X1 U13162 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10567) );
  MUX2_X1 U13163 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10567), .S(n10670), .Z(
        n10568) );
  INV_X1 U13164 ( .A(n10568), .ZN(n10569) );
  AOI211_X1 U13165 ( .C1(n10570), .C2(n10569), .A(n15120), .B(n10664), .ZN(
        n10583) );
  AOI21_X1 U13166 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n10572), .A(n10571), .ZN(
        n10589) );
  INV_X1 U13167 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10573) );
  MUX2_X1 U13168 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10573), .S(n10592), .Z(
        n10588) );
  NOR2_X1 U13169 ( .A1(n10589), .A2(n10588), .ZN(n10587) );
  INV_X1 U13170 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10575) );
  MUX2_X1 U13171 ( .A(n10575), .B(P2_REG1_REG_5__SCAN_IN), .S(n10670), .Z(
        n10576) );
  NOR2_X1 U13172 ( .A1(n10577), .A2(n10576), .ZN(n10669) );
  AOI211_X1 U13173 ( .C1(n10577), .C2(n10576), .A(n15135), .B(n10669), .ZN(
        n10582) );
  INV_X1 U13174 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10580) );
  NAND2_X1 U13175 ( .A1(n15141), .A2(n10670), .ZN(n10579) );
  NAND2_X1 U13176 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10578) );
  OAI211_X1 U13177 ( .C1(n10580), .C2(n15144), .A(n10579), .B(n10578), .ZN(
        n10581) );
  OR3_X1 U13178 ( .A1(n10583), .A2(n10582), .A3(n10581), .ZN(P2_U3219) );
  AOI211_X1 U13179 ( .C1(n10586), .C2(n10585), .A(n15120), .B(n10584), .ZN(
        n10595) );
  AOI211_X1 U13180 ( .C1(n10589), .C2(n10588), .A(n15135), .B(n10587), .ZN(
        n10594) );
  NAND2_X1 U13181 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10591) );
  NAND2_X1 U13182 ( .A1(n15056), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10590) );
  OAI211_X1 U13183 ( .C1(n11968), .C2(n10592), .A(n10591), .B(n10590), .ZN(
        n10593) );
  OR3_X1 U13184 ( .A1(n10595), .A2(n10594), .A3(n10593), .ZN(P2_U3218) );
  INV_X1 U13185 ( .A(n10596), .ZN(n10663) );
  AOI22_X1 U13186 ( .A1(n15089), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n13922), .ZN(n10597) );
  OAI21_X1 U13187 ( .B1(n10663), .B2(n13920), .A(n10597), .ZN(P2_U3316) );
  MUX2_X1 U13188 ( .A(n11328), .B(P1_REG2_REG_2__SCAN_IN), .S(n14157), .Z(
        n14161) );
  MUX2_X1 U13189 ( .A(n8940), .B(P1_REG2_REG_1__SCAN_IN), .S(n10608), .Z(
        n14143) );
  AND2_X1 U13190 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14149) );
  NAND2_X1 U13191 ( .A1(n14143), .A2(n14149), .ZN(n14142) );
  INV_X1 U13192 ( .A(n10608), .ZN(n14144) );
  NAND2_X1 U13193 ( .A1(n14144), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10598) );
  NAND2_X1 U13194 ( .A1(n14142), .A2(n10598), .ZN(n14160) );
  NAND2_X1 U13195 ( .A1(n14161), .A2(n14160), .ZN(n14159) );
  OR2_X1 U13196 ( .A1(n14157), .A2(n11328), .ZN(n10599) );
  NAND2_X1 U13197 ( .A1(n14159), .A2(n10599), .ZN(n14172) );
  INV_X1 U13198 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n13071) );
  MUX2_X1 U13199 ( .A(n13071), .B(P1_REG2_REG_3__SCAN_IN), .S(n10611), .Z(
        n14173) );
  NAND2_X1 U13200 ( .A1(n14172), .A2(n14173), .ZN(n14171) );
  OR2_X1 U13201 ( .A1(n10611), .A2(n13071), .ZN(n10600) );
  NAND2_X1 U13202 ( .A1(n14171), .A2(n10600), .ZN(n14190) );
  MUX2_X1 U13203 ( .A(n9016), .B(P1_REG2_REG_4__SCAN_IN), .S(n14182), .Z(
        n14191) );
  AND2_X1 U13204 ( .A1(n14190), .A2(n14191), .ZN(n14188) );
  XNOR2_X1 U13205 ( .A(n10653), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n10657) );
  MUX2_X1 U13206 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9047), .S(n10625), .Z(
        n10601) );
  INV_X1 U13207 ( .A(n10601), .ZN(n10605) );
  NAND2_X1 U13208 ( .A1(n10603), .A2(n10602), .ZN(n14862) );
  OR2_X1 U13209 ( .A1(n9524), .A2(n14545), .ZN(n10604) );
  OR2_X1 U13210 ( .A1(n14862), .A2(n10604), .ZN(n14868) );
  AOI211_X1 U13211 ( .C1(n10606), .C2(n10605), .A(n14868), .B(n10621), .ZN(
        n10620) );
  INV_X1 U13212 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10607) );
  MUX2_X1 U13213 ( .A(n10607), .B(P1_REG1_REG_6__SCAN_IN), .S(n10625), .Z(
        n10616) );
  INV_X1 U13214 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15033) );
  MUX2_X1 U13215 ( .A(n15033), .B(P1_REG1_REG_2__SCAN_IN), .S(n14157), .Z(
        n14164) );
  INV_X1 U13216 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15031) );
  MUX2_X1 U13217 ( .A(n15031), .B(P1_REG1_REG_1__SCAN_IN), .S(n10608), .Z(
        n14141) );
  AND2_X1 U13218 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14140) );
  NAND2_X1 U13219 ( .A1(n14141), .A2(n14140), .ZN(n14139) );
  NAND2_X1 U13220 ( .A1(n14144), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U13221 ( .A1(n14139), .A2(n10609), .ZN(n14163) );
  NAND2_X1 U13222 ( .A1(n14164), .A2(n14163), .ZN(n14162) );
  OR2_X1 U13223 ( .A1(n14157), .A2(n15033), .ZN(n10610) );
  NAND2_X1 U13224 ( .A1(n14162), .A2(n10610), .ZN(n14175) );
  INV_X1 U13225 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n15035) );
  MUX2_X1 U13226 ( .A(n15035), .B(P1_REG1_REG_3__SCAN_IN), .S(n10611), .Z(
        n14176) );
  NAND2_X1 U13227 ( .A1(n14175), .A2(n14176), .ZN(n14174) );
  INV_X1 U13228 ( .A(n10611), .ZN(n14170) );
  NAND2_X1 U13229 ( .A1(n14170), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13230 ( .A1(n14174), .A2(n10612), .ZN(n14186) );
  INV_X1 U13231 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15037) );
  MUX2_X1 U13232 ( .A(n15037), .B(P1_REG1_REG_4__SCAN_IN), .S(n14182), .Z(
        n14187) );
  AND2_X1 U13233 ( .A1(n14186), .A2(n14187), .ZN(n14184) );
  XNOR2_X1 U13234 ( .A(n10653), .B(n10614), .ZN(n10652) );
  NAND2_X1 U13235 ( .A1(n10651), .A2(n10652), .ZN(n10650) );
  OAI21_X1 U13236 ( .B1(n10653), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10650), .ZN(
        n10615) );
  NOR2_X1 U13237 ( .A1(n10615), .A2(n10616), .ZN(n10624) );
  AOI211_X1 U13238 ( .C1(n10616), .C2(n10615), .A(n10624), .B(n14864), .ZN(
        n10619) );
  INV_X1 U13239 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14555) );
  INV_X1 U13240 ( .A(n14907), .ZN(n14875) );
  NAND2_X1 U13241 ( .A1(n14875), .A2(n10625), .ZN(n10617) );
  NAND2_X1 U13242 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11656) );
  OAI211_X1 U13243 ( .C1(n14555), .C2(n14912), .A(n10617), .B(n11656), .ZN(
        n10618) );
  OR3_X1 U13244 ( .A1(n10620), .A2(n10619), .A3(n10618), .ZN(P1_U3249) );
  AOI21_X1 U13245 ( .B1(n10625), .B2(P1_REG2_REG_6__SCAN_IN), .A(n10621), .ZN(
        n10623) );
  XNOR2_X1 U13246 ( .A(n10641), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n10622) );
  AOI211_X1 U13247 ( .C1(n10623), .C2(n10622), .A(n14868), .B(n10640), .ZN(
        n10632) );
  XNOR2_X1 U13248 ( .A(n10641), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n10626) );
  NOR2_X1 U13249 ( .A1(n10627), .A2(n10626), .ZN(n10635) );
  AOI211_X1 U13250 ( .C1(n10627), .C2(n10626), .A(n14864), .B(n10635), .ZN(
        n10631) );
  INV_X1 U13251 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14619) );
  NAND2_X1 U13252 ( .A1(n14875), .A2(n10641), .ZN(n10629) );
  NAND2_X1 U13253 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10628) );
  OAI211_X1 U13254 ( .C1(n14619), .C2(n14912), .A(n10629), .B(n10628), .ZN(
        n10630) );
  OR3_X1 U13255 ( .A1(n10632), .A2(n10631), .A3(n10630), .ZN(P1_U3250) );
  OAI222_X1 U13256 ( .A1(P3_U3151), .A2(n14701), .B1(n13423), .B2(n10634), 
        .C1(n13419), .C2(n10633), .ZN(P3_U3280) );
  MUX2_X1 U13257 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10636), .S(n10709), .Z(
        n10637) );
  NAND2_X1 U13258 ( .A1(n10638), .A2(n10637), .ZN(n10702) );
  OAI21_X1 U13259 ( .B1(n10638), .B2(n10637), .A(n10702), .ZN(n10648) );
  INV_X1 U13260 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14623) );
  NAND2_X1 U13261 ( .A1(n14875), .A2(n10709), .ZN(n10639) );
  NAND2_X1 U13262 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11875) );
  OAI211_X1 U13263 ( .C1(n14623), .C2(n14912), .A(n10639), .B(n11875), .ZN(
        n10647) );
  INV_X1 U13264 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10642) );
  MUX2_X1 U13265 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10642), .S(n10709), .Z(
        n10643) );
  INV_X1 U13266 ( .A(n10643), .ZN(n10644) );
  AOI211_X1 U13267 ( .C1(n10645), .C2(n10644), .A(n14868), .B(n10708), .ZN(
        n10646) );
  AOI211_X1 U13268 ( .C1(n14898), .C2(n10648), .A(n10647), .B(n10646), .ZN(
        n10649) );
  INV_X1 U13269 ( .A(n10649), .ZN(P1_U3251) );
  OAI21_X1 U13270 ( .B1(n10652), .B2(n10651), .A(n10650), .ZN(n10661) );
  INV_X1 U13271 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14567) );
  NAND2_X1 U13272 ( .A1(n14875), .A2(n10653), .ZN(n10655) );
  NAND2_X1 U13273 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10654) );
  OAI211_X1 U13274 ( .C1(n14567), .C2(n14912), .A(n10655), .B(n10654), .ZN(
        n10660) );
  AOI211_X1 U13275 ( .C1(n10658), .C2(n10657), .A(n10656), .B(n14868), .ZN(
        n10659) );
  AOI211_X1 U13276 ( .C1(n14898), .C2(n10661), .A(n10660), .B(n10659), .ZN(
        n10662) );
  INV_X1 U13277 ( .A(n10662), .ZN(P1_U3248) );
  INV_X1 U13278 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n13235) );
  INV_X1 U13279 ( .A(n11427), .ZN(n11114) );
  OAI222_X1 U13280 ( .A1(n14542), .A2(n13235), .B1(n14544), .B2(n10663), .C1(
        P1_U3086), .C2(n11114), .ZN(P1_U3344) );
  AOI21_X1 U13281 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n10670), .A(n10664), .ZN(
        n10668) );
  INV_X1 U13282 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10665) );
  MUX2_X1 U13283 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10665), .S(n10752), .Z(
        n10666) );
  INV_X1 U13284 ( .A(n10666), .ZN(n10667) );
  NOR2_X1 U13285 ( .A1(n10668), .A2(n10667), .ZN(n10746) );
  AOI211_X1 U13286 ( .C1(n10668), .C2(n10667), .A(n15120), .B(n10746), .ZN(
        n10679) );
  AOI21_X1 U13287 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n10670), .A(n10669), .ZN(
        n10673) );
  INV_X1 U13288 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10671) );
  MUX2_X1 U13289 ( .A(n10671), .B(P2_REG1_REG_6__SCAN_IN), .S(n10752), .Z(
        n10672) );
  AOI211_X1 U13290 ( .C1(n10673), .C2(n10672), .A(n15135), .B(n10751), .ZN(
        n10678) );
  NAND2_X1 U13291 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10675) );
  NAND2_X1 U13292 ( .A1(n15056), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10674) );
  OAI211_X1 U13293 ( .C1(n11968), .C2(n10676), .A(n10675), .B(n10674), .ZN(
        n10677) );
  OR3_X1 U13294 ( .A1(n10679), .A2(n10678), .A3(n10677), .ZN(P2_U3220) );
  INV_X1 U13295 ( .A(n14937), .ZN(n14917) );
  OAI22_X1 U13296 ( .A1(n11383), .A2(n14917), .B1(n8986), .B2(n14268), .ZN(
        n11379) );
  OR2_X1 U13297 ( .A1(n10682), .A2(n10681), .ZN(n15013) );
  OAI22_X1 U13298 ( .A1(n11383), .A2(n14825), .B1(n11720), .B2(n10683), .ZN(
        n10684) );
  NOR2_X1 U13299 ( .A1(n11379), .A2(n10684), .ZN(n10695) );
  AND2_X1 U13300 ( .A1(n10686), .A2(n10685), .ZN(n10693) );
  INV_X1 U13301 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10688) );
  OR2_X1 U13302 ( .A1(n15030), .A2(n10688), .ZN(n10689) );
  OAI21_X1 U13303 ( .B1(n10695), .B2(n15029), .A(n10689), .ZN(P1_U3459) );
  NOR2_X1 U13304 ( .A1(n10691), .A2(n10690), .ZN(n10692) );
  NAND2_X1 U13305 ( .A1(n15043), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10694) );
  OAI21_X1 U13306 ( .B1(n10695), .B2(n15043), .A(n10694), .ZN(P1_U3528) );
  OAI222_X1 U13307 ( .A1(n13423), .A2(n10697), .B1(n13419), .B2(n10696), .C1(
        n12825), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U13308 ( .A(n10698), .ZN(n10700) );
  AOI22_X1 U13309 ( .A1(n13560), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n13922), .ZN(n10699) );
  OAI21_X1 U13310 ( .B1(n10700), .B2(n13920), .A(n10699), .ZN(P2_U3315) );
  INV_X1 U13311 ( .A(n11622), .ZN(n11433) );
  OAI222_X1 U13312 ( .A1(P1_U3086), .A2(n11433), .B1(n14544), .B2(n10700), 
        .C1(n13062), .C2(n14542), .ZN(P1_U3343) );
  MUX2_X1 U13313 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10701), .S(n10813), .Z(
        n10704) );
  OAI21_X1 U13314 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10709), .A(n10702), .ZN(
        n10703) );
  NAND2_X1 U13315 ( .A1(n10703), .A2(n10704), .ZN(n10812) );
  OAI21_X1 U13316 ( .B1(n10704), .B2(n10703), .A(n10812), .ZN(n10714) );
  NOR2_X1 U13317 ( .A1(n10705), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12005) );
  AOI21_X1 U13318 ( .B1(n14860), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n12005), .ZN(
        n10706) );
  OAI21_X1 U13319 ( .B1(n14907), .B2(n10707), .A(n10706), .ZN(n10713) );
  XNOR2_X1 U13320 ( .A(n10813), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n10710) );
  NOR2_X1 U13321 ( .A1(n10711), .A2(n10710), .ZN(n10806) );
  AOI211_X1 U13322 ( .C1(n10711), .C2(n10710), .A(n14868), .B(n10806), .ZN(
        n10712) );
  AOI211_X1 U13323 ( .C1(n14898), .C2(n10714), .A(n10713), .B(n10712), .ZN(
        n10715) );
  INV_X1 U13324 ( .A(n10715), .ZN(P1_U3252) );
  INV_X1 U13325 ( .A(n13408), .ZN(n10717) );
  NOR2_X1 U13326 ( .A1(n10717), .A2(n10716), .ZN(n10720) );
  CLKBUF_X1 U13327 ( .A(n10720), .Z(n10735) );
  INV_X1 U13328 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10718) );
  NOR2_X1 U13329 ( .A1(n10735), .A2(n10718), .ZN(P3_U3257) );
  INV_X1 U13330 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10719) );
  NOR2_X1 U13331 ( .A1(n10735), .A2(n10719), .ZN(P3_U3263) );
  INV_X1 U13332 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10721) );
  NOR2_X1 U13333 ( .A1(n10735), .A2(n10721), .ZN(P3_U3262) );
  INV_X1 U13334 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10722) );
  NOR2_X1 U13335 ( .A1(n10720), .A2(n10722), .ZN(P3_U3260) );
  INV_X1 U13336 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10723) );
  NOR2_X1 U13337 ( .A1(n10735), .A2(n10723), .ZN(P3_U3259) );
  INV_X1 U13338 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10724) );
  NOR2_X1 U13339 ( .A1(n10720), .A2(n10724), .ZN(P3_U3258) );
  INV_X1 U13340 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10725) );
  NOR2_X1 U13341 ( .A1(n10735), .A2(n10725), .ZN(P3_U3261) );
  INV_X1 U13342 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10726) );
  NOR2_X1 U13343 ( .A1(n10720), .A2(n10726), .ZN(P3_U3234) );
  INV_X1 U13344 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n13222) );
  NOR2_X1 U13345 ( .A1(n10735), .A2(n13222), .ZN(P3_U3256) );
  INV_X1 U13346 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10727) );
  NOR2_X1 U13347 ( .A1(n10735), .A2(n10727), .ZN(P3_U3255) );
  INV_X1 U13348 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10728) );
  NOR2_X1 U13349 ( .A1(n10735), .A2(n10728), .ZN(P3_U3254) );
  INV_X1 U13350 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10729) );
  NOR2_X1 U13351 ( .A1(n10735), .A2(n10729), .ZN(P3_U3253) );
  INV_X1 U13352 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10730) );
  NOR2_X1 U13353 ( .A1(n10735), .A2(n10730), .ZN(P3_U3252) );
  INV_X1 U13354 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10731) );
  NOR2_X1 U13355 ( .A1(n10735), .A2(n10731), .ZN(P3_U3251) );
  INV_X1 U13356 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10732) );
  NOR2_X1 U13357 ( .A1(n10735), .A2(n10732), .ZN(P3_U3250) );
  INV_X1 U13358 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n13200) );
  NOR2_X1 U13359 ( .A1(n10735), .A2(n13200), .ZN(P3_U3249) );
  INV_X1 U13360 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10733) );
  NOR2_X1 U13361 ( .A1(n10735), .A2(n10733), .ZN(P3_U3248) );
  INV_X1 U13362 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10734) );
  NOR2_X1 U13363 ( .A1(n10735), .A2(n10734), .ZN(P3_U3247) );
  INV_X1 U13364 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n13172) );
  NOR2_X1 U13365 ( .A1(n10735), .A2(n13172), .ZN(P3_U3246) );
  INV_X1 U13366 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10736) );
  NOR2_X1 U13367 ( .A1(n10720), .A2(n10736), .ZN(P3_U3245) );
  INV_X1 U13368 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10737) );
  NOR2_X1 U13369 ( .A1(n10720), .A2(n10737), .ZN(P3_U3244) );
  INV_X1 U13370 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10738) );
  NOR2_X1 U13371 ( .A1(n10720), .A2(n10738), .ZN(P3_U3243) );
  INV_X1 U13372 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10739) );
  NOR2_X1 U13373 ( .A1(n10720), .A2(n10739), .ZN(P3_U3242) );
  INV_X1 U13374 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10740) );
  NOR2_X1 U13375 ( .A1(n10720), .A2(n10740), .ZN(P3_U3241) );
  INV_X1 U13376 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10741) );
  NOR2_X1 U13377 ( .A1(n10720), .A2(n10741), .ZN(P3_U3240) );
  INV_X1 U13378 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n13223) );
  NOR2_X1 U13379 ( .A1(n10720), .A2(n13223), .ZN(P3_U3239) );
  INV_X1 U13380 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10742) );
  NOR2_X1 U13381 ( .A1(n10720), .A2(n10742), .ZN(P3_U3238) );
  INV_X1 U13382 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10743) );
  NOR2_X1 U13383 ( .A1(n10735), .A2(n10743), .ZN(P3_U3237) );
  INV_X1 U13384 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10744) );
  NOR2_X1 U13385 ( .A1(n10735), .A2(n10744), .ZN(P3_U3236) );
  INV_X1 U13386 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10745) );
  NOR2_X1 U13387 ( .A1(n10735), .A2(n10745), .ZN(P3_U3235) );
  AOI21_X1 U13388 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n10752), .A(n10746), .ZN(
        n10750) );
  INV_X1 U13389 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10747) );
  MUX2_X1 U13390 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10747), .S(n10850), .Z(
        n10748) );
  INV_X1 U13391 ( .A(n10748), .ZN(n10749) );
  NOR2_X1 U13392 ( .A1(n10750), .A2(n10749), .ZN(n10844) );
  AOI211_X1 U13393 ( .C1(n10750), .C2(n10749), .A(n15120), .B(n10844), .ZN(
        n10761) );
  AOI21_X1 U13394 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n10752), .A(n10751), .ZN(
        n10755) );
  INV_X1 U13395 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10753) );
  MUX2_X1 U13396 ( .A(n10753), .B(P2_REG1_REG_7__SCAN_IN), .S(n10850), .Z(
        n10754) );
  NOR2_X1 U13397 ( .A1(n10755), .A2(n10754), .ZN(n10849) );
  AOI211_X1 U13398 ( .C1(n10755), .C2(n10754), .A(n15135), .B(n10849), .ZN(
        n10760) );
  NAND2_X1 U13399 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n10757) );
  NAND2_X1 U13400 ( .A1(n15056), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10756) );
  OAI211_X1 U13401 ( .C1(n11968), .C2(n10758), .A(n10757), .B(n10756), .ZN(
        n10759) );
  OR3_X1 U13402 ( .A1(n10761), .A2(n10760), .A3(n10759), .ZN(P2_U3221) );
  INV_X1 U13403 ( .A(SI_17_), .ZN(n10763) );
  OAI222_X1 U13404 ( .A1(P3_U3151), .A2(n12849), .B1(n13423), .B2(n10763), 
        .C1(n13419), .C2(n10762), .ZN(P3_U3278) );
  AND2_X1 U13405 ( .A1(n13769), .A2(n9942), .ZN(n10764) );
  OR2_X1 U13406 ( .A1(n10764), .A2(n11471), .ZN(n10765) );
  NAND2_X1 U13407 ( .A1(n13510), .A2(n13551), .ZN(n10797) );
  AND2_X1 U13408 ( .A1(n10765), .A2(n10797), .ZN(n11469) );
  INV_X1 U13409 ( .A(n10766), .ZN(n10767) );
  OAI22_X1 U13410 ( .A1(n11471), .A2(n15223), .B1(n10767), .B2(n9588), .ZN(
        n10768) );
  INV_X1 U13411 ( .A(n10768), .ZN(n10769) );
  AND2_X1 U13412 ( .A1(n11469), .A2(n10769), .ZN(n15189) );
  NAND2_X1 U13413 ( .A1(n9959), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10770) );
  OAI21_X1 U13414 ( .B1(n9959), .B2(n15189), .A(n10770), .ZN(P2_U3499) );
  MUX2_X1 U13415 ( .A(n11127), .B(n12161), .S(n14133), .Z(n10771) );
  INV_X1 U13416 ( .A(n10771), .ZN(P1_U3575) );
  INV_X1 U13417 ( .A(n11896), .ZN(n10774) );
  INV_X1 U13418 ( .A(n10772), .ZN(n10776) );
  OAI222_X1 U13419 ( .A1(P1_U3086), .A2(n10774), .B1(n14544), .B2(n10776), 
        .C1(n10773), .C2(n14542), .ZN(P1_U3342) );
  INV_X1 U13420 ( .A(n13573), .ZN(n11967) );
  OAI222_X1 U13421 ( .A1(P2_U3088), .A2(n11967), .B1(n13920), .B2(n10776), 
        .C1(n10775), .C2(n13928), .ZN(P2_U3314) );
  INV_X1 U13422 ( .A(n14103), .ZN(n14093) );
  XNOR2_X1 U13423 ( .A(n10778), .B(n10779), .ZN(n10780) );
  NAND2_X1 U13424 ( .A1(n10780), .A2(n14082), .ZN(n10784) );
  INV_X1 U13425 ( .A(n14135), .ZN(n11317) );
  OAI22_X1 U13426 ( .A1(n11317), .A2(n14268), .B1(n8986), .B2(n14085), .ZN(
        n11326) );
  NAND2_X1 U13427 ( .A1(n10782), .A2(n10781), .ZN(n10888) );
  AOI22_X1 U13428 ( .A1(n14097), .A2(n11326), .B1(n10888), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10783) );
  OAI211_X1 U13429 ( .C1(n14973), .C2(n14093), .A(n10784), .B(n10783), .ZN(
        P1_U3237) );
  INV_X1 U13430 ( .A(n13515), .ZN(n13493) );
  AOI22_X1 U13431 ( .A1(n13510), .A2(n13547), .B1(n13509), .B2(n13549), .ZN(
        n11566) );
  INV_X1 U13432 ( .A(n11566), .ZN(n10785) );
  AOI22_X1 U13433 ( .A1(n13513), .A2(n10785), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10786) );
  OAI21_X1 U13434 ( .B1(n8883), .B2(n15209), .A(n10786), .ZN(n10792) );
  INV_X1 U13435 ( .A(n10787), .ZN(n10788) );
  AOI211_X1 U13436 ( .C1(n10790), .C2(n10789), .A(n13520), .B(n10788), .ZN(
        n10791) );
  AOI211_X1 U13437 ( .C1(n11568), .C2(n13493), .A(n10792), .B(n10791), .ZN(
        n10793) );
  INV_X1 U13438 ( .A(n10793), .ZN(P2_U3190) );
  INV_X1 U13439 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n13189) );
  NAND2_X1 U13440 ( .A1(P3_U3897), .A2(n13010), .ZN(n10794) );
  OAI21_X1 U13441 ( .B1(P3_U3897), .B2(n13189), .A(n10794), .ZN(P3_U3509) );
  INV_X1 U13442 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n13063) );
  NAND2_X1 U13443 ( .A1(P3_U3897), .A2(n12407), .ZN(n10795) );
  OAI21_X1 U13444 ( .B1(P3_U3897), .B2(n13063), .A(n10795), .ZN(P3_U3504) );
  AOI21_X1 U13445 ( .B1(n13742), .B2(n12224), .A(n13518), .ZN(n10801) );
  INV_X1 U13446 ( .A(n11471), .ZN(n10799) );
  NOR2_X1 U13447 ( .A1(n13520), .A2(n13742), .ZN(n13484) );
  AND2_X1 U13448 ( .A1(n10796), .A2(n15187), .ZN(n10952) );
  INV_X1 U13449 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11468) );
  OAI22_X1 U13450 ( .A1(n13491), .A2(n10797), .B1(n10952), .B2(n11468), .ZN(
        n10798) );
  AOI21_X1 U13451 ( .B1(n10799), .B2(n13484), .A(n10798), .ZN(n10800) );
  OAI21_X1 U13452 ( .B1(n10801), .B2(n9588), .A(n10800), .ZN(P2_U3204) );
  INV_X1 U13453 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U13454 ( .A1(n13284), .A2(P3_U3897), .ZN(n10802) );
  OAI21_X1 U13455 ( .B1(P3_U3897), .B2(n13030), .A(n10802), .ZN(P3_U3510) );
  INV_X1 U13456 ( .A(n10803), .ZN(n10805) );
  OAI222_X1 U13457 ( .A1(n12863), .A2(P3_U3151), .B1(n13419), .B2(n10805), 
        .C1(n10804), .C2(n13423), .ZN(P3_U3277) );
  INV_X1 U13458 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10807) );
  MUX2_X1 U13459 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10807), .S(n11116), .Z(
        n10808) );
  INV_X1 U13460 ( .A(n10808), .ZN(n10809) );
  AOI211_X1 U13461 ( .C1(n10810), .C2(n10809), .A(n14868), .B(n11115), .ZN(
        n10820) );
  MUX2_X1 U13462 ( .A(n10811), .B(P1_REG1_REG_10__SCAN_IN), .S(n11116), .Z(
        n10815) );
  OAI21_X1 U13463 ( .B1(n10813), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10812), .ZN(
        n10814) );
  NOR2_X1 U13464 ( .A1(n10814), .A2(n10815), .ZN(n11109) );
  AOI211_X1 U13465 ( .C1(n10815), .C2(n10814), .A(n14864), .B(n11109), .ZN(
        n10819) );
  INV_X1 U13466 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10817) );
  NAND2_X1 U13467 ( .A1(n14875), .A2(n11116), .ZN(n10816) );
  NAND2_X1 U13468 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n12153)
         );
  OAI211_X1 U13469 ( .C1(n10817), .C2(n14912), .A(n10816), .B(n12153), .ZN(
        n10818) );
  OR3_X1 U13470 ( .A1(n10820), .A2(n10819), .A3(n10818), .ZN(P1_U3253) );
  XNOR2_X1 U13471 ( .A(n10822), .B(n10821), .ZN(n14150) );
  NAND2_X1 U13472 ( .A1(n14097), .A2(n14071), .ZN(n14088) );
  INV_X1 U13473 ( .A(n14088), .ZN(n10823) );
  NAND2_X1 U13474 ( .A1(n10823), .A2(n14137), .ZN(n10825) );
  AOI22_X1 U13475 ( .A1(n14103), .A2(n11380), .B1(n10888), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10824) );
  OAI211_X1 U13476 ( .C1(n14150), .C2(n14106), .A(n10825), .B(n10824), .ZN(
        P1_U3232) );
  OAI21_X1 U13477 ( .B1(n10827), .B2(n10787), .A(n10915), .ZN(n10837) );
  INV_X1 U13478 ( .A(n10827), .ZN(n10829) );
  NAND4_X1 U13479 ( .A1(n13484), .A2(n10829), .A3(n10828), .A4(n6898), .ZN(
        n10835) );
  NAND2_X1 U13480 ( .A1(n13509), .A2(n6898), .ZN(n10831) );
  NAND2_X1 U13481 ( .A1(n13510), .A2(n13546), .ZN(n10830) );
  NAND2_X1 U13482 ( .A1(n10831), .A2(n10830), .ZN(n11262) );
  AOI22_X1 U13483 ( .A1(n13513), .A2(n11262), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10834) );
  OR2_X1 U13484 ( .A1(n13515), .A2(n11257), .ZN(n10833) );
  NAND2_X1 U13485 ( .A1(n13518), .A2(n11259), .ZN(n10832) );
  NAND4_X1 U13486 ( .A1(n10835), .A2(n10834), .A3(n10833), .A4(n10832), .ZN(
        n10836) );
  AOI21_X1 U13487 ( .B1(n10837), .B2(n12224), .A(n10836), .ZN(n10838) );
  INV_X1 U13488 ( .A(n10838), .ZN(P2_U3202) );
  NOR2_X1 U13489 ( .A1(n12689), .A2(P3_U3151), .ZN(n10882) );
  INV_X1 U13490 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10843) );
  AND2_X1 U13491 ( .A1(n10839), .A2(n12328), .ZN(n12417) );
  NOR2_X1 U13492 ( .A1(n12416), .A2(n12417), .ZN(n12383) );
  INV_X1 U13493 ( .A(n12383), .ZN(n10841) );
  OAI22_X1 U13494 ( .A1(n12685), .A2(n8111), .B1(n12328), .B2(n12706), .ZN(
        n10840) );
  AOI21_X1 U13495 ( .B1(n12696), .B2(n10841), .A(n10840), .ZN(n10842) );
  OAI21_X1 U13496 ( .B1(n10882), .B2(n10843), .A(n10842), .ZN(P3_U3172) );
  INV_X1 U13497 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10845) );
  MUX2_X1 U13498 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10845), .S(n10966), .Z(
        n10846) );
  INV_X1 U13499 ( .A(n10846), .ZN(n10847) );
  AOI211_X1 U13500 ( .C1(n10848), .C2(n10847), .A(n15120), .B(n10959), .ZN(
        n10859) );
  INV_X1 U13501 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10851) );
  MUX2_X1 U13502 ( .A(n10851), .B(P2_REG1_REG_8__SCAN_IN), .S(n10966), .Z(
        n10852) );
  AOI211_X1 U13503 ( .C1(n10853), .C2(n10852), .A(n15135), .B(n10965), .ZN(
        n10858) );
  NAND2_X1 U13504 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10855) );
  NAND2_X1 U13505 ( .A1(n15056), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10854) );
  OAI211_X1 U13506 ( .C1(n11968), .C2(n10856), .A(n10855), .B(n10854), .ZN(
        n10857) );
  OR3_X1 U13507 ( .A1(n10859), .A2(n10858), .A3(n10857), .ZN(P2_U3222) );
  INV_X1 U13508 ( .A(n10860), .ZN(n10862) );
  OAI222_X1 U13509 ( .A1(P3_U3151), .A2(n12889), .B1(n13419), .B2(n10862), 
        .C1(n10861), .C2(n13423), .ZN(P3_U3276) );
  INV_X1 U13510 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11176) );
  OAI22_X1 U13511 ( .A1(n12296), .A2(n6506), .B1(n10863), .B2(n12706), .ZN(
        n10864) );
  AOI21_X1 U13512 ( .B1(n12703), .B2(n6803), .A(n10864), .ZN(n10872) );
  INV_X1 U13513 ( .A(n12416), .ZN(n10866) );
  NAND3_X1 U13514 ( .A1(n10866), .A2(n10087), .A3(n10865), .ZN(n10867) );
  OAI211_X1 U13515 ( .C1(n10869), .C2(n11209), .A(n10868), .B(n10867), .ZN(
        n10870) );
  NAND2_X1 U13516 ( .A1(n10870), .A2(n12696), .ZN(n10871) );
  OAI211_X1 U13517 ( .C1(n10882), .C2(n11176), .A(n10872), .B(n10871), .ZN(
        P3_U3162) );
  INV_X1 U13518 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10881) );
  OAI21_X1 U13519 ( .B1(n10875), .B2(n10874), .A(n10873), .ZN(n10876) );
  NAND2_X1 U13520 ( .A1(n10876), .A2(n12696), .ZN(n10880) );
  OAI22_X1 U13521 ( .A1(n12296), .A2(n8111), .B1(n10877), .B2(n12706), .ZN(
        n10878) );
  AOI21_X1 U13522 ( .B1(n12703), .B2(n12719), .A(n10878), .ZN(n10879) );
  OAI211_X1 U13523 ( .C1(n10882), .C2(n10881), .A(n10880), .B(n10879), .ZN(
        P3_U3177) );
  AOI21_X1 U13524 ( .B1(n10885), .B2(n10884), .A(n10883), .ZN(n10890) );
  NOR3_X1 U13525 ( .A1(n14073), .A2(n8938), .A3(n14085), .ZN(n10887) );
  INV_X1 U13526 ( .A(n14136), .ZN(n11371) );
  OAI22_X1 U13527 ( .A1(n14964), .A2(n14093), .B1(n14088), .B2(n11371), .ZN(
        n10886) );
  AOI211_X1 U13528 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n10888), .A(n10887), .B(
        n10886), .ZN(n10889) );
  OAI21_X1 U13529 ( .B1(n10890), .B2(n14106), .A(n10889), .ZN(P1_U3222) );
  INV_X1 U13530 ( .A(n15125), .ZN(n10892) );
  INV_X1 U13531 ( .A(n10891), .ZN(n10894) );
  OAI222_X1 U13532 ( .A1(P2_U3088), .A2(n10892), .B1(n13920), .B2(n10894), 
        .C1(n13109), .C2(n13928), .ZN(P2_U3311) );
  INV_X1 U13533 ( .A(n14874), .ZN(n10895) );
  OAI222_X1 U13534 ( .A1(P1_U3086), .A2(n10895), .B1(n14544), .B2(n10894), 
        .C1(n10893), .C2(n14542), .ZN(P1_U3339) );
  OAI22_X1 U13535 ( .A1(n10897), .A2(n13468), .B1(n13469), .B2(n10896), .ZN(
        n11674) );
  INV_X1 U13536 ( .A(n11674), .ZN(n10898) );
  INV_X1 U13537 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11681) );
  OAI22_X1 U13538 ( .A1(n13491), .A2(n10898), .B1(n11681), .B2(n10952), .ZN(
        n10904) );
  AOI22_X1 U13539 ( .A1(n13484), .A2(n13551), .B1(n12224), .B2(n10899), .ZN(
        n10902) );
  INV_X1 U13540 ( .A(n10900), .ZN(n10948) );
  NOR3_X1 U13541 ( .A1(n10902), .A2(n10948), .A3(n10901), .ZN(n10903) );
  AOI211_X1 U13542 ( .C1(n15199), .C2(n13518), .A(n10904), .B(n10903), .ZN(
        n10905) );
  OAI21_X1 U13543 ( .B1(n10906), .B2(n13520), .A(n10905), .ZN(P2_U3209) );
  INV_X1 U13544 ( .A(n9168), .ZN(n10910) );
  INV_X1 U13545 ( .A(n15101), .ZN(n10907) );
  OAI222_X1 U13546 ( .A1(n13928), .A2(n10908), .B1(n13920), .B2(n10910), .C1(
        n10907), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13547 ( .A(n12062), .ZN(n10911) );
  OAI222_X1 U13548 ( .A1(P1_U3086), .A2(n10911), .B1(n14544), .B2(n10910), 
        .C1(n10909), .C2(n14542), .ZN(P1_U3341) );
  OAI22_X1 U13549 ( .A1(n10913), .A2(n13469), .B1(n13468), .B2(n10912), .ZN(
        n11269) );
  AOI22_X1 U13550 ( .A1(n13513), .A2(n11269), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10914) );
  OAI21_X1 U13551 ( .B1(n8883), .B2(n15227), .A(n10914), .ZN(n10921) );
  INV_X1 U13552 ( .A(n10915), .ZN(n10919) );
  AOI22_X1 U13553 ( .A1(n13484), .A2(n13547), .B1(n12224), .B2(n10916), .ZN(
        n10918) );
  NOR3_X1 U13554 ( .A1(n10919), .A2(n10918), .A3(n10917), .ZN(n10920) );
  AOI211_X1 U13555 ( .C1(n13493), .C2(n11275), .A(n10921), .B(n10920), .ZN(
        n10922) );
  OAI21_X1 U13556 ( .B1(n10923), .B2(n13520), .A(n10922), .ZN(P2_U3199) );
  XNOR2_X1 U13557 ( .A(n10925), .B(n10924), .ZN(n11695) );
  AOI21_X1 U13558 ( .B1(n11271), .B2(n11689), .A(n11852), .ZN(n10926) );
  AND2_X1 U13559 ( .A1(n11086), .A2(n10926), .ZN(n11687) );
  INV_X1 U13560 ( .A(n10927), .ZN(n10928) );
  AOI21_X1 U13561 ( .B1(n10930), .B2(n10929), .A(n10928), .ZN(n10931) );
  AOI22_X1 U13562 ( .A1(n13510), .A2(n13544), .B1(n13509), .B2(n13546), .ZN(
        n10942) );
  OAI21_X1 U13563 ( .B1(n10931), .B2(n13769), .A(n10942), .ZN(n11692) );
  AOI211_X1 U13564 ( .C1(n15212), .C2(n11695), .A(n11687), .B(n11692), .ZN(
        n10936) );
  INV_X1 U13565 ( .A(n13850), .ZN(n11886) );
  AOI22_X1 U13566 ( .A1(n11886), .A2(n11689), .B1(n9959), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10932) );
  OAI21_X1 U13567 ( .B1(n10936), .B2(n9959), .A(n10932), .ZN(P2_U3505) );
  INV_X1 U13568 ( .A(n13903), .ZN(n11884) );
  INV_X1 U13569 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10933) );
  NOR2_X1 U13570 ( .A1(n15242), .A2(n10933), .ZN(n10934) );
  AOI21_X1 U13571 ( .B1(n11884), .B2(n11689), .A(n10934), .ZN(n10935) );
  OAI21_X1 U13572 ( .B1(n10936), .B2(n15240), .A(n10935), .ZN(P2_U3448) );
  INV_X1 U13573 ( .A(n11689), .ZN(n10946) );
  INV_X1 U13574 ( .A(n10937), .ZN(n10986) );
  AOI211_X1 U13575 ( .C1(n10939), .C2(n10938), .A(n13520), .B(n10986), .ZN(
        n10940) );
  INV_X1 U13576 ( .A(n10940), .ZN(n10945) );
  INV_X1 U13577 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10941) );
  OAI22_X1 U13578 ( .A1(n13491), .A2(n10942), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10941), .ZN(n10943) );
  AOI21_X1 U13579 ( .B1(n11688), .B2(n13493), .A(n10943), .ZN(n10944) );
  OAI211_X1 U13580 ( .C1(n10946), .C2(n8883), .A(n10945), .B(n10944), .ZN(
        P2_U3211) );
  INV_X1 U13581 ( .A(n10947), .ZN(n10950) );
  INV_X1 U13582 ( .A(n10954), .ZN(n10949) );
  AOI21_X1 U13583 ( .B1(n10950), .B2(n10949), .A(n10948), .ZN(n10958) );
  AOI22_X1 U13584 ( .A1(n13509), .A2(n9589), .B1(n13510), .B2(n13549), .ZN(
        n15159) );
  INV_X1 U13585 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10951) );
  OAI22_X1 U13586 ( .A1(n13491), .A2(n15159), .B1(n10952), .B2(n10951), .ZN(
        n10956) );
  INV_X1 U13587 ( .A(n13484), .ZN(n12342) );
  NOR3_X1 U13588 ( .A1(n12342), .A2(n10954), .A3(n10953), .ZN(n10955) );
  AOI211_X1 U13589 ( .C1(n15171), .C2(n13518), .A(n10956), .B(n10955), .ZN(
        n10957) );
  OAI21_X1 U13590 ( .B1(n10958), .B2(n13520), .A(n10957), .ZN(P2_U3194) );
  INV_X1 U13591 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10960) );
  MUX2_X1 U13592 ( .A(n10960), .B(P2_REG2_REG_9__SCAN_IN), .S(n11960), .Z(
        n10961) );
  INV_X1 U13593 ( .A(n10961), .ZN(n10962) );
  OAI21_X1 U13594 ( .B1(n10963), .B2(n10962), .A(n11948), .ZN(n10964) );
  NAND2_X1 U13595 ( .A1(n10964), .A2(n15129), .ZN(n10975) );
  INV_X1 U13596 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10967) );
  MUX2_X1 U13597 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10967), .S(n11960), .Z(
        n10968) );
  OAI21_X1 U13598 ( .B1(n10969), .B2(n10968), .A(n11959), .ZN(n10973) );
  NAND2_X1 U13599 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U13600 ( .A1(n15056), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10970) );
  OAI211_X1 U13601 ( .C1(n11968), .C2(n10971), .A(n11237), .B(n10970), .ZN(
        n10972) );
  AOI21_X1 U13602 ( .B1(n10973), .B2(n13605), .A(n10972), .ZN(n10974) );
  NAND2_X1 U13603 ( .A1(n10975), .A2(n10974), .ZN(P2_U3223) );
  AND2_X1 U13604 ( .A1(n10873), .A2(n10976), .ZN(n10979) );
  OAI211_X1 U13605 ( .C1(n10979), .C2(n10978), .A(n12696), .B(n10977), .ZN(
        n10983) );
  NOR2_X1 U13606 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7720), .ZN(n11137) );
  AOI21_X1 U13607 ( .B1(n12679), .B2(n15373), .A(n11137), .ZN(n10980) );
  OAI21_X1 U13608 ( .B1(n12296), .B2(n11103), .A(n10980), .ZN(n10981) );
  AOI21_X1 U13609 ( .B1(n12703), .B2(n12718), .A(n10981), .ZN(n10982) );
  OAI211_X1 U13610 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12700), .A(n10983), .B(
        n10982), .ZN(P3_U3158) );
  NAND3_X1 U13611 ( .A1(n13484), .A2(n10984), .A3(n13545), .ZN(n10988) );
  OAI21_X1 U13612 ( .B1(n10986), .B2(n10985), .A(n12224), .ZN(n10987) );
  AOI21_X1 U13613 ( .B1(n10988), .B2(n10987), .A(n6685), .ZN(n10995) );
  INV_X1 U13614 ( .A(n15148), .ZN(n10993) );
  NAND2_X1 U13615 ( .A1(n13509), .A2(n13545), .ZN(n10990) );
  NAND2_X1 U13616 ( .A1(n13510), .A2(n13543), .ZN(n10989) );
  NAND2_X1 U13617 ( .A1(n10990), .A2(n10989), .ZN(n11089) );
  AOI22_X1 U13618 ( .A1(n13513), .A2(n11089), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10992) );
  NAND2_X1 U13619 ( .A1(n15146), .A2(n13518), .ZN(n10991) );
  OAI211_X1 U13620 ( .C1(n13515), .C2(n10993), .A(n10992), .B(n10991), .ZN(
        n10994) );
  OR2_X1 U13621 ( .A1(n10995), .A2(n10994), .ZN(P2_U3185) );
  INV_X1 U13622 ( .A(n14211), .ZN(n14889) );
  INV_X1 U13623 ( .A(n10996), .ZN(n10999) );
  OAI222_X1 U13624 ( .A1(P1_U3086), .A2(n14889), .B1(n14544), .B2(n10999), 
        .C1(n10997), .C2(n14542), .ZN(P1_U3338) );
  OAI222_X1 U13625 ( .A1(P2_U3088), .A2(n13587), .B1(n13920), .B2(n10999), 
        .C1(n10998), .C2(n13928), .ZN(P2_U3310) );
  NAND2_X1 U13626 ( .A1(P3_U3897), .A2(n13420), .ZN(n15296) );
  MUX2_X1 U13627 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n15255), .Z(n11017) );
  INV_X1 U13628 ( .A(n11017), .ZN(n11018) );
  INV_X1 U13629 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11001) );
  MUX2_X1 U13630 ( .A(n11001), .B(n11000), .S(n15255), .Z(n11002) );
  NAND2_X1 U13631 ( .A1(n11002), .A2(n11027), .ZN(n11016) );
  INV_X1 U13632 ( .A(n11002), .ZN(n11003) );
  NAND2_X1 U13633 ( .A1(n11003), .A2(n11047), .ZN(n11004) );
  AND2_X1 U13634 ( .A1(n11016), .A2(n11004), .ZN(n11133) );
  INV_X1 U13635 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U13636 ( .A1(n11013), .A2(n11206), .ZN(n11015) );
  INV_X1 U13637 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11221) );
  INV_X1 U13638 ( .A(n11041), .ZN(n11187) );
  AND2_X1 U13639 ( .A1(n11008), .A2(n11187), .ZN(n11012) );
  INV_X1 U13640 ( .A(n11012), .ZN(n11007) );
  OAI21_X1 U13641 ( .B1(n11187), .B2(n11008), .A(n11007), .ZN(n11175) );
  INV_X1 U13642 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U13643 ( .A1(n11011), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15263) );
  OAI21_X1 U13644 ( .B1(n11013), .B2(n11206), .A(n11015), .ZN(n11194) );
  NAND2_X1 U13645 ( .A1(n11015), .A2(n11014), .ZN(n11132) );
  XNOR2_X1 U13646 ( .A(n11017), .B(n12722), .ZN(n12732) );
  AOI21_X1 U13647 ( .B1(n12722), .B2(n11018), .A(n12735), .ZN(n11293) );
  MUX2_X1 U13648 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n15255), .Z(n11019) );
  OR2_X1 U13649 ( .A1(n11019), .A2(n11054), .ZN(n11292) );
  INV_X1 U13650 ( .A(n11292), .ZN(n11020) );
  AND2_X1 U13651 ( .A1(n11019), .A2(n11054), .ZN(n11294) );
  NOR2_X1 U13652 ( .A1(n11020), .A2(n11294), .ZN(n11021) );
  XNOR2_X1 U13653 ( .A(n11293), .B(n11021), .ZN(n11066) );
  OR2_X1 U13654 ( .A1(n11023), .A2(P3_U3151), .ZN(n12558) );
  INV_X1 U13655 ( .A(n12558), .ZN(n11022) );
  OR2_X1 U13656 ( .A1(n11219), .A2(n11022), .ZN(n11060) );
  AOI21_X1 U13657 ( .B1(n12530), .B2(n11023), .A(n6848), .ZN(n11058) );
  INV_X1 U13658 ( .A(n11038), .ZN(n11024) );
  MUX2_X1 U13659 ( .A(n12710), .B(n11024), .S(n13420), .Z(n15290) );
  INV_X1 U13660 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11035) );
  NOR2_X1 U13661 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11010), .ZN(n15253) );
  NAND2_X1 U13662 ( .A1(n11026), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11025) );
  OAI21_X1 U13663 ( .B1(n15253), .B2(n11041), .A(n11025), .ZN(n11173) );
  NOR2_X1 U13664 ( .A1(n11173), .A2(n11221), .ZN(n11172) );
  AOI21_X1 U13665 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n11026), .A(n11172), .ZN(
        n11191) );
  NOR2_X1 U13666 ( .A1(n11027), .A2(n11028), .ZN(n11029) );
  NAND2_X1 U13667 ( .A1(n11050), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n11032) );
  INV_X1 U13668 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11030) );
  NAND2_X1 U13669 ( .A1(n12722), .A2(n11030), .ZN(n11031) );
  NAND2_X1 U13670 ( .A1(n11032), .A2(n11031), .ZN(n12725) );
  AOI21_X1 U13671 ( .B1(n11035), .B2(n11034), .A(n11300), .ZN(n11063) );
  INV_X1 U13672 ( .A(n11036), .ZN(n11037) );
  NOR2_X1 U13673 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11040), .ZN(n11042) );
  NOR2_X1 U13674 ( .A1(n11042), .A2(n11179), .ZN(n11199) );
  NAND2_X1 U13675 ( .A1(P3_REG1_REG_2__SCAN_IN), .A2(n11043), .ZN(n11044) );
  OAI21_X1 U13676 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(n11043), .A(n11044), .ZN(
        n11198) );
  INV_X1 U13677 ( .A(n11044), .ZN(n11045) );
  NOR2_X1 U13678 ( .A1(n11027), .A2(n11046), .ZN(n11049) );
  NAND2_X1 U13679 ( .A1(n11050), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U13680 ( .A1(n12722), .A2(n11051), .ZN(n11052) );
  AOI21_X1 U13681 ( .B1(n7668), .B2(n11055), .A(n11304), .ZN(n11056) );
  INV_X1 U13682 ( .A(n11056), .ZN(n11057) );
  NAND2_X1 U13683 ( .A1(n15252), .A2(n11057), .ZN(n11062) );
  INV_X1 U13684 ( .A(n11058), .ZN(n11059) );
  NOR2_X1 U13685 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7664), .ZN(n11340) );
  AOI21_X1 U13686 ( .B1(n15274), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11340), .ZN(
        n11061) );
  OAI211_X1 U13687 ( .C1(n11063), .C2(n15304), .A(n11062), .B(n11061), .ZN(
        n11064) );
  AOI21_X1 U13688 ( .B1(n15281), .B2(n11033), .A(n11064), .ZN(n11065) );
  OAI21_X1 U13689 ( .B1(n15296), .B2(n11066), .A(n11065), .ZN(P3_U3187) );
  NOR3_X1 U13690 ( .A1(n11068), .A2(n11067), .A3(n12342), .ZN(n11069) );
  AOI21_X1 U13691 ( .B1(n6685), .B2(n12224), .A(n11069), .ZN(n11079) );
  INV_X1 U13692 ( .A(n11070), .ZN(n11242) );
  NAND2_X1 U13693 ( .A1(n11712), .A2(n13518), .ZN(n11074) );
  NAND2_X1 U13694 ( .A1(n13509), .A2(n13544), .ZN(n11072) );
  NAND2_X1 U13695 ( .A1(n13510), .A2(n13542), .ZN(n11071) );
  NAND2_X1 U13696 ( .A1(n11072), .A2(n11071), .ZN(n11162) );
  AOI22_X1 U13697 ( .A1(n13513), .A2(n11162), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11073) );
  OAI211_X1 U13698 ( .C1(n13515), .C2(n11075), .A(n11074), .B(n11073), .ZN(
        n11076) );
  AOI21_X1 U13699 ( .B1(n11242), .B2(n12224), .A(n11076), .ZN(n11077) );
  OAI21_X1 U13700 ( .B1(n11079), .B2(n11078), .A(n11077), .ZN(P2_U3193) );
  INV_X1 U13701 ( .A(n11080), .ZN(n11082) );
  OAI222_X1 U13702 ( .A1(n13419), .A2(n11082), .B1(n13423), .B2(n13024), .C1(
        P3_U3151), .C2(n11081), .ZN(P3_U3275) );
  OAI21_X1 U13703 ( .B1(n11085), .B2(n11084), .A(n11083), .ZN(n15155) );
  AOI211_X1 U13704 ( .C1(n15146), .C2(n11086), .A(n11852), .B(n11164), .ZN(
        n15147) );
  XNOR2_X1 U13705 ( .A(n11088), .B(n11087), .ZN(n11090) );
  AOI21_X1 U13706 ( .B1(n11090), .B2(n15161), .A(n11089), .ZN(n15157) );
  INV_X1 U13707 ( .A(n15157), .ZN(n11091) );
  AOI211_X1 U13708 ( .C1(n15212), .C2(n15155), .A(n15147), .B(n11091), .ZN(
        n11096) );
  AOI22_X1 U13709 ( .A1(n11886), .A2(n15146), .B1(n9959), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11092) );
  OAI21_X1 U13710 ( .B1(n11096), .B2(n9959), .A(n11092), .ZN(P2_U3506) );
  INV_X1 U13711 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11093) );
  NOR2_X1 U13712 ( .A1(n15242), .A2(n11093), .ZN(n11094) );
  AOI21_X1 U13713 ( .B1(n11884), .B2(n15146), .A(n11094), .ZN(n11095) );
  OAI21_X1 U13714 ( .B1(n11096), .B2(n15240), .A(n11095), .ZN(P2_U3451) );
  OAI21_X1 U13715 ( .B1(n11098), .B2(n8114), .A(n11097), .ZN(n11099) );
  INV_X1 U13716 ( .A(n11099), .ZN(n15370) );
  INV_X1 U13717 ( .A(n15411), .ZN(n11416) );
  NAND2_X1 U13718 ( .A1(n11100), .A2(n11101), .ZN(n11102) );
  AOI21_X1 U13719 ( .B1(n11102), .B2(n8114), .A(n15388), .ZN(n11106) );
  OAI22_X1 U13720 ( .A1(n11342), .A2(n15382), .B1(n11103), .B2(n15381), .ZN(
        n11104) );
  AOI21_X1 U13721 ( .B1(n11106), .B2(n11105), .A(n11104), .ZN(n15368) );
  OAI21_X1 U13722 ( .B1(n15370), .B2(n11416), .A(n15368), .ZN(n11563) );
  INV_X1 U13723 ( .A(n11563), .ZN(n11108) );
  INV_X1 U13724 ( .A(n13392), .ZN(n13401) );
  AOI22_X1 U13725 ( .A1(n13401), .A2(n15373), .B1(n15428), .B2(
        P3_REG0_REG_3__SCAN_IN), .ZN(n11107) );
  OAI21_X1 U13726 ( .B1(n11108), .B2(n15428), .A(n11107), .ZN(P3_U3399) );
  MUX2_X1 U13727 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11110), .S(n11427), .Z(
        n11111) );
  NAND2_X1 U13728 ( .A1(n11112), .A2(n11111), .ZN(n11423) );
  OAI21_X1 U13729 ( .B1(n11112), .B2(n11111), .A(n11423), .ZN(n11123) );
  AND2_X1 U13730 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12208) );
  AOI21_X1 U13731 ( .B1(n14860), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n12208), 
        .ZN(n11113) );
  OAI21_X1 U13732 ( .B1(n14907), .B2(n11114), .A(n11113), .ZN(n11122) );
  INV_X1 U13733 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11117) );
  MUX2_X1 U13734 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11117), .S(n11427), .Z(
        n11118) );
  INV_X1 U13735 ( .A(n11118), .ZN(n11119) );
  AOI211_X1 U13736 ( .C1(n11120), .C2(n11119), .A(n14868), .B(n11426), .ZN(
        n11121) );
  AOI211_X1 U13737 ( .C1(n14898), .C2(n11123), .A(n11122), .B(n11121), .ZN(
        n11124) );
  INV_X1 U13738 ( .A(n11124), .ZN(P1_U3254) );
  INV_X1 U13739 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n13185) );
  NAND2_X1 U13740 ( .A1(n12920), .A2(P3_U3897), .ZN(n11125) );
  OAI21_X1 U13741 ( .B1(P3_U3897), .B2(n13185), .A(n11125), .ZN(P3_U3516) );
  INV_X1 U13742 ( .A(n11126), .ZN(n11129) );
  INV_X1 U13743 ( .A(n15112), .ZN(n13580) );
  OAI222_X1 U13744 ( .A1(n13928), .A2(n11127), .B1(n13920), .B2(n11129), .C1(
        n13580), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI222_X1 U13745 ( .A1(P1_U3086), .A2(n12058), .B1(n14544), .B2(n11129), 
        .C1(n11128), .C2(n14542), .ZN(P1_U3340) );
  AOI21_X1 U13746 ( .B1(n11001), .B2(n11131), .A(n11130), .ZN(n11147) );
  INV_X1 U13747 ( .A(n11132), .ZN(n11136) );
  INV_X1 U13748 ( .A(n11133), .ZN(n11135) );
  AOI21_X1 U13749 ( .B1(n11136), .B2(n11135), .A(n11134), .ZN(n11139) );
  INV_X1 U13750 ( .A(n11137), .ZN(n11138) );
  OAI21_X1 U13751 ( .B1(n15296), .B2(n11139), .A(n11138), .ZN(n11144) );
  AOI21_X1 U13752 ( .B1(n11000), .B2(n11141), .A(n11140), .ZN(n11142) );
  NOR2_X1 U13753 ( .A1(n15298), .A2(n11142), .ZN(n11143) );
  AOI211_X1 U13754 ( .C1(n15274), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n11144), .B(
        n11143), .ZN(n11146) );
  NAND2_X1 U13755 ( .A1(n15281), .A2(n11027), .ZN(n11145) );
  OAI211_X1 U13756 ( .C1(n11147), .C2(n15304), .A(n11146), .B(n11145), .ZN(
        P3_U3185) );
  INV_X1 U13757 ( .A(n11148), .ZN(n11149) );
  AOI21_X1 U13758 ( .B1(n11151), .B2(n11150), .A(n11149), .ZN(n11157) );
  AND2_X1 U13759 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n12723) );
  NOR2_X1 U13760 ( .A1(n12706), .A2(n11577), .ZN(n11152) );
  AOI211_X1 U13761 ( .C1(n12698), .C2(n12719), .A(n12723), .B(n11152), .ZN(
        n11153) );
  OAI21_X1 U13762 ( .B1(n11454), .B2(n12685), .A(n11153), .ZN(n11154) );
  AOI21_X1 U13763 ( .B1(n11155), .B2(n12689), .A(n11154), .ZN(n11156) );
  OAI21_X1 U13764 ( .B1(n11157), .B2(n12691), .A(n11156), .ZN(P3_U3170) );
  INV_X1 U13765 ( .A(n11160), .ZN(n11159) );
  OAI21_X1 U13766 ( .B1(n6691), .B2(n11159), .A(n11158), .ZN(n11710) );
  XNOR2_X1 U13767 ( .A(n11161), .B(n11160), .ZN(n11163) );
  AOI21_X1 U13768 ( .B1(n11163), .B2(n15161), .A(n11162), .ZN(n11719) );
  OAI211_X1 U13769 ( .C1(n11168), .C2(n11164), .A(n13742), .B(n11351), .ZN(
        n11715) );
  OAI211_X1 U13770 ( .C1(n11710), .C2(n13861), .A(n11719), .B(n11715), .ZN(
        n11170) );
  OAI22_X1 U13771 ( .A1(n13850), .A2(n11168), .B1(n15250), .B2(n10851), .ZN(
        n11165) );
  AOI21_X1 U13772 ( .B1(n11170), .B2(n15250), .A(n11165), .ZN(n11166) );
  INV_X1 U13773 ( .A(n11166), .ZN(P2_U3507) );
  INV_X1 U13774 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11167) );
  OAI22_X1 U13775 ( .A1(n13903), .A2(n11168), .B1(n15242), .B2(n11167), .ZN(
        n11169) );
  AOI21_X1 U13776 ( .B1(n11170), .B2(n15242), .A(n11169), .ZN(n11171) );
  INV_X1 U13777 ( .A(n11171), .ZN(P2_U3454) );
  AOI21_X1 U13778 ( .B1(n11221), .B2(n11173), .A(n11172), .ZN(n11185) );
  AOI21_X1 U13779 ( .B1(n11175), .B2(n15263), .A(n11174), .ZN(n11177) );
  OAI22_X1 U13780 ( .A1(n15296), .A2(n11177), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11176), .ZN(n11178) );
  AOI21_X1 U13781 ( .B1(n15274), .B2(P3_ADDR_REG_1__SCAN_IN), .A(n11178), .ZN(
        n11184) );
  AOI21_X1 U13782 ( .B1(n15431), .B2(n11180), .A(n11179), .ZN(n11181) );
  INV_X1 U13783 ( .A(n11181), .ZN(n11182) );
  NAND2_X1 U13784 ( .A1(n15252), .A2(n11182), .ZN(n11183) );
  OAI211_X1 U13785 ( .C1(n11185), .C2(n15304), .A(n11184), .B(n11183), .ZN(
        n11186) );
  AOI21_X1 U13786 ( .B1(n15281), .B2(n11187), .A(n11186), .ZN(n11188) );
  INV_X1 U13787 ( .A(n11188), .ZN(P3_U3183) );
  AOI21_X1 U13788 ( .B1(n11191), .B2(n11190), .A(n11189), .ZN(n11204) );
  AOI21_X1 U13789 ( .B1(n11194), .B2(n11193), .A(n11192), .ZN(n11195) );
  OAI22_X1 U13790 ( .A1(n15296), .A2(n11195), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10881), .ZN(n11196) );
  AOI21_X1 U13791 ( .B1(n15274), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n11196), .ZN(
        n11203) );
  AOI21_X1 U13792 ( .B1(n11199), .B2(n11198), .A(n11197), .ZN(n11200) );
  INV_X1 U13793 ( .A(n11200), .ZN(n11201) );
  NAND2_X1 U13794 ( .A1(n15252), .A2(n11201), .ZN(n11202) );
  OAI211_X1 U13795 ( .C1(n11204), .C2(n15304), .A(n11203), .B(n11202), .ZN(
        n11205) );
  AOI21_X1 U13796 ( .B1(n15281), .B2(n11206), .A(n11205), .ZN(n11207) );
  INV_X1 U13797 ( .A(n11207), .ZN(P3_U3184) );
  AND2_X1 U13798 ( .A1(n15410), .A2(n11208), .ZN(n15400) );
  XNOR2_X1 U13799 ( .A(n10087), .B(n11209), .ZN(n11210) );
  NAND2_X1 U13800 ( .A1(n11210), .A2(n15341), .ZN(n11212) );
  AOI22_X1 U13801 ( .A1(n15326), .A2(n10839), .B1(n15324), .B2(n6803), .ZN(
        n11211) );
  NAND2_X1 U13802 ( .A1(n11212), .A2(n11211), .ZN(n15399) );
  AOI21_X1 U13803 ( .B1(n15400), .B2(n12551), .A(n15399), .ZN(n11220) );
  INV_X1 U13804 ( .A(n13407), .ZN(n11213) );
  XNOR2_X1 U13805 ( .A(n11214), .B(n11213), .ZN(n11215) );
  NAND3_X1 U13806 ( .A1(n11217), .A2(n11216), .A3(n11215), .ZN(n11704) );
  NOR2_X1 U13807 ( .A1(n15346), .A2(n12551), .ZN(n11218) );
  MUX2_X1 U13808 ( .A(n11221), .B(n11220), .S(n15396), .Z(n11223) );
  AND2_X1 U13809 ( .A1(n12414), .A2(n15392), .ZN(n15390) );
  INV_X1 U13810 ( .A(n10087), .ZN(n12384) );
  XNOR2_X1 U13811 ( .A(n12416), .B(n12384), .ZN(n15401) );
  INV_X2 U13812 ( .A(n15376), .ZN(n15395) );
  AOI22_X1 U13813 ( .A1(n13306), .A2(n15401), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15395), .ZN(n11222) );
  NAND2_X1 U13814 ( .A1(n11223), .A2(n11222), .ZN(P3_U3232) );
  OAI21_X1 U13815 ( .B1(n11225), .B2(n12435), .A(n11224), .ZN(n11226) );
  INV_X1 U13816 ( .A(n11226), .ZN(n15362) );
  OAI211_X1 U13817 ( .C1(n11229), .C2(n11228), .A(n11227), .B(n15341), .ZN(
        n11231) );
  AOI22_X1 U13818 ( .A1(n15326), .A2(n12719), .B1(n15324), .B2(n12717), .ZN(
        n11230) );
  AND2_X1 U13819 ( .A1(n11231), .A2(n11230), .ZN(n15361) );
  OAI21_X1 U13820 ( .B1(n15362), .B2(n11416), .A(n15361), .ZN(n11579) );
  INV_X1 U13821 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n11232) );
  OAI22_X1 U13822 ( .A1(n11577), .A2(n13392), .B1(n15430), .B2(n11232), .ZN(
        n11233) );
  AOI21_X1 U13823 ( .B1(n11579), .B2(n15430), .A(n11233), .ZN(n11234) );
  INV_X1 U13824 ( .A(n11234), .ZN(P3_U3402) );
  NAND2_X1 U13825 ( .A1(n13509), .A2(n13543), .ZN(n11236) );
  NAND2_X1 U13826 ( .A1(n13510), .A2(n13541), .ZN(n11235) );
  AND2_X1 U13827 ( .A1(n11236), .A2(n11235), .ZN(n11349) );
  NAND2_X1 U13828 ( .A1(n13493), .A2(n11354), .ZN(n11238) );
  OAI211_X1 U13829 ( .C1(n13491), .C2(n11349), .A(n11238), .B(n11237), .ZN(
        n11244) );
  AOI22_X1 U13830 ( .A1(n11239), .A2(n12224), .B1(n13484), .B2(n13543), .ZN(
        n11241) );
  NOR3_X1 U13831 ( .A1(n11242), .A2(n11241), .A3(n11240), .ZN(n11243) );
  AOI211_X1 U13832 ( .C1(n11443), .C2(n13518), .A(n11244), .B(n11243), .ZN(
        n11245) );
  OAI21_X1 U13833 ( .B1(n11246), .B2(n13520), .A(n11245), .ZN(P2_U3203) );
  INV_X1 U13834 ( .A(n11250), .ZN(n11470) );
  AND2_X1 U13835 ( .A1(n9942), .A2(n11470), .ZN(n11251) );
  XNOR2_X1 U13836 ( .A(n11252), .B(n11260), .ZN(n15218) );
  NOR2_X2 U13837 ( .A1(n11254), .A2(n13700), .ZN(n15169) );
  INV_X1 U13838 ( .A(n15169), .ZN(n13747) );
  INV_X1 U13839 ( .A(n11571), .ZN(n11256) );
  INV_X1 U13840 ( .A(n11255), .ZN(n11273) );
  OAI211_X1 U13841 ( .C1(n15217), .C2(n11256), .A(n11273), .B(n13742), .ZN(
        n15215) );
  OAI22_X1 U13842 ( .A1(n13747), .A2(n15215), .B1(n11257), .B2(n13774), .ZN(
        n11258) );
  AOI21_X1 U13843 ( .B1(n15170), .B2(n11259), .A(n11258), .ZN(n11265) );
  XNOR2_X1 U13844 ( .A(n11261), .B(n11260), .ZN(n11263) );
  AOI21_X1 U13845 ( .B1(n11263), .B2(n15161), .A(n11262), .ZN(n15216) );
  MUX2_X1 U13846 ( .A(n15216), .B(n10565), .S(n15174), .Z(n11264) );
  OAI211_X1 U13847 ( .C1(n13793), .C2(n15218), .A(n11265), .B(n11264), .ZN(
        P2_U3261) );
  XOR2_X1 U13848 ( .A(n11267), .B(n11266), .Z(n15222) );
  XOR2_X1 U13849 ( .A(n11268), .B(n11267), .Z(n11270) );
  AOI21_X1 U13850 ( .B1(n11270), .B2(n15161), .A(n11269), .ZN(n15226) );
  MUX2_X1 U13851 ( .A(n10567), .B(n15226), .S(n11353), .Z(n11279) );
  INV_X1 U13852 ( .A(n11271), .ZN(n11272) );
  AOI211_X1 U13853 ( .C1(n11274), .C2(n11273), .A(n11852), .B(n11272), .ZN(
        n15224) );
  INV_X1 U13854 ( .A(n11275), .ZN(n11276) );
  OAI22_X1 U13855 ( .A1(n15152), .A2(n15227), .B1(n13774), .B2(n11276), .ZN(
        n11277) );
  AOI21_X1 U13856 ( .B1(n15224), .B2(n15169), .A(n11277), .ZN(n11278) );
  OAI211_X1 U13857 ( .C1(n13793), .C2(n15222), .A(n11279), .B(n11278), .ZN(
        P2_U3260) );
  XNOR2_X1 U13858 ( .A(n11281), .B(n11280), .ZN(n11282) );
  XNOR2_X1 U13859 ( .A(n11283), .B(n11282), .ZN(n11289) );
  AOI22_X1 U13860 ( .A1(n14052), .A2(n14134), .B1(n14131), .B2(n14071), .ZN(
        n11388) );
  OAI22_X1 U13861 ( .A1(n14073), .A2(n11388), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11284), .ZN(n11286) );
  NOR2_X1 U13862 ( .A1(n14101), .A2(n11391), .ZN(n11285) );
  AOI211_X1 U13863 ( .C1(n14103), .C2(n11287), .A(n11286), .B(n11285), .ZN(
        n11288) );
  OAI21_X1 U13864 ( .B1(n11289), .B2(n14106), .A(n11288), .ZN(P1_U3227) );
  INV_X1 U13865 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11290) );
  NOR2_X1 U13866 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11290), .ZN(n11451) );
  MUX2_X1 U13867 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n15255), .Z(n11593) );
  INV_X1 U13868 ( .A(n11592), .ZN(n11291) );
  XNOR2_X1 U13869 ( .A(n11593), .B(n11291), .ZN(n11296) );
  OAI21_X1 U13870 ( .B1(n11294), .B2(n11293), .A(n11292), .ZN(n11295) );
  NAND2_X1 U13871 ( .A1(n11296), .A2(n11295), .ZN(n11594) );
  OAI21_X1 U13872 ( .B1(n11296), .B2(n11295), .A(n11594), .ZN(n11297) );
  AND2_X1 U13873 ( .A1(n15279), .A2(n11297), .ZN(n11298) );
  AOI211_X1 U13874 ( .C1(n15274), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n11451), .B(
        n11298), .ZN(n11310) );
  INV_X1 U13875 ( .A(n15304), .ZN(n15254) );
  NAND2_X1 U13876 ( .A1(n11592), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n11585) );
  OR2_X1 U13877 ( .A1(n11592), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n11302) );
  OAI21_X1 U13878 ( .B1(n6700), .B2(n6704), .A(n11586), .ZN(n11308) );
  NOR2_X1 U13879 ( .A1(n11033), .A2(n11303), .ZN(n11305) );
  NAND2_X1 U13880 ( .A1(n11592), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11604) );
  OR2_X1 U13881 ( .A1(n11592), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11306) );
  OAI21_X1 U13882 ( .B1(n7315), .B2(n6705), .A(n11605), .ZN(n11307) );
  AOI22_X1 U13883 ( .A1(n15254), .A2(n11308), .B1(n11307), .B2(n15252), .ZN(
        n11309) );
  OAI211_X1 U13884 ( .C1(n11592), .C2(n15290), .A(n11310), .B(n11309), .ZN(
        P3_U3188) );
  INV_X1 U13885 ( .A(n11311), .ZN(n11312) );
  AOI211_X1 U13886 ( .C1(n11314), .C2(n11313), .A(n14106), .B(n11312), .ZN(
        n11315) );
  INV_X1 U13887 ( .A(n11315), .ZN(n11320) );
  OAI22_X1 U13888 ( .A1(n11317), .A2(n14085), .B1(n11316), .B2(n14268), .ZN(
        n14936) );
  AND2_X1 U13889 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14180) );
  NOR2_X1 U13890 ( .A1(n14093), .A2(n14988), .ZN(n11318) );
  AOI211_X1 U13891 ( .C1(n14097), .C2(n14936), .A(n14180), .B(n11318), .ZN(
        n11319) );
  OAI211_X1 U13892 ( .C1(n14101), .C2(n14939), .A(n11320), .B(n11319), .ZN(
        P1_U3230) );
  XNOR2_X1 U13893 ( .A(n11321), .B(n11324), .ZN(n14971) );
  OR2_X1 U13894 ( .A1(n14942), .A2(n14674), .ZN(n14926) );
  OAI21_X1 U13895 ( .B1(n11324), .B2(n11323), .A(n11322), .ZN(n11327) );
  NOR2_X1 U13896 ( .A1(n14971), .A2(n14966), .ZN(n11325) );
  AOI211_X1 U13897 ( .C1(n14937), .C2(n11327), .A(n11326), .B(n11325), .ZN(
        n14974) );
  MUX2_X1 U13898 ( .A(n11328), .B(n14974), .S(n14427), .Z(n11335) );
  INV_X1 U13899 ( .A(n11721), .ZN(n11330) );
  INV_X1 U13900 ( .A(n11329), .ZN(n11365) );
  OAI211_X1 U13901 ( .C1(n14973), .C2(n11330), .A(n11365), .B(n14948), .ZN(
        n14972) );
  OAI22_X1 U13902 ( .A1(n14334), .A2(n14972), .B1(n11331), .B2(n14940), .ZN(
        n11332) );
  AOI21_X1 U13903 ( .B1(n14417), .B2(n11333), .A(n11332), .ZN(n11334) );
  OAI211_X1 U13904 ( .C1(n14971), .C2(n14926), .A(n11335), .B(n11334), .ZN(
        P1_U3291) );
  OAI21_X1 U13905 ( .B1(n11338), .B2(n11337), .A(n11336), .ZN(n11339) );
  NAND2_X1 U13906 ( .A1(n11339), .A2(n12696), .ZN(n11345) );
  AOI21_X1 U13907 ( .B1(n12679), .B2(n15358), .A(n11340), .ZN(n11341) );
  OAI21_X1 U13908 ( .B1(n12296), .B2(n11342), .A(n11341), .ZN(n11343) );
  AOI21_X1 U13909 ( .B1(n12703), .B2(n12716), .A(n11343), .ZN(n11344) );
  OAI211_X1 U13910 ( .C1(n15360), .C2(n12700), .A(n11345), .B(n11344), .ZN(
        P3_U3167) );
  XOR2_X1 U13911 ( .A(n11347), .B(n11346), .Z(n11439) );
  INV_X1 U13912 ( .A(n11439), .ZN(n11360) );
  OAI211_X1 U13913 ( .C1(n6849), .C2(n9850), .A(n15161), .B(n11348), .ZN(
        n11350) );
  NAND2_X1 U13914 ( .A1(n11350), .A2(n11349), .ZN(n11437) );
  INV_X1 U13915 ( .A(n11443), .ZN(n11357) );
  NAND2_X1 U13916 ( .A1(n11443), .A2(n11351), .ZN(n11352) );
  AND3_X1 U13917 ( .A1(n11496), .A2(n13742), .A3(n11352), .ZN(n11438) );
  NAND2_X1 U13918 ( .A1(n11438), .A2(n15169), .ZN(n11356) );
  AOI22_X1 U13919 ( .A1(n15149), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11354), 
        .B2(n15163), .ZN(n11355) );
  OAI211_X1 U13920 ( .C1(n11357), .C2(n15152), .A(n11356), .B(n11355), .ZN(
        n11358) );
  AOI21_X1 U13921 ( .B1(n11437), .B2(n11353), .A(n11358), .ZN(n11359) );
  OAI21_X1 U13922 ( .B1(n11360), .B2(n13793), .A(n11359), .ZN(P2_U3256) );
  INV_X1 U13923 ( .A(n11361), .ZN(n11363) );
  OAI22_X1 U13924 ( .A1(n12555), .A2(P3_U3151), .B1(SI_22_), .B2(n13423), .ZN(
        n11362) );
  AOI21_X1 U13925 ( .B1(n11363), .B2(n13410), .A(n11362), .ZN(P3_U3273) );
  XNOR2_X1 U13926 ( .A(n11369), .B(n11364), .ZN(n14983) );
  AOI211_X1 U13927 ( .C1(n14980), .C2(n11365), .A(n14829), .B(n14949), .ZN(
        n14978) );
  INV_X1 U13928 ( .A(n14978), .ZN(n11366) );
  OAI22_X1 U13929 ( .A1(n11366), .A2(n14334), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14940), .ZN(n11367) );
  AOI21_X1 U13930 ( .B1(n14417), .B2(n14980), .A(n11367), .ZN(n11375) );
  OAI21_X1 U13931 ( .B1(n11370), .B2(n11369), .A(n11368), .ZN(n11373) );
  OAI22_X1 U13932 ( .A1(n11372), .A2(n14268), .B1(n11371), .B2(n14085), .ZN(
        n13964) );
  AOI21_X1 U13933 ( .B1(n11373), .B2(n14937), .A(n13964), .ZN(n14982) );
  MUX2_X1 U13934 ( .A(n13071), .B(n14982), .S(n14427), .Z(n11374) );
  OAI211_X1 U13935 ( .C1(n14432), .C2(n14983), .A(n11375), .B(n11374), .ZN(
        P1_U3290) );
  OAI22_X1 U13936 ( .A1(n14427), .A2(n11377), .B1(n11376), .B2(n14940), .ZN(
        n11378) );
  AOI21_X1 U13937 ( .B1(n14427), .B2(n11379), .A(n11378), .ZN(n11382) );
  NOR2_X1 U13938 ( .A1(n14334), .A2(n14829), .ZN(n14263) );
  OAI21_X1 U13939 ( .B1(n14417), .B2(n14263), .A(n11380), .ZN(n11381) );
  OAI211_X1 U13940 ( .C1(n14432), .C2(n11383), .A(n11382), .B(n11381), .ZN(
        P1_U3293) );
  XNOR2_X1 U13941 ( .A(n11384), .B(n11387), .ZN(n14991) );
  OAI21_X1 U13942 ( .B1(n11387), .B2(n11386), .A(n11385), .ZN(n11390) );
  INV_X1 U13943 ( .A(n11388), .ZN(n11389) );
  AOI21_X1 U13944 ( .B1(n11390), .B2(n14937), .A(n11389), .ZN(n14993) );
  INV_X1 U13945 ( .A(n14993), .ZN(n11396) );
  OAI211_X1 U13946 ( .C1(n14951), .C2(n14994), .A(n14948), .B(n14927), .ZN(
        n14992) );
  NOR2_X1 U13947 ( .A1(n14992), .A2(n14334), .ZN(n11395) );
  NOR2_X1 U13948 ( .A1(n14940), .A2(n11391), .ZN(n11392) );
  AOI21_X1 U13949 ( .B1(n14942), .B2(P1_REG2_REG_5__SCAN_IN), .A(n11392), .ZN(
        n11393) );
  OAI21_X1 U13950 ( .B1(n14944), .B2(n14994), .A(n11393), .ZN(n11394) );
  AOI211_X1 U13951 ( .C1(n11396), .C2(n14427), .A(n11395), .B(n11394), .ZN(
        n11397) );
  OAI21_X1 U13952 ( .B1(n14432), .B2(n14991), .A(n11397), .ZN(P1_U3288) );
  XOR2_X1 U13953 ( .A(n11398), .B(n11399), .Z(n11549) );
  AOI21_X1 U13954 ( .B1(n11400), .B2(n11399), .A(n14917), .ZN(n11404) );
  OR2_X1 U13955 ( .A1(n11769), .A2(n14268), .ZN(n11402) );
  NAND2_X1 U13956 ( .A1(n14130), .A2(n14052), .ZN(n11401) );
  NAND2_X1 U13957 ( .A1(n11402), .A2(n11401), .ZN(n11873) );
  AOI21_X1 U13958 ( .B1(n11404), .B2(n11403), .A(n11873), .ZN(n11546) );
  INV_X1 U13959 ( .A(n11516), .ZN(n11405) );
  AOI21_X1 U13960 ( .B1(n11878), .B2(n11405), .A(n11530), .ZN(n11544) );
  AOI22_X1 U13961 ( .A1(n11544), .A2(n14948), .B1(n11878), .B2(n14979), .ZN(
        n11406) );
  OAI211_X1 U13962 ( .C1(n11549), .C2(n14825), .A(n11546), .B(n11406), .ZN(
        n11408) );
  NAND2_X1 U13963 ( .A1(n11408), .A2(n15045), .ZN(n11407) );
  OAI21_X1 U13964 ( .B1(n15045), .B2(n10636), .A(n11407), .ZN(P1_U3536) );
  NAND2_X1 U13965 ( .A1(n11408), .A2(n15030), .ZN(n11409) );
  OAI21_X1 U13966 ( .B1(n15030), .B2(n9082), .A(n11409), .ZN(P1_U3483) );
  OAI21_X1 U13967 ( .B1(n11411), .B2(n12382), .A(n11410), .ZN(n11412) );
  INV_X1 U13968 ( .A(n11412), .ZN(n15355) );
  OAI21_X1 U13969 ( .B1(n11414), .B2(n8119), .A(n11413), .ZN(n11415) );
  AOI222_X1 U13970 ( .A1(n15341), .A2(n11415), .B1(n12716), .B2(n15324), .C1(
        n12718), .C2(n15326), .ZN(n15354) );
  OAI21_X1 U13971 ( .B1(n11416), .B2(n15355), .A(n15354), .ZN(n11583) );
  INV_X1 U13972 ( .A(n11583), .ZN(n11418) );
  AOI22_X1 U13973 ( .A1(n13401), .A2(n15358), .B1(n15428), .B2(
        P3_REG0_REG_5__SCAN_IN), .ZN(n11417) );
  OAI21_X1 U13974 ( .B1(n11418), .B2(n15428), .A(n11417), .ZN(P3_U3405) );
  INV_X1 U13975 ( .A(n11419), .ZN(n11421) );
  OAI222_X1 U13976 ( .A1(n14906), .A2(P1_U3086), .B1(n14544), .B2(n11421), 
        .C1(n11420), .C2(n14542), .ZN(P1_U3337) );
  INV_X1 U13977 ( .A(n13596), .ZN(n13569) );
  OAI222_X1 U13978 ( .A1(n13928), .A2(n13234), .B1(n13920), .B2(n11421), .C1(
        P2_U3088), .C2(n13569), .ZN(P2_U3309) );
  MUX2_X1 U13979 ( .A(n9155), .B(P1_REG1_REG_12__SCAN_IN), .S(n11622), .Z(
        n11422) );
  INV_X1 U13980 ( .A(n11422), .ZN(n11425) );
  OAI21_X1 U13981 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n11427), .A(n11423), 
        .ZN(n11424) );
  OAI21_X1 U13982 ( .B1(n11425), .B2(n11424), .A(n11621), .ZN(n11435) );
  XOR2_X1 U13983 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11622), .Z(n11429) );
  AOI21_X1 U13984 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n11427), .A(n11426), 
        .ZN(n11428) );
  NAND2_X1 U13985 ( .A1(n11428), .A2(n11429), .ZN(n11617) );
  OAI21_X1 U13986 ( .B1(n11429), .B2(n11428), .A(n11617), .ZN(n11430) );
  NAND2_X1 U13987 ( .A1(n11430), .A2(n14903), .ZN(n11432) );
  NOR2_X1 U13988 ( .A1(n13041), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13995) );
  AOI21_X1 U13989 ( .B1(n14860), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n13995), 
        .ZN(n11431) );
  OAI211_X1 U13990 ( .C1(n14907), .C2(n11433), .A(n11432), .B(n11431), .ZN(
        n11434) );
  AOI21_X1 U13991 ( .B1(n14898), .B2(n11435), .A(n11434), .ZN(n11436) );
  INV_X1 U13992 ( .A(n11436), .ZN(P1_U3255) );
  AOI211_X1 U13993 ( .C1(n15212), .C2(n11439), .A(n11438), .B(n11437), .ZN(
        n11445) );
  INV_X1 U13994 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11440) );
  NOR2_X1 U13995 ( .A1(n15242), .A2(n11440), .ZN(n11441) );
  AOI21_X1 U13996 ( .B1(n11884), .B2(n11443), .A(n11441), .ZN(n11442) );
  OAI21_X1 U13997 ( .B1(n11445), .B2(n15240), .A(n11442), .ZN(P2_U3457) );
  AOI22_X1 U13998 ( .A1(n11886), .A2(n11443), .B1(n9959), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11444) );
  OAI21_X1 U13999 ( .B1(n11445), .B2(n9959), .A(n11444), .ZN(P2_U3508) );
  INV_X1 U14000 ( .A(n11446), .ZN(n11747) );
  AOI21_X1 U14001 ( .B1(n11448), .B2(n11447), .A(n12691), .ZN(n11450) );
  NAND2_X1 U14002 ( .A1(n11450), .A2(n11449), .ZN(n11457) );
  AOI21_X1 U14003 ( .B1(n12679), .B2(n11452), .A(n11451), .ZN(n11453) );
  OAI21_X1 U14004 ( .B1(n12296), .B2(n11454), .A(n11453), .ZN(n11455) );
  AOI21_X1 U14005 ( .B1(n12703), .B2(n12715), .A(n11455), .ZN(n11456) );
  OAI211_X1 U14006 ( .C1(n11747), .C2(n12700), .A(n11457), .B(n11456), .ZN(
        P3_U3179) );
  OAI211_X1 U14007 ( .C1(n11461), .C2(n11460), .A(n11459), .B(n15341), .ZN(
        n11463) );
  AOI22_X1 U14008 ( .A1(n15326), .A2(n12717), .B1(n15324), .B2(n12715), .ZN(
        n11462) );
  NAND2_X1 U14009 ( .A1(n11463), .A2(n11462), .ZN(n11749) );
  AOI21_X1 U14010 ( .B1(n15411), .B2(n11752), .A(n11749), .ZN(n11543) );
  INV_X1 U14011 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11464) );
  OAI22_X1 U14012 ( .A1(n11748), .A2(n13392), .B1(n15430), .B2(n11464), .ZN(
        n11465) );
  INV_X1 U14013 ( .A(n11465), .ZN(n11466) );
  OAI21_X1 U14014 ( .B1(n11543), .B2(n15428), .A(n11466), .ZN(P3_U3408) );
  AOI21_X1 U14015 ( .B1(n15169), .B2(n13742), .A(n15170), .ZN(n11475) );
  OAI22_X1 U14016 ( .A1(n15174), .A2(n11469), .B1(n11468), .B2(n13774), .ZN(
        n11473) );
  OR2_X1 U14017 ( .A1(n15174), .A2(n11470), .ZN(n13706) );
  NOR2_X1 U14018 ( .A1(n13706), .A2(n11471), .ZN(n11472) );
  AOI211_X1 U14019 ( .C1(n15174), .C2(P2_REG2_REG_0__SCAN_IN), .A(n11473), .B(
        n11472), .ZN(n11474) );
  OAI21_X1 U14020 ( .B1(n11475), .B2(n9588), .A(n11474), .ZN(P2_U3265) );
  INV_X1 U14021 ( .A(n11476), .ZN(n11646) );
  NOR3_X1 U14022 ( .A1(n11478), .A2(n11477), .A3(n12342), .ZN(n11479) );
  AOI21_X1 U14023 ( .B1(n11646), .B2(n12224), .A(n11479), .ZN(n11487) );
  INV_X1 U14024 ( .A(n11480), .ZN(n11637) );
  NAND2_X1 U14025 ( .A1(n11637), .A2(n12224), .ZN(n11485) );
  AOI22_X1 U14026 ( .A1(n13509), .A2(n13541), .B1(n13510), .B2(n13539), .ZN(
        n11788) );
  OAI22_X1 U14027 ( .A1(n13491), .A2(n11788), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11481), .ZN(n11483) );
  INV_X1 U14028 ( .A(n11887), .ZN(n11794) );
  NOR2_X1 U14029 ( .A1(n11794), .A2(n8883), .ZN(n11482) );
  AOI211_X1 U14030 ( .C1(n13493), .C2(n11792), .A(n11483), .B(n11482), .ZN(
        n11484) );
  OAI211_X1 U14031 ( .C1(n11487), .C2(n11486), .A(n11485), .B(n11484), .ZN(
        P2_U3208) );
  NAND2_X1 U14032 ( .A1(n12710), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11488) );
  OAI21_X1 U14033 ( .B1(n6543), .B2(n12710), .A(n11488), .ZN(P3_U3519) );
  XNOR2_X1 U14034 ( .A(n11490), .B(n11491), .ZN(n15231) );
  AOI21_X1 U14035 ( .B1(n6690), .B2(n11491), .A(n13769), .ZN(n11495) );
  NAND2_X1 U14036 ( .A1(n13509), .A2(n13542), .ZN(n11493) );
  NAND2_X1 U14037 ( .A1(n13510), .A2(n13540), .ZN(n11492) );
  NAND2_X1 U14038 ( .A1(n11493), .A2(n11492), .ZN(n11643) );
  AOI21_X1 U14039 ( .B1(n11495), .B2(n11494), .A(n11643), .ZN(n15234) );
  INV_X1 U14040 ( .A(n15234), .ZN(n11501) );
  AOI21_X1 U14041 ( .B1(n15232), .B2(n11496), .A(n11852), .ZN(n11497) );
  NAND2_X1 U14042 ( .A1(n11497), .A2(n11781), .ZN(n15233) );
  AOI22_X1 U14043 ( .A1(n15149), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11642), 
        .B2(n15163), .ZN(n11499) );
  NAND2_X1 U14044 ( .A1(n15232), .A2(n15170), .ZN(n11498) );
  OAI211_X1 U14045 ( .C1(n15233), .C2(n13747), .A(n11499), .B(n11498), .ZN(
        n11500) );
  AOI21_X1 U14046 ( .B1(n11501), .B2(n11353), .A(n11500), .ZN(n11502) );
  OAI21_X1 U14047 ( .B1(n15231), .B2(n13793), .A(n11502), .ZN(P2_U3255) );
  INV_X1 U14048 ( .A(n9256), .ZN(n11504) );
  OAI222_X1 U14049 ( .A1(n14218), .A2(P1_U3086), .B1(n14544), .B2(n11504), 
        .C1(n11503), .C2(n14542), .ZN(P1_U3336) );
  OAI222_X1 U14050 ( .A1(n13928), .A2(n11505), .B1(n13920), .B2(n11504), .C1(
        n13607), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U14051 ( .A(n11506), .B(n7572), .ZN(n15005) );
  INV_X1 U14052 ( .A(n15005), .ZN(n11523) );
  OAI21_X1 U14053 ( .B1(n11509), .B2(n11508), .A(n11507), .ZN(n11510) );
  NAND2_X1 U14054 ( .A1(n11510), .A2(n14937), .ZN(n11514) );
  OR2_X1 U14055 ( .A1(n11528), .A2(n14268), .ZN(n11512) );
  NAND2_X1 U14056 ( .A1(n14131), .A2(n14052), .ZN(n11511) );
  NAND2_X1 U14057 ( .A1(n11512), .A2(n11511), .ZN(n11666) );
  INV_X1 U14058 ( .A(n11666), .ZN(n11513) );
  NAND2_X1 U14059 ( .A1(n11514), .A2(n11513), .ZN(n15010) );
  NAND2_X1 U14060 ( .A1(n14928), .A2(n15006), .ZN(n11515) );
  NAND2_X1 U14061 ( .A1(n11515), .A2(n14948), .ZN(n11517) );
  OR2_X1 U14062 ( .A1(n11517), .A2(n11516), .ZN(n15007) );
  INV_X1 U14063 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11518) );
  OAI22_X1 U14064 ( .A1(n14427), .A2(n11518), .B1(n11668), .B2(n14940), .ZN(
        n11519) );
  AOI21_X1 U14065 ( .B1(n14417), .B2(n15006), .A(n11519), .ZN(n11520) );
  OAI21_X1 U14066 ( .B1(n15007), .B2(n14334), .A(n11520), .ZN(n11521) );
  AOI21_X1 U14067 ( .B1(n15010), .B2(n14427), .A(n11521), .ZN(n11522) );
  OAI21_X1 U14068 ( .B1(n14432), .B2(n11523), .A(n11522), .ZN(P1_U3286) );
  XNOR2_X1 U14069 ( .A(n11524), .B(n11526), .ZN(n15014) );
  OAI21_X1 U14070 ( .B1(n11527), .B2(n11526), .A(n11525), .ZN(n11529) );
  OAI22_X1 U14071 ( .A1(n11528), .A2(n14085), .B1(n11737), .B2(n14268), .ZN(
        n12006) );
  AOI21_X1 U14072 ( .B1(n11529), .B2(n14937), .A(n12006), .ZN(n15016) );
  INV_X1 U14073 ( .A(n15016), .ZN(n11535) );
  OAI211_X1 U14074 ( .C1(n11530), .C2(n15017), .A(n14948), .B(n11774), .ZN(
        n15015) );
  NAND2_X1 U14075 ( .A1(n14942), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11531) );
  OAI21_X1 U14076 ( .B1(n14940), .B2(n12008), .A(n11531), .ZN(n11532) );
  AOI21_X1 U14077 ( .B1(n12010), .B2(n14417), .A(n11532), .ZN(n11533) );
  OAI21_X1 U14078 ( .B1(n15015), .B2(n14334), .A(n11533), .ZN(n11534) );
  AOI21_X1 U14079 ( .B1(n11535), .B2(n14427), .A(n11534), .ZN(n11536) );
  OAI21_X1 U14080 ( .B1(n14432), .B2(n15014), .A(n11536), .ZN(P1_U3284) );
  NAND2_X1 U14081 ( .A1(n11537), .A2(n13410), .ZN(n11538) );
  OAI211_X1 U14082 ( .C1(n11539), .C2(n13423), .A(n11538), .B(n12558), .ZN(
        P3_U3272) );
  INV_X1 U14083 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n13032) );
  NAND2_X1 U14084 ( .A1(n12381), .A2(P3_U3897), .ZN(n11540) );
  OAI21_X1 U14085 ( .B1(P3_U3897), .B2(n13032), .A(n11540), .ZN(P3_U3521) );
  OAI22_X1 U14086 ( .A1(n13339), .A2(n11748), .B1(n15438), .B2(n7756), .ZN(
        n11541) );
  INV_X1 U14087 ( .A(n11541), .ZN(n11542) );
  OAI21_X1 U14088 ( .B1(n11543), .B2(n15439), .A(n11542), .ZN(P3_U3465) );
  INV_X1 U14089 ( .A(n14682), .ZN(n14361) );
  NAND2_X1 U14090 ( .A1(n11544), .A2(n14361), .ZN(n11545) );
  OAI211_X1 U14091 ( .C1(n14940), .C2(n11876), .A(n11546), .B(n11545), .ZN(
        n11547) );
  MUX2_X1 U14092 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11547), .S(n14427), .Z(
        n11551) );
  OAI22_X1 U14093 ( .A1(n11549), .A2(n14432), .B1(n11548), .B2(n14944), .ZN(
        n11550) );
  OR2_X1 U14094 ( .A1(n11551), .A2(n11550), .ZN(P1_U3285) );
  XNOR2_X1 U14095 ( .A(n11553), .B(n11552), .ZN(n11560) );
  AND2_X1 U14096 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n15273) );
  NOR2_X1 U14097 ( .A1(n12706), .A2(n11554), .ZN(n11555) );
  AOI211_X1 U14098 ( .C1(n12703), .C2(n15325), .A(n15273), .B(n11555), .ZN(
        n11556) );
  OAI21_X1 U14099 ( .B1(n11557), .B2(n12296), .A(n11556), .ZN(n11558) );
  AOI21_X1 U14100 ( .B1(n11705), .B2(n12689), .A(n11558), .ZN(n11559) );
  OAI21_X1 U14101 ( .B1(n11560), .B2(n12691), .A(n11559), .ZN(P3_U3153) );
  OAI22_X1 U14102 ( .A1(n13339), .A2(n11561), .B1(n15438), .B2(n11000), .ZN(
        n11562) );
  AOI21_X1 U14103 ( .B1(n11563), .B2(n15438), .A(n11562), .ZN(n11564) );
  INV_X1 U14104 ( .A(n11564), .ZN(P3_U3462) );
  XNOR2_X1 U14105 ( .A(n11565), .B(n6879), .ZN(n11567) );
  OAI21_X1 U14106 ( .B1(n11567), .B2(n13769), .A(n11566), .ZN(n15210) );
  AOI21_X1 U14107 ( .B1(n15163), .B2(n11568), .A(n15210), .ZN(n11576) );
  XNOR2_X1 U14108 ( .A(n11570), .B(n9840), .ZN(n15207) );
  NOR2_X1 U14109 ( .A1(n13793), .A2(n15207), .ZN(n11573) );
  OAI211_X1 U14110 ( .C1(n11680), .C2(n15209), .A(n13742), .B(n11571), .ZN(
        n15208) );
  OAI22_X1 U14111 ( .A1(n11353), .A2(n10550), .B1(n13747), .B2(n15208), .ZN(
        n11572) );
  AOI211_X1 U14112 ( .C1(n15170), .C2(n11574), .A(n11573), .B(n11572), .ZN(
        n11575) );
  OAI21_X1 U14113 ( .B1(n15174), .B2(n11576), .A(n11575), .ZN(P2_U3262) );
  OAI22_X1 U14114 ( .A1(n13339), .A2(n11577), .B1(n15438), .B2(n11051), .ZN(
        n11578) );
  AOI21_X1 U14115 ( .B1(n11579), .B2(n15438), .A(n11578), .ZN(n11580) );
  INV_X1 U14116 ( .A(n11580), .ZN(P3_U3463) );
  OAI22_X1 U14117 ( .A1(n13339), .A2(n11581), .B1(n15438), .B2(n7668), .ZN(
        n11582) );
  AOI21_X1 U14118 ( .B1(n11583), .B2(n15438), .A(n11582), .ZN(n11584) );
  INV_X1 U14119 ( .A(n11584), .ZN(P3_U3464) );
  INV_X1 U14120 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15267) );
  NOR2_X1 U14121 ( .A1(n15280), .A2(n11587), .ZN(n11588) );
  INV_X1 U14122 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n15351) );
  AOI22_X1 U14123 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11614), .B1(n11812), 
        .B2(n15351), .ZN(n11589) );
  AOI21_X1 U14124 ( .B1(n6699), .B2(n11589), .A(n11798), .ZN(n11616) );
  INV_X1 U14125 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11603) );
  MUX2_X1 U14126 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n15255), .Z(n11801) );
  XNOR2_X1 U14127 ( .A(n11801), .B(n11614), .ZN(n11598) );
  MUX2_X1 U14128 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n15255), .Z(n11591) );
  INV_X1 U14129 ( .A(n11591), .ZN(n11590) );
  NAND2_X1 U14130 ( .A1(n15280), .A2(n11590), .ZN(n11596) );
  XNOR2_X1 U14131 ( .A(n11591), .B(n15280), .ZN(n15277) );
  OR2_X1 U14132 ( .A1(n11593), .A2(n11592), .ZN(n11595) );
  NAND2_X1 U14133 ( .A1(n11595), .A2(n11594), .ZN(n15276) );
  NAND2_X1 U14134 ( .A1(n15277), .A2(n15276), .ZN(n15275) );
  NAND2_X1 U14135 ( .A1(n11596), .A2(n15275), .ZN(n11597) );
  NAND2_X1 U14136 ( .A1(n11598), .A2(n11597), .ZN(n11800) );
  OAI21_X1 U14137 ( .B1(n11598), .B2(n11597), .A(n11800), .ZN(n11599) );
  NAND2_X1 U14138 ( .A1(n15279), .A2(n11599), .ZN(n11602) );
  NOR2_X1 U14139 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11600), .ZN(n11757) );
  INV_X1 U14140 ( .A(n11757), .ZN(n11601) );
  OAI211_X1 U14141 ( .C1(n15287), .C2(n11603), .A(n11602), .B(n11601), .ZN(
        n11613) );
  XNOR2_X1 U14142 ( .A(n15280), .B(n11606), .ZN(n15269) );
  NOR2_X1 U14143 ( .A1(n15280), .A2(n11606), .ZN(n11607) );
  NAND2_X1 U14144 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11812), .ZN(n11608) );
  OAI21_X1 U14145 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n11812), .A(n11608), .ZN(
        n11609) );
  AOI21_X1 U14146 ( .B1(n11610), .B2(n11609), .A(n11811), .ZN(n11611) );
  NOR2_X1 U14147 ( .A1(n11611), .A2(n15298), .ZN(n11612) );
  AOI211_X1 U14148 ( .C1(n15281), .C2(n11614), .A(n11613), .B(n11612), .ZN(
        n11615) );
  OAI21_X1 U14149 ( .B1(n11616), .B2(n15304), .A(n11615), .ZN(P3_U3190) );
  XNOR2_X1 U14150 ( .A(n11896), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n11619) );
  OAI21_X1 U14151 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n11622), .A(n11617), 
        .ZN(n11618) );
  NOR2_X1 U14152 ( .A1(n11618), .A2(n11619), .ZN(n11895) );
  AOI211_X1 U14153 ( .C1(n11619), .C2(n11618), .A(n14868), .B(n11895), .ZN(
        n11629) );
  MUX2_X1 U14154 ( .A(n11620), .B(P1_REG1_REG_13__SCAN_IN), .S(n11896), .Z(
        n11624) );
  NOR2_X1 U14155 ( .A1(n11623), .A2(n11624), .ZN(n11890) );
  AOI211_X1 U14156 ( .C1(n11624), .C2(n11623), .A(n14864), .B(n11890), .ZN(
        n11628) );
  INV_X1 U14157 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14550) );
  NAND2_X1 U14158 ( .A1(n14875), .A2(n11896), .ZN(n11626) );
  NAND2_X1 U14159 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11625)
         );
  OAI211_X1 U14160 ( .C1(n14550), .C2(n14912), .A(n11626), .B(n11625), .ZN(
        n11627) );
  OR3_X1 U14161 ( .A1(n11629), .A2(n11628), .A3(n11627), .ZN(P1_U3256) );
  INV_X1 U14162 ( .A(n11854), .ZN(n11633) );
  NAND2_X1 U14163 ( .A1(n13509), .A2(n13540), .ZN(n11631) );
  NAND2_X1 U14164 ( .A1(n13510), .A2(n13538), .ZN(n11630) );
  NAND2_X1 U14165 ( .A1(n11631), .A2(n11630), .ZN(n11849) );
  NAND2_X1 U14166 ( .A1(n13513), .A2(n11849), .ZN(n11632) );
  NAND2_X1 U14167 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n13563)
         );
  OAI211_X1 U14168 ( .C1(n13515), .C2(n11633), .A(n11632), .B(n13563), .ZN(
        n11639) );
  AOI22_X1 U14169 ( .A1(n11634), .A2(n12224), .B1(n13484), .B2(n13540), .ZN(
        n11636) );
  NOR3_X1 U14170 ( .A1(n11637), .A2(n11636), .A3(n11635), .ZN(n11638) );
  AOI211_X1 U14171 ( .C1(n11855), .C2(n13518), .A(n11639), .B(n11638), .ZN(
        n11640) );
  OAI21_X1 U14172 ( .B1(n11641), .B2(n13520), .A(n11640), .ZN(P2_U3196) );
  INV_X1 U14173 ( .A(n11642), .ZN(n11645) );
  AOI22_X1 U14174 ( .A1(n13513), .A2(n11643), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11644) );
  OAI21_X1 U14175 ( .B1(n11645), .B2(n13515), .A(n11644), .ZN(n11650) );
  AOI211_X1 U14176 ( .C1(n11648), .C2(n11647), .A(n13520), .B(n11646), .ZN(
        n11649) );
  AOI211_X1 U14177 ( .C1(n15232), .C2(n13518), .A(n11650), .B(n11649), .ZN(
        n11651) );
  INV_X1 U14178 ( .A(n11651), .ZN(P2_U3189) );
  XOR2_X1 U14179 ( .A(n11652), .B(n11653), .Z(n11662) );
  NAND2_X1 U14180 ( .A1(n14130), .A2(n14071), .ZN(n11655) );
  NAND2_X1 U14181 ( .A1(n14132), .A2(n14052), .ZN(n11654) );
  NAND2_X1 U14182 ( .A1(n11655), .A2(n11654), .ZN(n14921) );
  INV_X1 U14183 ( .A(n11656), .ZN(n11657) );
  AOI21_X1 U14184 ( .B1(n14097), .B2(n14921), .A(n11657), .ZN(n11660) );
  NAND2_X1 U14185 ( .A1(n11658), .A2(n14103), .ZN(n11659) );
  OAI211_X1 U14186 ( .C1(n14101), .C2(n14922), .A(n11660), .B(n11659), .ZN(
        n11661) );
  AOI21_X1 U14187 ( .B1(n11662), .B2(n14082), .A(n11661), .ZN(n11663) );
  INV_X1 U14188 ( .A(n11663), .ZN(P1_U3239) );
  XNOR2_X1 U14189 ( .A(n11665), .B(n11664), .ZN(n11671) );
  AOI22_X1 U14190 ( .A1(n14097), .A2(n11666), .B1(P1_REG3_REG_7__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11667) );
  OAI21_X1 U14191 ( .B1(n14101), .B2(n11668), .A(n11667), .ZN(n11669) );
  AOI21_X1 U14192 ( .B1(n14103), .B2(n15006), .A(n11669), .ZN(n11670) );
  OAI21_X1 U14193 ( .B1(n11671), .B2(n14106), .A(n11670), .ZN(P1_U3213) );
  XNOR2_X1 U14194 ( .A(n11672), .B(n11673), .ZN(n11675) );
  AOI21_X1 U14195 ( .B1(n11675), .B2(n15161), .A(n11674), .ZN(n15205) );
  XNOR2_X1 U14196 ( .A(n11676), .B(n11677), .ZN(n15201) );
  NAND2_X1 U14197 ( .A1(n15164), .A2(n15199), .ZN(n11678) );
  NAND2_X1 U14198 ( .A1(n11678), .A2(n13742), .ZN(n11679) );
  NOR2_X1 U14199 ( .A1(n11680), .A2(n11679), .ZN(n15198) );
  AOI22_X1 U14200 ( .A1(n15169), .A2(n15198), .B1(n15163), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n11683) );
  NAND2_X1 U14201 ( .A1(n15149), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n11682) );
  OAI211_X1 U14202 ( .C1(n15152), .C2(n11684), .A(n11683), .B(n11682), .ZN(
        n11685) );
  AOI21_X1 U14203 ( .B1(n15168), .B2(n15201), .A(n11685), .ZN(n11686) );
  OAI21_X1 U14204 ( .B1(n15149), .B2(n15205), .A(n11686), .ZN(P2_U3263) );
  INV_X1 U14205 ( .A(n11687), .ZN(n11691) );
  AOI22_X1 U14206 ( .A1(n15170), .A2(n11689), .B1(n15163), .B2(n11688), .ZN(
        n11690) );
  OAI21_X1 U14207 ( .B1(n13747), .B2(n11691), .A(n11690), .ZN(n11694) );
  MUX2_X1 U14208 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11692), .S(n11353), .Z(
        n11693) );
  AOI211_X1 U14209 ( .C1(n15168), .C2(n11695), .A(n11694), .B(n11693), .ZN(
        n11696) );
  INV_X1 U14210 ( .A(n11696), .ZN(P2_U3259) );
  OAI21_X1 U14211 ( .B1(n11698), .B2(n12454), .A(n11697), .ZN(n15412) );
  INV_X1 U14212 ( .A(n15412), .ZN(n11709) );
  INV_X1 U14213 ( .A(n13306), .ZN(n11708) );
  OAI211_X1 U14214 ( .C1(n11701), .C2(n11700), .A(n11699), .B(n15341), .ZN(
        n11703) );
  AOI22_X1 U14215 ( .A1(n15326), .A2(n12716), .B1(n15324), .B2(n15325), .ZN(
        n11702) );
  AND2_X1 U14216 ( .A1(n11703), .A2(n11702), .ZN(n15414) );
  MUX2_X1 U14217 ( .A(n15414), .B(n15267), .S(n15398), .Z(n11707) );
  INV_X1 U14218 ( .A(n13304), .ZN(n15374) );
  AOI22_X1 U14219 ( .A1(n15374), .A2(n15409), .B1(n15395), .B2(n11705), .ZN(
        n11706) );
  OAI211_X1 U14220 ( .C1(n11709), .C2(n11708), .A(n11707), .B(n11706), .ZN(
        P3_U3226) );
  INV_X1 U14221 ( .A(n11710), .ZN(n11717) );
  AOI22_X1 U14222 ( .A1(n15149), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11711), 
        .B2(n15163), .ZN(n11714) );
  NAND2_X1 U14223 ( .A1(n15170), .A2(n11712), .ZN(n11713) );
  OAI211_X1 U14224 ( .C1(n11715), .C2(n13747), .A(n11714), .B(n11713), .ZN(
        n11716) );
  AOI21_X1 U14225 ( .B1(n11717), .B2(n15168), .A(n11716), .ZN(n11718) );
  OAI21_X1 U14226 ( .B1(n15174), .B2(n11719), .A(n11718), .ZN(P2_U3257) );
  OAI21_X1 U14227 ( .B1(n9960), .B2(n8938), .A(n14937), .ZN(n11726) );
  OR2_X1 U14228 ( .A1(n14964), .A2(n11720), .ZN(n11722) );
  AND2_X1 U14229 ( .A1(n11722), .A2(n11721), .ZN(n11729) );
  INV_X1 U14230 ( .A(n11729), .ZN(n11723) );
  XNOR2_X1 U14231 ( .A(n14137), .B(n11723), .ZN(n11724) );
  AOI21_X1 U14232 ( .B1(n11724), .B2(n14937), .A(n14138), .ZN(n11725) );
  AOI21_X1 U14233 ( .B1(n14085), .B2(n11726), .A(n11725), .ZN(n11727) );
  AOI21_X1 U14234 ( .B1(n14071), .B2(n14136), .A(n11727), .ZN(n14965) );
  XNOR2_X1 U14235 ( .A(n9960), .B(n11728), .ZN(n14970) );
  NAND2_X1 U14236 ( .A1(n11729), .A2(n14948), .ZN(n14963) );
  OAI22_X1 U14237 ( .A1(n14334), .A2(n14963), .B1(n11730), .B2(n14940), .ZN(
        n11731) );
  INV_X1 U14238 ( .A(n11731), .ZN(n11733) );
  NAND2_X1 U14239 ( .A1(n14942), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n11732) );
  OAI211_X1 U14240 ( .C1(n14944), .C2(n14964), .A(n11733), .B(n11732), .ZN(
        n11734) );
  AOI21_X1 U14241 ( .B1(n14954), .B2(n14970), .A(n11734), .ZN(n11735) );
  OAI21_X1 U14242 ( .B1(n14942), .B2(n14965), .A(n11735), .ZN(P1_U3292) );
  XNOR2_X1 U14243 ( .A(n11736), .B(n11743), .ZN(n11739) );
  OAI22_X1 U14244 ( .A1(n11738), .A2(n14268), .B1(n11737), .B2(n14085), .ZN(
        n12209) );
  AOI21_X1 U14245 ( .B1(n11739), .B2(n14937), .A(n12209), .ZN(n14836) );
  AOI211_X1 U14246 ( .C1(n11740), .C2(n11775), .A(n14829), .B(n11991), .ZN(
        n14834) );
  NOR2_X1 U14247 ( .A1(n7189), .A2(n14944), .ZN(n11742) );
  OAI22_X1 U14248 ( .A1(n14427), .A2(n11117), .B1(n12206), .B2(n14940), .ZN(
        n11741) );
  AOI211_X1 U14249 ( .C1(n14834), .C2(n14953), .A(n11742), .B(n11741), .ZN(
        n11746) );
  XNOR2_X1 U14250 ( .A(n11744), .B(n11743), .ZN(n14839) );
  NAND2_X1 U14251 ( .A1(n14839), .A2(n14954), .ZN(n11745) );
  OAI211_X1 U14252 ( .C1(n14836), .C2(n14942), .A(n11746), .B(n11745), .ZN(
        P1_U3282) );
  OAI22_X1 U14253 ( .A1(n13304), .A2(n11748), .B1(n11747), .B2(n15376), .ZN(
        n11751) );
  MUX2_X1 U14254 ( .A(n11749), .B(P3_REG2_REG_6__SCAN_IN), .S(n15398), .Z(
        n11750) );
  AOI211_X1 U14255 ( .C1(n13306), .C2(n11752), .A(n11751), .B(n11750), .ZN(
        n11753) );
  INV_X1 U14256 ( .A(n11753), .ZN(P3_U3227) );
  XNOR2_X1 U14257 ( .A(n11755), .B(n11754), .ZN(n11761) );
  NOR2_X1 U14258 ( .A1(n12706), .A2(n15347), .ZN(n11756) );
  AOI211_X1 U14259 ( .C1(n12698), .C2(n12715), .A(n11757), .B(n11756), .ZN(
        n11758) );
  OAI21_X1 U14260 ( .B1(n15339), .B2(n12685), .A(n11758), .ZN(n11759) );
  AOI21_X1 U14261 ( .B1(n15348), .B2(n12689), .A(n11759), .ZN(n11760) );
  OAI21_X1 U14262 ( .B1(n11761), .B2(n12691), .A(n11760), .ZN(P3_U3161) );
  INV_X1 U14263 ( .A(n11762), .ZN(n11765) );
  OAI222_X1 U14264 ( .A1(P1_U3086), .A2(n11764), .B1(n14544), .B2(n11765), 
        .C1(n11763), .C2(n14542), .ZN(P1_U3335) );
  OAI222_X1 U14265 ( .A1(n13928), .A2(n11767), .B1(P2_U3088), .B2(n11766), 
        .C1(n13920), .C2(n11765), .ZN(P2_U3307) );
  AOI21_X1 U14266 ( .B1(n11768), .B2(n11773), .A(n14917), .ZN(n11771) );
  NOR2_X1 U14267 ( .A1(n11769), .A2(n14085), .ZN(n12151) );
  AOI21_X1 U14268 ( .B1(n11771), .B2(n11770), .A(n12151), .ZN(n15024) );
  XNOR2_X1 U14269 ( .A(n11772), .B(n11773), .ZN(n15028) );
  AOI21_X1 U14270 ( .B1(n11774), .B2(n15022), .A(n14829), .ZN(n11776) );
  AOI22_X1 U14271 ( .A1(n11776), .A2(n11775), .B1(n14071), .B2(n14126), .ZN(
        n15023) );
  OAI22_X1 U14272 ( .A1(n14427), .A2(n10807), .B1(n12150), .B2(n14940), .ZN(
        n11777) );
  AOI21_X1 U14273 ( .B1(n15022), .B2(n14417), .A(n11777), .ZN(n11778) );
  OAI21_X1 U14274 ( .B1(n15023), .B2(n14334), .A(n11778), .ZN(n11779) );
  AOI21_X1 U14275 ( .B1(n15028), .B2(n14954), .A(n11779), .ZN(n11780) );
  OAI21_X1 U14276 ( .B1(n15024), .B2(n14942), .A(n11780), .ZN(P1_U3283) );
  NAND2_X1 U14277 ( .A1(n11887), .A2(n11781), .ZN(n11782) );
  NAND2_X1 U14278 ( .A1(n11782), .A2(n13742), .ZN(n11783) );
  NOR2_X1 U14279 ( .A1(n11853), .A2(n11783), .ZN(n11882) );
  INV_X1 U14280 ( .A(n11784), .ZN(n11785) );
  AOI21_X1 U14281 ( .B1(n11787), .B2(n11786), .A(n11785), .ZN(n11789) );
  OAI21_X1 U14282 ( .B1(n11789), .B2(n13769), .A(n11788), .ZN(n11881) );
  AOI21_X1 U14283 ( .B1(n11882), .B2(n13607), .A(n11881), .ZN(n11797) );
  XNOR2_X1 U14284 ( .A(n11791), .B(n11790), .ZN(n11883) );
  AOI22_X1 U14285 ( .A1(n15174), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11792), 
        .B2(n15163), .ZN(n11793) );
  OAI21_X1 U14286 ( .B1(n11794), .B2(n15152), .A(n11793), .ZN(n11795) );
  AOI21_X1 U14287 ( .B1(n11883), .B2(n15168), .A(n11795), .ZN(n11796) );
  OAI21_X1 U14288 ( .B1(n11797), .B2(n15149), .A(n11796), .ZN(P2_U3254) );
  INV_X1 U14289 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15333) );
  XNOR2_X1 U14290 ( .A(n11829), .B(n11825), .ZN(n11799) );
  AOI21_X1 U14291 ( .B1(n15333), .B2(n11799), .A(n11826), .ZN(n11818) );
  OAI21_X1 U14292 ( .B1(n11801), .B2(n11812), .A(n11800), .ZN(n11804) );
  MUX2_X1 U14293 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n15255), .Z(n11802) );
  NAND2_X1 U14294 ( .A1(n11802), .A2(n7302), .ZN(n11805) );
  NAND2_X1 U14295 ( .A1(n11804), .A2(n11805), .ZN(n11835) );
  INV_X1 U14296 ( .A(n11835), .ZN(n11807) );
  INV_X1 U14297 ( .A(n11802), .ZN(n11803) );
  NAND2_X1 U14298 ( .A1(n11803), .A2(n11829), .ZN(n11836) );
  AOI21_X1 U14299 ( .B1(n11836), .B2(n11805), .A(n11804), .ZN(n11806) );
  AOI21_X1 U14300 ( .B1(n11807), .B2(n11836), .A(n11806), .ZN(n11810) );
  NAND2_X1 U14301 ( .A1(n15274), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11809) );
  AND2_X1 U14302 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11913) );
  INV_X1 U14303 ( .A(n11913), .ZN(n11808) );
  OAI211_X1 U14304 ( .C1(n11810), .C2(n15296), .A(n11809), .B(n11808), .ZN(
        n11816) );
  AOI21_X1 U14305 ( .B1(n7805), .B2(n11813), .A(n11830), .ZN(n11814) );
  NOR2_X1 U14306 ( .A1(n11814), .A2(n15298), .ZN(n11815) );
  AOI211_X1 U14307 ( .C1(n15281), .C2(n11829), .A(n11816), .B(n11815), .ZN(
        n11817) );
  OAI21_X1 U14308 ( .B1(n11818), .B2(n15304), .A(n11817), .ZN(P3_U3191) );
  INV_X1 U14309 ( .A(n11819), .ZN(n11823) );
  OAI222_X1 U14310 ( .A1(n13928), .A2(n11821), .B1(n13920), .B2(n11823), .C1(
        n11820), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U14311 ( .A1(n11824), .A2(P1_U3086), .B1(n14544), .B2(n11823), 
        .C1(n11822), .C2(n14542), .ZN(P1_U3334) );
  INV_X1 U14312 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12041) );
  MUX2_X1 U14313 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n12041), .S(n12042), .Z(
        n11828) );
  INV_X1 U14314 ( .A(n12044), .ZN(n11827) );
  AOI21_X1 U14315 ( .B1(n6698), .B2(n11828), .A(n11827), .ZN(n11845) );
  MUX2_X1 U14316 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n12028), .S(n12042), .Z(
        n11831) );
  OAI21_X1 U14317 ( .B1(n6841), .B2(n6840), .A(n12030), .ZN(n11843) );
  INV_X1 U14318 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11832) );
  NOR2_X1 U14319 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11832), .ZN(n11940) );
  AOI21_X1 U14320 ( .B1(n15274), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11940), 
        .ZN(n11840) );
  MUX2_X1 U14321 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n15255), .Z(n11833) );
  NOR2_X1 U14322 ( .A1(n11833), .A2(n11841), .ZN(n12037) );
  AOI21_X1 U14323 ( .B1(n11833), .B2(n11841), .A(n12037), .ZN(n11834) );
  INV_X1 U14324 ( .A(n11834), .ZN(n11837) );
  AOI21_X1 U14325 ( .B1(n11836), .B2(n11835), .A(n11837), .ZN(n12036) );
  AND3_X1 U14326 ( .A1(n11837), .A2(n11836), .A3(n11835), .ZN(n11838) );
  OAI21_X1 U14327 ( .B1(n12036), .B2(n11838), .A(n15279), .ZN(n11839) );
  OAI211_X1 U14328 ( .C1(n15290), .C2(n11841), .A(n11840), .B(n11839), .ZN(
        n11842) );
  AOI21_X1 U14329 ( .B1(n11843), .B2(n15252), .A(n11842), .ZN(n11844) );
  OAI21_X1 U14330 ( .B1(n11845), .B2(n15304), .A(n11844), .ZN(P3_U3192) );
  XOR2_X1 U14331 ( .A(n11847), .B(n11846), .Z(n14790) );
  AOI21_X1 U14332 ( .B1(n11848), .B2(n11847), .A(n13769), .ZN(n11851) );
  AOI21_X1 U14333 ( .B1(n11851), .B2(n11850), .A(n11849), .ZN(n14792) );
  INV_X1 U14334 ( .A(n14792), .ZN(n11859) );
  OAI211_X1 U14335 ( .C1(n14793), .C2(n11853), .A(n13742), .B(n12014), .ZN(
        n14791) );
  AOI22_X1 U14336 ( .A1(n15149), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11854), 
        .B2(n15163), .ZN(n11857) );
  NAND2_X1 U14337 ( .A1(n11855), .A2(n15170), .ZN(n11856) );
  OAI211_X1 U14338 ( .C1(n14791), .C2(n13747), .A(n11857), .B(n11856), .ZN(
        n11858) );
  AOI21_X1 U14339 ( .B1(n11859), .B2(n11353), .A(n11858), .ZN(n11860) );
  OAI21_X1 U14340 ( .B1(n13793), .B2(n14790), .A(n11860), .ZN(P2_U3253) );
  INV_X1 U14341 ( .A(n14782), .ZN(n11870) );
  AOI211_X1 U14342 ( .C1(n11862), .C2(n11861), .A(n13520), .B(n12306), .ZN(
        n11863) );
  INV_X1 U14343 ( .A(n11863), .ZN(n11869) );
  NAND2_X1 U14344 ( .A1(n13509), .A2(n13539), .ZN(n11865) );
  NAND2_X1 U14345 ( .A1(n13510), .A2(n13537), .ZN(n11864) );
  AND2_X1 U14346 ( .A1(n11865), .A2(n11864), .ZN(n12023) );
  INV_X1 U14347 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11866) );
  OAI22_X1 U14348 ( .A1(n13491), .A2(n12023), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11866), .ZN(n11867) );
  AOI21_X1 U14349 ( .B1(n12017), .B2(n13493), .A(n11867), .ZN(n11868) );
  OAI211_X1 U14350 ( .C1(n11870), .C2(n8883), .A(n11869), .B(n11868), .ZN(
        P2_U3206) );
  AOI21_X1 U14351 ( .B1(n11872), .B2(n11871), .A(n6693), .ZN(n11880) );
  NAND2_X1 U14352 ( .A1(n14097), .A2(n11873), .ZN(n11874) );
  OAI211_X1 U14353 ( .C1(n14101), .C2(n11876), .A(n11875), .B(n11874), .ZN(
        n11877) );
  AOI21_X1 U14354 ( .B1(n14103), .B2(n11878), .A(n11877), .ZN(n11879) );
  OAI21_X1 U14355 ( .B1(n11880), .B2(n14106), .A(n11879), .ZN(P1_U3221) );
  AOI211_X1 U14356 ( .C1(n15212), .C2(n11883), .A(n11882), .B(n11881), .ZN(
        n11889) );
  AOI22_X1 U14357 ( .A1(n11887), .A2(n11884), .B1(n15240), .B2(
        P2_REG0_REG_11__SCAN_IN), .ZN(n11885) );
  OAI21_X1 U14358 ( .B1(n11889), .B2(n15240), .A(n11885), .ZN(P2_U3463) );
  INV_X1 U14359 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U14360 ( .A1(n11887), .A2(n11886), .B1(n9959), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11888) );
  OAI21_X1 U14361 ( .B1(n11889), .B2(n9959), .A(n11888), .ZN(P2_U3510) );
  MUX2_X1 U14362 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11891), .S(n12062), .Z(
        n11892) );
  NAND2_X1 U14363 ( .A1(n11893), .A2(n11892), .ZN(n12061) );
  OAI21_X1 U14364 ( .B1(n11893), .B2(n11892), .A(n12061), .ZN(n11903) );
  INV_X1 U14365 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14640) );
  NAND2_X1 U14366 ( .A1(n14875), .A2(n12062), .ZN(n11894) );
  NAND2_X1 U14367 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13944)
         );
  OAI211_X1 U14368 ( .C1(n14640), .C2(n14912), .A(n11894), .B(n13944), .ZN(
        n11902) );
  INV_X1 U14369 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11897) );
  MUX2_X1 U14370 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11897), .S(n12062), .Z(
        n11898) );
  INV_X1 U14371 ( .A(n11898), .ZN(n11899) );
  AOI211_X1 U14372 ( .C1(n11900), .C2(n11899), .A(n14868), .B(n12055), .ZN(
        n11901) );
  AOI211_X1 U14373 ( .C1(n14898), .C2(n11903), .A(n11902), .B(n11901), .ZN(
        n11904) );
  INV_X1 U14374 ( .A(n11904), .ZN(P1_U3257) );
  INV_X1 U14375 ( .A(n11905), .ZN(n11907) );
  OAI222_X1 U14376 ( .A1(n11908), .A2(P3_U3151), .B1(n13419), .B2(n11907), 
        .C1(n11906), .C2(n13423), .ZN(P3_U3271) );
  INV_X1 U14377 ( .A(n11935), .ZN(n11909) );
  AOI21_X1 U14378 ( .B1(n11911), .B2(n11910), .A(n11909), .ZN(n11917) );
  NOR2_X1 U14379 ( .A1(n12706), .A2(n12458), .ZN(n11912) );
  AOI211_X1 U14380 ( .C1(n12698), .C2(n15325), .A(n11913), .B(n11912), .ZN(
        n11914) );
  OAI21_X1 U14381 ( .B1(n14740), .B2(n12685), .A(n11914), .ZN(n11915) );
  AOI21_X1 U14382 ( .B1(n15331), .B2(n12689), .A(n11915), .ZN(n11916) );
  OAI21_X1 U14383 ( .B1(n11917), .B2(n12691), .A(n11916), .ZN(P3_U3171) );
  XNOR2_X1 U14384 ( .A(n11918), .B(n11922), .ZN(n11920) );
  OAI22_X1 U14385 ( .A1(n12107), .A2(n13468), .B1(n13469), .B2(n11919), .ZN(
        n12309) );
  AOI21_X1 U14386 ( .B1(n11920), .B2(n15161), .A(n12309), .ZN(n14777) );
  XNOR2_X1 U14387 ( .A(n11922), .B(n11921), .ZN(n14780) );
  INV_X1 U14388 ( .A(n12015), .ZN(n11924) );
  OAI211_X1 U14389 ( .C1(n14776), .C2(n11924), .A(n13742), .B(n12098), .ZN(
        n14775) );
  AOI22_X1 U14390 ( .A1(n15149), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11925), 
        .B2(n15163), .ZN(n11928) );
  NAND2_X1 U14391 ( .A1(n11926), .A2(n15170), .ZN(n11927) );
  OAI211_X1 U14392 ( .C1(n14775), .C2(n13747), .A(n11928), .B(n11927), .ZN(
        n11929) );
  AOI21_X1 U14393 ( .B1(n14780), .B2(n15168), .A(n11929), .ZN(n11930) );
  OAI21_X1 U14394 ( .B1(n14777), .B2(n15174), .A(n11930), .ZN(P2_U3251) );
  INV_X1 U14395 ( .A(n11931), .ZN(n11932) );
  OAI222_X1 U14396 ( .A1(n11933), .A2(P3_U3151), .B1(n13419), .B2(n11932), 
        .C1(n13160), .C2(n13423), .ZN(P3_U3270) );
  INV_X1 U14397 ( .A(n15315), .ZN(n11943) );
  AND2_X1 U14398 ( .A1(n11935), .A2(n11934), .ZN(n11938) );
  OAI211_X1 U14399 ( .C1(n11938), .C2(n11937), .A(n12696), .B(n11936), .ZN(
        n11942) );
  INV_X1 U14400 ( .A(n15314), .ZN(n12464) );
  OAI22_X1 U14401 ( .A1(n12685), .A2(n14728), .B1(n12706), .B2(n12464), .ZN(
        n11939) );
  AOI211_X1 U14402 ( .C1(n12698), .C2(n15310), .A(n11940), .B(n11939), .ZN(
        n11941) );
  OAI211_X1 U14403 ( .C1(n11943), .C2(n12700), .A(n11942), .B(n11941), .ZN(
        P3_U3157) );
  INV_X1 U14404 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11945) );
  NAND2_X1 U14405 ( .A1(n13573), .A2(n11945), .ZN(n11944) );
  OAI21_X1 U14406 ( .B1(n13573), .B2(n11945), .A(n11944), .ZN(n11946) );
  INV_X1 U14407 ( .A(n11946), .ZN(n11956) );
  INV_X1 U14408 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11947) );
  MUX2_X1 U14409 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11947), .S(n13560), .Z(
        n13556) );
  OAI21_X1 U14410 ( .B1(n11960), .B2(P2_REG2_REG_9__SCAN_IN), .A(n11948), .ZN(
        n15072) );
  INV_X1 U14411 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11949) );
  MUX2_X1 U14412 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n11949), .S(n15076), .Z(
        n11950) );
  INV_X1 U14413 ( .A(n11950), .ZN(n15073) );
  NOR2_X1 U14414 ( .A1(n15072), .A2(n15073), .ZN(n15071) );
  INV_X1 U14415 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11951) );
  MUX2_X1 U14416 ( .A(n11951), .B(P2_REG2_REG_11__SCAN_IN), .S(n15089), .Z(
        n11952) );
  INV_X1 U14417 ( .A(n11952), .ZN(n15084) );
  OR2_X1 U14418 ( .A1(n13560), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11953) );
  NAND2_X1 U14419 ( .A1(n13555), .A2(n11953), .ZN(n11955) );
  INV_X1 U14420 ( .A(n13575), .ZN(n11954) );
  AOI211_X1 U14421 ( .C1(n11956), .C2(n11955), .A(n11954), .B(n15120), .ZN(
        n11971) );
  INV_X1 U14422 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14789) );
  NOR2_X1 U14423 ( .A1(n13573), .A2(n14789), .ZN(n11957) );
  AOI21_X1 U14424 ( .B1(n13573), .B2(n14789), .A(n11957), .ZN(n11964) );
  INV_X1 U14425 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11958) );
  MUX2_X1 U14426 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11958), .S(n13560), .Z(
        n13553) );
  OAI21_X1 U14427 ( .B1(n11960), .B2(P2_REG1_REG_9__SCAN_IN), .A(n11959), .ZN(
        n15069) );
  INV_X1 U14428 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11961) );
  MUX2_X1 U14429 ( .A(n11961), .B(P2_REG1_REG_10__SCAN_IN), .S(n15076), .Z(
        n15070) );
  NOR2_X1 U14430 ( .A1(n15069), .A2(n15070), .ZN(n15068) );
  MUX2_X1 U14431 ( .A(n11962), .B(P2_REG1_REG_11__SCAN_IN), .S(n15089), .Z(
        n15081) );
  OAI21_X1 U14432 ( .B1(n13560), .B2(P2_REG1_REG_12__SCAN_IN), .A(n13552), 
        .ZN(n11963) );
  AOI211_X1 U14433 ( .C1(n11964), .C2(n11963), .A(n13565), .B(n15135), .ZN(
        n11970) );
  NAND2_X1 U14434 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n11966)
         );
  NAND2_X1 U14435 ( .A1(n15056), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n11965) );
  OAI211_X1 U14436 ( .C1(n11968), .C2(n11967), .A(n11966), .B(n11965), .ZN(
        n11969) );
  OR3_X1 U14437 ( .A1(n11971), .A2(n11970), .A3(n11969), .ZN(P2_U3227) );
  XNOR2_X1 U14438 ( .A(n11973), .B(n11972), .ZN(n14826) );
  XNOR2_X1 U14439 ( .A(n11974), .B(n11975), .ZN(n11976) );
  NAND2_X1 U14440 ( .A1(n11976), .A2(n14937), .ZN(n11979) );
  NAND2_X1 U14441 ( .A1(n14123), .A2(n14071), .ZN(n11978) );
  NAND2_X1 U14442 ( .A1(n14125), .A2(n14052), .ZN(n11977) );
  AND2_X1 U14443 ( .A1(n11978), .A2(n11977), .ZN(n14047) );
  NAND2_X1 U14444 ( .A1(n11979), .A2(n14047), .ZN(n14833) );
  NAND2_X1 U14445 ( .A1(n14827), .A2(n11990), .ZN(n11981) );
  NAND2_X1 U14446 ( .A1(n12079), .A2(n11981), .ZN(n14830) );
  OAI22_X1 U14447 ( .A1(n14830), .A2(n14682), .B1(n14046), .B2(n14940), .ZN(
        n11982) );
  OAI21_X1 U14448 ( .B1(n14833), .B2(n11982), .A(n14427), .ZN(n11984) );
  AOI22_X1 U14449 ( .A1(n14827), .A2(n14417), .B1(n14942), .B2(
        P1_REG2_REG_13__SCAN_IN), .ZN(n11983) );
  OAI211_X1 U14450 ( .C1(n14432), .C2(n14826), .A(n11984), .B(n11983), .ZN(
        P1_U3280) );
  INV_X1 U14451 ( .A(n11985), .ZN(n11986) );
  OAI222_X1 U14452 ( .A1(n13928), .A2(n11987), .B1(n13920), .B2(n11986), .C1(
        n9586), .C2(P2_U3088), .ZN(P2_U3305) );
  XNOR2_X1 U14453 ( .A(n11988), .B(n11989), .ZN(n14675) );
  OAI21_X1 U14454 ( .B1(n13999), .B2(n11991), .A(n11990), .ZN(n14683) );
  OAI22_X1 U14455 ( .A1(n14683), .A2(n14829), .B1(n13999), .B2(n15025), .ZN(
        n11998) );
  XNOR2_X1 U14456 ( .A(n11992), .B(n11993), .ZN(n11997) );
  NAND2_X1 U14457 ( .A1(n14124), .A2(n14071), .ZN(n11995) );
  NAND2_X1 U14458 ( .A1(n14126), .A2(n14052), .ZN(n11994) );
  NAND2_X1 U14459 ( .A1(n11995), .A2(n11994), .ZN(n13996) );
  INV_X1 U14460 ( .A(n13996), .ZN(n11996) );
  OAI21_X1 U14461 ( .B1(n11997), .B2(n14917), .A(n11996), .ZN(n14685) );
  AOI211_X1 U14462 ( .C1(n14675), .C2(n14442), .A(n11998), .B(n14685), .ZN(
        n12001) );
  NAND2_X1 U14463 ( .A1(n15029), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11999) );
  OAI21_X1 U14464 ( .B1(n12001), .B2(n15029), .A(n11999), .ZN(P1_U3495) );
  NAND2_X1 U14465 ( .A1(n15043), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n12000) );
  OAI21_X1 U14466 ( .B1(n12001), .B2(n15043), .A(n12000), .ZN(P1_U3540) );
  XNOR2_X1 U14467 ( .A(n12004), .B(n12003), .ZN(n12012) );
  AOI21_X1 U14468 ( .B1(n12006), .B2(n14097), .A(n12005), .ZN(n12007) );
  OAI21_X1 U14469 ( .B1(n14101), .B2(n12008), .A(n12007), .ZN(n12009) );
  AOI21_X1 U14470 ( .B1(n12010), .B2(n14103), .A(n12009), .ZN(n12011) );
  OAI21_X1 U14471 ( .B1(n12012), .B2(n14106), .A(n12011), .ZN(P1_U3231) );
  XNOR2_X1 U14472 ( .A(n12013), .B(n12021), .ZN(n14785) );
  AOI21_X1 U14473 ( .B1(n12014), .B2(n14782), .A(n11852), .ZN(n12016) );
  NAND2_X1 U14474 ( .A1(n12016), .A2(n12015), .ZN(n14784) );
  AOI22_X1 U14475 ( .A1(n15149), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12017), 
        .B2(n15163), .ZN(n12019) );
  NAND2_X1 U14476 ( .A1(n14782), .A2(n15170), .ZN(n12018) );
  OAI211_X1 U14477 ( .C1(n14784), .C2(n13747), .A(n12019), .B(n12018), .ZN(
        n12026) );
  OAI211_X1 U14478 ( .C1(n12022), .C2(n12021), .A(n12020), .B(n15161), .ZN(
        n12024) );
  AND2_X1 U14479 ( .A1(n12024), .A2(n12023), .ZN(n14788) );
  NOR2_X1 U14480 ( .A1(n14788), .A2(n15149), .ZN(n12025) );
  AOI211_X1 U14481 ( .C1(n14785), .C2(n15168), .A(n12026), .B(n12025), .ZN(
        n12027) );
  INV_X1 U14482 ( .A(n12027), .ZN(P2_U3252) );
  OR2_X1 U14483 ( .A1(n12042), .A2(n12028), .ZN(n12029) );
  NAND2_X1 U14484 ( .A1(n12755), .A2(n12033), .ZN(n12032) );
  OAI21_X1 U14485 ( .B1(n12755), .B2(n12033), .A(n12032), .ZN(n12034) );
  OAI21_X1 U14486 ( .B1(n7290), .B2(n12034), .A(n12757), .ZN(n12035) );
  NAND2_X1 U14487 ( .A1(n12035), .A2(n15252), .ZN(n12054) );
  MUX2_X1 U14488 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n15255), .Z(n12038) );
  NOR2_X1 U14489 ( .A1(n12038), .A2(n15289), .ZN(n12040) );
  AOI21_X1 U14490 ( .B1(n12038), .B2(n15289), .A(n12040), .ZN(n12039) );
  INV_X1 U14491 ( .A(n12039), .ZN(n15295) );
  MUX2_X1 U14492 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n15255), .Z(n12745) );
  XNOR2_X1 U14493 ( .A(n12745), .B(n12755), .ZN(n12746) );
  XNOR2_X1 U14494 ( .A(n12747), .B(n12746), .ZN(n12052) );
  INV_X1 U14495 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14552) );
  OR2_X1 U14496 ( .A1(n12042), .A2(n12041), .ZN(n12043) );
  NOR2_X1 U14497 ( .A1(n12045), .A2(n12046), .ZN(n12047) );
  INV_X1 U14498 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n15286) );
  NAND2_X1 U14499 ( .A1(n12755), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12742) );
  OAI21_X1 U14500 ( .B1(n12755), .B2(P3_REG2_REG_12__SCAN_IN), .A(n12742), 
        .ZN(n12740) );
  XNOR2_X1 U14501 ( .A(n12741), .B(n12740), .ZN(n12048) );
  NAND2_X1 U14502 ( .A1(n15254), .A2(n12048), .ZN(n12050) );
  INV_X1 U14503 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12049) );
  OR2_X1 U14504 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12049), .ZN(n12232) );
  OAI211_X1 U14505 ( .C1(n14552), .C2(n15287), .A(n12050), .B(n12232), .ZN(
        n12051) );
  AOI21_X1 U14506 ( .B1(n15279), .B2(n12052), .A(n12051), .ZN(n12053) );
  OAI211_X1 U14507 ( .C1(n15290), .C2(n12755), .A(n12054), .B(n12053), .ZN(
        P3_U3194) );
  NAND2_X1 U14508 ( .A1(n12056), .A2(n12125), .ZN(n14199) );
  OAI21_X1 U14509 ( .B1(n12056), .B2(n12125), .A(n14199), .ZN(n12060) );
  NAND2_X1 U14510 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14099)
         );
  NAND2_X1 U14511 ( .A1(n14860), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n12057) );
  OAI211_X1 U14512 ( .C1(n14907), .C2(n12058), .A(n14099), .B(n12057), .ZN(
        n12059) );
  AOI21_X1 U14513 ( .B1(n12060), .B2(n14903), .A(n12059), .ZN(n12066) );
  OAI21_X1 U14514 ( .B1(n12062), .B2(P1_REG1_REG_14__SCAN_IN), .A(n12061), 
        .ZN(n14206) );
  XNOR2_X1 U14515 ( .A(n14206), .B(n14208), .ZN(n12063) );
  INV_X1 U14516 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14818) );
  NAND2_X1 U14517 ( .A1(n12063), .A2(n14818), .ZN(n14207) );
  OAI21_X1 U14518 ( .B1(n12063), .B2(n14818), .A(n14207), .ZN(n12064) );
  NAND2_X1 U14519 ( .A1(n12064), .A2(n14898), .ZN(n12065) );
  NAND2_X1 U14520 ( .A1(n12066), .A2(n12065), .ZN(P1_U3258) );
  INV_X1 U14521 ( .A(n12070), .ZN(n12069) );
  NAND2_X1 U14522 ( .A1(n13922), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12068) );
  OAI211_X1 U14523 ( .C1(n12069), .C2(n13920), .A(n12068), .B(n12067), .ZN(
        P2_U3304) );
  NAND2_X1 U14524 ( .A1(n12070), .A2(n14536), .ZN(n12072) );
  OAI211_X1 U14525 ( .C1(n12073), .C2(n14542), .A(n12072), .B(n12071), .ZN(
        P1_U3332) );
  INV_X1 U14526 ( .A(n12074), .ZN(n12075) );
  OAI222_X1 U14527 ( .A1(P3_U3151), .A2(n12077), .B1(n13423), .B2(n12076), 
        .C1(n13419), .C2(n12075), .ZN(P3_U3269) );
  INV_X1 U14528 ( .A(n12078), .ZN(n12126) );
  AOI211_X1 U14529 ( .C1(n14820), .C2(n12079), .A(n14829), .B(n12126), .ZN(
        n14823) );
  XNOR2_X1 U14530 ( .A(n12080), .B(n12086), .ZN(n12083) );
  OAI22_X1 U14531 ( .A1(n12081), .A2(n14085), .B1(n12161), .B2(n14268), .ZN(
        n13942) );
  INV_X1 U14532 ( .A(n13942), .ZN(n12082) );
  OAI21_X1 U14533 ( .B1(n12083), .B2(n14917), .A(n12082), .ZN(n14824) );
  AOI21_X1 U14534 ( .B1(n14823), .B2(n14218), .A(n14824), .ZN(n12090) );
  OAI22_X1 U14535 ( .A1(n14427), .A2(n11897), .B1(n13945), .B2(n14940), .ZN(
        n12084) );
  AOI21_X1 U14536 ( .B1(n14820), .B2(n14417), .A(n12084), .ZN(n12089) );
  NAND2_X1 U14537 ( .A1(n12087), .A2(n12086), .ZN(n14819) );
  NAND3_X1 U14538 ( .A1(n12085), .A2(n14819), .A3(n14954), .ZN(n12088) );
  OAI211_X1 U14539 ( .C1(n12090), .C2(n14942), .A(n12089), .B(n12088), .ZN(
        P1_U3279) );
  XOR2_X1 U14540 ( .A(n12092), .B(n12091), .Z(n12181) );
  XNOR2_X1 U14541 ( .A(n12093), .B(n12092), .ZN(n12094) );
  NOR2_X1 U14542 ( .A1(n12094), .A2(n13769), .ZN(n12184) );
  NAND2_X1 U14543 ( .A1(n13535), .A2(n13510), .ZN(n12096) );
  NAND2_X1 U14544 ( .A1(n13509), .A2(n13537), .ZN(n12095) );
  NAND2_X1 U14545 ( .A1(n12096), .A2(n12095), .ZN(n12182) );
  OAI21_X1 U14546 ( .B1(n12184), .B2(n12182), .A(n11353), .ZN(n12103) );
  INV_X1 U14547 ( .A(n12135), .ZN(n12097) );
  AOI211_X1 U14548 ( .C1(n12109), .C2(n12098), .A(n11852), .B(n12097), .ZN(
        n12183) );
  INV_X1 U14549 ( .A(n12112), .ZN(n12099) );
  AOI22_X1 U14550 ( .A1(n15149), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12099), 
        .B2(n15163), .ZN(n12100) );
  OAI21_X1 U14551 ( .B1(n9944), .B2(n15152), .A(n12100), .ZN(n12101) );
  AOI21_X1 U14552 ( .B1(n12183), .B2(n15169), .A(n12101), .ZN(n12102) );
  OAI211_X1 U14553 ( .C1(n12181), .C2(n13793), .A(n12103), .B(n12102), .ZN(
        P2_U3250) );
  INV_X1 U14554 ( .A(n12104), .ZN(n12603) );
  AOI22_X1 U14555 ( .A1(n12105), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n13922), .ZN(n12106) );
  OAI21_X1 U14556 ( .B1(n12603), .B2(n13920), .A(n12106), .ZN(P2_U3303) );
  OAI22_X1 U14557 ( .A1(n12108), .A2(n13520), .B1(n12107), .B2(n12342), .ZN(
        n12115) );
  NAND2_X1 U14558 ( .A1(n12109), .A2(n13518), .ZN(n12111) );
  AOI22_X1 U14559 ( .A1(n13513), .A2(n12182), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12110) );
  OAI211_X1 U14560 ( .C1(n13515), .C2(n12112), .A(n12111), .B(n12110), .ZN(
        n12113) );
  AOI21_X1 U14561 ( .B1(n12115), .B2(n12114), .A(n12113), .ZN(n12116) );
  INV_X1 U14562 ( .A(n12116), .ZN(P2_U3213) );
  INV_X1 U14563 ( .A(n12117), .ZN(n12118) );
  AOI21_X1 U14564 ( .B1(n12121), .B2(n12119), .A(n12118), .ZN(n14810) );
  XNOR2_X1 U14565 ( .A(n12120), .B(n12121), .ZN(n12122) );
  NOR2_X1 U14566 ( .A1(n12122), .A2(n14917), .ZN(n14815) );
  OR2_X1 U14567 ( .A1(n14011), .A2(n14268), .ZN(n12124) );
  NAND2_X1 U14568 ( .A1(n14123), .A2(n14052), .ZN(n12123) );
  NAND2_X1 U14569 ( .A1(n12124), .A2(n12123), .ZN(n14811) );
  OAI21_X1 U14570 ( .B1(n14815), .B2(n14811), .A(n14427), .ZN(n12130) );
  OAI22_X1 U14571 ( .A1(n14427), .A2(n12125), .B1(n14100), .B2(n14940), .ZN(
        n12128) );
  OAI211_X1 U14572 ( .C1(n14814), .C2(n12126), .A(n14948), .B(n12168), .ZN(
        n14813) );
  NOR2_X1 U14573 ( .A1(n14813), .A2(n14334), .ZN(n12127) );
  AOI211_X1 U14574 ( .C1(n14417), .C2(n14104), .A(n12128), .B(n12127), .ZN(
        n12129) );
  OAI211_X1 U14575 ( .C1(n14810), .C2(n14432), .A(n12130), .B(n12129), .ZN(
        P1_U3278) );
  XOR2_X1 U14576 ( .A(n12131), .B(n12142), .Z(n12134) );
  AND2_X1 U14577 ( .A1(n13536), .A2(n13509), .ZN(n12132) );
  AOI21_X1 U14578 ( .B1(n13534), .B2(n13510), .A(n12132), .ZN(n12226) );
  INV_X1 U14579 ( .A(n12226), .ZN(n12133) );
  AOI21_X1 U14580 ( .B1(n12134), .B2(n15161), .A(n12133), .ZN(n13874) );
  NAND2_X1 U14581 ( .A1(n12135), .A2(n13869), .ZN(n12136) );
  NAND2_X1 U14582 ( .A1(n12136), .A2(n13742), .ZN(n12137) );
  NOR2_X1 U14583 ( .A1(n6568), .A2(n12137), .ZN(n13868) );
  NAND2_X1 U14584 ( .A1(n13869), .A2(n15170), .ZN(n12140) );
  INV_X1 U14585 ( .A(n12138), .ZN(n12228) );
  AOI22_X1 U14586 ( .A1(n15174), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12228), 
        .B2(n15163), .ZN(n12139) );
  NAND2_X1 U14587 ( .A1(n12140), .A2(n12139), .ZN(n12141) );
  AOI21_X1 U14588 ( .B1(n13868), .B2(n15169), .A(n12141), .ZN(n12145) );
  NAND2_X1 U14589 ( .A1(n12143), .A2(n12142), .ZN(n13870) );
  NAND3_X1 U14590 ( .A1(n13871), .A2(n15168), .A3(n13870), .ZN(n12144) );
  OAI211_X1 U14591 ( .C1(n13874), .C2(n15149), .A(n12145), .B(n12144), .ZN(
        P2_U3249) );
  INV_X1 U14592 ( .A(n12146), .ZN(n12147) );
  AOI21_X1 U14593 ( .B1(n12149), .B2(n6919), .A(n12147), .ZN(n12158) );
  NOR2_X1 U14594 ( .A1(n14101), .A2(n12150), .ZN(n12156) );
  NAND2_X1 U14595 ( .A1(n14097), .A2(n12151), .ZN(n12152) );
  OAI211_X1 U14596 ( .C1(n14088), .C2(n12154), .A(n12153), .B(n12152), .ZN(
        n12155) );
  AOI211_X1 U14597 ( .C1(n15022), .C2(n14103), .A(n12156), .B(n12155), .ZN(
        n12157) );
  OAI21_X1 U14598 ( .B1(n12158), .B2(n14106), .A(n12157), .ZN(P1_U3217) );
  XNOR2_X1 U14599 ( .A(n12159), .B(n12166), .ZN(n12160) );
  NAND2_X1 U14600 ( .A1(n12160), .A2(n14937), .ZN(n12165) );
  OR2_X1 U14601 ( .A1(n14072), .A2(n14268), .ZN(n12163) );
  OR2_X1 U14602 ( .A1(n12161), .A2(n14085), .ZN(n12162) );
  NAND2_X1 U14603 ( .A1(n12163), .A2(n12162), .ZN(n14004) );
  INV_X1 U14604 ( .A(n14004), .ZN(n12164) );
  NAND2_X1 U14605 ( .A1(n12165), .A2(n12164), .ZN(n14809) );
  INV_X1 U14606 ( .A(n14809), .ZN(n12174) );
  XNOR2_X1 U14607 ( .A(n12167), .B(n12166), .ZN(n14803) );
  AOI21_X1 U14608 ( .B1(n12168), .B2(n14804), .A(n14829), .ZN(n12169) );
  NAND2_X1 U14609 ( .A1(n12169), .A2(n6676), .ZN(n14805) );
  INV_X1 U14610 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14196) );
  OAI22_X1 U14611 ( .A1(n14427), .A2(n14196), .B1(n14006), .B2(n14940), .ZN(
        n12170) );
  AOI21_X1 U14612 ( .B1(n14804), .B2(n14417), .A(n12170), .ZN(n12171) );
  OAI21_X1 U14613 ( .B1(n14805), .B2(n14334), .A(n12171), .ZN(n12172) );
  AOI21_X1 U14614 ( .B1(n14803), .B2(n14954), .A(n12172), .ZN(n12173) );
  OAI21_X1 U14615 ( .B1(n12174), .B2(n14942), .A(n12173), .ZN(P1_U3277) );
  INV_X1 U14616 ( .A(n12175), .ZN(n12179) );
  INV_X1 U14617 ( .A(n12176), .ZN(n12177) );
  OAI222_X1 U14618 ( .A1(n13928), .A2(n12178), .B1(n13920), .B2(n12179), .C1(
        n12177), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U14619 ( .A1(n12180), .A2(P1_U3086), .B1(n14544), .B2(n12179), 
        .C1(n6736), .C2(n14542), .ZN(P1_U3330) );
  INV_X1 U14620 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15108) );
  NOR2_X1 U14621 ( .A1(n12181), .A2(n13861), .ZN(n12185) );
  NOR4_X1 U14622 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12187) );
  MUX2_X1 U14623 ( .A(n15108), .B(n12187), .S(n15250), .Z(n12186) );
  OAI21_X1 U14624 ( .B1(n9944), .B2(n13850), .A(n12186), .ZN(P2_U3514) );
  INV_X1 U14625 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13045) );
  MUX2_X1 U14626 ( .A(n13045), .B(n12187), .S(n15242), .Z(n12188) );
  OAI21_X1 U14627 ( .B1(n9944), .B2(n13903), .A(n12188), .ZN(P2_U3475) );
  OR2_X1 U14628 ( .A1(n12189), .A2(n12192), .ZN(n12190) );
  NAND2_X1 U14629 ( .A1(n12191), .A2(n12190), .ZN(n13862) );
  XNOR2_X1 U14630 ( .A(n12193), .B(n12192), .ZN(n12194) );
  NAND2_X1 U14631 ( .A1(n12194), .A2(n15161), .ZN(n12196) );
  AND2_X1 U14632 ( .A1(n13535), .A2(n13509), .ZN(n12195) );
  AOI21_X1 U14633 ( .B1(n13533), .B2(n13510), .A(n12195), .ZN(n12337) );
  NAND2_X1 U14634 ( .A1(n12196), .A2(n12337), .ZN(n13867) );
  NAND2_X1 U14635 ( .A1(n13867), .A2(n11353), .ZN(n12201) );
  INV_X1 U14636 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12197) );
  OAI22_X1 U14637 ( .A1(n11353), .A2(n12197), .B1(n12335), .B2(n13774), .ZN(
        n12199) );
  OAI211_X1 U14638 ( .C1(n6568), .C2(n13864), .A(n13785), .B(n13742), .ZN(
        n13863) );
  NOR2_X1 U14639 ( .A1(n13863), .A2(n13747), .ZN(n12198) );
  AOI211_X1 U14640 ( .C1(n15170), .C2(n12340), .A(n12199), .B(n12198), .ZN(
        n12200) );
  OAI211_X1 U14641 ( .C1(n13862), .C2(n13793), .A(n12201), .B(n12200), .ZN(
        P2_U3248) );
  OAI21_X1 U14642 ( .B1(n12204), .B2(n12203), .A(n13990), .ZN(n12205) );
  NAND2_X1 U14643 ( .A1(n12205), .A2(n14082), .ZN(n12211) );
  NOR2_X1 U14644 ( .A1(n14101), .A2(n12206), .ZN(n12207) );
  AOI211_X1 U14645 ( .C1(n14097), .C2(n12209), .A(n12208), .B(n12207), .ZN(
        n12210) );
  OAI211_X1 U14646 ( .C1(n7189), .C2(n14093), .A(n12211), .B(n12210), .ZN(
        P1_U3236) );
  XNOR2_X1 U14647 ( .A(n12212), .B(n12391), .ZN(n12213) );
  OAI222_X1 U14648 ( .A1(n15382), .A2(n12271), .B1(n15381), .B2(n14739), .C1(
        n12213), .C2(n15388), .ZN(n14754) );
  INV_X1 U14649 ( .A(n14754), .ZN(n12220) );
  XNOR2_X1 U14650 ( .A(n12214), .B(n12475), .ZN(n14756) );
  NOR2_X1 U14651 ( .A1(n12405), .A2(n15346), .ZN(n14755) );
  INV_X1 U14652 ( .A(n14755), .ZN(n12217) );
  AOI22_X1 U14653 ( .A1(n15398), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15395), 
        .B2(n12215), .ZN(n12216) );
  OAI21_X1 U14654 ( .B1(n12250), .B2(n12217), .A(n12216), .ZN(n12218) );
  AOI21_X1 U14655 ( .B1(n14756), .B2(n13306), .A(n12218), .ZN(n12219) );
  OAI21_X1 U14656 ( .B1(n12220), .B2(n15398), .A(n12219), .ZN(P3_U3220) );
  INV_X1 U14657 ( .A(n13869), .ZN(n12231) );
  OAI21_X1 U14658 ( .B1(n12223), .B2(n12222), .A(n12221), .ZN(n12225) );
  NAND2_X1 U14659 ( .A1(n12225), .A2(n12224), .ZN(n12230) );
  NAND2_X1 U14660 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n15126)
         );
  OAI21_X1 U14661 ( .B1(n13491), .B2(n12226), .A(n15126), .ZN(n12227) );
  AOI21_X1 U14662 ( .B1(n12228), .B2(n13493), .A(n12227), .ZN(n12229) );
  OAI211_X1 U14663 ( .C1(n12231), .C2(n8883), .A(n12230), .B(n12229), .ZN(
        P2_U3198) );
  NAND2_X1 U14664 ( .A1(n12703), .A2(n12407), .ZN(n12235) );
  NAND2_X1 U14665 ( .A1(n12698), .A2(n15309), .ZN(n12234) );
  NAND2_X1 U14666 ( .A1(n12689), .A2(n14731), .ZN(n12233) );
  NAND4_X1 U14667 ( .A1(n12235), .A2(n12234), .A3(n12233), .A4(n12232), .ZN(
        n12241) );
  NOR2_X1 U14668 ( .A1(n12237), .A2(n6687), .ZN(n12238) );
  XNOR2_X1 U14669 ( .A(n12236), .B(n12238), .ZN(n12239) );
  NOR2_X1 U14670 ( .A1(n12239), .A2(n12691), .ZN(n12240) );
  AOI211_X1 U14671 ( .C1(n12679), .C2(n14730), .A(n12241), .B(n12240), .ZN(
        n12242) );
  INV_X1 U14672 ( .A(n12242), .ZN(P3_U3164) );
  XNOR2_X1 U14673 ( .A(n12243), .B(n12408), .ZN(n12244) );
  OAI222_X1 U14674 ( .A1(n15382), .A2(n12245), .B1(n15381), .B2(n14729), .C1(
        n12244), .C2(n15388), .ZN(n14751) );
  INV_X1 U14675 ( .A(n14751), .ZN(n12254) );
  XNOR2_X1 U14676 ( .A(n12246), .B(n12476), .ZN(n14753) );
  NOR2_X1 U14677 ( .A1(n12247), .A2(n15346), .ZN(n14752) );
  INV_X1 U14678 ( .A(n14752), .ZN(n12251) );
  AOI22_X1 U14679 ( .A1(n15398), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15395), 
        .B2(n12248), .ZN(n12249) );
  OAI21_X1 U14680 ( .B1(n12251), .B2(n12250), .A(n12249), .ZN(n12252) );
  AOI21_X1 U14681 ( .B1(n14753), .B2(n13306), .A(n12252), .ZN(n12253) );
  OAI21_X1 U14682 ( .B1(n12254), .B2(n15398), .A(n12253), .ZN(P3_U3219) );
  INV_X1 U14683 ( .A(n12255), .ZN(n12260) );
  OAI222_X1 U14684 ( .A1(P1_U3086), .A2(n12257), .B1(n14544), .B2(n12260), 
        .C1(n12256), .C2(n14542), .ZN(P1_U3329) );
  INV_X1 U14685 ( .A(n12258), .ZN(n12261) );
  OAI222_X1 U14686 ( .A1(n12261), .A2(P2_U3088), .B1(n13920), .B2(n12260), 
        .C1(n12259), .C2(n13928), .ZN(P2_U3301) );
  XNOR2_X1 U14687 ( .A(n12262), .B(n12482), .ZN(n12263) );
  AOI222_X1 U14688 ( .A1(n15341), .A2(n12263), .B1(n12713), .B2(n15326), .C1(
        n12711), .C2(n15324), .ZN(n13364) );
  XNOR2_X1 U14689 ( .A(n12264), .B(n12482), .ZN(n13362) );
  AOI22_X1 U14690 ( .A1(n15398), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15395), 
        .B2(n12274), .ZN(n12265) );
  OAI21_X1 U14691 ( .B1(n13365), .B2(n13304), .A(n12265), .ZN(n12266) );
  AOI21_X1 U14692 ( .B1(n13362), .B2(n13306), .A(n12266), .ZN(n12267) );
  OAI21_X1 U14693 ( .B1(n13364), .B2(n15398), .A(n12267), .ZN(P3_U3218) );
  XNOR2_X1 U14694 ( .A(n12269), .B(n12268), .ZN(n12276) );
  AND2_X1 U14695 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14713) );
  AOI21_X1 U14696 ( .B1(n12703), .B2(n12711), .A(n14713), .ZN(n12270) );
  OAI21_X1 U14697 ( .B1(n12271), .B2(n12296), .A(n12270), .ZN(n12273) );
  NOR2_X1 U14698 ( .A1(n13365), .A2(n12706), .ZN(n12272) );
  AOI211_X1 U14699 ( .C1(n12274), .C2(n12689), .A(n12273), .B(n12272), .ZN(
        n12275) );
  OAI21_X1 U14700 ( .B1(n12276), .B2(n12691), .A(n12275), .ZN(P3_U3181) );
  XNOR2_X1 U14701 ( .A(n12278), .B(n12392), .ZN(n12279) );
  AOI222_X1 U14702 ( .A1(n15341), .A2(n12279), .B1(n13283), .B2(n15324), .C1(
        n12712), .C2(n15326), .ZN(n13361) );
  OAI21_X1 U14703 ( .B1(n12281), .B2(n12392), .A(n12280), .ZN(n13359) );
  AOI22_X1 U14704 ( .A1(n15398), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15395), 
        .B2(n12641), .ZN(n12282) );
  OAI21_X1 U14705 ( .B1(n7601), .B2(n13304), .A(n12282), .ZN(n12283) );
  AOI21_X1 U14706 ( .B1(n13359), .B2(n13306), .A(n12283), .ZN(n12284) );
  OAI21_X1 U14707 ( .B1(n13361), .B2(n15398), .A(n12284), .ZN(P3_U3217) );
  INV_X1 U14708 ( .A(n12285), .ZN(n12287) );
  INV_X1 U14709 ( .A(n12290), .ZN(n13924) );
  OAI222_X1 U14710 ( .A1(n9524), .A2(P1_U3086), .B1(n14544), .B2(n13924), .C1(
        n13127), .C2(n14542), .ZN(P1_U3327) );
  XNOR2_X1 U14711 ( .A(n12399), .B(n10865), .ZN(n12298) );
  INV_X1 U14712 ( .A(n12298), .ZN(n12291) );
  NAND2_X1 U14713 ( .A1(n12291), .A2(n12696), .ZN(n12305) );
  INV_X1 U14714 ( .A(n12292), .ZN(n12293) );
  NAND4_X1 U14715 ( .A1(n12304), .A2(n12696), .A3(n12293), .A4(n12298), .ZN(
        n12303) );
  AOI22_X1 U14716 ( .A1(n12898), .A2(n12689), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12295) );
  NAND2_X1 U14717 ( .A1(n12707), .A2(n12703), .ZN(n12294) );
  OAI211_X1 U14718 ( .C1(n12529), .C2(n12296), .A(n12295), .B(n12294), .ZN(
        n12300) );
  NOR4_X1 U14719 ( .A1(n12298), .A2(n12297), .A3(n12691), .A4(n12921), .ZN(
        n12299) );
  AOI211_X1 U14720 ( .C1(n12679), .C2(n12301), .A(n12300), .B(n12299), .ZN(
        n12302) );
  OAI211_X1 U14721 ( .C1(n12305), .C2(n12304), .A(n12303), .B(n12302), .ZN(
        P3_U3160) );
  NAND3_X1 U14722 ( .A1(n12307), .A2(n13484), .A3(n13538), .ZN(n12308) );
  OAI21_X1 U14723 ( .B1(n6940), .B2(n13520), .A(n12308), .ZN(n12315) );
  NOR2_X1 U14724 ( .A1(n14776), .A2(n8883), .ZN(n12313) );
  NAND2_X1 U14725 ( .A1(n13513), .A2(n12309), .ZN(n12310) );
  NAND2_X1 U14726 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15102)
         );
  OAI211_X1 U14727 ( .C1(n13515), .C2(n12311), .A(n12310), .B(n15102), .ZN(
        n12312) );
  AOI211_X1 U14728 ( .C1(n12315), .C2(n12314), .A(n12313), .B(n12312), .ZN(
        n12316) );
  OAI21_X1 U14729 ( .B1(n12317), .B2(n13520), .A(n12316), .ZN(P2_U3187) );
  OR3_X1 U14730 ( .A1(n12383), .A2(n15410), .A3(n12318), .ZN(n12319) );
  OAI21_X1 U14731 ( .B1(n8111), .B2(n15382), .A(n12319), .ZN(n12325) );
  INV_X1 U14732 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n12320) );
  NOR2_X1 U14733 ( .A1(n15430), .A2(n12320), .ZN(n12321) );
  AOI21_X1 U14734 ( .B1(n15430), .B2(n12325), .A(n12321), .ZN(n12322) );
  OAI21_X1 U14735 ( .B1(n12328), .B2(n13392), .A(n12322), .ZN(P3_U3390) );
  NOR2_X1 U14736 ( .A1(n15438), .A2(n11009), .ZN(n12323) );
  AOI21_X1 U14737 ( .B1(n15438), .B2(n12325), .A(n12323), .ZN(n12324) );
  OAI21_X1 U14738 ( .B1(n12328), .B2(n13339), .A(n12324), .ZN(P3_U3459) );
  AOI21_X1 U14739 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15395), .A(n12325), .ZN(
        n12326) );
  MUX2_X1 U14740 ( .A(n11010), .B(n12326), .S(n15396), .Z(n12327) );
  OAI21_X1 U14741 ( .B1(n12328), .B2(n13304), .A(n12327), .ZN(P3_U3233) );
  INV_X1 U14742 ( .A(n12329), .ZN(n12331) );
  OAI222_X1 U14743 ( .A1(n13419), .A2(n12331), .B1(n13423), .B2(n12330), .C1(
        P3_U3151), .C2(n15255), .ZN(P3_U3268) );
  INV_X1 U14744 ( .A(n12332), .ZN(n13919) );
  OAI222_X1 U14745 ( .A1(P1_U3086), .A2(n12334), .B1(n14544), .B2(n13919), 
        .C1(n12333), .C2(n14542), .ZN(P1_U3326) );
  NOR2_X1 U14746 ( .A1(n13515), .A2(n12335), .ZN(n12339) );
  OAI22_X1 U14747 ( .A1(n13491), .A2(n12337), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12336), .ZN(n12338) );
  AOI211_X1 U14748 ( .C1(n12340), .C2(n13518), .A(n12339), .B(n12338), .ZN(
        n12348) );
  INV_X1 U14749 ( .A(n12341), .ZN(n12346) );
  OAI22_X1 U14750 ( .A1(n12344), .A2(n13520), .B1(n12343), .B2(n12342), .ZN(
        n12345) );
  NAND3_X1 U14751 ( .A1(n12221), .A2(n12346), .A3(n12345), .ZN(n12347) );
  OAI211_X1 U14752 ( .C1(n12349), .C2(n13520), .A(n12348), .B(n12347), .ZN(
        P2_U3200) );
  OAI222_X1 U14753 ( .A1(n13419), .A2(n12351), .B1(n13423), .B2(n13055), .C1(
        P3_U3151), .C2(n12350), .ZN(P3_U3274) );
  OAI22_X1 U14754 ( .A1(n14539), .A2(n13914), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12368) );
  NAND2_X1 U14755 ( .A1(n12368), .A2(n12367), .ZN(n12354) );
  OAI21_X1 U14756 ( .B1(n13914), .B2(P2_DATAO_REG_30__SCAN_IN), .A(n12354), 
        .ZN(n12357) );
  INV_X1 U14757 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12355) );
  INV_X1 U14758 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14532) );
  AOI22_X1 U14759 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n12355), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n14532), .ZN(n12356) );
  XOR2_X1 U14760 ( .A(n12357), .B(n12356), .Z(n13411) );
  INV_X1 U14761 ( .A(SI_31_), .ZN(n13416) );
  NOR2_X1 U14762 ( .A1(n12358), .A2(n13416), .ZN(n12359) );
  INV_X1 U14763 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14748) );
  NAND2_X1 U14764 ( .A1(n12360), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12362) );
  NAND2_X1 U14765 ( .A1(n9570), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12361) );
  OAI211_X1 U14766 ( .C1(n14748), .C2(n12363), .A(n12362), .B(n12361), .ZN(
        n12364) );
  INV_X1 U14767 ( .A(n12364), .ZN(n12365) );
  NAND2_X1 U14768 ( .A1(n12366), .A2(n12365), .ZN(n14718) );
  NAND2_X1 U14769 ( .A1(n14745), .A2(n14718), .ZN(n12549) );
  INV_X1 U14770 ( .A(n14718), .ZN(n12373) );
  INV_X1 U14771 ( .A(n12367), .ZN(n12369) );
  XNOR2_X1 U14772 ( .A(n12369), .B(n12368), .ZN(n12559) );
  NAND2_X1 U14773 ( .A1(n12370), .A2(n12559), .ZN(n12372) );
  INV_X1 U14774 ( .A(SI_30_), .ZN(n12561) );
  OR2_X1 U14775 ( .A1(n12358), .A2(n12561), .ZN(n12371) );
  OAI21_X1 U14776 ( .B1(n12546), .B2(n12373), .A(n12380), .ZN(n12374) );
  NAND3_X1 U14777 ( .A1(n12549), .A2(n12374), .A3(n12540), .ZN(n12378) );
  INV_X1 U14778 ( .A(n12380), .ZN(n12375) );
  NAND2_X1 U14779 ( .A1(n12381), .A2(n12375), .ZN(n12545) );
  NOR2_X1 U14780 ( .A1(n12545), .A2(n14745), .ZN(n12376) );
  NOR2_X1 U14781 ( .A1(n14745), .A2(n14718), .ZN(n12548) );
  NAND2_X1 U14782 ( .A1(n12514), .A2(n12513), .ZN(n12978) );
  INV_X1 U14783 ( .A(n12978), .ZN(n12972) );
  INV_X1 U14784 ( .A(n12519), .ZN(n12397) );
  XNOR2_X1 U14785 ( .A(n12381), .B(n12380), .ZN(n12541) );
  XNOR2_X1 U14786 ( .A(n15325), .B(n15347), .ZN(n15336) );
  NAND4_X1 U14787 ( .A1(n15379), .A2(n12435), .A3(n12382), .A4(n12454), .ZN(
        n12387) );
  NAND4_X1 U14788 ( .A1(n8114), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        n12386) );
  NOR4_X1 U14789 ( .A1(n15336), .A2(n6505), .A3(n12387), .A4(n12386), .ZN(
        n12388) );
  NAND4_X1 U14790 ( .A1(n14737), .A2(n12463), .A3(n12388), .A4(n14725), .ZN(
        n12389) );
  NOR4_X1 U14791 ( .A1(n12391), .A2(n12408), .A3(n12390), .A4(n12389), .ZN(
        n12393) );
  AND3_X1 U14792 ( .A1(n13300), .A2(n12393), .A3(n12392), .ZN(n12394) );
  INV_X1 U14793 ( .A(n12989), .ZN(n12396) );
  INV_X1 U14794 ( .A(n12401), .ZN(n12404) );
  INV_X1 U14795 ( .A(n12402), .ZN(n12403) );
  MUX2_X1 U14796 ( .A(n12404), .B(n12403), .S(n12530), .Z(n12532) );
  INV_X1 U14797 ( .A(n13383), .ZN(n13329) );
  INV_X1 U14798 ( .A(n12405), .ZN(n12406) );
  MUX2_X1 U14799 ( .A(n12407), .B(n12406), .S(n12530), .Z(n12409) );
  AOI21_X1 U14800 ( .B1(n12410), .B2(n12409), .A(n12408), .ZN(n12479) );
  INV_X1 U14801 ( .A(n12411), .ZN(n12413) );
  MUX2_X1 U14802 ( .A(n12413), .B(n6503), .S(n12547), .Z(n12478) );
  NOR2_X1 U14803 ( .A1(n12417), .A2(n12555), .ZN(n12415) );
  MUX2_X1 U14804 ( .A(n12416), .B(n12415), .S(n12414), .Z(n12420) );
  INV_X1 U14805 ( .A(n8109), .ZN(n12422) );
  INV_X1 U14806 ( .A(n12417), .ZN(n12418) );
  AOI21_X1 U14807 ( .B1(n12421), .B2(n12418), .A(n12547), .ZN(n12419) );
  NOR3_X1 U14808 ( .A1(n12420), .A2(n12422), .A3(n12419), .ZN(n12426) );
  INV_X1 U14809 ( .A(n12421), .ZN(n12423) );
  MUX2_X1 U14810 ( .A(n12423), .B(n12422), .S(n12530), .Z(n12425) );
  INV_X1 U14811 ( .A(n15379), .ZN(n12424) );
  NOR3_X1 U14812 ( .A1(n12426), .A2(n12425), .A3(n12424), .ZN(n12434) );
  NAND2_X1 U14813 ( .A1(n7735), .A2(n12427), .ZN(n12430) );
  NAND2_X1 U14814 ( .A1(n12431), .A2(n12428), .ZN(n12429) );
  MUX2_X1 U14815 ( .A(n12430), .B(n12429), .S(n12530), .Z(n12433) );
  MUX2_X1 U14816 ( .A(n12431), .B(n7735), .S(n12530), .Z(n12432) );
  OAI21_X1 U14817 ( .B1(n12434), .B2(n12433), .A(n12432), .ZN(n12436) );
  NAND2_X1 U14818 ( .A1(n12436), .A2(n12435), .ZN(n12440) );
  MUX2_X1 U14819 ( .A(n12438), .B(n12437), .S(n12530), .Z(n12439) );
  NAND2_X1 U14820 ( .A1(n12446), .A2(n12441), .ZN(n12444) );
  NAND2_X1 U14821 ( .A1(n12445), .A2(n12442), .ZN(n12443) );
  MUX2_X1 U14822 ( .A(n12444), .B(n12443), .S(n12530), .Z(n12448) );
  MUX2_X1 U14823 ( .A(n12446), .B(n12445), .S(n12547), .Z(n12447) );
  INV_X1 U14824 ( .A(n12449), .ZN(n12452) );
  INV_X1 U14825 ( .A(n12450), .ZN(n12451) );
  MUX2_X1 U14826 ( .A(n12452), .B(n12451), .S(n12547), .Z(n12453) );
  MUX2_X1 U14827 ( .A(n12456), .B(n12455), .S(n12547), .Z(n12457) );
  NAND2_X1 U14828 ( .A1(n12458), .A2(n15310), .ZN(n12460) );
  MUX2_X1 U14829 ( .A(n12460), .B(n12459), .S(n12530), .Z(n12461) );
  AND2_X1 U14830 ( .A1(n12462), .A2(n12461), .ZN(n12468) );
  NAND2_X1 U14831 ( .A1(n12464), .A2(n15323), .ZN(n12466) );
  MUX2_X1 U14832 ( .A(n12466), .B(n12465), .S(n12530), .Z(n12467) );
  INV_X1 U14833 ( .A(n12473), .ZN(n12470) );
  OAI21_X1 U14834 ( .B1(n6504), .B2(n12470), .A(n12547), .ZN(n12471) );
  AOI21_X1 U14835 ( .B1(n6674), .B2(n12472), .A(n12547), .ZN(n12474) );
  OAI21_X1 U14836 ( .B1(n12479), .B2(n12478), .A(n12477), .ZN(n12483) );
  OAI21_X1 U14837 ( .B1(n13358), .B2(n13296), .A(n12480), .ZN(n12481) );
  AOI22_X1 U14838 ( .A1(n12483), .A2(n12482), .B1(n12547), .B2(n12481), .ZN(
        n12487) );
  AND2_X1 U14839 ( .A1(n12485), .A2(n12484), .ZN(n12486) );
  OAI22_X1 U14840 ( .A1(n12487), .A2(n7226), .B1(n12486), .B2(n12547), .ZN(
        n12490) );
  NAND3_X1 U14841 ( .A1(n7601), .A2(n12530), .A3(n12711), .ZN(n12489) );
  INV_X1 U14842 ( .A(n13300), .ZN(n12488) );
  AOI211_X1 U14843 ( .C1(n12490), .C2(n12489), .A(n12488), .B(n6502), .ZN(
        n12502) );
  INV_X1 U14844 ( .A(n12494), .ZN(n12493) );
  OAI211_X1 U14845 ( .C1(n12493), .C2(n12492), .A(n12498), .B(n12491), .ZN(
        n12497) );
  OAI211_X1 U14846 ( .C1(n6502), .C2(n12495), .A(n12499), .B(n12494), .ZN(
        n12496) );
  MUX2_X1 U14847 ( .A(n12497), .B(n12496), .S(n12547), .Z(n12501) );
  MUX2_X1 U14848 ( .A(n12499), .B(n12498), .S(n12547), .Z(n12500) );
  OAI211_X1 U14849 ( .C1(n12502), .C2(n12501), .A(n13001), .B(n12500), .ZN(
        n12512) );
  NOR2_X1 U14850 ( .A1(n12615), .A2(n12547), .ZN(n12504) );
  NOR2_X1 U14851 ( .A1(n13011), .A2(n12530), .ZN(n12503) );
  MUX2_X1 U14852 ( .A(n12504), .B(n12503), .S(n13396), .Z(n12505) );
  NOR2_X1 U14853 ( .A1(n12989), .A2(n12505), .ZN(n12511) );
  INV_X1 U14854 ( .A(n12506), .ZN(n12509) );
  INV_X1 U14855 ( .A(n12507), .ZN(n12508) );
  MUX2_X1 U14856 ( .A(n12509), .B(n12508), .S(n12547), .Z(n12510) );
  AOI211_X1 U14857 ( .C1(n12512), .C2(n12511), .A(n12510), .B(n12978), .ZN(
        n12518) );
  INV_X1 U14858 ( .A(n12513), .ZN(n12516) );
  INV_X1 U14859 ( .A(n12514), .ZN(n12515) );
  MUX2_X1 U14860 ( .A(n12516), .B(n12515), .S(n12530), .Z(n12517) );
  OAI33_X1 U14861 ( .A1(n12709), .A2(n13329), .A3(n12547), .B1(n12519), .B2(
        n12518), .B3(n12517), .ZN(n12520) );
  INV_X1 U14862 ( .A(n12521), .ZN(n12523) );
  OAI21_X1 U14863 ( .B1(n12523), .B2(n8053), .A(n12525), .ZN(n12524) );
  MUX2_X1 U14864 ( .A(n12525), .B(n12524), .S(n12547), .Z(n12526) );
  MUX2_X1 U14865 ( .A(n12913), .B(n12527), .S(n12530), .Z(n12528) );
  XNOR2_X1 U14866 ( .A(n12534), .B(n12547), .ZN(n12535) );
  AOI21_X1 U14867 ( .B1(n9537), .B2(n12536), .A(n12535), .ZN(n12537) );
  AOI21_X1 U14868 ( .B1(n9537), .B2(n12538), .A(n12537), .ZN(n12544) );
  MUX2_X1 U14869 ( .A(n12540), .B(n12539), .S(n12547), .Z(n12542) );
  NOR3_X1 U14870 ( .A1(n12554), .A2(n12553), .A3(n13420), .ZN(n12557) );
  OAI21_X1 U14871 ( .B1(n12558), .B2(n12555), .A(P3_B_REG_SCAN_IN), .ZN(n12556) );
  INV_X1 U14872 ( .A(n12559), .ZN(n12560) );
  OAI222_X1 U14873 ( .A1(n12562), .A2(P3_U3151), .B1(n13423), .B2(n12561), 
        .C1(n13419), .C2(n12560), .ZN(P3_U3265) );
  AND2_X1 U14874 ( .A1(n14029), .A2(n12566), .ZN(n12565) );
  NAND2_X1 U14875 ( .A1(n14030), .A2(n12565), .ZN(n14078) );
  INV_X1 U14876 ( .A(n12566), .ZN(n12568) );
  NAND2_X1 U14877 ( .A1(n14455), .A2(n12588), .ZN(n12570) );
  NAND2_X1 U14878 ( .A1(n14112), .A2(n12591), .ZN(n12569) );
  NAND2_X1 U14879 ( .A1(n12570), .A2(n12569), .ZN(n12571) );
  XNOR2_X1 U14880 ( .A(n12571), .B(n12589), .ZN(n12575) );
  NAND2_X1 U14881 ( .A1(n14455), .A2(n12591), .ZN(n12573) );
  NAND2_X1 U14882 ( .A1(n10196), .A2(n14112), .ZN(n12572) );
  NAND2_X1 U14883 ( .A1(n12573), .A2(n12572), .ZN(n12574) );
  NOR2_X1 U14884 ( .A1(n12575), .A2(n12574), .ZN(n12577) );
  AOI21_X1 U14885 ( .B1(n12575), .B2(n12574), .A(n12577), .ZN(n14081) );
  AND2_X1 U14886 ( .A1(n14077), .A2(n14081), .ZN(n12576) );
  INV_X1 U14887 ( .A(n12577), .ZN(n12578) );
  NAND2_X1 U14888 ( .A1(n14450), .A2(n12588), .ZN(n12580) );
  NAND2_X1 U14889 ( .A1(n14111), .A2(n12591), .ZN(n12579) );
  NAND2_X1 U14890 ( .A1(n12580), .A2(n12579), .ZN(n12581) );
  XNOR2_X1 U14891 ( .A(n12581), .B(n12589), .ZN(n12585) );
  NAND2_X1 U14892 ( .A1(n14450), .A2(n12591), .ZN(n12583) );
  NAND2_X1 U14893 ( .A1(n10196), .A2(n14111), .ZN(n12582) );
  NAND2_X1 U14894 ( .A1(n12583), .A2(n12582), .ZN(n12584) );
  NOR2_X1 U14895 ( .A1(n12585), .A2(n12584), .ZN(n12586) );
  AOI21_X1 U14896 ( .B1(n12585), .B2(n12584), .A(n12586), .ZN(n13932) );
  AOI22_X1 U14897 ( .A1(n14446), .A2(n12588), .B1(n12591), .B2(n14110), .ZN(
        n12590) );
  XNOR2_X1 U14898 ( .A(n12590), .B(n12589), .ZN(n12593) );
  AOI22_X1 U14899 ( .A1(n14446), .A2(n12591), .B1(n10196), .B2(n14110), .ZN(
        n12592) );
  XNOR2_X1 U14900 ( .A(n12593), .B(n12592), .ZN(n12594) );
  XNOR2_X1 U14901 ( .A(n12595), .B(n12594), .ZN(n12601) );
  NAND2_X1 U14902 ( .A1(n14109), .A2(n14071), .ZN(n12597) );
  NAND2_X1 U14903 ( .A1(n14111), .A2(n14052), .ZN(n12596) );
  NAND2_X1 U14904 ( .A1(n12597), .A2(n12596), .ZN(n14237) );
  AOI22_X1 U14905 ( .A1(n14097), .A2(n14237), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12598) );
  OAI21_X1 U14906 ( .B1(n14101), .B2(n14240), .A(n12598), .ZN(n12599) );
  AOI21_X1 U14907 ( .B1(n14446), .B2(n14103), .A(n12599), .ZN(n12600) );
  OAI21_X1 U14908 ( .B1(n12601), .B2(n14106), .A(n12600), .ZN(P1_U3220) );
  OAI222_X1 U14909 ( .A1(n12604), .A2(P1_U3086), .B1(n14544), .B2(n12603), 
        .C1(n12602), .C2(n14542), .ZN(P1_U3331) );
  NOR2_X1 U14910 ( .A1(n6579), .A2(n12605), .ZN(n12656) );
  AOI21_X1 U14911 ( .B1(n6579), .B2(n12605), .A(n12656), .ZN(n12606) );
  NAND2_X1 U14912 ( .A1(n12606), .A2(n12976), .ZN(n12659) );
  OAI21_X1 U14913 ( .B1(n12976), .B2(n12606), .A(n12659), .ZN(n12607) );
  NAND2_X1 U14914 ( .A1(n12607), .A2(n12696), .ZN(n12611) );
  AOI22_X1 U14915 ( .A1(n12698), .A2(n12987), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12608) );
  OAI21_X1 U14916 ( .B1(n12933), .B2(n12685), .A(n12608), .ZN(n12609) );
  AOI21_X1 U14917 ( .B1(n12964), .B2(n12689), .A(n12609), .ZN(n12610) );
  OAI211_X1 U14918 ( .C1(n13329), .C2(n12706), .A(n12611), .B(n12610), .ZN(
        P3_U3156) );
  XNOR2_X1 U14919 ( .A(n12613), .B(n12612), .ZN(n12619) );
  NAND2_X1 U14920 ( .A1(n12698), .A2(n13010), .ZN(n12614) );
  NAND2_X1 U14921 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12888)
         );
  OAI211_X1 U14922 ( .C1(n12615), .C2(n12685), .A(n12614), .B(n12888), .ZN(
        n12617) );
  INV_X1 U14923 ( .A(n13400), .ZN(n13018) );
  NOR2_X1 U14924 ( .A1(n13018), .A2(n12706), .ZN(n12616) );
  AOI211_X1 U14925 ( .C1(n13016), .C2(n12689), .A(n12617), .B(n12616), .ZN(
        n12618) );
  OAI21_X1 U14926 ( .B1(n12619), .B2(n12691), .A(n12618), .ZN(P3_U3159) );
  OAI21_X1 U14927 ( .B1(n12622), .B2(n12621), .A(n12620), .ZN(n12623) );
  NAND2_X1 U14928 ( .A1(n12623), .A2(n12696), .ZN(n12628) );
  AOI22_X1 U14929 ( .A1(n12698), .A2(n13011), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12624) );
  OAI21_X1 U14930 ( .B1(n12625), .B2(n12685), .A(n12624), .ZN(n12626) );
  AOI21_X1 U14931 ( .B1(n12991), .B2(n12689), .A(n12626), .ZN(n12627) );
  OAI211_X1 U14932 ( .C1(n13393), .C2(n12706), .A(n12628), .B(n12627), .ZN(
        P3_U3163) );
  INV_X1 U14933 ( .A(n13375), .ZN(n13318) );
  INV_X1 U14934 ( .A(n12629), .ZN(n12633) );
  NOR3_X1 U14935 ( .A1(n12660), .A2(n12631), .A3(n12630), .ZN(n12632) );
  OAI21_X1 U14936 ( .B1(n12633), .B2(n12632), .A(n12696), .ZN(n12637) );
  AOI22_X1 U14937 ( .A1(n12960), .A2(n12698), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12634) );
  OAI21_X1 U14938 ( .B1(n12934), .B2(n12685), .A(n12634), .ZN(n12635) );
  AOI21_X1 U14939 ( .B1(n12941), .B2(n12689), .A(n12635), .ZN(n12636) );
  OAI211_X1 U14940 ( .C1(n13318), .C2(n12706), .A(n12637), .B(n12636), .ZN(
        P3_U3165) );
  XNOR2_X1 U14941 ( .A(n12639), .B(n12638), .ZN(n12647) );
  NOR2_X1 U14942 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12640), .ZN(n12806) );
  AOI21_X1 U14943 ( .B1(n12698), .B2(n12712), .A(n12806), .ZN(n12643) );
  NAND2_X1 U14944 ( .A1(n12689), .A2(n12641), .ZN(n12642) );
  OAI211_X1 U14945 ( .C1(n12644), .C2(n12685), .A(n12643), .B(n12642), .ZN(
        n12645) );
  AOI21_X1 U14946 ( .B1(n13358), .B2(n12679), .A(n12645), .ZN(n12646) );
  OAI21_X1 U14947 ( .B1(n12647), .B2(n12691), .A(n12646), .ZN(P3_U3166) );
  XNOR2_X1 U14948 ( .A(n12649), .B(n12648), .ZN(n12654) );
  NAND2_X1 U14949 ( .A1(n12698), .A2(n12711), .ZN(n12650) );
  NAND2_X1 U14950 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12832)
         );
  OAI211_X1 U14951 ( .C1(n13295), .C2(n12685), .A(n12650), .B(n12832), .ZN(
        n12652) );
  NOR2_X1 U14952 ( .A1(n13357), .A2(n12706), .ZN(n12651) );
  AOI211_X1 U14953 ( .C1(n13302), .C2(n12689), .A(n12652), .B(n12651), .ZN(
        n12653) );
  OAI21_X1 U14954 ( .B1(n12654), .B2(n12691), .A(n12653), .ZN(P3_U3168) );
  INV_X1 U14955 ( .A(n12655), .ZN(n13380) );
  INV_X1 U14956 ( .A(n12656), .ZN(n12657) );
  AND3_X1 U14957 ( .A1(n12659), .A2(n12658), .A3(n12657), .ZN(n12661) );
  OAI21_X1 U14958 ( .B1(n12661), .B2(n12660), .A(n12696), .ZN(n12665) );
  AOI22_X1 U14959 ( .A1(n12709), .A2(n12698), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12662) );
  OAI21_X1 U14960 ( .B1(n12949), .B2(n12685), .A(n12662), .ZN(n12663) );
  AOI21_X1 U14961 ( .B1(n12953), .B2(n12689), .A(n12663), .ZN(n12664) );
  OAI211_X1 U14962 ( .C1(n13380), .C2(n12706), .A(n12665), .B(n12664), .ZN(
        P3_U3169) );
  XNOR2_X1 U14963 ( .A(n12666), .B(n12667), .ZN(n12672) );
  AOI22_X1 U14964 ( .A1(n12698), .A2(n13284), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12669) );
  NAND2_X1 U14965 ( .A1(n12689), .A2(n13003), .ZN(n12668) );
  OAI211_X1 U14966 ( .C1(n12975), .C2(n12685), .A(n12669), .B(n12668), .ZN(
        n12670) );
  AOI21_X1 U14967 ( .B1(n13396), .B2(n12679), .A(n12670), .ZN(n12671) );
  OAI21_X1 U14968 ( .B1(n12672), .B2(n12691), .A(n12671), .ZN(P3_U3173) );
  INV_X1 U14969 ( .A(n12673), .ZN(n12674) );
  AOI21_X1 U14970 ( .B1(n12987), .B2(n12675), .A(n12674), .ZN(n12681) );
  AOI22_X1 U14971 ( .A1(n12698), .A2(n12998), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12677) );
  NAND2_X1 U14972 ( .A1(n12689), .A2(n12980), .ZN(n12676) );
  OAI211_X1 U14973 ( .C1(n12976), .C2(n12685), .A(n12677), .B(n12676), .ZN(
        n12678) );
  AOI21_X1 U14974 ( .B1(n12979), .B2(n12679), .A(n12678), .ZN(n12680) );
  OAI21_X1 U14975 ( .B1(n12681), .B2(n12691), .A(n12680), .ZN(P3_U3175) );
  XNOR2_X1 U14976 ( .A(n12683), .B(n12682), .ZN(n12692) );
  NAND2_X1 U14977 ( .A1(n12698), .A2(n13283), .ZN(n12684) );
  NAND2_X1 U14978 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12858)
         );
  OAI211_X1 U14979 ( .C1(n12686), .C2(n12685), .A(n12684), .B(n12858), .ZN(
        n12688) );
  INV_X1 U14980 ( .A(n13350), .ZN(n13291) );
  NOR2_X1 U14981 ( .A1(n13291), .A2(n12706), .ZN(n12687) );
  AOI211_X1 U14982 ( .C1(n13289), .C2(n12689), .A(n12688), .B(n12687), .ZN(
        n12690) );
  OAI21_X1 U14983 ( .B1(n12692), .B2(n12691), .A(n12690), .ZN(P3_U3178) );
  OAI21_X1 U14984 ( .B1(n12695), .B2(n12694), .A(n12693), .ZN(n12697) );
  NAND2_X1 U14985 ( .A1(n12697), .A2(n12696), .ZN(n12705) );
  INV_X1 U14986 ( .A(n12925), .ZN(n12701) );
  AOI22_X1 U14987 ( .A1(n12920), .A2(n12698), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12699) );
  OAI21_X1 U14988 ( .B1(n12701), .B2(n12700), .A(n12699), .ZN(n12702) );
  AOI21_X1 U14989 ( .B1(n12703), .B2(n12921), .A(n12702), .ZN(n12704) );
  OAI211_X1 U14990 ( .C1(n13372), .C2(n12706), .A(n12705), .B(n12704), .ZN(
        P3_U3180) );
  MUX2_X1 U14991 ( .A(n14718), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12710), .Z(
        P3_U3522) );
  MUX2_X1 U14992 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12707), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14993 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12921), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14994 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12708), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14995 ( .A(n12960), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12710), .Z(
        P3_U3515) );
  MUX2_X1 U14996 ( .A(n12709), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12710), .Z(
        P3_U3514) );
  MUX2_X1 U14997 ( .A(n12987), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12710), .Z(
        P3_U3513) );
  MUX2_X1 U14998 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12998), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14999 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13011), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15000 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13283), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15001 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12711), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15002 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12712), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15003 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12713), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15004 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12714), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15005 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n15309), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15006 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n15323), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15007 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n15310), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15008 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n15325), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15009 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12715), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15010 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12716), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15011 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12717), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15012 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12718), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15013 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12719), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15014 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n6803), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15015 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12721), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15016 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n10839), .S(P3_U3897), .Z(
        P3_U3491) );
  NAND2_X1 U15017 ( .A1(n15281), .A2(n12722), .ZN(n12739) );
  AOI21_X1 U15018 ( .B1(n15274), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n12723), .ZN(
        n12738) );
  INV_X1 U15019 ( .A(n12724), .ZN(n12728) );
  INV_X1 U15020 ( .A(n12725), .ZN(n12727) );
  OAI21_X1 U15021 ( .B1(n12728), .B2(n12727), .A(n12726), .ZN(n12731) );
  OAI21_X1 U15022 ( .B1(n6574), .B2(n6706), .A(n12729), .ZN(n12730) );
  AOI22_X1 U15023 ( .A1(n15254), .A2(n12731), .B1(n15252), .B2(n12730), .ZN(
        n12737) );
  NOR2_X1 U15024 ( .A1(n12733), .A2(n12732), .ZN(n12734) );
  OAI21_X1 U15025 ( .B1(n12735), .B2(n12734), .A(n15279), .ZN(n12736) );
  NAND4_X1 U15026 ( .A1(n12739), .A2(n12738), .A3(n12737), .A4(n12736), .ZN(
        P3_U3186) );
  INV_X1 U15027 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12744) );
  AOI21_X1 U15028 ( .B1(n12744), .B2(n12743), .A(n12769), .ZN(n12763) );
  MUX2_X1 U15029 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n15255), .Z(n12773) );
  XNOR2_X1 U15030 ( .A(n12773), .B(n12772), .ZN(n12751) );
  NAND2_X1 U15031 ( .A1(n12745), .A2(n12755), .ZN(n12749) );
  NAND2_X1 U15032 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  AOI21_X1 U15033 ( .B1(n12751), .B2(n12750), .A(n12776), .ZN(n12754) );
  AOI21_X1 U15034 ( .B1(n15274), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12752), 
        .ZN(n12753) );
  OAI21_X1 U15035 ( .B1(n12754), .B2(n15296), .A(n12753), .ZN(n12761) );
  NAND2_X1 U15036 ( .A1(n12755), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12756) );
  AOI21_X1 U15037 ( .B1(n7883), .B2(n12758), .A(n12764), .ZN(n12759) );
  NOR2_X1 U15038 ( .A1(n12759), .A2(n15298), .ZN(n12760) );
  AOI211_X1 U15039 ( .C1(n15281), .C2(n12768), .A(n12761), .B(n12760), .ZN(
        n12762) );
  OAI21_X1 U15040 ( .B1(n12763), .B2(n15304), .A(n12762), .ZN(P3_U3195) );
  NAND2_X1 U15041 ( .A1(n12771), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12808) );
  OAI21_X1 U15042 ( .B1(n12771), .B2(P3_REG1_REG_14__SCAN_IN), .A(n12808), 
        .ZN(n12774) );
  AOI21_X1 U15043 ( .B1(n6684), .B2(n12774), .A(n12809), .ZN(n12785) );
  NOR2_X1 U15044 ( .A1(n12768), .A2(n12767), .ZN(n12770) );
  NAND2_X1 U15045 ( .A1(n12771), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12795) );
  OAI21_X1 U15046 ( .B1(n12771), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12795), 
        .ZN(n12788) );
  XNOR2_X1 U15047 ( .A(n12789), .B(n12788), .ZN(n12783) );
  NOR2_X1 U15048 ( .A1(n15290), .A2(n12771), .ZN(n12782) );
  INV_X1 U15049 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n13043) );
  NOR2_X1 U15050 ( .A1(n12773), .A2(n12772), .ZN(n12777) );
  MUX2_X1 U15051 ( .A(n12788), .B(n12774), .S(n15255), .Z(n12775) );
  OAI21_X1 U15052 ( .B1(n12777), .B2(n12776), .A(n12775), .ZN(n12778) );
  NAND3_X1 U15053 ( .A1(n15279), .A2(n12797), .A3(n12778), .ZN(n12779) );
  OAI211_X1 U15054 ( .C1(n15287), .C2(n13043), .A(n12780), .B(n12779), .ZN(
        n12781) );
  AOI211_X1 U15055 ( .C1(n12783), .C2(n15254), .A(n12782), .B(n12781), .ZN(
        n12784) );
  OAI21_X1 U15056 ( .B1(n12785), .B2(n15298), .A(n12784), .ZN(P3_U3196) );
  INV_X1 U15057 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U15058 ( .A1(n12825), .A2(n12801), .ZN(n12786) );
  OAI21_X1 U15059 ( .B1(n12825), .B2(n12801), .A(n12786), .ZN(n12787) );
  INV_X1 U15060 ( .A(n12787), .ZN(n12794) );
  AND2_X1 U15061 ( .A1(n14701), .A2(n12790), .ZN(n12791) );
  INV_X1 U15062 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14699) );
  NOR2_X1 U15063 ( .A1(n14699), .A2(n14698), .ZN(n14697) );
  INV_X1 U15064 ( .A(n12827), .ZN(n12792) );
  AOI21_X1 U15065 ( .B1(n12794), .B2(n12793), .A(n12792), .ZN(n12820) );
  MUX2_X1 U15066 ( .A(n12795), .B(n12808), .S(n15255), .Z(n12796) );
  AOI21_X1 U15067 ( .B1(n14701), .B2(n12798), .A(n12799), .ZN(n14706) );
  MUX2_X1 U15068 ( .A(n14699), .B(n14704), .S(n15255), .Z(n14705) );
  AND2_X1 U15069 ( .A1(n14706), .A2(n14705), .ZN(n14708) );
  NOR2_X1 U15070 ( .A1(n12799), .A2(n14708), .ZN(n12835) );
  MUX2_X1 U15071 ( .A(n12801), .B(n12800), .S(n15255), .Z(n12803) );
  INV_X1 U15072 ( .A(n12825), .ZN(n12802) );
  NAND2_X1 U15073 ( .A1(n12803), .A2(n12802), .ZN(n12834) );
  MUX2_X1 U15074 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n15255), .Z(n12804) );
  AND2_X1 U15075 ( .A1(n12804), .A2(n12825), .ZN(n12836) );
  NAND2_X1 U15076 ( .A1(n12834), .A2(n7004), .ZN(n12805) );
  XNOR2_X1 U15077 ( .A(n12835), .B(n12805), .ZN(n12818) );
  AOI21_X1 U15078 ( .B1(n15274), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12806), 
        .ZN(n12807) );
  OAI21_X1 U15079 ( .B1(n15290), .B2(n12825), .A(n12807), .ZN(n12817) );
  NOR2_X1 U15080 ( .A1(n12811), .A2(n12810), .ZN(n12812) );
  NOR2_X1 U15081 ( .A1(n14704), .A2(n14703), .ZN(n14702) );
  NAND2_X1 U15082 ( .A1(n12825), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12821) );
  OAI21_X1 U15083 ( .B1(n12825), .B2(P3_REG1_REG_16__SCAN_IN), .A(n12821), 
        .ZN(n12813) );
  NAND2_X1 U15084 ( .A1(n12814), .A2(n12813), .ZN(n12815) );
  AOI21_X1 U15085 ( .B1(n12822), .B2(n12815), .A(n15298), .ZN(n12816) );
  AOI211_X1 U15086 ( .C1(n15279), .C2(n12818), .A(n12817), .B(n12816), .ZN(
        n12819) );
  OAI21_X1 U15087 ( .B1(n12820), .B2(n15304), .A(n12819), .ZN(P3_U3198) );
  AOI21_X1 U15088 ( .B1(n12824), .B2(n12823), .A(n12861), .ZN(n12842) );
  INV_X1 U15089 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U15090 ( .A1(n12825), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U15091 ( .A1(n15274), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12831) );
  OAI211_X1 U15092 ( .C1(n15304), .C2(n12833), .A(n12832), .B(n12831), .ZN(
        n12840) );
  MUX2_X1 U15093 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n15255), .Z(n12850) );
  XNOR2_X1 U15094 ( .A(n12850), .B(n12849), .ZN(n12837) );
  AOI211_X1 U15095 ( .C1(n12838), .C2(n12837), .A(n6665), .B(n15296), .ZN(
        n12839) );
  AOI211_X1 U15096 ( .C1(n15281), .C2(n12860), .A(n12840), .B(n12839), .ZN(
        n12841) );
  OAI21_X1 U15097 ( .B1(n12842), .B2(n15298), .A(n12841), .ZN(P3_U3199) );
  NOR2_X1 U15098 ( .A1(n12860), .A2(n12843), .ZN(n12845) );
  NAND2_X1 U15099 ( .A1(n12863), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12870) );
  OAI21_X1 U15100 ( .B1(n12863), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12870), 
        .ZN(n12847) );
  INV_X1 U15101 ( .A(n12871), .ZN(n12846) );
  AOI21_X1 U15102 ( .B1(n12848), .B2(n12847), .A(n12846), .ZN(n12869) );
  INV_X1 U15103 ( .A(n12863), .ZN(n12880) );
  INV_X1 U15104 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14656) );
  NAND2_X1 U15105 ( .A1(n12850), .A2(n12849), .ZN(n12851) );
  XNOR2_X1 U15106 ( .A(n12878), .B(n12880), .ZN(n12855) );
  INV_X1 U15107 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12853) );
  MUX2_X1 U15108 ( .A(n12853), .B(n12852), .S(n15255), .Z(n12854) );
  AND2_X1 U15109 ( .A1(n12855), .A2(n12854), .ZN(n12879) );
  NOR2_X1 U15110 ( .A1(n12855), .A2(n12854), .ZN(n12856) );
  OAI21_X1 U15111 ( .B1(n12879), .B2(n12856), .A(n15279), .ZN(n12857) );
  OAI211_X1 U15112 ( .C1(n15287), .C2(n14656), .A(n12858), .B(n12857), .ZN(
        n12867) );
  NOR2_X1 U15113 ( .A1(n12860), .A2(n12859), .ZN(n12862) );
  NAND2_X1 U15114 ( .A1(n12863), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12875) );
  OAI21_X1 U15115 ( .B1(n12863), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12875), 
        .ZN(n12864) );
  AOI21_X1 U15116 ( .B1(n12865), .B2(n12864), .A(n12877), .ZN(n12866) );
  OAI21_X1 U15117 ( .B1(n12869), .B2(n15304), .A(n12868), .ZN(P3_U3200) );
  NAND2_X1 U15118 ( .A1(n12871), .A2(n12870), .ZN(n12874) );
  XNOR2_X1 U15119 ( .A(n12872), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12883) );
  INV_X1 U15120 ( .A(n12883), .ZN(n12873) );
  XNOR2_X1 U15121 ( .A(n12874), .B(n12873), .ZN(n12891) );
  INV_X1 U15122 ( .A(n12875), .ZN(n12876) );
  XNOR2_X1 U15123 ( .A(n12889), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12882) );
  INV_X1 U15124 ( .A(n12878), .ZN(n12881) );
  AOI21_X1 U15125 ( .B1(n12881), .B2(n12880), .A(n12879), .ZN(n12886) );
  INV_X1 U15126 ( .A(n12882), .ZN(n12884) );
  MUX2_X1 U15127 ( .A(n12884), .B(n12883), .S(n12553), .Z(n12885) );
  NAND2_X1 U15128 ( .A1(n15274), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12887) );
  OAI211_X1 U15129 ( .C1(n15290), .C2(n12889), .A(n12888), .B(n12887), .ZN(
        n12890) );
  INV_X1 U15130 ( .A(n12892), .ZN(n12897) );
  AOI22_X1 U15131 ( .A1(n14719), .A2(n15395), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15398), .ZN(n12893) );
  OAI21_X1 U15132 ( .B1(n12894), .B2(n13304), .A(n12893), .ZN(n12895) );
  OAI21_X1 U15133 ( .B1(n12897), .B2(n15398), .A(n12896), .ZN(P3_U3204) );
  AOI22_X1 U15134 ( .A1(n12898), .A2(n15395), .B1(n15398), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12899) );
  OAI21_X1 U15135 ( .B1(n12900), .B2(n13304), .A(n12899), .ZN(n12901) );
  AOI21_X1 U15136 ( .B1(n12902), .B2(n13306), .A(n12901), .ZN(n12903) );
  OAI21_X1 U15137 ( .B1(n12904), .B2(n15398), .A(n12903), .ZN(P3_U3205) );
  INV_X1 U15138 ( .A(n12905), .ZN(n12911) );
  AND2_X1 U15139 ( .A1(n15396), .A2(n15390), .ZN(n12968) );
  AOI22_X1 U15140 ( .A1(n12906), .A2(n15395), .B1(n15398), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12907) );
  OAI21_X1 U15141 ( .B1(n13368), .B2(n13304), .A(n12907), .ZN(n12908) );
  AOI21_X1 U15142 ( .B1(n12909), .B2(n12968), .A(n12908), .ZN(n12910) );
  OAI21_X1 U15143 ( .B1(n12911), .B2(n15398), .A(n12910), .ZN(P3_U3206) );
  INV_X1 U15144 ( .A(n15385), .ZN(n15345) );
  NAND2_X1 U15145 ( .A1(n12912), .A2(n12913), .ZN(n12914) );
  NAND2_X1 U15146 ( .A1(n12914), .A2(n12917), .ZN(n12916) );
  NAND2_X1 U15147 ( .A1(n12916), .A2(n12915), .ZN(n12924) );
  XOR2_X1 U15148 ( .A(n12918), .B(n12917), .Z(n12919) );
  NAND2_X1 U15149 ( .A1(n12919), .A2(n15341), .ZN(n12923) );
  AOI22_X1 U15150 ( .A1(n12921), .A2(n15324), .B1(n15326), .B2(n12920), .ZN(
        n12922) );
  OAI211_X1 U15151 ( .C1(n15345), .C2(n12924), .A(n12923), .B(n12922), .ZN(
        n13308) );
  INV_X1 U15152 ( .A(n13308), .ZN(n12929) );
  INV_X1 U15153 ( .A(n12924), .ZN(n13309) );
  AOI22_X1 U15154 ( .A1(n12925), .A2(n15395), .B1(n15398), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12926) );
  OAI21_X1 U15155 ( .B1(n13372), .B2(n13304), .A(n12926), .ZN(n12927) );
  AOI21_X1 U15156 ( .B1(n13309), .B2(n12968), .A(n12927), .ZN(n12928) );
  OAI21_X1 U15157 ( .B1(n12929), .B2(n15398), .A(n12928), .ZN(P3_U3207) );
  NAND2_X1 U15158 ( .A1(n12930), .A2(n12938), .ZN(n12931) );
  NAND3_X1 U15159 ( .A1(n12932), .A2(n15341), .A3(n12931), .ZN(n12937) );
  OAI22_X1 U15160 ( .A1(n12934), .A2(n15382), .B1(n12933), .B2(n15381), .ZN(
        n12935) );
  INV_X1 U15161 ( .A(n12935), .ZN(n12936) );
  OR2_X1 U15162 ( .A1(n12939), .A2(n12938), .ZN(n12940) );
  NAND2_X1 U15163 ( .A1(n12912), .A2(n12940), .ZN(n13312) );
  AOI22_X1 U15164 ( .A1(n15398), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12941), 
        .B2(n15395), .ZN(n12942) );
  OAI21_X1 U15165 ( .B1(n13318), .B2(n13304), .A(n12942), .ZN(n12943) );
  AOI21_X1 U15166 ( .B1(n13312), .B2(n13306), .A(n12943), .ZN(n12944) );
  OAI21_X1 U15167 ( .B1(n13314), .B2(n15398), .A(n12944), .ZN(P3_U3208) );
  XNOR2_X1 U15168 ( .A(n12946), .B(n12945), .ZN(n12952) );
  OAI21_X1 U15169 ( .B1(n12948), .B2(n7070), .A(n12947), .ZN(n13320) );
  OAI22_X1 U15170 ( .A1(n12949), .A2(n15382), .B1(n12976), .B2(n15381), .ZN(
        n12950) );
  AOI21_X1 U15171 ( .B1(n13320), .B2(n15385), .A(n12950), .ZN(n12951) );
  OAI21_X1 U15172 ( .B1(n12952), .B2(n15388), .A(n12951), .ZN(n13319) );
  INV_X1 U15173 ( .A(n13319), .ZN(n12957) );
  AOI22_X1 U15174 ( .A1(n15398), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12953), 
        .B2(n15395), .ZN(n12954) );
  OAI21_X1 U15175 ( .B1(n13380), .B2(n13304), .A(n12954), .ZN(n12955) );
  AOI21_X1 U15176 ( .B1(n13320), .B2(n12968), .A(n12955), .ZN(n12956) );
  OAI21_X1 U15177 ( .B1(n12957), .B2(n15398), .A(n12956), .ZN(P3_U3209) );
  XNOR2_X1 U15178 ( .A(n12958), .B(n12397), .ZN(n12963) );
  XNOR2_X1 U15179 ( .A(n12959), .B(n12397), .ZN(n13323) );
  AOI22_X1 U15180 ( .A1(n12960), .A2(n15324), .B1(n15326), .B2(n12987), .ZN(
        n12961) );
  OAI21_X1 U15181 ( .B1(n13323), .B2(n15345), .A(n12961), .ZN(n12962) );
  AOI21_X1 U15182 ( .B1(n12963), .B2(n15341), .A(n12962), .ZN(n13326) );
  INV_X1 U15183 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12966) );
  INV_X1 U15184 ( .A(n12964), .ZN(n12965) );
  OAI22_X1 U15185 ( .A1(n15396), .A2(n12966), .B1(n12965), .B2(n15376), .ZN(
        n12967) );
  AOI21_X1 U15186 ( .B1(n13383), .B2(n15374), .A(n12967), .ZN(n12971) );
  INV_X1 U15187 ( .A(n12968), .ZN(n12969) );
  OR2_X1 U15188 ( .A1(n13323), .A2(n12969), .ZN(n12970) );
  OAI211_X1 U15189 ( .C1(n13326), .C2(n15398), .A(n12971), .B(n12970), .ZN(
        P3_U3210) );
  XNOR2_X1 U15190 ( .A(n12973), .B(n12972), .ZN(n12974) );
  OAI222_X1 U15191 ( .A1(n15382), .A2(n12976), .B1(n15381), .B2(n12975), .C1(
        n15388), .C2(n12974), .ZN(n13330) );
  INV_X1 U15192 ( .A(n13330), .ZN(n12984) );
  XNOR2_X1 U15193 ( .A(n12977), .B(n12978), .ZN(n13331) );
  INV_X1 U15194 ( .A(n12979), .ZN(n13388) );
  AOI22_X1 U15195 ( .A1(n15398), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15395), 
        .B2(n12980), .ZN(n12981) );
  OAI21_X1 U15196 ( .B1(n13388), .B2(n13304), .A(n12981), .ZN(n12982) );
  AOI21_X1 U15197 ( .B1(n13331), .B2(n13306), .A(n12982), .ZN(n12983) );
  OAI21_X1 U15198 ( .B1(n12984), .B2(n15398), .A(n12983), .ZN(P3_U3211) );
  OAI21_X1 U15199 ( .B1(n12986), .B2(n12989), .A(n12985), .ZN(n12988) );
  AOI222_X1 U15200 ( .A1(n15341), .A2(n12988), .B1(n12987), .B2(n15324), .C1(
        n13011), .C2(n15326), .ZN(n13334) );
  XNOR2_X1 U15201 ( .A(n12990), .B(n12989), .ZN(n13336) );
  AOI22_X1 U15202 ( .A1(n15398), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15395), 
        .B2(n12991), .ZN(n12992) );
  OAI21_X1 U15203 ( .B1(n13393), .B2(n13304), .A(n12992), .ZN(n12993) );
  AOI21_X1 U15204 ( .B1(n13336), .B2(n13306), .A(n12993), .ZN(n12994) );
  OAI21_X1 U15205 ( .B1(n13334), .B2(n15398), .A(n12994), .ZN(P3_U3212) );
  OAI211_X1 U15206 ( .C1(n12997), .C2(n12996), .A(n6839), .B(n15341), .ZN(
        n13000) );
  AOI22_X1 U15207 ( .A1(n12998), .A2(n15324), .B1(n13284), .B2(n15326), .ZN(
        n12999) );
  AND2_X1 U15208 ( .A1(n13000), .A2(n12999), .ZN(n13342) );
  XNOR2_X1 U15209 ( .A(n13002), .B(n13001), .ZN(n13340) );
  AOI22_X1 U15210 ( .A1(n15398), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15395), 
        .B2(n13003), .ZN(n13004) );
  OAI21_X1 U15211 ( .B1(n6500), .B2(n13304), .A(n13004), .ZN(n13005) );
  AOI21_X1 U15212 ( .B1(n13340), .B2(n13306), .A(n13005), .ZN(n13006) );
  OAI21_X1 U15213 ( .B1(n13342), .B2(n15398), .A(n13006), .ZN(P3_U3213) );
  NAND2_X1 U15214 ( .A1(n13007), .A2(n13014), .ZN(n13008) );
  NAND3_X1 U15215 ( .A1(n13009), .A2(n15341), .A3(n13008), .ZN(n13013) );
  AOI22_X1 U15216 ( .A1(n13011), .A2(n15324), .B1(n15326), .B2(n13010), .ZN(
        n13012) );
  AND2_X1 U15217 ( .A1(n13013), .A2(n13012), .ZN(n13347) );
  XNOR2_X1 U15218 ( .A(n13015), .B(n6861), .ZN(n13345) );
  AOI22_X1 U15219 ( .A1(n15398), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15395), 
        .B2(n13016), .ZN(n13017) );
  OAI21_X1 U15220 ( .B1(n13018), .B2(n13304), .A(n13017), .ZN(n13019) );
  AOI21_X1 U15221 ( .B1(n13345), .B2(n13306), .A(n13019), .ZN(n13020) );
  OAI21_X1 U15222 ( .B1(n13347), .B2(n15398), .A(n13020), .ZN(n13280) );
  INV_X1 U15223 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U15224 ( .A1(n13022), .A2(keyinput91), .B1(keyinput89), .B2(n13244), 
        .ZN(n13021) );
  OAI221_X1 U15225 ( .B1(n13022), .B2(keyinput91), .C1(n13244), .C2(keyinput89), .A(n13021), .ZN(n13028) );
  INV_X1 U15226 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U15227 ( .A1(n13024), .A2(keyinput93), .B1(keyinput12), .B2(n13833), 
        .ZN(n13023) );
  OAI221_X1 U15228 ( .B1(n13024), .B2(keyinput93), .C1(n13833), .C2(keyinput12), .A(n13023), .ZN(n13027) );
  XNOR2_X1 U15229 ( .A(keyinput76), .B(n11377), .ZN(n13026) );
  INV_X1 U15230 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14551) );
  XNOR2_X1 U15231 ( .A(keyinput40), .B(n14551), .ZN(n13025) );
  OR4_X1 U15232 ( .A1(n13028), .A2(n13027), .A3(n13026), .A4(n13025), .ZN(
        n13036) );
  AOI22_X1 U15233 ( .A1(n13030), .A2(keyinput53), .B1(n7664), .B2(keyinput111), 
        .ZN(n13029) );
  OAI221_X1 U15234 ( .B1(n13030), .B2(keyinput53), .C1(n7664), .C2(keyinput111), .A(n13029), .ZN(n13035) );
  AOI22_X1 U15235 ( .A1(n13033), .A2(keyinput71), .B1(keyinput78), .B2(n13032), 
        .ZN(n13031) );
  OAI221_X1 U15236 ( .B1(n13033), .B2(keyinput71), .C1(n13032), .C2(keyinput78), .A(n13031), .ZN(n13034) );
  NOR3_X1 U15237 ( .A1(n13036), .A2(n13035), .A3(n13034), .ZN(n13078) );
  INV_X1 U15238 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n13038) );
  AOI22_X1 U15239 ( .A1(n14556), .A2(keyinput70), .B1(n13038), .B2(keyinput17), 
        .ZN(n13037) );
  OAI221_X1 U15240 ( .B1(n14556), .B2(keyinput70), .C1(n13038), .C2(keyinput17), .A(n13037), .ZN(n13050) );
  INV_X1 U15241 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U15242 ( .A1(n13041), .A2(keyinput41), .B1(n13040), .B2(keyinput19), 
        .ZN(n13039) );
  OAI221_X1 U15243 ( .B1(n13041), .B2(keyinput41), .C1(n13040), .C2(keyinput19), .A(n13039), .ZN(n13049) );
  INV_X1 U15244 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U15245 ( .A1(n13043), .A2(keyinput22), .B1(n14801), .B2(keyinput98), 
        .ZN(n13042) );
  OAI221_X1 U15246 ( .B1(n13043), .B2(keyinput22), .C1(n14801), .C2(keyinput98), .A(n13042), .ZN(n13048) );
  INV_X1 U15247 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U15248 ( .A1(n13046), .A2(keyinput65), .B1(n13045), .B2(keyinput16), 
        .ZN(n13044) );
  OAI221_X1 U15249 ( .B1(n13046), .B2(keyinput65), .C1(n13045), .C2(keyinput16), .A(n13044), .ZN(n13047) );
  NOR4_X1 U15250 ( .A1(n13050), .A2(n13049), .A3(n13048), .A4(n13047), .ZN(
        n13077) );
  INV_X1 U15251 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U15252 ( .A1(n15128), .A2(keyinput99), .B1(n7832), .B2(keyinput46), 
        .ZN(n13051) );
  OAI221_X1 U15253 ( .B1(n15128), .B2(keyinput99), .C1(n7832), .C2(keyinput46), 
        .A(n13051), .ZN(n13060) );
  INV_X1 U15254 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U15255 ( .A1(n15431), .A2(keyinput5), .B1(keyinput11), .B2(n13053), 
        .ZN(n13052) );
  OAI221_X1 U15256 ( .B1(n15431), .B2(keyinput5), .C1(n13053), .C2(keyinput11), 
        .A(n13052), .ZN(n13059) );
  AOI22_X1 U15257 ( .A1(n13055), .A2(keyinput56), .B1(n13223), .B2(keyinput58), 
        .ZN(n13054) );
  OAI221_X1 U15258 ( .B1(n13055), .B2(keyinput56), .C1(n13223), .C2(keyinput58), .A(n13054), .ZN(n13058) );
  INV_X1 U15259 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15177) );
  AOI22_X1 U15260 ( .A1(P1_U3086), .A2(keyinput7), .B1(n15177), .B2(keyinput14), .ZN(n13056) );
  OAI221_X1 U15261 ( .B1(P1_U3086), .B2(keyinput7), .C1(n15177), .C2(
        keyinput14), .A(n13056), .ZN(n13057) );
  NOR4_X1 U15262 ( .A1(n13060), .A2(n13059), .A3(n13058), .A4(n13057), .ZN(
        n13076) );
  AOI22_X1 U15263 ( .A1(n13063), .A2(keyinput105), .B1(n13062), .B2(keyinput38), .ZN(n13061) );
  OAI221_X1 U15264 ( .B1(n13063), .B2(keyinput105), .C1(n13062), .C2(
        keyinput38), .A(n13061), .ZN(n13068) );
  INV_X1 U15265 ( .A(P2_B_REG_SCAN_IN), .ZN(n13065) );
  AOI22_X1 U15266 ( .A1(n13235), .A2(keyinput103), .B1(keyinput116), .B2(
        n13065), .ZN(n13064) );
  OAI221_X1 U15267 ( .B1(n13235), .B2(keyinput103), .C1(n13065), .C2(
        keyinput116), .A(n13064), .ZN(n13067) );
  XNOR2_X1 U15268 ( .A(n14640), .B(keyinput67), .ZN(n13066) );
  OR3_X1 U15269 ( .A1(n13068), .A2(n13067), .A3(n13066), .ZN(n13074) );
  AOI22_X1 U15270 ( .A1(n13233), .A2(keyinput54), .B1(keyinput88), .B2(n10636), 
        .ZN(n13069) );
  OAI221_X1 U15271 ( .B1(n13233), .B2(keyinput54), .C1(n10636), .C2(keyinput88), .A(n13069), .ZN(n13073) );
  INV_X1 U15272 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13232) );
  AOI22_X1 U15273 ( .A1(n13232), .A2(keyinput118), .B1(keyinput104), .B2(
        n13071), .ZN(n13070) );
  OAI221_X1 U15274 ( .B1(n13232), .B2(keyinput118), .C1(n13071), .C2(
        keyinput104), .A(n13070), .ZN(n13072) );
  NOR3_X1 U15275 ( .A1(n13074), .A2(n13073), .A3(n13072), .ZN(n13075) );
  NAND4_X1 U15276 ( .A1(n13078), .A2(n13077), .A3(n13076), .A4(n13075), .ZN(
        n13146) );
  AOI22_X1 U15277 ( .A1(n13080), .A2(keyinput13), .B1(n7731), .B2(keyinput66), 
        .ZN(n13079) );
  OAI221_X1 U15278 ( .B1(n13080), .B2(keyinput13), .C1(n7731), .C2(keyinput66), 
        .A(n13079), .ZN(n13089) );
  AOI22_X1 U15279 ( .A1(n13082), .A2(keyinput108), .B1(n8161), .B2(keyinput114), .ZN(n13081) );
  OAI221_X1 U15280 ( .B1(n13082), .B2(keyinput108), .C1(n8161), .C2(
        keyinput114), .A(n13081), .ZN(n13088) );
  AOI22_X1 U15281 ( .A1(n13084), .A2(keyinput32), .B1(n9401), .B2(keyinput1), 
        .ZN(n13083) );
  OAI221_X1 U15282 ( .B1(n13084), .B2(keyinput32), .C1(n9401), .C2(keyinput1), 
        .A(n13083), .ZN(n13087) );
  INV_X1 U15283 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13589) );
  AOI22_X1 U15284 ( .A1(n13589), .A2(keyinput115), .B1(n13221), .B2(keyinput96), .ZN(n13085) );
  OAI221_X1 U15285 ( .B1(n13589), .B2(keyinput115), .C1(n13221), .C2(
        keyinput96), .A(n13085), .ZN(n13086) );
  NOR4_X1 U15286 ( .A1(n13089), .A2(n13088), .A3(n13087), .A4(n13086), .ZN(
        n13092) );
  INV_X1 U15287 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14957) );
  XOR2_X1 U15288 ( .A(n14957), .B(keyinput59), .Z(n13091) );
  INV_X1 U15289 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14960) );
  XOR2_X1 U15290 ( .A(n14960), .B(keyinput74), .Z(n13090) );
  NAND3_X1 U15291 ( .A1(n13092), .A2(n13091), .A3(n13090), .ZN(n13145) );
  INV_X1 U15292 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15188) );
  AOI22_X1 U15293 ( .A1(n11009), .A2(keyinput3), .B1(keyinput122), .B2(n15188), 
        .ZN(n13093) );
  OAI221_X1 U15294 ( .B1(n11009), .B2(keyinput3), .C1(n15188), .C2(keyinput122), .A(n13093), .ZN(n13103) );
  AOI22_X1 U15295 ( .A1(n9370), .A2(keyinput90), .B1(n10881), .B2(keyinput123), 
        .ZN(n13094) );
  OAI221_X1 U15296 ( .B1(n9370), .B2(keyinput90), .C1(n10881), .C2(keyinput123), .A(n13094), .ZN(n13102) );
  INV_X1 U15297 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14553) );
  AOI22_X1 U15298 ( .A1(n14553), .A2(keyinput92), .B1(n13096), .B2(keyinput80), 
        .ZN(n13095) );
  OAI221_X1 U15299 ( .B1(n14553), .B2(keyinput92), .C1(n13096), .C2(keyinput80), .A(n13095), .ZN(n13101) );
  INV_X1 U15300 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U15301 ( .A1(n13099), .A2(keyinput52), .B1(keyinput43), .B2(n13098), 
        .ZN(n13097) );
  OAI221_X1 U15302 ( .B1(n13099), .B2(keyinput52), .C1(n13098), .C2(keyinput43), .A(n13097), .ZN(n13100) );
  OR4_X1 U15303 ( .A1(n13103), .A2(n13102), .A3(n13101), .A4(n13100), .ZN(
        n13144) );
  XOR2_X1 U15304 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput81), .Z(n13107) );
  XOR2_X1 U15305 ( .A(P3_IR_REG_31__SCAN_IN), .B(keyinput126), .Z(n13106) );
  XOR2_X1 U15306 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput61), .Z(n13105) );
  XOR2_X1 U15307 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput69), .Z(n13104) );
  NOR4_X1 U15308 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13142) );
  AOI22_X1 U15309 ( .A1(n10671), .A2(keyinput82), .B1(n13109), .B2(keyinput87), 
        .ZN(n13108) );
  OAI221_X1 U15310 ( .B1(n10671), .B2(keyinput82), .C1(n13109), .C2(keyinput87), .A(n13108), .ZN(n13125) );
  XOR2_X1 U15311 ( .A(keyinput63), .B(n8719), .Z(n13113) );
  XOR2_X1 U15312 ( .A(keyinput77), .B(n14204), .Z(n13112) );
  XNOR2_X1 U15313 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput124), .ZN(n13111) );
  XNOR2_X1 U15314 ( .A(P3_IR_REG_25__SCAN_IN), .B(keyinput39), .ZN(n13110) );
  NAND4_X1 U15315 ( .A1(n13113), .A2(n13112), .A3(n13111), .A4(n13110), .ZN(
        n13124) );
  XNOR2_X1 U15316 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput34), .ZN(n13117) );
  XNOR2_X1 U15317 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput125), .ZN(n13116)
         );
  XNOR2_X1 U15318 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(keyinput49), .ZN(n13115)
         );
  XNOR2_X1 U15319 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput85), .ZN(n13114) );
  NAND4_X1 U15320 ( .A1(n13117), .A2(n13116), .A3(n13115), .A4(n13114), .ZN(
        n13123) );
  XNOR2_X1 U15321 ( .A(P1_REG2_REG_21__SCAN_IN), .B(keyinput102), .ZN(n13121)
         );
  XNOR2_X1 U15322 ( .A(P3_D_REG_1__SCAN_IN), .B(keyinput101), .ZN(n13120) );
  XNOR2_X1 U15323 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput44), .ZN(n13119)
         );
  XNOR2_X1 U15324 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput31), .ZN(n13118) );
  NAND4_X1 U15325 ( .A1(n13121), .A2(n13120), .A3(n13119), .A4(n13118), .ZN(
        n13122) );
  NOR4_X1 U15326 ( .A1(n13125), .A2(n13124), .A3(n13123), .A4(n13122), .ZN(
        n13141) );
  INV_X1 U15327 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U15328 ( .A1(n13128), .A2(keyinput109), .B1(n13127), .B2(keyinput75), .ZN(n13126) );
  OAI221_X1 U15329 ( .B1(n13128), .B2(keyinput109), .C1(n13127), .C2(
        keyinput75), .A(n13126), .ZN(n13132) );
  XOR2_X1 U15330 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput35), .Z(n13131) );
  XOR2_X1 U15331 ( .A(SI_22_), .B(keyinput42), .Z(n13130) );
  XNOR2_X1 U15332 ( .A(keyinput36), .B(n11568), .ZN(n13129) );
  NOR4_X1 U15333 ( .A1(n13132), .A2(n13131), .A3(n13130), .A4(n13129), .ZN(
        n13140) );
  XOR2_X1 U15334 ( .A(P3_IR_REG_14__SCAN_IN), .B(keyinput15), .Z(n13138) );
  XOR2_X1 U15335 ( .A(P3_IR_REG_24__SCAN_IN), .B(keyinput64), .Z(n13137) );
  XNOR2_X1 U15336 ( .A(n13133), .B(keyinput97), .ZN(n13136) );
  XNOR2_X1 U15337 ( .A(n13134), .B(keyinput8), .ZN(n13135) );
  NOR4_X1 U15338 ( .A1(n13138), .A2(n13137), .A3(n13136), .A4(n13135), .ZN(
        n13139) );
  NAND4_X1 U15339 ( .A1(n13142), .A2(n13141), .A3(n13140), .A4(n13139), .ZN(
        n13143) );
  NOR4_X1 U15340 ( .A1(n13146), .A2(n13145), .A3(n13144), .A4(n13143), .ZN(
        n13182) );
  AOI22_X1 U15341 ( .A1(n7883), .A2(keyinput26), .B1(keyinput79), .B2(n9137), 
        .ZN(n13147) );
  OAI221_X1 U15342 ( .B1(n7883), .B2(keyinput26), .C1(n9137), .C2(keyinput79), 
        .A(n13147), .ZN(n13155) );
  INV_X1 U15343 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15092) );
  AOI22_X1 U15344 ( .A1(n15092), .A2(keyinput55), .B1(n14070), .B2(keyinput6), 
        .ZN(n13148) );
  OAI221_X1 U15345 ( .B1(n15092), .B2(keyinput55), .C1(n14070), .C2(keyinput6), 
        .A(n13148), .ZN(n13154) );
  INV_X1 U15346 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U15347 ( .A1(n13150), .A2(keyinput47), .B1(n12028), .B2(keyinput112), .ZN(n13149) );
  OAI221_X1 U15348 ( .B1(n13150), .B2(keyinput47), .C1(n12028), .C2(
        keyinput112), .A(n13149), .ZN(n13153) );
  AOI22_X1 U15349 ( .A1(n7419), .A2(keyinput120), .B1(keyinput4), .B2(n13234), 
        .ZN(n13151) );
  OAI221_X1 U15350 ( .B1(n7419), .B2(keyinput120), .C1(n13234), .C2(keyinput4), 
        .A(n13151), .ZN(n13152) );
  NOR4_X1 U15351 ( .A1(n13155), .A2(n13154), .A3(n13153), .A4(n13152), .ZN(
        n13181) );
  INV_X1 U15352 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U15353 ( .A1(n13157), .A2(keyinput48), .B1(n7720), .B2(keyinput117), 
        .ZN(n13156) );
  OAI221_X1 U15354 ( .B1(n13157), .B2(keyinput48), .C1(n7720), .C2(keyinput117), .A(n13156), .ZN(n13166) );
  AOI22_X1 U15355 ( .A1(n14567), .A2(keyinput119), .B1(n11006), .B2(keyinput23), .ZN(n13158) );
  OAI221_X1 U15356 ( .B1(n14567), .B2(keyinput119), .C1(n11006), .C2(
        keyinput23), .A(n13158), .ZN(n13165) );
  AOI22_X1 U15357 ( .A1(n13160), .A2(keyinput20), .B1(keyinput45), .B2(n9328), 
        .ZN(n13159) );
  OAI221_X1 U15358 ( .B1(n13160), .B2(keyinput20), .C1(n9328), .C2(keyinput45), 
        .A(n13159), .ZN(n13164) );
  INV_X1 U15359 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13889) );
  AOI22_X1 U15360 ( .A1(n13162), .A2(keyinput95), .B1(keyinput10), .B2(n13889), 
        .ZN(n13161) );
  OAI221_X1 U15361 ( .B1(n13162), .B2(keyinput95), .C1(n13889), .C2(keyinput10), .A(n13161), .ZN(n13163) );
  NOR4_X1 U15362 ( .A1(n13166), .A2(n13165), .A3(n13164), .A4(n13163), .ZN(
        n13180) );
  INV_X1 U15363 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14577) );
  AOI22_X1 U15364 ( .A1(n13168), .A2(keyinput27), .B1(keyinput127), .B2(n14577), .ZN(n13167) );
  OAI221_X1 U15365 ( .B1(n13168), .B2(keyinput27), .C1(n14577), .C2(
        keyinput127), .A(n13167), .ZN(n13178) );
  INV_X1 U15366 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14913) );
  INV_X1 U15367 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n13170) );
  AOI22_X1 U15368 ( .A1(n14913), .A2(keyinput106), .B1(n13170), .B2(keyinput9), 
        .ZN(n13169) );
  OAI221_X1 U15369 ( .B1(n14913), .B2(keyinput106), .C1(n13170), .C2(keyinput9), .A(n13169), .ZN(n13177) );
  AOI22_X1 U15370 ( .A1(n8973), .A2(keyinput0), .B1(n13172), .B2(keyinput121), 
        .ZN(n13171) );
  OAI221_X1 U15371 ( .B1(n8973), .B2(keyinput0), .C1(n13172), .C2(keyinput121), 
        .A(n13171), .ZN(n13176) );
  INV_X1 U15372 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n13174) );
  AOI22_X1 U15373 ( .A1(n11891), .A2(keyinput107), .B1(n13174), .B2(keyinput50), .ZN(n13173) );
  OAI221_X1 U15374 ( .B1(n11891), .B2(keyinput107), .C1(n13174), .C2(
        keyinput50), .A(n13173), .ZN(n13175) );
  NOR4_X1 U15375 ( .A1(n13178), .A2(n13177), .A3(n13176), .A4(n13175), .ZN(
        n13179) );
  AND4_X1 U15376 ( .A1(n13182), .A2(n13181), .A3(n13180), .A4(n13179), .ZN(
        n13220) );
  AOI22_X1 U15377 ( .A1(n13185), .A2(keyinput62), .B1(n13184), .B2(keyinput33), 
        .ZN(n13183) );
  OAI221_X1 U15378 ( .B1(n13185), .B2(keyinput62), .C1(n13184), .C2(keyinput33), .A(n13183), .ZN(n13194) );
  INV_X1 U15379 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14958) );
  AOI22_X1 U15380 ( .A1(n13187), .A2(keyinput60), .B1(keyinput83), .B2(n14958), 
        .ZN(n13186) );
  OAI221_X1 U15381 ( .B1(n13187), .B2(keyinput60), .C1(n14958), .C2(keyinput83), .A(n13186), .ZN(n13193) );
  AOI22_X1 U15382 ( .A1(n13222), .A2(keyinput24), .B1(keyinput25), .B2(n13189), 
        .ZN(n13188) );
  OAI221_X1 U15383 ( .B1(n13222), .B2(keyinput24), .C1(n13189), .C2(keyinput25), .A(n13188), .ZN(n13192) );
  AOI22_X1 U15384 ( .A1(n15351), .A2(keyinput73), .B1(keyinput84), .B2(n15108), 
        .ZN(n13190) );
  OAI221_X1 U15385 ( .B1(n15351), .B2(keyinput73), .C1(n15108), .C2(keyinput84), .A(n13190), .ZN(n13191) );
  NOR4_X1 U15386 ( .A1(n13194), .A2(n13193), .A3(n13192), .A4(n13191), .ZN(
        n13219) );
  INV_X1 U15387 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U15388 ( .A1(n13893), .A2(keyinput2), .B1(n12033), .B2(keyinput28), 
        .ZN(n13195) );
  OAI221_X1 U15389 ( .B1(n13893), .B2(keyinput2), .C1(n12033), .C2(keyinput28), 
        .A(n13195), .ZN(n13206) );
  INV_X1 U15390 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14878) );
  AOI22_X1 U15391 ( .A1(n13197), .A2(keyinput29), .B1(keyinput21), .B2(n14878), 
        .ZN(n13196) );
  OAI221_X1 U15392 ( .B1(n13197), .B2(keyinput29), .C1(n14878), .C2(keyinput21), .A(n13196), .ZN(n13205) );
  INV_X1 U15393 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U15394 ( .A1(n13200), .A2(keyinput94), .B1(keyinput86), .B2(n13199), 
        .ZN(n13198) );
  OAI221_X1 U15395 ( .B1(n13200), .B2(keyinput94), .C1(n13199), .C2(keyinput86), .A(n13198), .ZN(n13204) );
  INV_X1 U15396 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13202) );
  AOI22_X1 U15397 ( .A1(n13202), .A2(keyinput110), .B1(n13459), .B2(keyinput18), .ZN(n13201) );
  OAI221_X1 U15398 ( .B1(n13202), .B2(keyinput110), .C1(n13459), .C2(
        keyinput18), .A(n13201), .ZN(n13203) );
  NOR4_X1 U15399 ( .A1(n13206), .A2(n13205), .A3(n13204), .A4(n13203), .ZN(
        n13218) );
  AOI22_X1 U15400 ( .A1(n13208), .A2(keyinput113), .B1(n14532), .B2(keyinput57), .ZN(n13207) );
  OAI221_X1 U15401 ( .B1(n13208), .B2(keyinput113), .C1(n14532), .C2(
        keyinput57), .A(n13207), .ZN(n13216) );
  INV_X1 U15402 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15178) );
  AOI22_X1 U15403 ( .A1(n15178), .A2(keyinput30), .B1(n6720), .B2(keyinput72), 
        .ZN(n13209) );
  OAI221_X1 U15404 ( .B1(n15178), .B2(keyinput30), .C1(n6720), .C2(keyinput72), 
        .A(n13209), .ZN(n13215) );
  AOI22_X1 U15405 ( .A1(n13927), .A2(keyinput68), .B1(keyinput100), .B2(n13211), .ZN(n13210) );
  OAI221_X1 U15406 ( .B1(n13927), .B2(keyinput68), .C1(n13211), .C2(
        keyinput100), .A(n13210), .ZN(n13214) );
  INV_X1 U15407 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14959) );
  AOI22_X1 U15408 ( .A1(n14959), .A2(keyinput51), .B1(n13224), .B2(keyinput37), 
        .ZN(n13212) );
  OAI221_X1 U15409 ( .B1(n14959), .B2(keyinput51), .C1(n13224), .C2(keyinput37), .A(n13212), .ZN(n13213) );
  NOR4_X1 U15410 ( .A1(n13216), .A2(n13215), .A3(n13214), .A4(n13213), .ZN(
        n13217) );
  NAND4_X1 U15411 ( .A1(n13220), .A2(n13219), .A3(n13218), .A4(n13217), .ZN(
        n13278) );
  NOR4_X1 U15412 ( .A1(P3_REG1_REG_1__SCAN_IN), .A2(P3_REG1_REG_20__SCAN_IN), 
        .A3(n13221), .A4(n11009), .ZN(n13229) );
  NOR4_X1 U15413 ( .A1(SI_4_), .A2(P3_REG0_REG_3__SCAN_IN), .A3(
        P3_REG3_REG_2__SCAN_IN), .A4(n11006), .ZN(n13228) );
  NOR4_X1 U15414 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P3_DATAO_REG_30__SCAN_IN), 
        .A3(P3_DATAO_REG_25__SCAN_IN), .A4(P3_DATAO_REG_19__SCAN_IN), .ZN(
        n13227) );
  NOR4_X1 U15415 ( .A1(n13225), .A2(n13224), .A3(n13223), .A4(n13222), .ZN(
        n13226) );
  NAND4_X1 U15416 ( .A1(n13229), .A2(n13228), .A3(n13227), .A4(n13226), .ZN(
        n13261) );
  INV_X1 U15417 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n13230) );
  NOR4_X1 U15418 ( .A1(n13231), .A2(n13230), .A3(P3_IR_REG_25__SCAN_IN), .A4(
        P3_IR_REG_24__SCAN_IN), .ZN(n13256) );
  NOR4_X1 U15419 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(SI_14_), .A3(n13232), 
        .A4(n12033), .ZN(n13239) );
  NOR4_X1 U15420 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(P3_REG2_REG_8__SCAN_IN), 
        .A3(P3_REG0_REG_5__SCAN_IN), .A4(n13233), .ZN(n13238) );
  NOR4_X1 U15421 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .A3(n13234), .A4(n14567), .ZN(n13237) );
  NOR4_X1 U15422 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P2_DATAO_REG_12__SCAN_IN), 
        .A3(P2_DATAO_REG_1__SCAN_IN), .A4(n13235), .ZN(n13236) );
  NAND4_X1 U15423 ( .A1(n13239), .A2(n13238), .A3(n13237), .A4(n13236), .ZN(
        n13250) );
  NAND4_X1 U15424 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_REG2_REG_18__SCAN_IN), 
        .A3(P2_REG1_REG_6__SCAN_IN), .A4(P1_IR_REG_24__SCAN_IN), .ZN(n13243)
         );
  NAND4_X1 U15425 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .A3(P1_REG2_REG_26__SCAN_IN), .A4(P1_ADDR_REG_11__SCAN_IN), .ZN(n13242) );
  NAND4_X1 U15426 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), .A3(P2_REG2_REG_23__SCAN_IN), .A4(P1_REG1_REG_31__SCAN_IN), .ZN(n13241) );
  NAND4_X1 U15427 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(P1_REG2_REG_23__SCAN_IN), 
        .A3(P1_REG1_REG_21__SCAN_IN), .A4(P1_REG1_REG_8__SCAN_IN), .ZN(n13240)
         );
  NOR4_X1 U15428 ( .A1(n13243), .A2(n13242), .A3(n13241), .A4(n13240), .ZN(
        n13248) );
  NAND4_X1 U15429 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(P3_REG0_REG_25__SCAN_IN), .A3(P2_B_REG_SCAN_IN), .A4(P2_REG0_REG_12__SCAN_IN), .ZN(n13246) );
  NAND4_X1 U15430 ( .A1(SI_22_), .A2(P2_REG3_REG_25__SCAN_IN), .A3(
        P2_REG1_REG_28__SCAN_IN), .A4(P2_REG2_REG_30__SCAN_IN), .ZN(n13245) );
  NOR4_X1 U15431 ( .A1(n13246), .A2(n13245), .A3(n7832), .A4(n13244), .ZN(
        n13247) );
  NAND2_X1 U15432 ( .A1(n13248), .A2(n13247), .ZN(n13249) );
  NOR4_X1 U15433 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_1__SCAN_IN), 
        .A3(n13250), .A4(n13249), .ZN(n13254) );
  NAND4_X1 U15434 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(P1_REG0_REG_21__SCAN_IN), 
        .A3(P1_REG2_REG_0__SCAN_IN), .A4(P3_DATAO_REG_13__SCAN_IN), .ZN(n13252) );
  NAND4_X1 U15435 ( .A1(P3_REG1_REG_29__SCAN_IN), .A2(P2_REG1_REG_15__SCAN_IN), 
        .A3(P1_IR_REG_6__SCAN_IN), .A4(P3_DATAO_REG_18__SCAN_IN), .ZN(n13251)
         );
  NOR2_X1 U15436 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  NAND4_X1 U15437 ( .A1(n13256), .A2(n13255), .A3(n13254), .A4(n13253), .ZN(
        n13260) );
  NAND4_X1 U15438 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .A3(P1_D_REG_1__SCAN_IN), .A4(P1_ADDR_REG_16__SCAN_IN), .ZN(n13257) );
  NOR3_X1 U15439 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(P1_REG1_REG_14__SCAN_IN), 
        .A3(n13257), .ZN(n13258) );
  NAND3_X1 U15440 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .A3(n13258), .ZN(n13259) );
  NOR3_X1 U15441 ( .A1(n13261), .A2(n13260), .A3(n13259), .ZN(n13276) );
  NOR4_X1 U15442 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .A3(n6720), .A4(n7664), .ZN(n13275) );
  NOR4_X1 U15443 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_REG0_REG_11__SCAN_IN), .A4(P2_REG0_REG_23__SCAN_IN), .ZN(n13265) );
  NOR4_X1 U15444 ( .A1(P3_REG0_REG_28__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .A3(P2_REG1_REG_23__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n13264)
         );
  NOR4_X1 U15445 ( .A1(SI_21_), .A2(P2_REG2_REG_21__SCAN_IN), .A3(
        P2_REG0_REG_15__SCAN_IN), .A4(P2_DATAO_REG_31__SCAN_IN), .ZN(n13263)
         );
  NOR4_X1 U15446 ( .A1(SI_20_), .A2(P2_REG3_REG_3__SCAN_IN), .A3(
        P2_REG0_REG_0__SCAN_IN), .A4(P2_ADDR_REG_16__SCAN_IN), .ZN(n13262) );
  NAND4_X1 U15447 ( .A1(n13265), .A2(n13264), .A3(n13263), .A4(n13262), .ZN(
        n13268) );
  NAND2_X1 U15448 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n14640), .ZN(n14639) );
  NAND4_X1 U15449 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .A3(P1_REG0_REG_27__SCAN_IN), .A4(P1_REG2_REG_3__SCAN_IN), .ZN(n13267)
         );
  NAND4_X1 U15450 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P1_REG0_REG_3__SCAN_IN), 
        .A3(P1_REG1_REG_0__SCAN_IN), .A4(P1_ADDR_REG_18__SCAN_IN), .ZN(n13266)
         );
  NOR4_X1 U15451 ( .A1(n13268), .A2(n14639), .A3(n13267), .A4(n13266), .ZN(
        n13274) );
  NOR4_X1 U15452 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG1_REG_24__SCAN_IN), 
        .A3(P1_REG0_REG_20__SCAN_IN), .A4(P1_REG1_REG_29__SCAN_IN), .ZN(n13272) );
  NOR4_X1 U15453 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(P1_REG0_REG_30__SCAN_IN), 
        .A3(P2_ADDR_REG_8__SCAN_IN), .A4(P1_U3086), .ZN(n13271) );
  NOR4_X1 U15454 ( .A1(SI_25_), .A2(P1_IR_REG_16__SCAN_IN), .A3(
        P1_ADDR_REG_12__SCAN_IN), .A4(P3_ADDR_REG_9__SCAN_IN), .ZN(n13270) );
  NOR4_X1 U15455 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_REG3_REG_7__SCAN_IN), .A4(P1_REG0_REG_11__SCAN_IN), .ZN(n13269) );
  AND4_X1 U15456 ( .A1(n13272), .A2(n13271), .A3(n13270), .A4(n13269), .ZN(
        n13273) );
  NAND4_X1 U15457 ( .A1(n13276), .A2(n13275), .A3(n13274), .A4(n13273), .ZN(
        n13277) );
  XNOR2_X1 U15458 ( .A(n13278), .B(n13277), .ZN(n13279) );
  XNOR2_X1 U15459 ( .A(n13280), .B(n13279), .ZN(P3_U3214) );
  OAI21_X1 U15460 ( .B1(n13282), .B2(n6502), .A(n13281), .ZN(n13285) );
  AOI222_X1 U15461 ( .A1(n15341), .A2(n13285), .B1(n13284), .B2(n15324), .C1(
        n13283), .C2(n15326), .ZN(n13353) );
  INV_X1 U15462 ( .A(n13286), .ZN(n13287) );
  AOI21_X1 U15463 ( .B1(n6502), .B2(n13288), .A(n13287), .ZN(n13351) );
  AOI22_X1 U15464 ( .A1(n15398), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15395), 
        .B2(n13289), .ZN(n13290) );
  OAI21_X1 U15465 ( .B1(n13291), .B2(n13304), .A(n13290), .ZN(n13292) );
  AOI21_X1 U15466 ( .B1(n13351), .B2(n13306), .A(n13292), .ZN(n13293) );
  OAI21_X1 U15467 ( .B1(n13353), .B2(n15398), .A(n13293), .ZN(P3_U3215) );
  AOI21_X1 U15468 ( .B1(n13294), .B2(n13300), .A(n15388), .ZN(n13299) );
  OAI22_X1 U15469 ( .A1(n13296), .A2(n15381), .B1(n13295), .B2(n15382), .ZN(
        n13297) );
  AOI21_X1 U15470 ( .B1(n13299), .B2(n13298), .A(n13297), .ZN(n13356) );
  XNOR2_X1 U15471 ( .A(n13301), .B(n13300), .ZN(n13354) );
  AOI22_X1 U15472 ( .A1(n15398), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15395), 
        .B2(n13302), .ZN(n13303) );
  OAI21_X1 U15473 ( .B1(n13357), .B2(n13304), .A(n13303), .ZN(n13305) );
  AOI21_X1 U15474 ( .B1(n13354), .B2(n13306), .A(n13305), .ZN(n13307) );
  OAI21_X1 U15475 ( .B1(n13356), .B2(n15398), .A(n13307), .ZN(P3_U3216) );
  INV_X1 U15476 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13310) );
  AOI21_X1 U15477 ( .B1(n15426), .B2(n13309), .A(n13308), .ZN(n13369) );
  MUX2_X1 U15478 ( .A(n13310), .B(n13369), .S(n15438), .Z(n13311) );
  OAI21_X1 U15479 ( .B1(n13372), .B2(n13339), .A(n13311), .ZN(P3_U3485) );
  NAND2_X1 U15480 ( .A1(n13312), .A2(n15411), .ZN(n13313) );
  NAND2_X1 U15481 ( .A1(n13314), .A2(n13313), .ZN(n13373) );
  INV_X1 U15482 ( .A(n13373), .ZN(n13316) );
  MUX2_X1 U15483 ( .A(n13316), .B(n13315), .S(n15439), .Z(n13317) );
  OAI21_X1 U15484 ( .B1(n13318), .B2(n13339), .A(n13317), .ZN(P3_U3484) );
  INV_X1 U15485 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13321) );
  AOI21_X1 U15486 ( .B1(n15426), .B2(n13320), .A(n13319), .ZN(n13377) );
  MUX2_X1 U15487 ( .A(n13321), .B(n13377), .S(n15438), .Z(n13322) );
  OAI21_X1 U15488 ( .B1(n13380), .B2(n13339), .A(n13322), .ZN(P3_U3483) );
  INV_X1 U15489 ( .A(n13323), .ZN(n13324) );
  NAND2_X1 U15490 ( .A1(n13324), .A2(n15426), .ZN(n13325) );
  NAND2_X1 U15491 ( .A1(n13326), .A2(n13325), .ZN(n13381) );
  MUX2_X1 U15492 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13381), .S(n15438), .Z(
        n13327) );
  INV_X1 U15493 ( .A(n13327), .ZN(n13328) );
  OAI21_X1 U15494 ( .B1(n13329), .B2(n13339), .A(n13328), .ZN(P3_U3482) );
  INV_X1 U15495 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13332) );
  AOI21_X1 U15496 ( .B1(n15411), .B2(n13331), .A(n13330), .ZN(n13385) );
  MUX2_X1 U15497 ( .A(n13332), .B(n13385), .S(n15438), .Z(n13333) );
  OAI21_X1 U15498 ( .B1(n13388), .B2(n13339), .A(n13333), .ZN(P3_U3481) );
  INV_X1 U15499 ( .A(n13334), .ZN(n13335) );
  AOI21_X1 U15500 ( .B1(n15411), .B2(n13336), .A(n13335), .ZN(n13389) );
  MUX2_X1 U15501 ( .A(n13337), .B(n13389), .S(n15438), .Z(n13338) );
  OAI21_X1 U15502 ( .B1(n13393), .B2(n13339), .A(n13338), .ZN(P3_U3480) );
  NAND2_X1 U15503 ( .A1(n13340), .A2(n15411), .ZN(n13341) );
  NAND2_X1 U15504 ( .A1(n13342), .A2(n13341), .ZN(n13394) );
  MUX2_X1 U15505 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13394), .S(n15438), .Z(
        n13343) );
  AOI21_X1 U15506 ( .B1(n10409), .B2(n13396), .A(n13343), .ZN(n13344) );
  INV_X1 U15507 ( .A(n13344), .ZN(P3_U3479) );
  NAND2_X1 U15508 ( .A1(n13345), .A2(n15411), .ZN(n13346) );
  NAND2_X1 U15509 ( .A1(n13347), .A2(n13346), .ZN(n13398) );
  MUX2_X1 U15510 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13398), .S(n15438), .Z(
        n13348) );
  AOI21_X1 U15511 ( .B1(n10409), .B2(n13400), .A(n13348), .ZN(n13349) );
  INV_X1 U15512 ( .A(n13349), .ZN(P3_U3478) );
  AOI22_X1 U15513 ( .A1(n13351), .A2(n15411), .B1(n15410), .B2(n13350), .ZN(
        n13352) );
  NAND2_X1 U15514 ( .A1(n13353), .A2(n13352), .ZN(n13403) );
  MUX2_X1 U15515 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13403), .S(n15438), .Z(
        P3_U3477) );
  NAND2_X1 U15516 ( .A1(n13354), .A2(n15411), .ZN(n13355) );
  OAI211_X1 U15517 ( .C1(n13357), .C2(n15346), .A(n13356), .B(n13355), .ZN(
        n13404) );
  MUX2_X1 U15518 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13404), .S(n15438), .Z(
        P3_U3476) );
  AOI22_X1 U15519 ( .A1(n13359), .A2(n15411), .B1(n15410), .B2(n13358), .ZN(
        n13360) );
  NAND2_X1 U15520 ( .A1(n13361), .A2(n13360), .ZN(n13405) );
  MUX2_X1 U15521 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13405), .S(n15438), .Z(
        P3_U3475) );
  NAND2_X1 U15522 ( .A1(n13362), .A2(n15411), .ZN(n13363) );
  OAI211_X1 U15523 ( .C1(n13365), .C2(n15346), .A(n13364), .B(n13363), .ZN(
        n13406) );
  MUX2_X1 U15524 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13406), .S(n15438), .Z(
        P3_U3474) );
  MUX2_X1 U15525 ( .A(n13370), .B(n13369), .S(n15430), .Z(n13371) );
  OAI21_X1 U15526 ( .B1(n13372), .B2(n13392), .A(n13371), .ZN(P3_U3453) );
  MUX2_X1 U15527 ( .A(n13373), .B(P3_REG0_REG_25__SCAN_IN), .S(n15428), .Z(
        n13374) );
  AOI21_X1 U15528 ( .B1(n13401), .B2(n13375), .A(n13374), .ZN(n13376) );
  INV_X1 U15529 ( .A(n13376), .ZN(P3_U3452) );
  MUX2_X1 U15530 ( .A(n13378), .B(n13377), .S(n15430), .Z(n13379) );
  OAI21_X1 U15531 ( .B1(n13380), .B2(n13392), .A(n13379), .ZN(P3_U3451) );
  MUX2_X1 U15532 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13381), .S(n15430), .Z(
        n13382) );
  AOI21_X1 U15533 ( .B1(n13401), .B2(n13383), .A(n13382), .ZN(n13384) );
  INV_X1 U15534 ( .A(n13384), .ZN(P3_U3450) );
  MUX2_X1 U15535 ( .A(n13386), .B(n13385), .S(n15430), .Z(n13387) );
  OAI21_X1 U15536 ( .B1(n13388), .B2(n13392), .A(n13387), .ZN(P3_U3449) );
  INV_X1 U15537 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13390) );
  MUX2_X1 U15538 ( .A(n13390), .B(n13389), .S(n15430), .Z(n13391) );
  OAI21_X1 U15539 ( .B1(n13393), .B2(n13392), .A(n13391), .ZN(P3_U3448) );
  MUX2_X1 U15540 ( .A(n13394), .B(P3_REG0_REG_20__SCAN_IN), .S(n15428), .Z(
        n13395) );
  AOI21_X1 U15541 ( .B1(n13401), .B2(n13396), .A(n13395), .ZN(n13397) );
  INV_X1 U15542 ( .A(n13397), .ZN(P3_U3447) );
  MUX2_X1 U15543 ( .A(n13398), .B(P3_REG0_REG_19__SCAN_IN), .S(n15428), .Z(
        n13399) );
  AOI21_X1 U15544 ( .B1(n13401), .B2(n13400), .A(n13399), .ZN(n13402) );
  INV_X1 U15545 ( .A(n13402), .ZN(P3_U3446) );
  MUX2_X1 U15546 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13403), .S(n15430), .Z(
        P3_U3444) );
  MUX2_X1 U15547 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13404), .S(n15430), .Z(
        P3_U3441) );
  MUX2_X1 U15548 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13405), .S(n15430), .Z(
        P3_U3438) );
  MUX2_X1 U15549 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13406), .S(n15430), .Z(
        P3_U3435) );
  MUX2_X1 U15550 ( .A(P3_D_REG_1__SCAN_IN), .B(n13407), .S(n13408), .Z(
        P3_U3377) );
  MUX2_X1 U15551 ( .A(P3_D_REG_0__SCAN_IN), .B(n13409), .S(n13408), .Z(
        P3_U3376) );
  NAND2_X1 U15552 ( .A1(n13411), .A2(n13410), .ZN(n13415) );
  INV_X1 U15553 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13413) );
  NAND4_X1 U15554 ( .A1(n6707), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n13413), .ZN(n13414) );
  OAI211_X1 U15555 ( .C1(n13416), .C2(n13423), .A(n13415), .B(n13414), .ZN(
        P3_U3264) );
  INV_X1 U15556 ( .A(n13417), .ZN(n13418) );
  OAI222_X1 U15557 ( .A1(n13423), .A2(n13422), .B1(P3_U3151), .B2(n13420), 
        .C1(n13419), .C2(n13418), .ZN(P3_U3267) );
  XNOR2_X1 U15558 ( .A(n13425), .B(n13424), .ZN(n13430) );
  AOI22_X1 U15559 ( .A1(n13525), .A2(n13509), .B1(n13510), .B2(n13523), .ZN(
        n13648) );
  OAI22_X1 U15560 ( .A1(n13491), .A2(n13648), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13426), .ZN(n13427) );
  AOI21_X1 U15561 ( .B1(n13652), .B2(n13493), .A(n13427), .ZN(n13429) );
  NAND2_X1 U15562 ( .A1(n13809), .A2(n13518), .ZN(n13428) );
  OAI211_X1 U15563 ( .C1(n13430), .C2(n13520), .A(n13429), .B(n13428), .ZN(
        P2_U3186) );
  NAND2_X1 U15564 ( .A1(n13484), .A2(n13528), .ZN(n13434) );
  OR2_X1 U15565 ( .A1(n13520), .A2(n13431), .ZN(n13433) );
  MUX2_X1 U15566 ( .A(n13434), .B(n13433), .S(n13432), .Z(n13438) );
  AOI22_X1 U15567 ( .A1(n13527), .A2(n13510), .B1(n13509), .B2(n13529), .ZN(
        n13708) );
  OAI22_X1 U15568 ( .A1(n13491), .A2(n13708), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13435), .ZN(n13436) );
  AOI21_X1 U15569 ( .B1(n13714), .B2(n13493), .A(n13436), .ZN(n13437) );
  OAI211_X1 U15570 ( .C1(n7264), .C2(n8883), .A(n13438), .B(n13437), .ZN(
        P2_U3188) );
  NAND2_X1 U15571 ( .A1(n13440), .A2(n13439), .ZN(n13442) );
  XOR2_X1 U15572 ( .A(n13442), .B(n13441), .Z(n13447) );
  NOR2_X1 U15573 ( .A1(n13515), .A2(n13775), .ZN(n13445) );
  AND2_X1 U15574 ( .A1(n13533), .A2(n13509), .ZN(n13443) );
  AOI21_X1 U15575 ( .B1(n13531), .B2(n13510), .A(n13443), .ZN(n13768) );
  NAND2_X1 U15576 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13609)
         );
  OAI21_X1 U15577 ( .B1(n13768), .B2(n13491), .A(n13609), .ZN(n13444) );
  AOI211_X1 U15578 ( .C1(n13853), .C2(n13518), .A(n13445), .B(n13444), .ZN(
        n13446) );
  OAI21_X1 U15579 ( .B1(n13447), .B2(n13520), .A(n13446), .ZN(P2_U3191) );
  XNOR2_X1 U15580 ( .A(n13448), .B(n13449), .ZN(n13456) );
  INV_X1 U15581 ( .A(n13743), .ZN(n13453) );
  OAI22_X1 U15582 ( .A1(n13451), .A2(n13469), .B1(n13450), .B2(n13468), .ZN(
        n13739) );
  AOI22_X1 U15583 ( .A1(n13739), .A2(n13513), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13452) );
  OAI21_X1 U15584 ( .B1(n13453), .B2(n13515), .A(n13452), .ZN(n13454) );
  AOI21_X1 U15585 ( .B1(n13744), .B2(n13518), .A(n13454), .ZN(n13455) );
  OAI21_X1 U15586 ( .B1(n13456), .B2(n13520), .A(n13455), .ZN(P2_U3195) );
  XNOR2_X1 U15587 ( .A(n13457), .B(n13458), .ZN(n13463) );
  AOI22_X1 U15588 ( .A1(n13509), .A2(n13527), .B1(n13525), .B2(n13510), .ZN(
        n13680) );
  OAI22_X1 U15589 ( .A1(n13491), .A2(n13680), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13459), .ZN(n13460) );
  AOI21_X1 U15590 ( .B1(n13685), .B2(n13493), .A(n13460), .ZN(n13462) );
  NAND2_X1 U15591 ( .A1(n13682), .A2(n13518), .ZN(n13461) );
  OAI211_X1 U15592 ( .C1(n13463), .C2(n13520), .A(n13462), .B(n13461), .ZN(
        P2_U3197) );
  XNOR2_X1 U15593 ( .A(n13465), .B(n13464), .ZN(n13474) );
  INV_X1 U15594 ( .A(n13466), .ZN(n13699) );
  OAI22_X1 U15595 ( .A1(n13470), .A2(n13469), .B1(n13468), .B2(n13467), .ZN(
        n13694) );
  AOI22_X1 U15596 ( .A1(n13513), .A2(n13694), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13471) );
  OAI21_X1 U15597 ( .B1(n13699), .B2(n13515), .A(n13471), .ZN(n13472) );
  AOI21_X1 U15598 ( .B1(n13703), .B2(n13518), .A(n13472), .ZN(n13473) );
  OAI21_X1 U15599 ( .B1(n13474), .B2(n13520), .A(n13473), .ZN(P2_U3201) );
  INV_X1 U15600 ( .A(n13475), .ZN(n13476) );
  AOI21_X1 U15601 ( .B1(n13478), .B2(n13477), .A(n13476), .ZN(n13483) );
  AOI22_X1 U15602 ( .A1(n13530), .A2(n13510), .B1(n13509), .B2(n13532), .ZN(
        n13752) );
  INV_X1 U15603 ( .A(n13752), .ZN(n13479) );
  AOI22_X1 U15604 ( .A1(n13479), .A2(n13513), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13480) );
  OAI21_X1 U15605 ( .B1(n13758), .B2(n13515), .A(n13480), .ZN(n13481) );
  AOI21_X1 U15606 ( .B1(n13757), .B2(n13518), .A(n13481), .ZN(n13482) );
  OAI21_X1 U15607 ( .B1(n13483), .B2(n13520), .A(n13482), .ZN(P2_U3205) );
  INV_X1 U15608 ( .A(n13836), .ZN(n13728) );
  NAND2_X1 U15609 ( .A1(n13484), .A2(n13529), .ZN(n13488) );
  OR2_X1 U15610 ( .A1(n13520), .A2(n13485), .ZN(n13487) );
  MUX2_X1 U15611 ( .A(n13488), .B(n13487), .S(n13486), .Z(n13495) );
  AND2_X1 U15612 ( .A1(n13510), .A2(n13528), .ZN(n13489) );
  AOI21_X1 U15613 ( .B1(n13530), .B2(n13509), .A(n13489), .ZN(n13721) );
  OAI22_X1 U15614 ( .A1(n13721), .A2(n13491), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13490), .ZN(n13492) );
  AOI21_X1 U15615 ( .B1(n13726), .B2(n13493), .A(n13492), .ZN(n13494) );
  OAI211_X1 U15616 ( .C1(n13728), .C2(n8883), .A(n13495), .B(n13494), .ZN(
        P2_U3207) );
  AOI21_X1 U15617 ( .B1(n13497), .B2(n13496), .A(n13520), .ZN(n13499) );
  NAND2_X1 U15618 ( .A1(n13499), .A2(n13498), .ZN(n13504) );
  NAND2_X1 U15619 ( .A1(n13532), .A2(n13510), .ZN(n13501) );
  NAND2_X1 U15620 ( .A1(n13534), .A2(n13509), .ZN(n13500) );
  NAND2_X1 U15621 ( .A1(n13501), .A2(n13500), .ZN(n13782) );
  AND2_X1 U15622 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13572) );
  NOR2_X1 U15623 ( .A1(n13515), .A2(n13786), .ZN(n13502) );
  AOI211_X1 U15624 ( .C1(n13513), .C2(n13782), .A(n13572), .B(n13502), .ZN(
        n13503) );
  OAI211_X1 U15625 ( .C1(n6988), .C2(n8883), .A(n13504), .B(n13503), .ZN(
        P2_U3210) );
  INV_X1 U15626 ( .A(n13505), .ZN(n13506) );
  AOI21_X1 U15627 ( .B1(n13508), .B2(n13507), .A(n13506), .ZN(n13521) );
  INV_X1 U15628 ( .A(n13666), .ZN(n13516) );
  NAND2_X1 U15629 ( .A1(n13509), .A2(n13526), .ZN(n13512) );
  NAND2_X1 U15630 ( .A1(n13510), .A2(n13524), .ZN(n13511) );
  NAND2_X1 U15631 ( .A1(n13512), .A2(n13511), .ZN(n13661) );
  AOI22_X1 U15632 ( .A1(n13513), .A2(n13661), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13514) );
  OAI21_X1 U15633 ( .B1(n13516), .B2(n13515), .A(n13514), .ZN(n13517) );
  AOI21_X1 U15634 ( .B1(n13815), .B2(n13518), .A(n13517), .ZN(n13519) );
  OAI21_X1 U15635 ( .B1(n13521), .B2(n13520), .A(n13519), .ZN(P2_U3212) );
  MUX2_X1 U15636 ( .A(n13614), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13550), .Z(
        P2_U3562) );
  MUX2_X1 U15637 ( .A(n9894), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13550), .Z(
        P2_U3561) );
  MUX2_X1 U15638 ( .A(n13522), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13550), .Z(
        P2_U3560) );
  MUX2_X1 U15639 ( .A(n13523), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13550), .Z(
        P2_U3559) );
  MUX2_X1 U15640 ( .A(n13524), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13550), .Z(
        P2_U3558) );
  MUX2_X1 U15641 ( .A(n13525), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13550), .Z(
        P2_U3557) );
  MUX2_X1 U15642 ( .A(n13526), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13550), .Z(
        P2_U3556) );
  MUX2_X1 U15643 ( .A(n13527), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13550), .Z(
        P2_U3555) );
  MUX2_X1 U15644 ( .A(n13528), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13550), .Z(
        P2_U3554) );
  MUX2_X1 U15645 ( .A(n13529), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13550), .Z(
        P2_U3553) );
  MUX2_X1 U15646 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13530), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15647 ( .A(n13531), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13550), .Z(
        P2_U3551) );
  MUX2_X1 U15648 ( .A(n13532), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13550), .Z(
        P2_U3550) );
  MUX2_X1 U15649 ( .A(n13533), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13550), .Z(
        P2_U3549) );
  MUX2_X1 U15650 ( .A(n13534), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13550), .Z(
        P2_U3548) );
  MUX2_X1 U15651 ( .A(n13535), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13550), .Z(
        P2_U3547) );
  MUX2_X1 U15652 ( .A(n13536), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13550), .Z(
        P2_U3546) );
  MUX2_X1 U15653 ( .A(n13537), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13550), .Z(
        P2_U3545) );
  MUX2_X1 U15654 ( .A(n13538), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13550), .Z(
        P2_U3544) );
  MUX2_X1 U15655 ( .A(n13539), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13550), .Z(
        P2_U3543) );
  MUX2_X1 U15656 ( .A(n13540), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13550), .Z(
        P2_U3542) );
  MUX2_X1 U15657 ( .A(n13541), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13550), .Z(
        P2_U3541) );
  MUX2_X1 U15658 ( .A(n13542), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13550), .Z(
        P2_U3540) );
  MUX2_X1 U15659 ( .A(n13543), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13550), .Z(
        P2_U3539) );
  MUX2_X1 U15660 ( .A(n13544), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13550), .Z(
        P2_U3538) );
  MUX2_X1 U15661 ( .A(n13545), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13550), .Z(
        P2_U3537) );
  MUX2_X1 U15662 ( .A(n13546), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13550), .Z(
        P2_U3536) );
  MUX2_X1 U15663 ( .A(n13547), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13550), .Z(
        P2_U3535) );
  MUX2_X1 U15664 ( .A(n6898), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13550), .Z(
        P2_U3534) );
  MUX2_X1 U15665 ( .A(n13549), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13550), .Z(
        P2_U3533) );
  MUX2_X1 U15666 ( .A(n13551), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13550), .Z(
        P2_U3532) );
  OAI21_X1 U15667 ( .B1(n13554), .B2(n13553), .A(n13552), .ZN(n13559) );
  OAI21_X1 U15668 ( .B1(n13557), .B2(n13556), .A(n13555), .ZN(n13558) );
  AOI22_X1 U15669 ( .A1(n13605), .A2(n13559), .B1(n15129), .B2(n13558), .ZN(
        n13564) );
  NAND2_X1 U15670 ( .A1(n15141), .A2(n13560), .ZN(n13562) );
  NAND2_X1 U15671 ( .A1(n15056), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n13561) );
  NAND4_X1 U15672 ( .A1(n13564), .A2(n13563), .A3(n13562), .A4(n13561), .ZN(
        P2_U3226) );
  INV_X1 U15673 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14781) );
  NOR2_X1 U15674 ( .A1(n15101), .A2(n14781), .ZN(n13566) );
  AOI21_X1 U15675 ( .B1(n15101), .B2(n14781), .A(n13566), .ZN(n15095) );
  NOR2_X1 U15676 ( .A1(n13567), .A2(n13580), .ZN(n13568) );
  XNOR2_X1 U15677 ( .A(n15125), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15116) );
  XNOR2_X1 U15678 ( .A(n15140), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15136) );
  NOR2_X1 U15679 ( .A1(n15137), .A2(n15136), .ZN(n15134) );
  INV_X1 U15680 ( .A(n13602), .ZN(n13570) );
  OAI211_X1 U15681 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13571), .A(n13570), 
        .B(n13605), .ZN(n13595) );
  AOI21_X1 U15682 ( .B1(n15056), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n13572), 
        .ZN(n13594) );
  NAND2_X1 U15683 ( .A1(n13573), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n13574) );
  NAND2_X1 U15684 ( .A1(n13575), .A2(n13574), .ZN(n13576) );
  NOR2_X1 U15685 ( .A1(n13576), .A2(n15101), .ZN(n13577) );
  INV_X1 U15686 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n15098) );
  NOR2_X1 U15687 ( .A1(n13579), .A2(n13580), .ZN(n13581) );
  INV_X1 U15688 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n15105) );
  NOR2_X1 U15689 ( .A1(n13581), .A2(n15104), .ZN(n15122) );
  INV_X1 U15690 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13583) );
  NAND2_X1 U15691 ( .A1(n15125), .A2(n13583), .ZN(n13582) );
  OAI21_X1 U15692 ( .B1(n15125), .B2(n13583), .A(n13582), .ZN(n13584) );
  INV_X1 U15693 ( .A(n13584), .ZN(n15121) );
  NAND2_X1 U15694 ( .A1(n15125), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13585) );
  NAND2_X1 U15695 ( .A1(n15118), .A2(n13585), .ZN(n15132) );
  NAND2_X1 U15696 ( .A1(n13587), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13586) );
  OAI21_X1 U15697 ( .B1(n13587), .B2(P2_REG2_REG_17__SCAN_IN), .A(n13586), 
        .ZN(n15131) );
  NAND2_X1 U15698 ( .A1(n15132), .A2(n15131), .ZN(n15130) );
  NAND2_X1 U15699 ( .A1(n15140), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13588) );
  NAND2_X1 U15700 ( .A1(n15130), .A2(n13588), .ZN(n13597) );
  XOR2_X1 U15701 ( .A(n13596), .B(n13597), .Z(n13590) );
  NAND2_X1 U15702 ( .A1(n13590), .A2(n13589), .ZN(n13599) );
  OAI21_X1 U15703 ( .B1(n13590), .B2(n13589), .A(n13599), .ZN(n13591) );
  NAND2_X1 U15704 ( .A1(n13591), .A2(n15129), .ZN(n13593) );
  NAND2_X1 U15705 ( .A1(n15141), .A2(n13596), .ZN(n13592) );
  NAND4_X1 U15706 ( .A1(n13595), .A2(n13594), .A3(n13593), .A4(n13592), .ZN(
        P2_U3232) );
  OR2_X1 U15707 ( .A1(n13597), .A2(n13596), .ZN(n13598) );
  NAND2_X1 U15708 ( .A1(n13599), .A2(n13598), .ZN(n13600) );
  XNOR2_X1 U15709 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13600), .ZN(n13606) );
  XNOR2_X1 U15710 ( .A(n13603), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13604) );
  AOI22_X1 U15711 ( .A1(n13606), .A2(n15129), .B1(n13605), .B2(n13604), .ZN(
        n13608) );
  NAND2_X1 U15712 ( .A1(n7632), .A2(n13614), .ZN(n13800) );
  NOR2_X1 U15713 ( .A1(n15174), .A2(n13800), .ZN(n13620) );
  NOR2_X1 U15714 ( .A1(n13612), .A2(n15152), .ZN(n13615) );
  AOI211_X1 U15715 ( .C1(n15149), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13620), 
        .B(n13615), .ZN(n13616) );
  OAI21_X1 U15716 ( .B1(n13797), .B2(n13747), .A(n13616), .ZN(P2_U3234) );
  OAI211_X1 U15717 ( .C1(n13880), .C2(n13618), .A(n13742), .B(n13617), .ZN(
        n13801) );
  NOR2_X1 U15718 ( .A1(n13880), .A2(n15152), .ZN(n13619) );
  AOI211_X1 U15719 ( .C1(n15174), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13620), 
        .B(n13619), .ZN(n13621) );
  OAI21_X1 U15720 ( .B1(n13747), .B2(n13801), .A(n13621), .ZN(P2_U3235) );
  AOI22_X1 U15721 ( .A1(n15149), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n13624), 
        .B2(n15163), .ZN(n13625) );
  OAI21_X1 U15722 ( .B1(n6993), .B2(n15152), .A(n13625), .ZN(n13626) );
  AOI21_X1 U15723 ( .B1(n13627), .B2(n15169), .A(n13626), .ZN(n13628) );
  OR2_X1 U15724 ( .A1(n13630), .A2(n13629), .ZN(n13631) );
  NAND2_X1 U15725 ( .A1(n13632), .A2(n13631), .ZN(n13806) );
  INV_X1 U15726 ( .A(n13636), .ZN(n13637) );
  INV_X1 U15727 ( .A(n13805), .ZN(n13642) );
  AOI21_X1 U15728 ( .B1(n13643), .B2(n6610), .A(n11852), .ZN(n13639) );
  NAND2_X1 U15729 ( .A1(n13639), .A2(n13638), .ZN(n13804) );
  OAI22_X1 U15730 ( .A1(n13804), .A2(n13700), .B1(n13774), .B2(n13640), .ZN(
        n13641) );
  OAI21_X1 U15731 ( .B1(n13642), .B2(n13641), .A(n11353), .ZN(n13645) );
  AOI22_X1 U15732 ( .A1(n13643), .A2(n15170), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n15174), .ZN(n13644) );
  OAI211_X1 U15733 ( .C1(n13793), .C2(n13806), .A(n13645), .B(n13644), .ZN(
        P2_U3237) );
  XNOR2_X1 U15734 ( .A(n13647), .B(n13646), .ZN(n13650) );
  INV_X1 U15735 ( .A(n13648), .ZN(n13649) );
  AOI21_X1 U15736 ( .B1(n13650), .B2(n15161), .A(n13649), .ZN(n13812) );
  AOI21_X1 U15737 ( .B1(n13809), .B2(n13664), .A(n11852), .ZN(n13651) );
  NAND2_X1 U15738 ( .A1(n13651), .A2(n6610), .ZN(n13810) );
  AOI22_X1 U15739 ( .A1(n15149), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13652), 
        .B2(n15163), .ZN(n13654) );
  NAND2_X1 U15740 ( .A1(n13809), .A2(n15170), .ZN(n13653) );
  OAI211_X1 U15741 ( .C1(n13810), .C2(n13747), .A(n13654), .B(n13653), .ZN(
        n13655) );
  INV_X1 U15742 ( .A(n13655), .ZN(n13659) );
  OR2_X1 U15743 ( .A1(n13657), .A2(n13656), .ZN(n13808) );
  NAND3_X1 U15744 ( .A1(n13808), .A2(n15168), .A3(n13807), .ZN(n13658) );
  OAI211_X1 U15745 ( .C1(n13812), .C2(n15174), .A(n13659), .B(n13658), .ZN(
        P2_U3238) );
  XNOR2_X1 U15746 ( .A(n13660), .B(n13669), .ZN(n13662) );
  AOI21_X1 U15747 ( .B1(n13662), .B2(n15161), .A(n13661), .ZN(n13817) );
  INV_X1 U15748 ( .A(n13663), .ZN(n13684) );
  INV_X1 U15749 ( .A(n13664), .ZN(n13665) );
  AOI211_X1 U15750 ( .C1(n13815), .C2(n13684), .A(n11852), .B(n13665), .ZN(
        n13814) );
  AOI22_X1 U15751 ( .A1(n15174), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13666), 
        .B2(n15163), .ZN(n13667) );
  OAI21_X1 U15752 ( .B1(n13668), .B2(n15152), .A(n13667), .ZN(n13673) );
  INV_X1 U15753 ( .A(n13669), .ZN(n13670) );
  XNOR2_X1 U15754 ( .A(n13671), .B(n13670), .ZN(n13818) );
  NOR2_X1 U15755 ( .A1(n13818), .A2(n13793), .ZN(n13672) );
  AOI211_X1 U15756 ( .C1(n13814), .C2(n15169), .A(n13673), .B(n13672), .ZN(
        n13674) );
  OAI21_X1 U15757 ( .B1(n15174), .B2(n13817), .A(n13674), .ZN(P2_U3239) );
  XNOR2_X1 U15758 ( .A(n13675), .B(n13677), .ZN(n13821) );
  INV_X1 U15759 ( .A(n13821), .ZN(n13690) );
  OAI21_X1 U15760 ( .B1(n13678), .B2(n13677), .A(n13676), .ZN(n13679) );
  NAND2_X1 U15761 ( .A1(n13679), .A2(n15161), .ZN(n13681) );
  NAND2_X1 U15762 ( .A1(n13681), .A2(n13680), .ZN(n13819) );
  INV_X1 U15763 ( .A(n13682), .ZN(n13887) );
  NAND2_X1 U15764 ( .A1(n13682), .A2(n13697), .ZN(n13683) );
  NAND2_X1 U15765 ( .A1(n13820), .A2(n15169), .ZN(n13687) );
  AOI22_X1 U15766 ( .A1(n15174), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13685), 
        .B2(n15163), .ZN(n13686) );
  OAI211_X1 U15767 ( .C1(n13887), .C2(n15152), .A(n13687), .B(n13686), .ZN(
        n13688) );
  AOI21_X1 U15768 ( .B1(n13819), .B2(n11353), .A(n13688), .ZN(n13689) );
  OAI21_X1 U15769 ( .B1(n13690), .B2(n13793), .A(n13689), .ZN(P2_U3240) );
  XNOR2_X1 U15770 ( .A(n13691), .B(n13693), .ZN(n13824) );
  OAI21_X1 U15771 ( .B1(n6654), .B2(n13693), .A(n13692), .ZN(n13695) );
  AOI21_X1 U15772 ( .B1(n13695), .B2(n15161), .A(n13694), .ZN(n13696) );
  OAI21_X1 U15773 ( .B1(n13824), .B2(n9942), .A(n13696), .ZN(n13825) );
  INV_X1 U15774 ( .A(n13697), .ZN(n13698) );
  AOI211_X1 U15775 ( .C1(n13703), .C2(n6985), .A(n11852), .B(n13698), .ZN(
        n13826) );
  INV_X1 U15776 ( .A(n13826), .ZN(n13701) );
  OAI22_X1 U15777 ( .A1(n13701), .A2(n13700), .B1(n13774), .B2(n13699), .ZN(
        n13702) );
  OAI21_X1 U15778 ( .B1(n13825), .B2(n13702), .A(n11353), .ZN(n13705) );
  AOI22_X1 U15779 ( .A1(n13703), .A2(n15170), .B1(n15149), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n13704) );
  OAI211_X1 U15780 ( .C1(n13824), .C2(n13706), .A(n13705), .B(n13704), .ZN(
        P2_U3241) );
  XNOR2_X1 U15781 ( .A(n13707), .B(n13710), .ZN(n13709) );
  OAI21_X1 U15782 ( .B1(n13709), .B2(n13769), .A(n13708), .ZN(n13830) );
  INV_X1 U15783 ( .A(n13830), .ZN(n13719) );
  XNOR2_X1 U15784 ( .A(n13711), .B(n13710), .ZN(n13832) );
  AOI211_X1 U15785 ( .C1(n13713), .C2(n13724), .A(n11852), .B(n13712), .ZN(
        n13831) );
  NAND2_X1 U15786 ( .A1(n13831), .A2(n15169), .ZN(n13716) );
  AOI22_X1 U15787 ( .A1(n15174), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13714), 
        .B2(n15163), .ZN(n13715) );
  OAI211_X1 U15788 ( .C1(n7264), .C2(n15152), .A(n13716), .B(n13715), .ZN(
        n13717) );
  AOI21_X1 U15789 ( .B1(n15168), .B2(n13832), .A(n13717), .ZN(n13718) );
  OAI21_X1 U15790 ( .B1(n13719), .B2(n15149), .A(n13718), .ZN(P2_U3242) );
  XNOR2_X1 U15791 ( .A(n13720), .B(n13730), .ZN(n13723) );
  INV_X1 U15792 ( .A(n13721), .ZN(n13722) );
  AOI21_X1 U15793 ( .B1(n13723), .B2(n15161), .A(n13722), .ZN(n13838) );
  INV_X1 U15794 ( .A(n13724), .ZN(n13725) );
  AOI211_X1 U15795 ( .C1(n13836), .C2(n13741), .A(n11852), .B(n13725), .ZN(
        n13835) );
  AOI22_X1 U15796 ( .A1(n15174), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13726), 
        .B2(n15163), .ZN(n13727) );
  OAI21_X1 U15797 ( .B1(n13728), .B2(n15152), .A(n13727), .ZN(n13733) );
  OAI21_X1 U15798 ( .B1(n13731), .B2(n13730), .A(n13729), .ZN(n13839) );
  NOR2_X1 U15799 ( .A1(n13839), .A2(n13793), .ZN(n13732) );
  AOI211_X1 U15800 ( .C1(n13835), .C2(n15169), .A(n13733), .B(n13732), .ZN(
        n13734) );
  OAI21_X1 U15801 ( .B1(n15149), .B2(n13838), .A(n13734), .ZN(P2_U3243) );
  XNOR2_X1 U15802 ( .A(n13735), .B(n13737), .ZN(n13842) );
  AOI21_X1 U15803 ( .B1(n13751), .B2(n13754), .A(n13736), .ZN(n13738) );
  XNOR2_X1 U15804 ( .A(n13738), .B(n13737), .ZN(n13740) );
  AOI21_X1 U15805 ( .B1(n13740), .B2(n15161), .A(n13739), .ZN(n13841) );
  INV_X1 U15806 ( .A(n13841), .ZN(n13749) );
  OAI211_X1 U15807 ( .C1(n13756), .C2(n13899), .A(n13742), .B(n13741), .ZN(
        n13840) );
  AOI22_X1 U15808 ( .A1(n15149), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13743), 
        .B2(n15163), .ZN(n13746) );
  NAND2_X1 U15809 ( .A1(n13744), .A2(n15170), .ZN(n13745) );
  OAI211_X1 U15810 ( .C1(n13840), .C2(n13747), .A(n13746), .B(n13745), .ZN(
        n13748) );
  AOI21_X1 U15811 ( .B1(n13749), .B2(n11353), .A(n13748), .ZN(n13750) );
  OAI21_X1 U15812 ( .B1(n13842), .B2(n13793), .A(n13750), .ZN(P2_U3244) );
  XOR2_X1 U15813 ( .A(n13751), .B(n13754), .Z(n13753) );
  OAI21_X1 U15814 ( .B1(n13753), .B2(n13769), .A(n13752), .ZN(n13845) );
  INV_X1 U15815 ( .A(n13845), .ZN(n13764) );
  XNOR2_X1 U15816 ( .A(n13755), .B(n13754), .ZN(n13847) );
  INV_X1 U15817 ( .A(n13757), .ZN(n13904) );
  AOI211_X1 U15818 ( .C1(n13757), .C2(n13772), .A(n11852), .B(n13756), .ZN(
        n13846) );
  NAND2_X1 U15819 ( .A1(n13846), .A2(n15169), .ZN(n13761) );
  INV_X1 U15820 ( .A(n13758), .ZN(n13759) );
  AOI22_X1 U15821 ( .A1(n15149), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13759), 
        .B2(n15163), .ZN(n13760) );
  OAI211_X1 U15822 ( .C1(n13904), .C2(n15152), .A(n13761), .B(n13760), .ZN(
        n13762) );
  AOI21_X1 U15823 ( .B1(n15168), .B2(n13847), .A(n13762), .ZN(n13763) );
  OAI21_X1 U15824 ( .B1(n13764), .B2(n15174), .A(n13763), .ZN(P2_U3245) );
  XOR2_X1 U15825 ( .A(n13765), .B(n13766), .Z(n13855) );
  XOR2_X1 U15826 ( .A(n13767), .B(n13766), .Z(n13770) );
  OAI21_X1 U15827 ( .B1(n13770), .B2(n13769), .A(n13768), .ZN(n13851) );
  NAND2_X1 U15828 ( .A1(n13851), .A2(n11353), .ZN(n13780) );
  INV_X1 U15829 ( .A(n13771), .ZN(n13784) );
  INV_X1 U15830 ( .A(n13772), .ZN(n13773) );
  AOI211_X1 U15831 ( .C1(n13853), .C2(n13784), .A(n11852), .B(n13773), .ZN(
        n13852) );
  NOR2_X1 U15832 ( .A1(n9945), .A2(n15152), .ZN(n13778) );
  OAI22_X1 U15833 ( .A1(n11353), .A2(n13776), .B1(n13775), .B2(n13774), .ZN(
        n13777) );
  AOI211_X1 U15834 ( .C1(n13852), .C2(n15169), .A(n13778), .B(n13777), .ZN(
        n13779) );
  OAI211_X1 U15835 ( .C1(n13793), .C2(n13855), .A(n13780), .B(n13779), .ZN(
        P2_U3246) );
  XNOR2_X1 U15836 ( .A(n13781), .B(n13792), .ZN(n13783) );
  AOI21_X1 U15837 ( .B1(n13783), .B2(n15161), .A(n13782), .ZN(n13859) );
  AOI211_X1 U15838 ( .C1(n13857), .C2(n13785), .A(n11852), .B(n13771), .ZN(
        n13856) );
  INV_X1 U15839 ( .A(n13786), .ZN(n13787) );
  AOI22_X1 U15840 ( .A1(n15149), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13787), 
        .B2(n15163), .ZN(n13788) );
  OAI21_X1 U15841 ( .B1(n6988), .B2(n15152), .A(n13788), .ZN(n13795) );
  INV_X1 U15842 ( .A(n13789), .ZN(n13790) );
  AOI21_X1 U15843 ( .B1(n13792), .B2(n13791), .A(n13790), .ZN(n13860) );
  NOR2_X1 U15844 ( .A1(n13860), .A2(n13793), .ZN(n13794) );
  AOI211_X1 U15845 ( .C1(n13856), .C2(n15169), .A(n13795), .B(n13794), .ZN(
        n13796) );
  OAI21_X1 U15846 ( .B1(n15149), .B2(n13859), .A(n13796), .ZN(P2_U3247) );
  INV_X1 U15847 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13798) );
  OAI21_X1 U15848 ( .B1(n13612), .B2(n13850), .A(n13799), .ZN(P2_U3530) );
  INV_X1 U15849 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13802) );
  AND2_X1 U15850 ( .A1(n13801), .A2(n13800), .ZN(n13877) );
  MUX2_X1 U15851 ( .A(n13802), .B(n13877), .S(n15250), .Z(n13803) );
  OAI21_X1 U15852 ( .B1(n13880), .B2(n13850), .A(n13803), .ZN(P2_U3529) );
  NAND3_X1 U15853 ( .A1(n13808), .A2(n15212), .A3(n13807), .ZN(n13813) );
  NAND2_X1 U15854 ( .A1(n13809), .A2(n15200), .ZN(n13811) );
  NAND4_X1 U15855 ( .A1(n13813), .A2(n13812), .A3(n13811), .A4(n13810), .ZN(
        n13882) );
  MUX2_X1 U15856 ( .A(n13882), .B(P2_REG1_REG_27__SCAN_IN), .S(n9959), .Z(
        P2_U3526) );
  AOI21_X1 U15857 ( .B1(n15200), .B2(n13815), .A(n13814), .ZN(n13816) );
  OAI211_X1 U15858 ( .C1(n13818), .C2(n13861), .A(n13817), .B(n13816), .ZN(
        n13883) );
  MUX2_X1 U15859 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13883), .S(n15250), .Z(
        P2_U3525) );
  INV_X1 U15860 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13822) );
  AOI211_X1 U15861 ( .C1(n15212), .C2(n13821), .A(n13820), .B(n13819), .ZN(
        n13884) );
  MUX2_X1 U15862 ( .A(n13822), .B(n13884), .S(n15250), .Z(n13823) );
  OAI21_X1 U15863 ( .B1(n13887), .B2(n13850), .A(n13823), .ZN(P2_U3524) );
  INV_X1 U15864 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13828) );
  INV_X1 U15865 ( .A(n13824), .ZN(n13827) );
  AOI211_X1 U15866 ( .C1(n13827), .C2(n15239), .A(n13826), .B(n13825), .ZN(
        n13888) );
  MUX2_X1 U15867 ( .A(n13828), .B(n13888), .S(n15250), .Z(n13829) );
  OAI21_X1 U15868 ( .B1(n13891), .B2(n13850), .A(n13829), .ZN(P2_U3523) );
  AOI211_X1 U15869 ( .C1(n15212), .C2(n13832), .A(n13831), .B(n13830), .ZN(
        n13892) );
  MUX2_X1 U15870 ( .A(n13833), .B(n13892), .S(n15250), .Z(n13834) );
  OAI21_X1 U15871 ( .B1(n7264), .B2(n13850), .A(n13834), .ZN(P2_U3522) );
  AOI21_X1 U15872 ( .B1(n15200), .B2(n13836), .A(n13835), .ZN(n13837) );
  OAI211_X1 U15873 ( .C1(n13839), .C2(n13861), .A(n13838), .B(n13837), .ZN(
        n13895) );
  MUX2_X1 U15874 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13895), .S(n15250), .Z(
        P2_U3521) );
  OAI211_X1 U15875 ( .C1(n13861), .C2(n13842), .A(n13841), .B(n13840), .ZN(
        n13896) );
  MUX2_X1 U15876 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13896), .S(n15250), .Z(
        n13843) );
  INV_X1 U15877 ( .A(n13843), .ZN(n13844) );
  OAI21_X1 U15878 ( .B1(n13899), .B2(n13850), .A(n13844), .ZN(P2_U3520) );
  INV_X1 U15879 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n13848) );
  AOI211_X1 U15880 ( .C1(n13847), .C2(n15212), .A(n13846), .B(n13845), .ZN(
        n13900) );
  MUX2_X1 U15881 ( .A(n13848), .B(n13900), .S(n15250), .Z(n13849) );
  OAI21_X1 U15882 ( .B1(n13904), .B2(n13850), .A(n13849), .ZN(P2_U3519) );
  AOI211_X1 U15883 ( .C1(n15200), .C2(n13853), .A(n13852), .B(n13851), .ZN(
        n13854) );
  OAI21_X1 U15884 ( .B1(n13861), .B2(n13855), .A(n13854), .ZN(n13905) );
  MUX2_X1 U15885 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13905), .S(n15250), .Z(
        P2_U3518) );
  AOI21_X1 U15886 ( .B1(n15200), .B2(n13857), .A(n13856), .ZN(n13858) );
  OAI211_X1 U15887 ( .C1(n13860), .C2(n13861), .A(n13859), .B(n13858), .ZN(
        n13906) );
  MUX2_X1 U15888 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13906), .S(n15250), .Z(
        P2_U3517) );
  NOR2_X1 U15889 ( .A1(n13862), .A2(n13861), .ZN(n13866) );
  INV_X1 U15890 ( .A(n15200), .ZN(n15235) );
  OAI21_X1 U15891 ( .B1(n13864), .B2(n15235), .A(n13863), .ZN(n13865) );
  MUX2_X1 U15892 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13907), .S(n15250), .Z(
        P2_U3516) );
  AOI21_X1 U15893 ( .B1(n15200), .B2(n13869), .A(n13868), .ZN(n13873) );
  NAND3_X1 U15894 ( .A1(n13871), .A2(n15212), .A3(n13870), .ZN(n13872) );
  NAND3_X1 U15895 ( .A1(n13874), .A2(n13873), .A3(n13872), .ZN(n13908) );
  MUX2_X1 U15896 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13908), .S(n15250), .Z(
        P2_U3515) );
  INV_X1 U15897 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13876) );
  INV_X1 U15898 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13878) );
  MUX2_X1 U15899 ( .A(n13878), .B(n13877), .S(n15242), .Z(n13879) );
  OAI21_X1 U15900 ( .B1(n13880), .B2(n13903), .A(n13879), .ZN(P2_U3497) );
  MUX2_X1 U15901 ( .A(n13882), .B(P2_REG0_REG_27__SCAN_IN), .S(n15240), .Z(
        P2_U3494) );
  MUX2_X1 U15902 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13883), .S(n15242), .Z(
        P2_U3493) );
  INV_X1 U15903 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13885) );
  MUX2_X1 U15904 ( .A(n13885), .B(n13884), .S(n15242), .Z(n13886) );
  OAI21_X1 U15905 ( .B1(n13887), .B2(n13903), .A(n13886), .ZN(P2_U3492) );
  MUX2_X1 U15906 ( .A(n13889), .B(n13888), .S(n15242), .Z(n13890) );
  OAI21_X1 U15907 ( .B1(n13891), .B2(n13903), .A(n13890), .ZN(P2_U3491) );
  MUX2_X1 U15908 ( .A(n13893), .B(n13892), .S(n15242), .Z(n13894) );
  OAI21_X1 U15909 ( .B1(n7264), .B2(n13903), .A(n13894), .ZN(P2_U3490) );
  MUX2_X1 U15910 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13895), .S(n15242), .Z(
        P2_U3489) );
  MUX2_X1 U15911 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13896), .S(n15242), .Z(
        n13897) );
  INV_X1 U15912 ( .A(n13897), .ZN(n13898) );
  OAI21_X1 U15913 ( .B1(n13899), .B2(n13903), .A(n13898), .ZN(P2_U3488) );
  MUX2_X1 U15914 ( .A(n13901), .B(n13900), .S(n15242), .Z(n13902) );
  OAI21_X1 U15915 ( .B1(n13904), .B2(n13903), .A(n13902), .ZN(P2_U3487) );
  MUX2_X1 U15916 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13905), .S(n15242), .Z(
        P2_U3486) );
  MUX2_X1 U15917 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13906), .S(n15242), .Z(
        P2_U3484) );
  MUX2_X1 U15918 ( .A(n13907), .B(P2_REG0_REG_17__SCAN_IN), .S(n15240), .Z(
        P2_U3481) );
  MUX2_X1 U15919 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13908), .S(n15242), .Z(
        P2_U3478) );
  INV_X1 U15920 ( .A(n14537), .ZN(n13911) );
  NOR4_X1 U15921 ( .A1(n6777), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8519), .A4(
        P2_U3088), .ZN(n13909) );
  AOI21_X1 U15922 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13922), .A(n13909), 
        .ZN(n13910) );
  OAI21_X1 U15923 ( .B1(n13911), .B2(n13920), .A(n13910), .ZN(P2_U3296) );
  INV_X1 U15924 ( .A(n13912), .ZN(n14540) );
  INV_X1 U15925 ( .A(n13913), .ZN(n13915) );
  OAI222_X1 U15926 ( .A1(n13920), .A2(n14540), .B1(P2_U3088), .B2(n13915), 
        .C1(n13914), .C2(n13928), .ZN(P2_U3297) );
  OAI222_X1 U15927 ( .A1(n13920), .A2(n13919), .B1(P2_U3088), .B2(n13917), 
        .C1(n13916), .C2(n13928), .ZN(P2_U3298) );
  AOI21_X1 U15928 ( .B1(n13922), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13921), 
        .ZN(n13923) );
  OAI21_X1 U15929 ( .B1(n13924), .B2(n13920), .A(n13923), .ZN(P2_U3299) );
  INV_X1 U15930 ( .A(n13925), .ZN(n14543) );
  OAI222_X1 U15931 ( .A1(n13928), .A2(n13927), .B1(n13920), .B2(n14543), .C1(
        n13926), .C2(P2_U3088), .ZN(P2_U3300) );
  MUX2_X1 U15932 ( .A(n13929), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U15933 ( .B1(n13932), .B2(n13931), .A(n13930), .ZN(n13933) );
  INV_X1 U15934 ( .A(n13934), .ZN(n14257) );
  INV_X1 U15935 ( .A(n14101), .ZN(n14090) );
  AOI22_X1 U15936 ( .A1(n14052), .A2(n14112), .B1(n14110), .B2(n14071), .ZN(
        n14251) );
  OAI22_X1 U15937 ( .A1(n14073), .A2(n14251), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13935), .ZN(n13936) );
  AOI21_X1 U15938 ( .B1(n14257), .B2(n14090), .A(n13936), .ZN(n13937) );
  INV_X1 U15939 ( .A(n13938), .ZN(n13939) );
  AOI21_X1 U15940 ( .B1(n13941), .B2(n13940), .A(n13939), .ZN(n13948) );
  NAND2_X1 U15941 ( .A1(n13942), .A2(n14097), .ZN(n13943) );
  OAI211_X1 U15942 ( .C1(n14101), .C2(n13945), .A(n13944), .B(n13943), .ZN(
        n13946) );
  AOI21_X1 U15943 ( .B1(n14820), .B2(n14103), .A(n13946), .ZN(n13947) );
  OAI21_X1 U15944 ( .B1(n13948), .B2(n14106), .A(n13947), .ZN(P1_U3215) );
  OR2_X1 U15945 ( .A1(n13983), .A2(n14085), .ZN(n13951) );
  OR2_X1 U15946 ( .A1(n13949), .A2(n14268), .ZN(n13950) );
  NAND2_X1 U15947 ( .A1(n13951), .A2(n13950), .ZN(n14323) );
  AOI22_X1 U15948 ( .A1(n14097), .A2(n14323), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13952) );
  OAI21_X1 U15949 ( .B1(n14101), .B2(n14320), .A(n13952), .ZN(n13959) );
  INV_X1 U15950 ( .A(n13954), .ZN(n13955) );
  NAND3_X1 U15951 ( .A1(n14061), .A2(n13956), .A3(n13955), .ZN(n13957) );
  AOI21_X1 U15952 ( .B1(n14030), .B2(n13957), .A(n14106), .ZN(n13958) );
  AOI211_X1 U15953 ( .C1(n14103), .C2(n14472), .A(n13959), .B(n13958), .ZN(
        n13960) );
  INV_X1 U15954 ( .A(n13960), .ZN(P1_U3216) );
  OAI211_X1 U15955 ( .C1(n13963), .C2(n13962), .A(n13961), .B(n14082), .ZN(
        n13967) );
  AOI22_X1 U15956 ( .A1(n14103), .A2(n14980), .B1(n13964), .B2(n14097), .ZN(
        n13966) );
  MUX2_X1 U15957 ( .A(n14101), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n13965) );
  NAND3_X1 U15958 ( .A1(n13967), .A2(n13966), .A3(n13965), .ZN(P1_U3218) );
  INV_X1 U15959 ( .A(n14498), .ZN(n14399) );
  INV_X1 U15960 ( .A(n14065), .ZN(n13971) );
  OAI21_X1 U15961 ( .B1(n13971), .B2(n13970), .A(n13969), .ZN(n13973) );
  NAND3_X1 U15962 ( .A1(n13973), .A2(n14082), .A3(n13972), .ZN(n13979) );
  OR2_X1 U15963 ( .A1(n13984), .A2(n14268), .ZN(n13975) );
  NAND2_X1 U15964 ( .A1(n14120), .A2(n14052), .ZN(n13974) );
  NAND2_X1 U15965 ( .A1(n13975), .A2(n13974), .ZN(n14390) );
  NOR2_X1 U15966 ( .A1(n13976), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14220) );
  NOR2_X1 U15967 ( .A1(n14101), .A2(n14395), .ZN(n13977) );
  AOI211_X1 U15968 ( .C1(n14097), .C2(n14390), .A(n14220), .B(n13977), .ZN(
        n13978) );
  OAI211_X1 U15969 ( .C1(n14399), .C2(n14093), .A(n13979), .B(n13978), .ZN(
        P1_U3219) );
  INV_X1 U15970 ( .A(n14059), .ZN(n13980) );
  AOI21_X1 U15971 ( .B1(n13982), .B2(n13981), .A(n13980), .ZN(n13988) );
  OAI22_X1 U15972 ( .A1(n13984), .A2(n14085), .B1(n13983), .B2(n14268), .ZN(
        n14357) );
  AOI22_X1 U15973 ( .A1(n14357), .A2(n14097), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13985) );
  OAI21_X1 U15974 ( .B1(n14101), .B2(n14363), .A(n13985), .ZN(n13986) );
  AOI21_X1 U15975 ( .B1(n14486), .B2(n14103), .A(n13986), .ZN(n13987) );
  OAI21_X1 U15976 ( .B1(n13988), .B2(n14106), .A(n13987), .ZN(P1_U3223) );
  AND2_X1 U15977 ( .A1(n13990), .A2(n13989), .ZN(n13993) );
  OAI211_X1 U15978 ( .C1(n13993), .C2(n13992), .A(n14082), .B(n13991), .ZN(
        n13998) );
  NOR2_X1 U15979 ( .A1(n14101), .A2(n14687), .ZN(n13994) );
  AOI211_X1 U15980 ( .C1(n14097), .C2(n13996), .A(n13995), .B(n13994), .ZN(
        n13997) );
  OAI211_X1 U15981 ( .C1(n13999), .C2(n14093), .A(n13998), .B(n13997), .ZN(
        P1_U3224) );
  INV_X1 U15982 ( .A(n14019), .ZN(n14001) );
  AOI21_X1 U15983 ( .B1(n14003), .B2(n14002), .A(n14001), .ZN(n14009) );
  NAND2_X1 U15984 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14876)
         );
  NAND2_X1 U15985 ( .A1(n14097), .A2(n14004), .ZN(n14005) );
  OAI211_X1 U15986 ( .C1(n14101), .C2(n14006), .A(n14876), .B(n14005), .ZN(
        n14007) );
  AOI21_X1 U15987 ( .B1(n14804), .B2(n14103), .A(n14007), .ZN(n14008) );
  OAI21_X1 U15988 ( .B1(n14009), .B2(n14106), .A(n14008), .ZN(P1_U3226) );
  NAND2_X1 U15989 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14891)
         );
  OR2_X1 U15990 ( .A1(n14010), .A2(n14268), .ZN(n14013) );
  OR2_X1 U15991 ( .A1(n14011), .A2(n14085), .ZN(n14012) );
  NAND2_X1 U15992 ( .A1(n14013), .A2(n14012), .ZN(n14509) );
  NAND2_X1 U15993 ( .A1(n14097), .A2(n14509), .ZN(n14014) );
  OAI211_X1 U15994 ( .C1(n14101), .C2(n14425), .A(n14891), .B(n14014), .ZN(
        n14022) );
  INV_X1 U15995 ( .A(n14016), .ZN(n14017) );
  NAND3_X1 U15996 ( .A1(n14019), .A2(n14018), .A3(n14017), .ZN(n14020) );
  AOI21_X1 U15997 ( .B1(n14015), .B2(n14020), .A(n14106), .ZN(n14021) );
  AOI211_X1 U15998 ( .C1(n14103), .C2(n14510), .A(n14022), .B(n14021), .ZN(
        n14023) );
  INV_X1 U15999 ( .A(n14023), .ZN(P1_U3228) );
  NAND2_X1 U16000 ( .A1(n14115), .A2(n14052), .ZN(n14025) );
  NAND2_X1 U16001 ( .A1(n14113), .A2(n14071), .ZN(n14024) );
  NAND2_X1 U16002 ( .A1(n14025), .A2(n14024), .ZN(n14304) );
  AOI22_X1 U16003 ( .A1(n14097), .A2(n14304), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14026) );
  OAI21_X1 U16004 ( .B1(n14101), .B2(n14312), .A(n14026), .ZN(n14034) );
  INV_X1 U16005 ( .A(n14027), .ZN(n14028) );
  NAND3_X1 U16006 ( .A1(n14030), .A2(n14029), .A3(n14028), .ZN(n14031) );
  AOI21_X1 U16007 ( .B1(n14032), .B2(n14031), .A(n14106), .ZN(n14033) );
  XNOR2_X1 U16008 ( .A(n14035), .B(n14036), .ZN(n14043) );
  INV_X1 U16009 ( .A(n14378), .ZN(n14040) );
  OAI22_X1 U16010 ( .A1(n14038), .A2(n14085), .B1(n14037), .B2(n14268), .ZN(
        n14368) );
  AOI22_X1 U16011 ( .A1(n14368), .A2(n14097), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14039) );
  OAI21_X1 U16012 ( .B1(n14101), .B2(n14040), .A(n14039), .ZN(n14041) );
  AOI21_X1 U16013 ( .B1(n14492), .B2(n14103), .A(n14041), .ZN(n14042) );
  OAI21_X1 U16014 ( .B1(n14043), .B2(n14106), .A(n14042), .ZN(P1_U3233) );
  XNOR2_X1 U16015 ( .A(n14045), .B(n14044), .ZN(n14051) );
  NOR2_X1 U16016 ( .A1(n14101), .A2(n14046), .ZN(n14049) );
  OAI22_X1 U16017 ( .A1(n14073), .A2(n14047), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9184), .ZN(n14048) );
  AOI211_X1 U16018 ( .C1(n14827), .C2(n14103), .A(n14049), .B(n14048), .ZN(
        n14050) );
  OAI21_X1 U16019 ( .B1(n14051), .B2(n14106), .A(n14050), .ZN(P1_U3234) );
  NAND2_X1 U16020 ( .A1(n14117), .A2(n14052), .ZN(n14054) );
  NAND2_X1 U16021 ( .A1(n14115), .A2(n14071), .ZN(n14053) );
  NAND2_X1 U16022 ( .A1(n14054), .A2(n14053), .ZN(n14340) );
  AOI22_X1 U16023 ( .A1(n14097), .A2(n14340), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14055) );
  OAI21_X1 U16024 ( .B1(n14101), .B2(n14345), .A(n14055), .ZN(n14063) );
  INV_X1 U16025 ( .A(n14056), .ZN(n14057) );
  NAND3_X1 U16026 ( .A1(n14059), .A2(n14058), .A3(n14057), .ZN(n14060) );
  AOI21_X1 U16027 ( .B1(n14061), .B2(n14060), .A(n14106), .ZN(n14062) );
  AOI211_X1 U16028 ( .C1(n14103), .C2(n14482), .A(n14063), .B(n14062), .ZN(
        n14064) );
  INV_X1 U16029 ( .A(n14064), .ZN(P1_U3235) );
  OAI21_X1 U16030 ( .B1(n14067), .B2(n14066), .A(n14065), .ZN(n14068) );
  NAND2_X1 U16031 ( .A1(n14068), .A2(n14082), .ZN(n14076) );
  INV_X1 U16032 ( .A(n14069), .ZN(n14412) );
  NOR2_X1 U16033 ( .A1(n14070), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14909) );
  NAND2_X1 U16034 ( .A1(n14119), .A2(n14071), .ZN(n14411) );
  OR2_X1 U16035 ( .A1(n14072), .A2(n14085), .ZN(n14407) );
  AOI21_X1 U16036 ( .B1(n14411), .B2(n14407), .A(n14073), .ZN(n14074) );
  AOI211_X1 U16037 ( .C1(n14412), .C2(n14090), .A(n14909), .B(n14074), .ZN(
        n14075) );
  OAI211_X1 U16038 ( .C1(n14409), .C2(n14093), .A(n14076), .B(n14075), .ZN(
        P1_U3238) );
  AND2_X1 U16039 ( .A1(n14078), .A2(n14077), .ZN(n14080) );
  OAI21_X1 U16040 ( .B1(n14081), .B2(n14080), .A(n14079), .ZN(n14083) );
  NAND2_X1 U16041 ( .A1(n14083), .A2(n14082), .ZN(n14092) );
  INV_X1 U16042 ( .A(n14084), .ZN(n14277) );
  INV_X1 U16043 ( .A(n14111), .ZN(n14269) );
  NOR2_X1 U16044 ( .A1(n14086), .A2(n14085), .ZN(n14270) );
  AOI22_X1 U16045 ( .A1(n14097), .A2(n14270), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14087) );
  OAI21_X1 U16046 ( .B1(n14088), .B2(n14269), .A(n14087), .ZN(n14089) );
  AOI21_X1 U16047 ( .B1(n14277), .B2(n14090), .A(n14089), .ZN(n14091) );
  OAI211_X1 U16048 ( .C1(n14094), .C2(n14093), .A(n14092), .B(n14091), .ZN(
        P1_U3240) );
  XNOR2_X1 U16049 ( .A(n14096), .B(n14095), .ZN(n14107) );
  NAND2_X1 U16050 ( .A1(n14097), .A2(n14811), .ZN(n14098) );
  OAI211_X1 U16051 ( .C1(n14101), .C2(n14100), .A(n14099), .B(n14098), .ZN(
        n14102) );
  AOI21_X1 U16052 ( .B1(n14104), .B2(n14103), .A(n14102), .ZN(n14105) );
  OAI21_X1 U16053 ( .B1(n14107), .B2(n14106), .A(n14105), .ZN(P1_U3241) );
  MUX2_X1 U16054 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14224), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16055 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14108), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16056 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14109), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16057 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14110), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16058 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14111), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16059 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14112), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16060 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14113), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16061 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14114), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16062 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14115), .S(n14133), .Z(
        P1_U3583) );
  MUX2_X1 U16063 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14116), .S(n14133), .Z(
        P1_U3582) );
  MUX2_X1 U16064 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14117), .S(n14133), .Z(
        P1_U3581) );
  MUX2_X1 U16065 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14118), .S(n14133), .Z(
        P1_U3580) );
  MUX2_X1 U16066 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14119), .S(n14133), .Z(
        P1_U3579) );
  MUX2_X1 U16067 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14120), .S(n14133), .Z(
        P1_U3578) );
  MUX2_X1 U16068 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14121), .S(n14133), .Z(
        P1_U3577) );
  MUX2_X1 U16069 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14122), .S(n14133), .Z(
        P1_U3576) );
  MUX2_X1 U16070 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14123), .S(n14133), .Z(
        P1_U3574) );
  MUX2_X1 U16071 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14124), .S(n14133), .Z(
        P1_U3573) );
  MUX2_X1 U16072 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14125), .S(n14133), .Z(
        P1_U3572) );
  MUX2_X1 U16073 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14126), .S(n14133), .Z(
        P1_U3571) );
  MUX2_X1 U16074 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14127), .S(n14133), .Z(
        P1_U3570) );
  MUX2_X1 U16075 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14128), .S(n14133), .Z(
        P1_U3569) );
  MUX2_X1 U16076 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14129), .S(n14133), .Z(
        P1_U3568) );
  MUX2_X1 U16077 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14130), .S(n14133), .Z(
        P1_U3567) );
  MUX2_X1 U16078 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14131), .S(n14133), .Z(
        P1_U3566) );
  MUX2_X1 U16079 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14132), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16080 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14134), .S(n14133), .Z(
        P1_U3564) );
  MUX2_X1 U16081 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14135), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16082 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14136), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16083 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14137), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16084 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14138), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16085 ( .C1(n14141), .C2(n14140), .A(n14898), .B(n14139), .ZN(
        n14148) );
  OAI211_X1 U16086 ( .C1(n14143), .C2(n14149), .A(n14903), .B(n14142), .ZN(
        n14147) );
  AOI22_X1 U16087 ( .A1(n14860), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14146) );
  NAND2_X1 U16088 ( .A1(n14875), .A2(n14144), .ZN(n14145) );
  NAND4_X1 U16089 ( .A1(n14148), .A2(n14147), .A3(n14146), .A4(n14145), .ZN(
        P1_U3244) );
  AOI21_X1 U16090 ( .B1(n14857), .B2(n11377), .A(n9524), .ZN(n14856) );
  MUX2_X1 U16091 ( .A(n14150), .B(n14149), .S(n14857), .Z(n14152) );
  NAND2_X1 U16092 ( .A1(n14152), .A2(n14151), .ZN(n14154) );
  OAI211_X1 U16093 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14856), .A(n14154), .B(
        P1_U4016), .ZN(n14195) );
  NAND2_X1 U16094 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n14156) );
  NAND2_X1 U16095 ( .A1(n14860), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n14155) );
  OAI211_X1 U16096 ( .C1(n14907), .C2(n14157), .A(n14156), .B(n14155), .ZN(
        n14158) );
  INV_X1 U16097 ( .A(n14158), .ZN(n14167) );
  OAI211_X1 U16098 ( .C1(n14161), .C2(n14160), .A(n14903), .B(n14159), .ZN(
        n14166) );
  OAI211_X1 U16099 ( .C1(n14164), .C2(n14163), .A(n14898), .B(n14162), .ZN(
        n14165) );
  NAND4_X1 U16100 ( .A1(n14195), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        P1_U3245) );
  NAND2_X1 U16101 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n14168) );
  OAI21_X1 U16102 ( .B1(n14912), .B2(n14603), .A(n14168), .ZN(n14169) );
  AOI21_X1 U16103 ( .B1(n14170), .B2(n14875), .A(n14169), .ZN(n14179) );
  OAI211_X1 U16104 ( .C1(n14173), .C2(n14172), .A(n14903), .B(n14171), .ZN(
        n14178) );
  OAI211_X1 U16105 ( .C1(n14176), .C2(n14175), .A(n14898), .B(n14174), .ZN(
        n14177) );
  NAND3_X1 U16106 ( .A1(n14179), .A2(n14178), .A3(n14177), .ZN(P1_U3246) );
  AOI21_X1 U16107 ( .B1(n14860), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14180), .ZN(
        n14181) );
  OAI21_X1 U16108 ( .B1(n14907), .B2(n14182), .A(n14181), .ZN(n14183) );
  INV_X1 U16109 ( .A(n14183), .ZN(n14194) );
  INV_X1 U16110 ( .A(n14184), .ZN(n14185) );
  OAI211_X1 U16111 ( .C1(n14187), .C2(n14186), .A(n14898), .B(n14185), .ZN(
        n14193) );
  INV_X1 U16112 ( .A(n14188), .ZN(n14189) );
  OAI211_X1 U16113 ( .C1(n14191), .C2(n14190), .A(n14903), .B(n14189), .ZN(
        n14192) );
  NAND4_X1 U16114 ( .A1(n14195), .A2(n14194), .A3(n14193), .A4(n14192), .ZN(
        P1_U3247) );
  NOR2_X1 U16115 ( .A1(n14874), .A2(n14196), .ZN(n14197) );
  AOI21_X1 U16116 ( .B1(n14874), .B2(n14196), .A(n14197), .ZN(n14870) );
  INV_X1 U16117 ( .A(n14198), .ZN(n14200) );
  OAI21_X1 U16118 ( .B1(n14200), .B2(n14208), .A(n14199), .ZN(n14871) );
  NOR2_X1 U16119 ( .A1(n14870), .A2(n14871), .ZN(n14869) );
  AOI21_X1 U16120 ( .B1(n14874), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14869), 
        .ZN(n14884) );
  MUX2_X1 U16121 ( .A(n14426), .B(P1_REG2_REG_17__SCAN_IN), .S(n14211), .Z(
        n14885) );
  NOR2_X1 U16122 ( .A1(n14884), .A2(n14885), .ZN(n14883) );
  NOR2_X1 U16123 ( .A1(n14201), .A2(n14906), .ZN(n14202) );
  XNOR2_X1 U16124 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14203), .ZN(n14217) );
  INV_X1 U16125 ( .A(n14217), .ZN(n14215) );
  NOR2_X1 U16126 ( .A1(n14874), .A2(n14204), .ZN(n14205) );
  AOI21_X1 U16127 ( .B1(n14204), .B2(n14874), .A(n14205), .ZN(n14866) );
  INV_X1 U16128 ( .A(n14206), .ZN(n14209) );
  OAI21_X1 U16129 ( .B1(n14209), .B2(n14208), .A(n14207), .ZN(n14867) );
  NOR2_X1 U16130 ( .A1(n14866), .A2(n14867), .ZN(n14865) );
  MUX2_X1 U16131 ( .A(n14210), .B(P1_REG1_REG_17__SCAN_IN), .S(n14211), .Z(
        n14881) );
  NOR2_X1 U16132 ( .A1(n14880), .A2(n14881), .ZN(n14879) );
  NOR2_X1 U16133 ( .A1(n14212), .A2(n14906), .ZN(n14213) );
  XNOR2_X1 U16134 ( .A(n14906), .B(n14212), .ZN(n14896) );
  NOR2_X1 U16135 ( .A1(n14895), .A2(n14896), .ZN(n14894) );
  OAI21_X1 U16136 ( .B1(n14216), .B2(n14864), .A(n14907), .ZN(n14214) );
  AOI22_X1 U16137 ( .A1(n14217), .A2(n14903), .B1(n14216), .B2(n14898), .ZN(
        n14219) );
  AOI21_X1 U16138 ( .B1(n14860), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n14220), 
        .ZN(n14221) );
  NAND2_X1 U16139 ( .A1(n14222), .A2(n14221), .ZN(P1_U3262) );
  NAND2_X1 U16140 ( .A1(n14438), .A2(n14228), .ZN(n14227) );
  XNOR2_X1 U16141 ( .A(n14435), .B(n14227), .ZN(n14433) );
  NAND2_X1 U16142 ( .A1(n14433), .A2(n14263), .ZN(n14226) );
  NAND2_X1 U16143 ( .A1(n14224), .A2(n14223), .ZN(n14436) );
  NOR2_X1 U16144 ( .A1(n14942), .A2(n14436), .ZN(n14230) );
  AOI21_X1 U16145 ( .B1(n14942), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14230), 
        .ZN(n14225) );
  OAI211_X1 U16146 ( .C1(n14435), .C2(n14944), .A(n14226), .B(n14225), .ZN(
        P1_U3263) );
  OAI211_X1 U16147 ( .C1(n14438), .C2(n14228), .A(n14948), .B(n14227), .ZN(
        n14437) );
  AND2_X1 U16148 ( .A1(n14942), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14229) );
  NOR2_X1 U16149 ( .A1(n14230), .A2(n14229), .ZN(n14233) );
  NAND2_X1 U16150 ( .A1(n14231), .A2(n14417), .ZN(n14232) );
  OAI211_X1 U16151 ( .C1(n14437), .C2(n14334), .A(n14233), .B(n14232), .ZN(
        P1_U3264) );
  OAI21_X1 U16152 ( .B1(n14236), .B2(n14235), .A(n14234), .ZN(n14238) );
  AOI21_X1 U16153 ( .B1(n14238), .B2(n14937), .A(n14237), .ZN(n14448) );
  AOI211_X1 U16154 ( .C1(n14446), .C2(n14255), .A(n14829), .B(n14239), .ZN(
        n14445) );
  INV_X1 U16155 ( .A(n14240), .ZN(n14241) );
  INV_X1 U16156 ( .A(n14940), .ZN(n14413) );
  AOI22_X1 U16157 ( .A1(n14942), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14241), 
        .B2(n14413), .ZN(n14242) );
  OAI21_X1 U16158 ( .B1(n14243), .B2(n14944), .A(n14242), .ZN(n14247) );
  OAI21_X1 U16159 ( .B1(n14448), .B2(n14942), .A(n14248), .ZN(P1_U3265) );
  OAI21_X1 U16160 ( .B1(n14250), .B2(n14261), .A(n14249), .ZN(n14253) );
  INV_X1 U16161 ( .A(n14251), .ZN(n14252) );
  AOI21_X1 U16162 ( .B1(n14253), .B2(n14937), .A(n14252), .ZN(n14453) );
  INV_X1 U16163 ( .A(n14255), .ZN(n14256) );
  AOI21_X1 U16164 ( .B1(n14450), .B2(n7187), .A(n14256), .ZN(n14451) );
  AOI22_X1 U16165 ( .A1(n14942), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14257), 
        .B2(n14413), .ZN(n14258) );
  OAI21_X1 U16166 ( .B1(n14259), .B2(n14944), .A(n14258), .ZN(n14262) );
  AOI21_X1 U16167 ( .B1(n14261), .B2(n14260), .A(n6605), .ZN(n14454) );
  OAI21_X1 U16168 ( .B1(n14942), .B2(n14453), .A(n14264), .ZN(P1_U3266) );
  AOI21_X1 U16169 ( .B1(n14455), .B2(n14292), .A(n14254), .ZN(n14456) );
  INV_X1 U16170 ( .A(n14456), .ZN(n14273) );
  OAI21_X1 U16171 ( .B1(n14267), .B2(n14266), .A(n14265), .ZN(n14272) );
  NOR2_X1 U16172 ( .A1(n14269), .A2(n14268), .ZN(n14271) );
  AOI211_X1 U16173 ( .C1(n14272), .C2(n14937), .A(n14271), .B(n14270), .ZN(
        n14458) );
  OAI21_X1 U16174 ( .B1(n14682), .B2(n14273), .A(n14458), .ZN(n14281) );
  OAI21_X1 U16175 ( .B1(n14276), .B2(n14275), .A(n14274), .ZN(n14459) );
  AOI22_X1 U16176 ( .A1(n14942), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14277), 
        .B2(n14413), .ZN(n14279) );
  NAND2_X1 U16177 ( .A1(n14455), .A2(n14417), .ZN(n14278) );
  OAI211_X1 U16178 ( .C1(n14459), .C2(n14432), .A(n14279), .B(n14278), .ZN(
        n14280) );
  AOI21_X1 U16179 ( .B1(n14281), .B2(n14427), .A(n14280), .ZN(n14282) );
  INV_X1 U16180 ( .A(n14282), .ZN(P1_U3267) );
  OAI21_X1 U16181 ( .B1(n14283), .B2(n14285), .A(n14284), .ZN(n14287) );
  AOI21_X1 U16182 ( .B1(n14287), .B2(n14937), .A(n14286), .ZN(n14464) );
  OAI21_X1 U16183 ( .B1(n14288), .B2(n14940), .A(n14464), .ZN(n14297) );
  OAI21_X1 U16184 ( .B1(n14289), .B2(n14291), .A(n14290), .ZN(n14465) );
  NOR2_X1 U16185 ( .A1(n14465), .A2(n14432), .ZN(n14296) );
  OAI211_X1 U16186 ( .C1(n14293), .C2(n14311), .A(n14948), .B(n14292), .ZN(
        n14462) );
  AOI22_X1 U16187 ( .A1(n14460), .A2(n14417), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n14942), .ZN(n14294) );
  OAI21_X1 U16188 ( .B1(n14462), .B2(n14334), .A(n14294), .ZN(n14295) );
  AOI211_X1 U16189 ( .C1(n14297), .C2(n14427), .A(n14296), .B(n14295), .ZN(
        n14298) );
  INV_X1 U16190 ( .A(n14298), .ZN(P1_U3268) );
  NAND2_X1 U16191 ( .A1(n14300), .A2(n14299), .ZN(n14301) );
  NAND2_X1 U16192 ( .A1(n14301), .A2(n14937), .ZN(n14302) );
  OR2_X1 U16193 ( .A1(n14303), .A2(n14302), .ZN(n14306) );
  INV_X1 U16194 ( .A(n14304), .ZN(n14305) );
  NAND2_X1 U16195 ( .A1(n14306), .A2(n14305), .ZN(n14471) );
  INV_X1 U16196 ( .A(n14471), .ZN(n14319) );
  NAND2_X1 U16197 ( .A1(n14307), .A2(n7565), .ZN(n14308) );
  NAND2_X1 U16198 ( .A1(n6792), .A2(n14308), .ZN(n14466) );
  NAND2_X1 U16199 ( .A1(n14314), .A2(n14331), .ZN(n14309) );
  NAND2_X1 U16200 ( .A1(n14309), .A2(n14948), .ZN(n14310) );
  OR2_X1 U16201 ( .A1(n14311), .A2(n14310), .ZN(n14467) );
  INV_X1 U16202 ( .A(n14312), .ZN(n14313) );
  AOI22_X1 U16203 ( .A1(n14942), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14313), 
        .B2(n14413), .ZN(n14316) );
  NAND2_X1 U16204 ( .A1(n14314), .A2(n14417), .ZN(n14315) );
  OAI211_X1 U16205 ( .C1(n14467), .C2(n14334), .A(n14316), .B(n14315), .ZN(
        n14317) );
  AOI21_X1 U16206 ( .B1(n14466), .B2(n14954), .A(n14317), .ZN(n14318) );
  OAI21_X1 U16207 ( .B1(n14319), .B2(n14942), .A(n14318), .ZN(P1_U3269) );
  INV_X1 U16208 ( .A(n14320), .ZN(n14326) );
  OAI21_X1 U16209 ( .B1(n14322), .B2(n14327), .A(n14321), .ZN(n14324) );
  AOI21_X1 U16210 ( .B1(n14324), .B2(n14937), .A(n14323), .ZN(n14478) );
  INV_X1 U16211 ( .A(n14478), .ZN(n14325) );
  AOI21_X1 U16212 ( .B1(n14326), .B2(n14413), .A(n14325), .ZN(n14337) );
  NAND2_X1 U16213 ( .A1(n14328), .A2(n14327), .ZN(n14329) );
  AND2_X1 U16214 ( .A1(n14330), .A2(n14329), .ZN(n14476) );
  AOI21_X1 U16215 ( .B1(n14472), .B2(n14342), .A(n14829), .ZN(n14332) );
  NAND2_X1 U16216 ( .A1(n14332), .A2(n14331), .ZN(n14474) );
  AOI22_X1 U16217 ( .A1(n14472), .A2(n14417), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n14942), .ZN(n14333) );
  OAI21_X1 U16218 ( .B1(n14474), .B2(n14334), .A(n14333), .ZN(n14335) );
  AOI21_X1 U16219 ( .B1(n14476), .B2(n14954), .A(n14335), .ZN(n14336) );
  OAI21_X1 U16220 ( .B1(n14337), .B2(n14942), .A(n14336), .ZN(P1_U3270) );
  CLKBUF_X1 U16221 ( .A(n14338), .Z(n14339) );
  XNOR2_X1 U16222 ( .A(n14339), .B(n14350), .ZN(n14341) );
  AOI21_X1 U16223 ( .B1(n14341), .B2(n14937), .A(n14340), .ZN(n14484) );
  INV_X1 U16224 ( .A(n14360), .ZN(n14344) );
  INV_X1 U16225 ( .A(n14342), .ZN(n14343) );
  AOI211_X1 U16226 ( .C1(n14482), .C2(n14344), .A(n14829), .B(n14343), .ZN(
        n14481) );
  INV_X1 U16227 ( .A(n14345), .ZN(n14346) );
  AOI22_X1 U16228 ( .A1(n14942), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14346), 
        .B2(n14413), .ZN(n14347) );
  OAI21_X1 U16229 ( .B1(n14348), .B2(n14944), .A(n14347), .ZN(n14352) );
  XNOR2_X1 U16230 ( .A(n14349), .B(n14350), .ZN(n14485) );
  NOR2_X1 U16231 ( .A1(n14485), .A2(n14432), .ZN(n14351) );
  AOI211_X1 U16232 ( .C1(n14481), .C2(n14953), .A(n14352), .B(n14351), .ZN(
        n14353) );
  OAI21_X1 U16233 ( .B1(n14942), .B2(n14484), .A(n14353), .ZN(P1_U3271) );
  AOI21_X1 U16234 ( .B1(n14355), .B2(n14354), .A(n6617), .ZN(n14490) );
  XOR2_X1 U16235 ( .A(n14356), .B(n14355), .Z(n14358) );
  AOI21_X1 U16236 ( .B1(n14358), .B2(n14937), .A(n14357), .ZN(n14489) );
  AND2_X1 U16237 ( .A1(n14376), .A2(n14486), .ZN(n14359) );
  NOR2_X1 U16238 ( .A1(n14360), .A2(n14359), .ZN(n14487) );
  NAND2_X1 U16239 ( .A1(n14487), .A2(n14361), .ZN(n14362) );
  OAI211_X1 U16240 ( .C1(n14940), .C2(n14363), .A(n14489), .B(n14362), .ZN(
        n14364) );
  NAND2_X1 U16241 ( .A1(n14364), .A2(n14427), .ZN(n14366) );
  AOI22_X1 U16242 ( .A1(n14486), .A2(n14417), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n14942), .ZN(n14365) );
  OAI211_X1 U16243 ( .C1(n14490), .C2(n14432), .A(n14366), .B(n14365), .ZN(
        P1_U3272) );
  AOI21_X1 U16244 ( .B1(n14367), .B2(n14373), .A(n14917), .ZN(n14370) );
  AOI21_X1 U16245 ( .B1(n14370), .B2(n14369), .A(n14368), .ZN(n14494) );
  INV_X1 U16246 ( .A(n14371), .ZN(n14374) );
  OAI21_X1 U16247 ( .B1(n14374), .B2(n14373), .A(n14372), .ZN(n14495) );
  INV_X1 U16248 ( .A(n14495), .ZN(n14383) );
  INV_X1 U16249 ( .A(n14375), .ZN(n14393) );
  INV_X1 U16250 ( .A(n14376), .ZN(n14377) );
  AOI211_X1 U16251 ( .C1(n14492), .C2(n14393), .A(n14829), .B(n14377), .ZN(
        n14491) );
  NAND2_X1 U16252 ( .A1(n14491), .A2(n14953), .ZN(n14380) );
  AOI22_X1 U16253 ( .A1(n14942), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14378), 
        .B2(n14413), .ZN(n14379) );
  OAI211_X1 U16254 ( .C1(n14381), .C2(n14944), .A(n14380), .B(n14379), .ZN(
        n14382) );
  AOI21_X1 U16255 ( .B1(n14383), .B2(n14954), .A(n14382), .ZN(n14384) );
  OAI21_X1 U16256 ( .B1(n14494), .B2(n14942), .A(n14384), .ZN(P1_U3273) );
  XOR2_X1 U16257 ( .A(n14385), .B(n14389), .Z(n14500) );
  INV_X1 U16258 ( .A(n14386), .ZN(n14387) );
  AOI21_X1 U16259 ( .B1(n14389), .B2(n14388), .A(n14387), .ZN(n14392) );
  INV_X1 U16260 ( .A(n14390), .ZN(n14391) );
  OAI21_X1 U16261 ( .B1(n14392), .B2(n14917), .A(n14391), .ZN(n14496) );
  AOI21_X1 U16262 ( .B1(n6679), .B2(n14498), .A(n14829), .ZN(n14394) );
  AND2_X1 U16263 ( .A1(n14394), .A2(n14393), .ZN(n14497) );
  NAND2_X1 U16264 ( .A1(n14497), .A2(n14953), .ZN(n14398) );
  INV_X1 U16265 ( .A(n14395), .ZN(n14396) );
  AOI22_X1 U16266 ( .A1(n14942), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14396), 
        .B2(n14413), .ZN(n14397) );
  OAI211_X1 U16267 ( .C1(n14399), .C2(n14944), .A(n14398), .B(n14397), .ZN(
        n14400) );
  AOI21_X1 U16268 ( .B1(n14496), .B2(n14427), .A(n14400), .ZN(n14401) );
  OAI21_X1 U16269 ( .B1(n14500), .B2(n14432), .A(n14401), .ZN(P1_U3274) );
  INV_X1 U16270 ( .A(n14402), .ZN(n14405) );
  XNOR2_X1 U16271 ( .A(n14403), .B(n14405), .ZN(n14505) );
  XNOR2_X1 U16272 ( .A(n14404), .B(n14405), .ZN(n14406) );
  NAND2_X1 U16273 ( .A1(n14406), .A2(n14937), .ZN(n14408) );
  OAI211_X1 U16274 ( .C1(n14966), .C2(n14505), .A(n14408), .B(n14407), .ZN(
        n14507) );
  OR2_X1 U16275 ( .A1(n14409), .A2(n14423), .ZN(n14410) );
  NAND3_X1 U16276 ( .A1(n6679), .A2(n14410), .A3(n14948), .ZN(n14503) );
  INV_X1 U16277 ( .A(n14411), .ZN(n14501) );
  AOI21_X1 U16278 ( .B1(n14413), .B2(n14412), .A(n14501), .ZN(n14414) );
  OAI21_X1 U16279 ( .B1(n14503), .B2(n14415), .A(n14414), .ZN(n14416) );
  OAI21_X1 U16280 ( .B1(n14507), .B2(n14416), .A(n14427), .ZN(n14419) );
  AOI22_X1 U16281 ( .A1(n14502), .A2(n14417), .B1(n14942), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n14418) );
  OAI211_X1 U16282 ( .C1(n14505), .C2(n14926), .A(n14419), .B(n14418), .ZN(
        P1_U3275) );
  XNOR2_X1 U16283 ( .A(n14420), .B(n6553), .ZN(n14513) );
  OAI211_X1 U16284 ( .C1(n6681), .C2(n6553), .A(n14937), .B(n14421), .ZN(
        n14511) );
  INV_X1 U16285 ( .A(n14511), .ZN(n14422) );
  OAI21_X1 U16286 ( .B1(n14422), .B2(n14509), .A(n14427), .ZN(n14431) );
  AOI211_X1 U16287 ( .C1(n14510), .C2(n6676), .A(n14829), .B(n14423), .ZN(
        n14508) );
  INV_X1 U16288 ( .A(n14510), .ZN(n14424) );
  NOR2_X1 U16289 ( .A1(n14424), .A2(n14944), .ZN(n14429) );
  OAI22_X1 U16290 ( .A1(n14427), .A2(n14426), .B1(n14425), .B2(n14940), .ZN(
        n14428) );
  AOI211_X1 U16291 ( .C1(n14508), .C2(n14953), .A(n14429), .B(n14428), .ZN(
        n14430) );
  OAI211_X1 U16292 ( .C1(n14513), .C2(n14432), .A(n14431), .B(n14430), .ZN(
        P1_U3276) );
  NAND2_X1 U16293 ( .A1(n14433), .A2(n14948), .ZN(n14434) );
  OAI211_X1 U16294 ( .C1(n14435), .C2(n15025), .A(n14434), .B(n14436), .ZN(
        n14514) );
  MUX2_X1 U16295 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14514), .S(n15045), .Z(
        P1_U3559) );
  OAI211_X1 U16296 ( .C1(n14438), .C2(n15025), .A(n14437), .B(n14436), .ZN(
        n14515) );
  MUX2_X1 U16297 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14515), .S(n15045), .Z(
        P1_U3558) );
  INV_X1 U16298 ( .A(n14825), .ZN(n14442) );
  MUX2_X1 U16299 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14516), .S(n15045), .Z(
        P1_U3557) );
  AOI21_X1 U16300 ( .B1(n14446), .B2(n14979), .A(n14445), .ZN(n14447) );
  MUX2_X1 U16301 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14517), .S(n15045), .Z(
        P1_U3556) );
  AOI22_X1 U16302 ( .A1(n14451), .A2(n14948), .B1(n14450), .B2(n14979), .ZN(
        n14452) );
  OAI211_X1 U16303 ( .C1(n14825), .C2(n14454), .A(n14453), .B(n14452), .ZN(
        n14518) );
  MUX2_X1 U16304 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14518), .S(n15045), .Z(
        P1_U3555) );
  AOI22_X1 U16305 ( .A1(n14456), .A2(n14948), .B1(n14455), .B2(n14979), .ZN(
        n14457) );
  OAI211_X1 U16306 ( .C1(n14825), .C2(n14459), .A(n14458), .B(n14457), .ZN(
        n14519) );
  MUX2_X1 U16307 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14519), .S(n15045), .Z(
        P1_U3554) );
  NAND2_X1 U16308 ( .A1(n14460), .A2(n14979), .ZN(n14461) );
  AND2_X1 U16309 ( .A1(n14462), .A2(n14461), .ZN(n14463) );
  OAI211_X1 U16310 ( .C1(n14825), .C2(n14465), .A(n14464), .B(n14463), .ZN(
        n14520) );
  MUX2_X1 U16311 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14520), .S(n15045), .Z(
        P1_U3553) );
  NAND2_X1 U16312 ( .A1(n14466), .A2(n14442), .ZN(n14468) );
  OAI211_X1 U16313 ( .C1(n14469), .C2(n15025), .A(n14468), .B(n14467), .ZN(
        n14470) );
  MUX2_X1 U16314 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14521), .S(n15045), .Z(
        P1_U3552) );
  INV_X1 U16315 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n14479) );
  NAND2_X1 U16316 ( .A1(n14472), .A2(n14979), .ZN(n14473) );
  NAND2_X1 U16317 ( .A1(n14474), .A2(n14473), .ZN(n14475) );
  AOI21_X1 U16318 ( .B1(n14476), .B2(n14442), .A(n14475), .ZN(n14477) );
  AND2_X1 U16319 ( .A1(n14478), .A2(n14477), .ZN(n14522) );
  MUX2_X1 U16320 ( .A(n14479), .B(n14522), .S(n15045), .Z(n14480) );
  INV_X1 U16321 ( .A(n14480), .ZN(P1_U3551) );
  AOI21_X1 U16322 ( .B1(n14482), .B2(n14979), .A(n14481), .ZN(n14483) );
  OAI211_X1 U16323 ( .C1(n14825), .C2(n14485), .A(n14484), .B(n14483), .ZN(
        n14525) );
  MUX2_X1 U16324 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14525), .S(n15045), .Z(
        P1_U3550) );
  AOI22_X1 U16325 ( .A1(n14487), .A2(n14948), .B1(n14486), .B2(n14979), .ZN(
        n14488) );
  OAI211_X1 U16326 ( .C1(n14825), .C2(n14490), .A(n14489), .B(n14488), .ZN(
        n14526) );
  MUX2_X1 U16327 ( .A(n14526), .B(P1_REG1_REG_21__SCAN_IN), .S(n15043), .Z(
        P1_U3549) );
  AOI21_X1 U16328 ( .B1(n14492), .B2(n14979), .A(n14491), .ZN(n14493) );
  OAI211_X1 U16329 ( .C1(n14825), .C2(n14495), .A(n14494), .B(n14493), .ZN(
        n14527) );
  MUX2_X1 U16330 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14527), .S(n15045), .Z(
        P1_U3548) );
  AOI211_X1 U16331 ( .C1(n14498), .C2(n14979), .A(n14497), .B(n14496), .ZN(
        n14499) );
  OAI21_X1 U16332 ( .B1(n14825), .B2(n14500), .A(n14499), .ZN(n14528) );
  MUX2_X1 U16333 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14528), .S(n15045), .Z(
        P1_U3547) );
  AOI21_X1 U16334 ( .B1(n14502), .B2(n14979), .A(n14501), .ZN(n14504) );
  OAI211_X1 U16335 ( .C1(n14505), .C2(n15013), .A(n14504), .B(n14503), .ZN(
        n14506) );
  OR2_X1 U16336 ( .A1(n14507), .A2(n14506), .ZN(n14529) );
  MUX2_X1 U16337 ( .A(n14529), .B(P1_REG1_REG_18__SCAN_IN), .S(n15043), .Z(
        P1_U3546) );
  AOI211_X1 U16338 ( .C1(n14510), .C2(n14979), .A(n14509), .B(n14508), .ZN(
        n14512) );
  OAI211_X1 U16339 ( .C1(n14825), .C2(n14513), .A(n14512), .B(n14511), .ZN(
        n14530) );
  MUX2_X1 U16340 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14530), .S(n15045), .Z(
        P1_U3545) );
  MUX2_X1 U16341 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14514), .S(n15030), .Z(
        P1_U3527) );
  MUX2_X1 U16342 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14515), .S(n15030), .Z(
        P1_U3526) );
  MUX2_X1 U16343 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14516), .S(n15030), .Z(
        P1_U3525) );
  MUX2_X1 U16344 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14517), .S(n15030), .Z(
        P1_U3524) );
  MUX2_X1 U16345 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14518), .S(n15030), .Z(
        P1_U3523) );
  MUX2_X1 U16346 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14519), .S(n15030), .Z(
        P1_U3522) );
  MUX2_X1 U16347 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14520), .S(n15030), .Z(
        P1_U3521) );
  MUX2_X1 U16348 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14521), .S(n15030), .Z(
        P1_U3520) );
  MUX2_X1 U16349 ( .A(n14523), .B(n14522), .S(n15030), .Z(n14524) );
  INV_X1 U16350 ( .A(n14524), .ZN(P1_U3519) );
  MUX2_X1 U16351 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14525), .S(n15030), .Z(
        P1_U3518) );
  MUX2_X1 U16352 ( .A(n14526), .B(P1_REG0_REG_21__SCAN_IN), .S(n15029), .Z(
        P1_U3517) );
  MUX2_X1 U16353 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14527), .S(n15030), .Z(
        P1_U3516) );
  MUX2_X1 U16354 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14528), .S(n15030), .Z(
        P1_U3515) );
  MUX2_X1 U16355 ( .A(n14529), .B(P1_REG0_REG_18__SCAN_IN), .S(n15029), .Z(
        P1_U3513) );
  MUX2_X1 U16356 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14530), .S(n15030), .Z(
        P1_U3510) );
  NAND3_X1 U16357 ( .A1(n14531), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14533) );
  OAI22_X1 U16358 ( .A1(n14534), .A2(n14533), .B1(n14532), .B2(n14542), .ZN(
        n14535) );
  AOI21_X1 U16359 ( .B1(n14537), .B2(n14536), .A(n14535), .ZN(n14538) );
  INV_X1 U16360 ( .A(n14538), .ZN(P1_U3324) );
  OAI222_X1 U16361 ( .A1(P1_U3086), .A2(n14541), .B1(n14544), .B2(n14540), 
        .C1(n14539), .C2(n14542), .ZN(P1_U3325) );
  OAI222_X1 U16362 ( .A1(P1_U3086), .A2(n14545), .B1(n14544), .B2(n14543), 
        .C1(n7419), .C2(n14542), .ZN(P1_U3328) );
  MUX2_X1 U16363 ( .A(n14547), .B(n14546), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16364 ( .A(n14548), .ZN(n14549) );
  MUX2_X1 U16365 ( .A(n14549), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16366 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14700) );
  XNOR2_X1 U16367 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14644) );
  INV_X1 U16368 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14585) );
  XOR2_X1 U16369 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(n14550), .Z(n14635) );
  NAND2_X1 U16370 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n14551), .ZN(n14583) );
  AOI22_X1 U16371 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n14552), .B1(
        P3_ADDR_REG_12__SCAN_IN), .B2(n14551), .ZN(n14590) );
  NAND2_X1 U16372 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n14553), .ZN(n14581) );
  INV_X1 U16373 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15288) );
  AOI22_X1 U16374 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n15288), .B1(
        P3_ADDR_REG_11__SCAN_IN), .B2(n14553), .ZN(n14632) );
  INV_X1 U16375 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14579) );
  NAND2_X1 U16376 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n14577), .ZN(n14554) );
  OAI21_X1 U16377 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14577), .A(n14554), .ZN(
        n14626) );
  XOR2_X1 U16378 ( .A(n14570), .B(n14555), .Z(n14613) );
  XNOR2_X2 U16379 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14594) );
  NAND2_X1 U16380 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n14556), .ZN(n14557) );
  NAND2_X1 U16381 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14561), .ZN(n14563) );
  INV_X1 U16382 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14593) );
  NAND2_X1 U16383 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14564), .ZN(n14565) );
  NAND2_X1 U16384 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14566), .ZN(n14569) );
  NAND2_X1 U16385 ( .A1(n14571), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n14573) );
  NAND2_X1 U16386 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n14574), .ZN(n14575) );
  XNOR2_X1 U16387 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n14629) );
  NAND2_X1 U16388 ( .A1(n14630), .A2(n14629), .ZN(n14578) );
  NAND2_X1 U16389 ( .A1(n14632), .A2(n14633), .ZN(n14580) );
  NAND2_X1 U16390 ( .A1(n14581), .A2(n14580), .ZN(n14591) );
  NAND2_X1 U16391 ( .A1(n14590), .A2(n14591), .ZN(n14582) );
  NAND2_X1 U16392 ( .A1(n14583), .A2(n14582), .ZN(n14636) );
  NAND2_X1 U16393 ( .A1(n14635), .A2(n14636), .ZN(n14584) );
  OAI21_X1 U16394 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14640), .A(n14642), 
        .ZN(n14586) );
  NAND2_X1 U16395 ( .A1(n14639), .A2(n14586), .ZN(n14643) );
  NAND2_X1 U16396 ( .A1(n14644), .A2(n14643), .ZN(n14587) );
  NAND2_X1 U16397 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14878), .ZN(n14588) );
  OAI21_X1 U16398 ( .B1(P3_ADDR_REG_16__SCAN_IN), .B2(n14878), .A(n14588), 
        .ZN(n14589) );
  XOR2_X1 U16399 ( .A(n14650), .B(n14589), .Z(n14854) );
  XNOR2_X1 U16400 ( .A(n14591), .B(n14590), .ZN(n14634) );
  INV_X1 U16401 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15079) );
  NOR2_X1 U16402 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14606), .ZN(n14608) );
  INV_X1 U16403 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14662) );
  XNOR2_X1 U16404 ( .A(n14595), .B(n14594), .ZN(n14660) );
  XNOR2_X1 U16405 ( .A(n14596), .B(n14597), .ZN(n14598) );
  NAND2_X1 U16406 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14598), .ZN(n14600) );
  AOI21_X1 U16407 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15258), .A(n14597), .ZN(
        n15445) );
  INV_X1 U16408 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15444) );
  NOR2_X1 U16409 ( .A1(n15445), .A2(n15444), .ZN(n15453) );
  NAND2_X1 U16410 ( .A1(n14600), .A2(n14599), .ZN(n14661) );
  NAND2_X1 U16411 ( .A1(n14660), .A2(n14661), .ZN(n14601) );
  NOR2_X1 U16412 ( .A1(n14660), .A2(n14661), .ZN(n14659) );
  XNOR2_X1 U16413 ( .A(n14603), .B(n14602), .ZN(n15450) );
  NOR2_X1 U16414 ( .A1(n15449), .A2(n15450), .ZN(n14605) );
  INV_X1 U16415 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14604) );
  NAND2_X1 U16416 ( .A1(n15449), .A2(n15450), .ZN(n15448) );
  OAI21_X1 U16417 ( .B1(n14605), .B2(n14604), .A(n15448), .ZN(n15442) );
  NOR2_X1 U16418 ( .A1(n15442), .A2(n15441), .ZN(n14607) );
  XOR2_X1 U16419 ( .A(n14613), .B(n14612), .Z(n14664) );
  NAND2_X1 U16420 ( .A1(n14614), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14615) );
  NAND2_X1 U16421 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14617), .ZN(n14621) );
  INV_X1 U16422 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14616) );
  XNOR2_X1 U16423 ( .A(n14619), .B(n14618), .ZN(n15446) );
  NAND2_X1 U16424 ( .A1(n15447), .A2(n15446), .ZN(n14620) );
  XNOR2_X1 U16425 ( .A(n14623), .B(n14622), .ZN(n14624) );
  XNOR2_X1 U16426 ( .A(n14630), .B(n14629), .ZN(n14671) );
  NAND2_X1 U16427 ( .A1(n14672), .A2(n14671), .ZN(n14631) );
  XNOR2_X1 U16428 ( .A(n14633), .B(n14632), .ZN(n14846) );
  XNOR2_X1 U16429 ( .A(n14636), .B(n14635), .ZN(n14637) );
  OAI21_X1 U16430 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14640), .A(n14639), 
        .ZN(n14641) );
  XNOR2_X1 U16431 ( .A(n14644), .B(n14643), .ZN(n14645) );
  INV_X1 U16432 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14653) );
  INV_X1 U16433 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14648) );
  NAND2_X1 U16434 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14648), .ZN(n14649) );
  AOI22_X1 U16435 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14878), .B1(n14650), 
        .B2(n14649), .ZN(n14651) );
  XNOR2_X1 U16436 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14651), .ZN(n14652) );
  NOR2_X1 U16437 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14651), .ZN(n14655) );
  NOR2_X1 U16438 ( .A1(n14653), .A2(n14652), .ZN(n14654) );
  NOR2_X1 U16439 ( .A1(n14655), .A2(n14654), .ZN(n14691) );
  AOI22_X1 U16440 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(P3_ADDR_REG_18__SCAN_IN), 
        .B1(n14656), .B2(n14913), .ZN(n14690) );
  XNOR2_X1 U16441 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14689), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16442 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14657) );
  OAI21_X1 U16443 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14657), 
        .ZN(U28) );
  AOI21_X1 U16444 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14658) );
  OAI21_X1 U16445 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14658), 
        .ZN(U29) );
  AOI21_X1 U16446 ( .B1(n14661), .B2(n14660), .A(n14659), .ZN(n14663) );
  XNOR2_X1 U16447 ( .A(n14663), .B(n14662), .ZN(SUB_1596_U61) );
  XOR2_X1 U16448 ( .A(n14665), .B(n14664), .Z(SUB_1596_U57) );
  XNOR2_X1 U16449 ( .A(n14666), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  NOR2_X1 U16450 ( .A1(n14668), .A2(n14667), .ZN(n14669) );
  XOR2_X1 U16451 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14669), .Z(SUB_1596_U54) );
  AOI21_X1 U16452 ( .B1(n14672), .B2(n14671), .A(n14670), .ZN(n14673) );
  XNOR2_X1 U16453 ( .A(n14673), .B(n15079), .ZN(SUB_1596_U70) );
  INV_X1 U16454 ( .A(n14674), .ZN(n14676) );
  INV_X1 U16455 ( .A(n14966), .ZN(n15020) );
  OAI21_X1 U16456 ( .B1(n14676), .B2(n15020), .A(n14675), .ZN(n14681) );
  INV_X1 U16457 ( .A(n14677), .ZN(n14678) );
  AOI21_X1 U16458 ( .B1(n14679), .B2(n14678), .A(n14942), .ZN(n14680) );
  OAI211_X1 U16459 ( .C1(n14683), .C2(n14682), .A(n14681), .B(n14680), .ZN(
        n14684) );
  OAI22_X1 U16460 ( .A1(n14685), .A2(n14684), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14427), .ZN(n14686) );
  OAI21_X1 U16461 ( .B1(n14687), .B2(n14940), .A(n14686), .ZN(P1_U3281) );
  XNOR2_X1 U16462 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14688), .ZN(SUB_1596_U63)
         );
  NOR2_X1 U16463 ( .A1(n14691), .A2(n14690), .ZN(n14692) );
  AOI21_X1 U16464 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14913), .A(n14692), 
        .ZN(n14696) );
  XNOR2_X1 U16465 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14693) );
  XNOR2_X1 U16466 ( .A(n14694), .B(n14693), .ZN(n14695) );
  AOI21_X1 U16467 ( .B1(n14699), .B2(n14698), .A(n14697), .ZN(n14715) );
  OAI22_X1 U16468 ( .A1(n15290), .A2(n14701), .B1(n14700), .B2(n15287), .ZN(
        n14712) );
  AOI21_X1 U16469 ( .B1(n14704), .B2(n14703), .A(n14702), .ZN(n14710) );
  NOR2_X1 U16470 ( .A1(n14706), .A2(n14705), .ZN(n14707) );
  OAI21_X1 U16471 ( .B1(n14708), .B2(n14707), .A(n15279), .ZN(n14709) );
  OAI21_X1 U16472 ( .B1(n14710), .B2(n15298), .A(n14709), .ZN(n14711) );
  NOR3_X1 U16473 ( .A1(n14713), .A2(n14712), .A3(n14711), .ZN(n14714) );
  OAI21_X1 U16474 ( .B1(n14715), .B2(n15304), .A(n14714), .ZN(P3_U3197) );
  INV_X1 U16475 ( .A(n14716), .ZN(n14717) );
  AOI22_X1 U16476 ( .A1(n14719), .A2(n15395), .B1(n14749), .B2(n15396), .ZN(
        n14723) );
  INV_X1 U16477 ( .A(n14745), .ZN(n14720) );
  AOI22_X1 U16478 ( .A1(n14720), .A2(n15374), .B1(n15398), .B2(
        P3_REG2_REG_31__SCAN_IN), .ZN(n14721) );
  NAND2_X1 U16479 ( .A1(n14723), .A2(n14721), .ZN(P3_U3202) );
  AOI22_X1 U16480 ( .A1(n15374), .A2(n12380), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15398), .ZN(n14722) );
  NAND2_X1 U16481 ( .A1(n14723), .A2(n14722), .ZN(P3_U3203) );
  XNOR2_X1 U16482 ( .A(n14724), .B(n14725), .ZN(n14759) );
  XNOR2_X1 U16483 ( .A(n14726), .B(n14725), .ZN(n14727) );
  OAI222_X1 U16484 ( .A1(n15382), .A2(n14729), .B1(n15381), .B2(n14728), .C1(
        n14727), .C2(n15388), .ZN(n14757) );
  AOI21_X1 U16485 ( .B1(n15353), .B2(n14759), .A(n14757), .ZN(n14734) );
  INV_X1 U16486 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n14733) );
  AND2_X1 U16487 ( .A1(n14730), .A2(n15410), .ZN(n14758) );
  AOI22_X1 U16488 ( .A1(n15349), .A2(n14758), .B1(n15395), .B2(n14731), .ZN(
        n14732) );
  OAI221_X1 U16489 ( .B1(n15398), .B2(n14734), .C1(n15396), .C2(n14733), .A(
        n14732), .ZN(P3_U3221) );
  XNOR2_X1 U16490 ( .A(n14735), .B(n14737), .ZN(n14762) );
  XOR2_X1 U16491 ( .A(n14737), .B(n14736), .Z(n14738) );
  OAI222_X1 U16492 ( .A1(n15381), .A2(n14740), .B1(n15382), .B2(n14739), .C1(
        n14738), .C2(n15388), .ZN(n14760) );
  AOI21_X1 U16493 ( .B1(n14762), .B2(n15353), .A(n14760), .ZN(n14744) );
  AND2_X1 U16494 ( .A1(n14741), .A2(n15410), .ZN(n14761) );
  AOI22_X1 U16495 ( .A1(n15349), .A2(n14761), .B1(n15395), .B2(n14742), .ZN(
        n14743) );
  OAI221_X1 U16496 ( .B1(n15398), .B2(n14744), .C1(n15396), .C2(n15286), .A(
        n14743), .ZN(P3_U3222) );
  OR2_X1 U16497 ( .A1(n14745), .A2(n15346), .ZN(n14747) );
  INV_X1 U16498 ( .A(n14749), .ZN(n14746) );
  AOI22_X1 U16499 ( .A1(n15438), .A2(n14764), .B1(n14748), .B2(n15439), .ZN(
        P3_U3490) );
  AOI21_X1 U16500 ( .B1(n15410), .B2(n12380), .A(n14749), .ZN(n14766) );
  AOI22_X1 U16501 ( .A1(n15438), .A2(n14766), .B1(n14750), .B2(n15439), .ZN(
        P3_U3489) );
  AOI211_X1 U16502 ( .C1(n14753), .C2(n15411), .A(n14752), .B(n14751), .ZN(
        n14768) );
  AOI22_X1 U16503 ( .A1(n15438), .A2(n14768), .B1(n7900), .B2(n15439), .ZN(
        P3_U3473) );
  AOI211_X1 U16504 ( .C1(n14756), .C2(n15411), .A(n14755), .B(n14754), .ZN(
        n14770) );
  AOI22_X1 U16505 ( .A1(n15438), .A2(n14770), .B1(n7883), .B2(n15439), .ZN(
        P3_U3472) );
  AOI211_X1 U16506 ( .C1(n15411), .C2(n14759), .A(n14758), .B(n14757), .ZN(
        n14772) );
  AOI22_X1 U16507 ( .A1(n15438), .A2(n14772), .B1(n12033), .B2(n15439), .ZN(
        P3_U3471) );
  AOI211_X1 U16508 ( .C1(n14762), .C2(n15411), .A(n14761), .B(n14760), .ZN(
        n14774) );
  AOI22_X1 U16509 ( .A1(n15438), .A2(n14774), .B1(n7841), .B2(n15439), .ZN(
        P3_U3470) );
  INV_X1 U16510 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14763) );
  AOI22_X1 U16511 ( .A1(n15430), .A2(n14764), .B1(n14763), .B2(n15428), .ZN(
        P3_U3458) );
  INV_X1 U16512 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14765) );
  AOI22_X1 U16513 ( .A1(n15430), .A2(n14766), .B1(n14765), .B2(n15428), .ZN(
        P3_U3457) );
  INV_X1 U16514 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14767) );
  AOI22_X1 U16515 ( .A1(n15430), .A2(n14768), .B1(n14767), .B2(n15428), .ZN(
        P3_U3432) );
  INV_X1 U16516 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14769) );
  AOI22_X1 U16517 ( .A1(n15430), .A2(n14770), .B1(n14769), .B2(n15428), .ZN(
        P3_U3429) );
  INV_X1 U16518 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14771) );
  AOI22_X1 U16519 ( .A1(n15430), .A2(n14772), .B1(n14771), .B2(n15428), .ZN(
        P3_U3426) );
  INV_X1 U16520 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14773) );
  AOI22_X1 U16521 ( .A1(n15430), .A2(n14774), .B1(n14773), .B2(n15428), .ZN(
        P3_U3423) );
  OAI21_X1 U16522 ( .B1(n14776), .B2(n15235), .A(n14775), .ZN(n14779) );
  INV_X1 U16523 ( .A(n14777), .ZN(n14778) );
  AOI211_X1 U16524 ( .C1(n15212), .C2(n14780), .A(n14779), .B(n14778), .ZN(
        n14798) );
  AOI22_X1 U16525 ( .A1(n15250), .A2(n14798), .B1(n14781), .B2(n9959), .ZN(
        P2_U3513) );
  NAND2_X1 U16526 ( .A1(n14782), .A2(n15200), .ZN(n14783) );
  AND2_X1 U16527 ( .A1(n14784), .A2(n14783), .ZN(n14787) );
  NAND2_X1 U16528 ( .A1(n14785), .A2(n15212), .ZN(n14786) );
  AND3_X1 U16529 ( .A1(n14788), .A2(n14787), .A3(n14786), .ZN(n14800) );
  AOI22_X1 U16530 ( .A1(n15250), .A2(n14800), .B1(n14789), .B2(n9959), .ZN(
        P2_U3512) );
  INV_X1 U16531 ( .A(n14790), .ZN(n14796) );
  NOR2_X1 U16532 ( .A1(n14790), .A2(n9942), .ZN(n14795) );
  OAI211_X1 U16533 ( .C1(n14793), .C2(n15235), .A(n14792), .B(n14791), .ZN(
        n14794) );
  AOI211_X1 U16534 ( .C1(n15239), .C2(n14796), .A(n14795), .B(n14794), .ZN(
        n14802) );
  AOI22_X1 U16535 ( .A1(n15250), .A2(n14802), .B1(n11958), .B2(n9959), .ZN(
        P2_U3511) );
  INV_X1 U16536 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14797) );
  AOI22_X1 U16537 ( .A1(n15242), .A2(n14798), .B1(n14797), .B2(n15240), .ZN(
        P2_U3472) );
  INV_X1 U16538 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14799) );
  AOI22_X1 U16539 ( .A1(n15242), .A2(n14800), .B1(n14799), .B2(n15240), .ZN(
        P2_U3469) );
  AOI22_X1 U16540 ( .A1(n15242), .A2(n14802), .B1(n14801), .B2(n15240), .ZN(
        P2_U3466) );
  AND2_X1 U16541 ( .A1(n14803), .A2(n14442), .ZN(n14808) );
  INV_X1 U16542 ( .A(n14804), .ZN(n14806) );
  OAI21_X1 U16543 ( .B1(n14806), .B2(n15025), .A(n14805), .ZN(n14807) );
  NOR3_X1 U16544 ( .A1(n14809), .A2(n14808), .A3(n14807), .ZN(n14840) );
  AOI22_X1 U16545 ( .A1(n15045), .A2(n14840), .B1(n14204), .B2(n15043), .ZN(
        P1_U3544) );
  INV_X1 U16546 ( .A(n14810), .ZN(n14817) );
  INV_X1 U16547 ( .A(n14811), .ZN(n14812) );
  OAI211_X1 U16548 ( .C1(n14814), .C2(n15025), .A(n14813), .B(n14812), .ZN(
        n14816) );
  AOI211_X1 U16549 ( .C1(n14442), .C2(n14817), .A(n14816), .B(n14815), .ZN(
        n14841) );
  AOI22_X1 U16550 ( .A1(n15045), .A2(n14841), .B1(n14818), .B2(n15043), .ZN(
        P1_U3543) );
  AND3_X1 U16551 ( .A1(n12085), .A2(n14442), .A3(n14819), .ZN(n14822) );
  NOR2_X1 U16552 ( .A1(n10067), .A2(n15025), .ZN(n14821) );
  NOR4_X1 U16553 ( .A1(n14824), .A2(n14823), .A3(n14822), .A4(n14821), .ZN(
        n14842) );
  AOI22_X1 U16554 ( .A1(n15045), .A2(n14842), .B1(n11891), .B2(n15043), .ZN(
        P1_U3542) );
  NOR2_X1 U16555 ( .A1(n14826), .A2(n14825), .ZN(n14832) );
  INV_X1 U16556 ( .A(n14827), .ZN(n14828) );
  OAI22_X1 U16557 ( .A1(n14830), .A2(n14829), .B1(n14828), .B2(n15025), .ZN(
        n14831) );
  NOR3_X1 U16558 ( .A1(n14833), .A2(n14832), .A3(n14831), .ZN(n14843) );
  AOI22_X1 U16559 ( .A1(n15045), .A2(n14843), .B1(n11620), .B2(n15043), .ZN(
        P1_U3541) );
  INV_X1 U16560 ( .A(n14834), .ZN(n14835) );
  OAI21_X1 U16561 ( .B1(n7189), .B2(n15025), .A(n14835), .ZN(n14838) );
  INV_X1 U16562 ( .A(n14836), .ZN(n14837) );
  AOI211_X1 U16563 ( .C1(n14839), .C2(n14442), .A(n14838), .B(n14837), .ZN(
        n14844) );
  AOI22_X1 U16564 ( .A1(n15045), .A2(n14844), .B1(n11110), .B2(n15043), .ZN(
        P1_U3539) );
  AOI22_X1 U16565 ( .A1(n15030), .A2(n14840), .B1(n9229), .B2(n15029), .ZN(
        P1_U3507) );
  AOI22_X1 U16566 ( .A1(n15030), .A2(n14841), .B1(n9212), .B2(n15029), .ZN(
        P1_U3504) );
  AOI22_X1 U16567 ( .A1(n15030), .A2(n14842), .B1(n9179), .B2(n15029), .ZN(
        P1_U3501) );
  AOI22_X1 U16568 ( .A1(n15030), .A2(n14843), .B1(n9186), .B2(n15029), .ZN(
        P1_U3498) );
  AOI22_X1 U16569 ( .A1(n15030), .A2(n14844), .B1(n9137), .B2(n15029), .ZN(
        P1_U3492) );
  AOI21_X1 U16570 ( .B1(n14847), .B2(n14846), .A(n14845), .ZN(n14848) );
  XNOR2_X1 U16571 ( .A(n14848), .B(n15092), .ZN(SUB_1596_U69) );
  XNOR2_X1 U16572 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14849), .ZN(SUB_1596_U68)
         );
  XNOR2_X1 U16573 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n14850), .ZN(SUB_1596_U66)
         );
  XNOR2_X1 U16574 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14851), .ZN(SUB_1596_U65)
         );
  AOI21_X1 U16575 ( .B1(n14854), .B2(n14853), .A(n14852), .ZN(n14855) );
  XNOR2_X1 U16576 ( .A(n14855), .B(n15128), .ZN(SUB_1596_U64) );
  OAI21_X1 U16577 ( .B1(n14857), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14856), .ZN(
        n14859) );
  XNOR2_X1 U16578 ( .A(n14859), .B(n14858), .ZN(n14863) );
  AOI22_X1 U16579 ( .A1(n14860), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14861) );
  OAI21_X1 U16580 ( .B1(n14863), .B2(n14862), .A(n14861), .ZN(P1_U3243) );
  AOI211_X1 U16581 ( .C1(n14867), .C2(n14866), .A(n14865), .B(n14864), .ZN(
        n14873) );
  AOI211_X1 U16582 ( .C1(n14871), .C2(n14870), .A(n14869), .B(n14868), .ZN(
        n14872) );
  AOI211_X1 U16583 ( .C1(n14875), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n14877) );
  OAI211_X1 U16584 ( .C1(n14878), .C2(n14912), .A(n14877), .B(n14876), .ZN(
        P1_U3259) );
  INV_X1 U16585 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14893) );
  AOI21_X1 U16586 ( .B1(n14881), .B2(n14880), .A(n14879), .ZN(n14882) );
  NAND2_X1 U16587 ( .A1(n14898), .A2(n14882), .ZN(n14888) );
  AOI21_X1 U16588 ( .B1(n14885), .B2(n14884), .A(n14883), .ZN(n14886) );
  NAND2_X1 U16589 ( .A1(n14903), .A2(n14886), .ZN(n14887) );
  OAI211_X1 U16590 ( .C1(n14907), .C2(n14889), .A(n14888), .B(n14887), .ZN(
        n14890) );
  INV_X1 U16591 ( .A(n14890), .ZN(n14892) );
  OAI211_X1 U16592 ( .C1(n14893), .C2(n14912), .A(n14892), .B(n14891), .ZN(
        P1_U3260) );
  AOI21_X1 U16593 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14897) );
  NAND2_X1 U16594 ( .A1(n14898), .A2(n14897), .ZN(n14905) );
  AOI21_X1 U16595 ( .B1(n14901), .B2(n14900), .A(n14899), .ZN(n14902) );
  NAND2_X1 U16596 ( .A1(n14903), .A2(n14902), .ZN(n14904) );
  OAI211_X1 U16597 ( .C1(n14907), .C2(n14906), .A(n14905), .B(n14904), .ZN(
        n14908) );
  INV_X1 U16598 ( .A(n14908), .ZN(n14911) );
  INV_X1 U16599 ( .A(n14909), .ZN(n14910) );
  OAI211_X1 U16600 ( .C1(n14913), .C2(n14912), .A(n14911), .B(n14910), .ZN(
        P1_U3261) );
  XNOR2_X1 U16601 ( .A(n14914), .B(n14916), .ZN(n15003) );
  NAND3_X1 U16602 ( .A1(n11385), .A2(n14916), .A3(n14915), .ZN(n14918) );
  AOI21_X1 U16603 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(n14920) );
  AOI211_X1 U16604 ( .C1(n15020), .C2(n15003), .A(n14921), .B(n14920), .ZN(
        n15000) );
  NOR2_X1 U16605 ( .A1(n14940), .A2(n14922), .ZN(n14923) );
  AOI21_X1 U16606 ( .B1(n14942), .B2(P1_REG2_REG_6__SCAN_IN), .A(n14923), .ZN(
        n14924) );
  OAI21_X1 U16607 ( .B1(n14944), .B2(n14999), .A(n14924), .ZN(n14925) );
  INV_X1 U16608 ( .A(n14925), .ZN(n14933) );
  INV_X1 U16609 ( .A(n14926), .ZN(n14931) );
  INV_X1 U16610 ( .A(n14927), .ZN(n14929) );
  OAI211_X1 U16611 ( .C1(n14929), .C2(n14999), .A(n14948), .B(n14928), .ZN(
        n14998) );
  INV_X1 U16612 ( .A(n14998), .ZN(n14930) );
  AOI22_X1 U16613 ( .A1(n15003), .A2(n14931), .B1(n14953), .B2(n14930), .ZN(
        n14932) );
  OAI211_X1 U16614 ( .C1(n14942), .C2(n15000), .A(n14933), .B(n14932), .ZN(
        P1_U3287) );
  XNOR2_X1 U16615 ( .A(n14934), .B(n14935), .ZN(n14938) );
  AOI21_X1 U16616 ( .B1(n14938), .B2(n14937), .A(n14936), .ZN(n14987) );
  NOR2_X1 U16617 ( .A1(n14940), .A2(n14939), .ZN(n14941) );
  AOI21_X1 U16618 ( .B1(n14942), .B2(P1_REG2_REG_4__SCAN_IN), .A(n14941), .ZN(
        n14943) );
  OAI21_X1 U16619 ( .B1(n14944), .B2(n14988), .A(n14943), .ZN(n14945) );
  INV_X1 U16620 ( .A(n14945), .ZN(n14956) );
  XNOR2_X1 U16621 ( .A(n14947), .B(n14946), .ZN(n14990) );
  OAI21_X1 U16622 ( .B1(n14949), .B2(n14988), .A(n14948), .ZN(n14950) );
  OR2_X1 U16623 ( .A1(n14951), .A2(n14950), .ZN(n14986) );
  INV_X1 U16624 ( .A(n14986), .ZN(n14952) );
  AOI22_X1 U16625 ( .A1(n14990), .A2(n14954), .B1(n14953), .B2(n14952), .ZN(
        n14955) );
  OAI211_X1 U16626 ( .C1(n14942), .C2(n14987), .A(n14956), .B(n14955), .ZN(
        P1_U3289) );
  AND2_X1 U16627 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14962), .ZN(P1_U3294) );
  AND2_X1 U16628 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14962), .ZN(P1_U3295) );
  AND2_X1 U16629 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14962), .ZN(P1_U3296) );
  AND2_X1 U16630 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14962), .ZN(P1_U3297) );
  AND2_X1 U16631 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14962), .ZN(P1_U3298) );
  INV_X1 U16632 ( .A(n14962), .ZN(n14961) );
  NOR2_X1 U16633 ( .A1(n14961), .A2(n14957), .ZN(P1_U3299) );
  AND2_X1 U16634 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14962), .ZN(P1_U3300) );
  AND2_X1 U16635 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14962), .ZN(P1_U3301) );
  AND2_X1 U16636 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14962), .ZN(P1_U3302) );
  AND2_X1 U16637 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14962), .ZN(P1_U3303) );
  AND2_X1 U16638 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14962), .ZN(P1_U3304) );
  AND2_X1 U16639 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14962), .ZN(P1_U3305) );
  AND2_X1 U16640 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14962), .ZN(P1_U3306) );
  AND2_X1 U16641 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14962), .ZN(P1_U3307) );
  AND2_X1 U16642 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14962), .ZN(P1_U3308) );
  AND2_X1 U16643 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14962), .ZN(P1_U3309) );
  AND2_X1 U16644 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14962), .ZN(P1_U3310) );
  AND2_X1 U16645 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14962), .ZN(P1_U3311) );
  AND2_X1 U16646 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14962), .ZN(P1_U3312) );
  AND2_X1 U16647 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14962), .ZN(P1_U3313) );
  NOR2_X1 U16648 ( .A1(n14961), .A2(n14958), .ZN(P1_U3314) );
  AND2_X1 U16649 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14962), .ZN(P1_U3315) );
  NOR2_X1 U16650 ( .A1(n14961), .A2(n14959), .ZN(P1_U3316) );
  AND2_X1 U16651 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14962), .ZN(P1_U3317) );
  AND2_X1 U16652 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14962), .ZN(P1_U3318) );
  AND2_X1 U16653 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14962), .ZN(P1_U3319) );
  AND2_X1 U16654 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14962), .ZN(P1_U3320) );
  NOR2_X1 U16655 ( .A1(n14961), .A2(n14960), .ZN(P1_U3321) );
  AND2_X1 U16656 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14962), .ZN(P1_U3322) );
  AND2_X1 U16657 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14962), .ZN(P1_U3323) );
  INV_X1 U16658 ( .A(n15013), .ZN(n15004) );
  OAI21_X1 U16659 ( .B1(n14964), .B2(n15025), .A(n14963), .ZN(n14969) );
  INV_X1 U16660 ( .A(n14970), .ZN(n14967) );
  OAI21_X1 U16661 ( .B1(n14967), .B2(n14966), .A(n14965), .ZN(n14968) );
  AOI211_X1 U16662 ( .C1(n15004), .C2(n14970), .A(n14969), .B(n14968), .ZN(
        n15032) );
  AOI22_X1 U16663 ( .A1(n15030), .A2(n15032), .B1(n8939), .B2(n15029), .ZN(
        P1_U3462) );
  INV_X1 U16664 ( .A(n14971), .ZN(n14977) );
  OAI21_X1 U16665 ( .B1(n14973), .B2(n15025), .A(n14972), .ZN(n14976) );
  INV_X1 U16666 ( .A(n14974), .ZN(n14975) );
  AOI211_X1 U16667 ( .C1(n15004), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        n15034) );
  AOI22_X1 U16668 ( .A1(n15030), .A2(n15034), .B1(n8953), .B2(n15029), .ZN(
        P1_U3465) );
  INV_X1 U16669 ( .A(n14983), .ZN(n14985) );
  AOI21_X1 U16670 ( .B1(n14980), .B2(n14979), .A(n14978), .ZN(n14981) );
  OAI211_X1 U16671 ( .C1(n15013), .C2(n14983), .A(n14982), .B(n14981), .ZN(
        n14984) );
  AOI21_X1 U16672 ( .B1(n15020), .B2(n14985), .A(n14984), .ZN(n15036) );
  AOI22_X1 U16673 ( .A1(n15030), .A2(n15036), .B1(n8973), .B2(n15029), .ZN(
        P1_U3468) );
  OAI211_X1 U16674 ( .C1(n14988), .C2(n15025), .A(n14987), .B(n14986), .ZN(
        n14989) );
  AOI21_X1 U16675 ( .B1(n14990), .B2(n14442), .A(n14989), .ZN(n15038) );
  AOI22_X1 U16676 ( .A1(n15030), .A2(n15038), .B1(n9018), .B2(n15029), .ZN(
        P1_U3471) );
  INV_X1 U16677 ( .A(n14991), .ZN(n14997) );
  NOR2_X1 U16678 ( .A1(n14991), .A2(n15013), .ZN(n14996) );
  OAI211_X1 U16679 ( .C1(n14994), .C2(n15025), .A(n14993), .B(n14992), .ZN(
        n14995) );
  AOI211_X1 U16680 ( .C1(n15020), .C2(n14997), .A(n14996), .B(n14995), .ZN(
        n15039) );
  AOI22_X1 U16681 ( .A1(n15030), .A2(n15039), .B1(n9035), .B2(n15029), .ZN(
        P1_U3474) );
  OAI21_X1 U16682 ( .B1(n14999), .B2(n15025), .A(n14998), .ZN(n15002) );
  INV_X1 U16683 ( .A(n15000), .ZN(n15001) );
  AOI211_X1 U16684 ( .C1(n15004), .C2(n15003), .A(n15002), .B(n15001), .ZN(
        n15040) );
  AOI22_X1 U16685 ( .A1(n15030), .A2(n15040), .B1(n9050), .B2(n15029), .ZN(
        P1_U3477) );
  AND2_X1 U16686 ( .A1(n15005), .A2(n15020), .ZN(n15012) );
  AND2_X1 U16687 ( .A1(n15005), .A2(n15004), .ZN(n15011) );
  INV_X1 U16688 ( .A(n15006), .ZN(n15008) );
  OAI21_X1 U16689 ( .B1(n15008), .B2(n15025), .A(n15007), .ZN(n15009) );
  NOR4_X1 U16690 ( .A1(n15012), .A2(n15011), .A3(n15010), .A4(n15009), .ZN(
        n15041) );
  AOI22_X1 U16691 ( .A1(n15030), .A2(n15041), .B1(n9066), .B2(n15029), .ZN(
        P1_U3480) );
  INV_X1 U16692 ( .A(n15014), .ZN(n15021) );
  NOR2_X1 U16693 ( .A1(n15014), .A2(n15013), .ZN(n15019) );
  OAI211_X1 U16694 ( .C1(n15017), .C2(n15025), .A(n15016), .B(n15015), .ZN(
        n15018) );
  AOI211_X1 U16695 ( .C1(n15021), .C2(n15020), .A(n15019), .B(n15018), .ZN(
        n15042) );
  AOI22_X1 U16696 ( .A1(n15030), .A2(n15042), .B1(n9102), .B2(n15029), .ZN(
        P1_U3486) );
  INV_X1 U16697 ( .A(n15022), .ZN(n15026) );
  OAI211_X1 U16698 ( .C1(n15026), .C2(n15025), .A(n15024), .B(n15023), .ZN(
        n15027) );
  AOI21_X1 U16699 ( .B1(n14442), .B2(n15028), .A(n15027), .ZN(n15044) );
  AOI22_X1 U16700 ( .A1(n15030), .A2(n15044), .B1(n9113), .B2(n15029), .ZN(
        P1_U3489) );
  AOI22_X1 U16701 ( .A1(n15045), .A2(n15032), .B1(n15031), .B2(n15043), .ZN(
        P1_U3529) );
  AOI22_X1 U16702 ( .A1(n15045), .A2(n15034), .B1(n15033), .B2(n15043), .ZN(
        P1_U3530) );
  AOI22_X1 U16703 ( .A1(n15045), .A2(n15036), .B1(n15035), .B2(n15043), .ZN(
        P1_U3531) );
  AOI22_X1 U16704 ( .A1(n15045), .A2(n15038), .B1(n15037), .B2(n15043), .ZN(
        P1_U3532) );
  AOI22_X1 U16705 ( .A1(n15045), .A2(n15039), .B1(n10614), .B2(n15043), .ZN(
        P1_U3533) );
  AOI22_X1 U16706 ( .A1(n15045), .A2(n15040), .B1(n10607), .B2(n15043), .ZN(
        P1_U3534) );
  AOI22_X1 U16707 ( .A1(n15045), .A2(n15041), .B1(n9063), .B2(n15043), .ZN(
        P1_U3535) );
  AOI22_X1 U16708 ( .A1(n15045), .A2(n15042), .B1(n10701), .B2(n15043), .ZN(
        P1_U3537) );
  AOI22_X1 U16709 ( .A1(n15045), .A2(n15044), .B1(n10811), .B2(n15043), .ZN(
        P1_U3538) );
  NOR2_X1 U16710 ( .A1(n15056), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16711 ( .A1(n15056), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15055) );
  NAND2_X1 U16712 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15047) );
  AOI211_X1 U16713 ( .C1(n15047), .C2(n6703), .A(n15046), .B(n15135), .ZN(
        n15052) );
  AOI211_X1 U16714 ( .C1(n15050), .C2(n15049), .A(n15048), .B(n15120), .ZN(
        n15051) );
  AOI211_X1 U16715 ( .C1(n15141), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        n15054) );
  NAND2_X1 U16716 ( .A1(n15055), .A2(n15054), .ZN(P2_U3215) );
  AOI22_X1 U16717 ( .A1(n15056), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15067) );
  AOI211_X1 U16718 ( .C1(n15059), .C2(n15058), .A(n15057), .B(n15135), .ZN(
        n15064) );
  AOI211_X1 U16719 ( .C1(n15062), .C2(n15061), .A(n15060), .B(n15120), .ZN(
        n15063) );
  AOI211_X1 U16720 ( .C1(n15141), .C2(n15065), .A(n15064), .B(n15063), .ZN(
        n15066) );
  NAND2_X1 U16721 ( .A1(n15067), .A2(n15066), .ZN(P2_U3216) );
  AOI211_X1 U16722 ( .C1(n15070), .C2(n15069), .A(n15135), .B(n15068), .ZN(
        n15075) );
  AOI211_X1 U16723 ( .C1(n15073), .C2(n15072), .A(n15120), .B(n15071), .ZN(
        n15074) );
  AOI211_X1 U16724 ( .C1(n15141), .C2(n15076), .A(n15075), .B(n15074), .ZN(
        n15078) );
  NAND2_X1 U16725 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n15077)
         );
  OAI211_X1 U16726 ( .C1(n15079), .C2(n15144), .A(n15078), .B(n15077), .ZN(
        P2_U3224) );
  AOI211_X1 U16727 ( .C1(n15082), .C2(n15081), .A(n15135), .B(n15080), .ZN(
        n15088) );
  OAI21_X1 U16728 ( .B1(n15085), .B2(n15084), .A(n15083), .ZN(n15086) );
  AND2_X1 U16729 ( .A1(n15086), .A2(n15129), .ZN(n15087) );
  AOI211_X1 U16730 ( .C1(n15141), .C2(n15089), .A(n15088), .B(n15087), .ZN(
        n15091) );
  NAND2_X1 U16731 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n15090)
         );
  OAI211_X1 U16732 ( .C1(n15092), .C2(n15144), .A(n15091), .B(n15090), .ZN(
        P2_U3225) );
  AOI211_X1 U16733 ( .C1(n15095), .C2(n15094), .A(n15093), .B(n15135), .ZN(
        n15100) );
  AOI211_X1 U16734 ( .C1(n15098), .C2(n15097), .A(n15096), .B(n15120), .ZN(
        n15099) );
  AOI211_X1 U16735 ( .C1(n15141), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        n15103) );
  OAI211_X1 U16736 ( .C1(n7363), .C2(n15144), .A(n15103), .B(n15102), .ZN(
        P2_U3228) );
  AOI211_X1 U16737 ( .C1(n15106), .C2(n15105), .A(n15104), .B(n15120), .ZN(
        n15111) );
  AOI211_X1 U16738 ( .C1(n15109), .C2(n15108), .A(n15107), .B(n15135), .ZN(
        n15110) );
  AOI211_X1 U16739 ( .C1(n15141), .C2(n15112), .A(n15111), .B(n15110), .ZN(
        n15114) );
  NAND2_X1 U16740 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15113)
         );
  OAI211_X1 U16741 ( .C1(n7137), .C2(n15144), .A(n15114), .B(n15113), .ZN(
        P2_U3229) );
  AOI211_X1 U16742 ( .C1(n15117), .C2(n15116), .A(n15135), .B(n15115), .ZN(
        n15124) );
  INV_X1 U16743 ( .A(n15118), .ZN(n15119) );
  AOI211_X1 U16744 ( .C1(n15122), .C2(n15121), .A(n15120), .B(n15119), .ZN(
        n15123) );
  AOI211_X1 U16745 ( .C1(n15141), .C2(n15125), .A(n15124), .B(n15123), .ZN(
        n15127) );
  OAI211_X1 U16746 ( .C1(n15128), .C2(n15144), .A(n15127), .B(n15126), .ZN(
        P2_U3230) );
  INV_X1 U16747 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15145) );
  OAI211_X1 U16748 ( .C1(n15132), .C2(n15131), .A(n15130), .B(n15129), .ZN(
        n15133) );
  INV_X1 U16749 ( .A(n15133), .ZN(n15139) );
  AOI211_X1 U16750 ( .C1(n15137), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        n15138) );
  AOI211_X1 U16751 ( .C1(n15141), .C2(n15140), .A(n15139), .B(n15138), .ZN(
        n15143) );
  NAND2_X1 U16752 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n15142)
         );
  OAI211_X1 U16753 ( .C1(n15145), .C2(n15144), .A(n15143), .B(n15142), .ZN(
        P2_U3231) );
  INV_X1 U16754 ( .A(n15146), .ZN(n15153) );
  NAND2_X1 U16755 ( .A1(n15147), .A2(n15169), .ZN(n15151) );
  AOI22_X1 U16756 ( .A1(n15149), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n15148), 
        .B2(n15163), .ZN(n15150) );
  OAI211_X1 U16757 ( .C1(n15153), .C2(n15152), .A(n15151), .B(n15150), .ZN(
        n15154) );
  AOI21_X1 U16758 ( .B1(n15168), .B2(n15155), .A(n15154), .ZN(n15156) );
  OAI21_X1 U16759 ( .B1(n15174), .B2(n15157), .A(n15156), .ZN(P2_U3258) );
  INV_X1 U16760 ( .A(n15159), .ZN(n15160) );
  AOI21_X1 U16761 ( .B1(n15162), .B2(n15161), .A(n15160), .ZN(n15193) );
  AOI22_X1 U16762 ( .A1(n15163), .A2(P2_REG3_REG_1__SCAN_IN), .B1(
        P2_REG2_REG_1__SCAN_IN), .B2(n15174), .ZN(n15173) );
  INV_X1 U16763 ( .A(n15164), .ZN(n15165) );
  AOI211_X1 U16764 ( .C1(n15166), .C2(n15171), .A(n11852), .B(n15165), .ZN(
        n15190) );
  AOI222_X1 U16765 ( .A1(n15171), .A2(n15170), .B1(n15169), .B2(n15190), .C1(
        n15196), .C2(n15168), .ZN(n15172) );
  OAI211_X1 U16766 ( .C1(n15174), .C2(n15193), .A(n15173), .B(n15172), .ZN(
        P2_U3264) );
  INV_X1 U16767 ( .A(n15175), .ZN(n15176) );
  AND2_X1 U16768 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15180), .ZN(P2_U3266) );
  AND2_X1 U16769 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15180), .ZN(P2_U3267) );
  AND2_X1 U16770 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15180), .ZN(P2_U3268) );
  AND2_X1 U16771 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15180), .ZN(P2_U3269) );
  AND2_X1 U16772 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15180), .ZN(P2_U3270) );
  AND2_X1 U16773 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15180), .ZN(P2_U3271) );
  AND2_X1 U16774 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15180), .ZN(P2_U3272) );
  AND2_X1 U16775 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15180), .ZN(P2_U3273) );
  AND2_X1 U16776 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15180), .ZN(P2_U3274) );
  INV_X1 U16777 ( .A(n15180), .ZN(n15179) );
  NOR2_X1 U16778 ( .A1(n15179), .A2(n15177), .ZN(P2_U3275) );
  AND2_X1 U16779 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15180), .ZN(P2_U3276) );
  AND2_X1 U16780 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15180), .ZN(P2_U3277) );
  AND2_X1 U16781 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15180), .ZN(P2_U3278) );
  AND2_X1 U16782 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15180), .ZN(P2_U3279) );
  NOR2_X1 U16783 ( .A1(n15179), .A2(n15178), .ZN(P2_U3280) );
  AND2_X1 U16784 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15180), .ZN(P2_U3281) );
  AND2_X1 U16785 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15180), .ZN(P2_U3282) );
  AND2_X1 U16786 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15180), .ZN(P2_U3283) );
  AND2_X1 U16787 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15180), .ZN(P2_U3284) );
  AND2_X1 U16788 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15180), .ZN(P2_U3285) );
  AND2_X1 U16789 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15180), .ZN(P2_U3286) );
  AND2_X1 U16790 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15180), .ZN(P2_U3287) );
  AND2_X1 U16791 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15180), .ZN(P2_U3288) );
  AND2_X1 U16792 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15180), .ZN(P2_U3289) );
  AND2_X1 U16793 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15180), .ZN(P2_U3290) );
  AND2_X1 U16794 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15180), .ZN(P2_U3291) );
  AND2_X1 U16795 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15180), .ZN(P2_U3292) );
  AND2_X1 U16796 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15180), .ZN(P2_U3293) );
  AND2_X1 U16797 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15180), .ZN(P2_U3294) );
  AND2_X1 U16798 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15180), .ZN(P2_U3295) );
  INV_X1 U16799 ( .A(n15187), .ZN(n15184) );
  AOI22_X1 U16800 ( .A1(n15187), .A2(n15182), .B1(n15181), .B2(n15184), .ZN(
        P2_U3416) );
  INV_X1 U16801 ( .A(n15183), .ZN(n15186) );
  AOI22_X1 U16802 ( .A1(n15187), .A2(n15186), .B1(n15185), .B2(n15184), .ZN(
        P2_U3417) );
  AOI22_X1 U16803 ( .A1(n15242), .A2(n15189), .B1(n15188), .B2(n15240), .ZN(
        P2_U3430) );
  INV_X1 U16804 ( .A(n15190), .ZN(n15191) );
  OAI21_X1 U16805 ( .B1(n15192), .B2(n15235), .A(n15191), .ZN(n15195) );
  INV_X1 U16806 ( .A(n15193), .ZN(n15194) );
  AOI211_X1 U16807 ( .C1(n15196), .C2(n15212), .A(n15195), .B(n15194), .ZN(
        n15244) );
  INV_X1 U16808 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15197) );
  AOI22_X1 U16809 ( .A1(n15242), .A2(n15244), .B1(n15197), .B2(n15240), .ZN(
        P2_U3433) );
  AOI21_X1 U16810 ( .B1(n15200), .B2(n15199), .A(n15198), .ZN(n15204) );
  INV_X1 U16811 ( .A(n9942), .ZN(n15202) );
  OAI21_X1 U16812 ( .B1(n15202), .B2(n15239), .A(n15201), .ZN(n15203) );
  AND3_X1 U16813 ( .A1(n15205), .A2(n15204), .A3(n15203), .ZN(n15245) );
  INV_X1 U16814 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15206) );
  AOI22_X1 U16815 ( .A1(n15242), .A2(n15245), .B1(n15206), .B2(n15240), .ZN(
        P2_U3436) );
  INV_X1 U16816 ( .A(n15207), .ZN(n15213) );
  OAI21_X1 U16817 ( .B1(n15209), .B2(n15235), .A(n15208), .ZN(n15211) );
  AOI211_X1 U16818 ( .C1(n15213), .C2(n15212), .A(n15211), .B(n15210), .ZN(
        n15246) );
  INV_X1 U16819 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15214) );
  AOI22_X1 U16820 ( .A1(n15242), .A2(n15246), .B1(n15214), .B2(n15240), .ZN(
        P2_U3439) );
  OAI211_X1 U16821 ( .C1(n15217), .C2(n15235), .A(n15216), .B(n15215), .ZN(
        n15220) );
  AOI21_X1 U16822 ( .B1(n9942), .B2(n15223), .A(n15218), .ZN(n15219) );
  NOR2_X1 U16823 ( .A1(n15220), .A2(n15219), .ZN(n15247) );
  INV_X1 U16824 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15221) );
  AOI22_X1 U16825 ( .A1(n15242), .A2(n15247), .B1(n15221), .B2(n15240), .ZN(
        P2_U3442) );
  AOI21_X1 U16826 ( .B1(n9942), .B2(n15223), .A(n15222), .ZN(n15229) );
  INV_X1 U16827 ( .A(n15224), .ZN(n15225) );
  OAI211_X1 U16828 ( .C1(n15227), .C2(n15235), .A(n15226), .B(n15225), .ZN(
        n15228) );
  NOR2_X1 U16829 ( .A1(n15229), .A2(n15228), .ZN(n15248) );
  INV_X1 U16830 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U16831 ( .A1(n15242), .A2(n15248), .B1(n15230), .B2(n15240), .ZN(
        P2_U3445) );
  INV_X1 U16832 ( .A(n15231), .ZN(n15238) );
  NOR2_X1 U16833 ( .A1(n15231), .A2(n9942), .ZN(n15237) );
  OAI211_X1 U16834 ( .C1(n6967), .C2(n15235), .A(n15234), .B(n15233), .ZN(
        n15236) );
  AOI211_X1 U16835 ( .C1(n15239), .C2(n15238), .A(n15237), .B(n15236), .ZN(
        n15249) );
  INV_X1 U16836 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15241) );
  AOI22_X1 U16837 ( .A1(n15242), .A2(n15249), .B1(n15241), .B2(n15240), .ZN(
        P2_U3460) );
  AOI22_X1 U16838 ( .A1(n15250), .A2(n15244), .B1(n15243), .B2(n9959), .ZN(
        P2_U3500) );
  AOI22_X1 U16839 ( .A1(n15250), .A2(n15245), .B1(n10554), .B2(n9959), .ZN(
        P2_U3501) );
  AOI22_X1 U16840 ( .A1(n15250), .A2(n15246), .B1(n10555), .B2(n9959), .ZN(
        P2_U3502) );
  AOI22_X1 U16841 ( .A1(n15250), .A2(n15247), .B1(n10573), .B2(n9959), .ZN(
        P2_U3503) );
  AOI22_X1 U16842 ( .A1(n15250), .A2(n15248), .B1(n10575), .B2(n9959), .ZN(
        P2_U3504) );
  AOI22_X1 U16843 ( .A1(n15250), .A2(n15249), .B1(n11961), .B2(n9959), .ZN(
        P2_U3509) );
  NOR2_X1 U16844 ( .A1(P3_U3897), .A2(n15274), .ZN(P3_U3150) );
  NOR3_X1 U16845 ( .A1(n15254), .A2(n15252), .A3(n15279), .ZN(n15264) );
  AOI22_X1 U16846 ( .A1(n15254), .A2(n15253), .B1(n15252), .B2(n15251), .ZN(
        n15262) );
  MUX2_X1 U16847 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n15255), .Z(n15256) );
  AND2_X1 U16848 ( .A1(n15279), .A2(n15256), .ZN(n15257) );
  MUX2_X1 U16849 ( .A(n15257), .B(n15281), .S(P3_IR_REG_0__SCAN_IN), .Z(n15260) );
  OAI22_X1 U16850 ( .A1(n15287), .A2(n15258), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10843), .ZN(n15259) );
  NOR2_X1 U16851 ( .A1(n15260), .A2(n15259), .ZN(n15261) );
  OAI211_X1 U16852 ( .C1(n15264), .C2(n15263), .A(n15262), .B(n15261), .ZN(
        P3_U3182) );
  AOI21_X1 U16853 ( .B1(n15267), .B2(n15266), .A(n15265), .ZN(n15271) );
  AOI21_X1 U16854 ( .B1(n7771), .B2(n15269), .A(n15268), .ZN(n15270) );
  OAI22_X1 U16855 ( .A1(n15271), .A2(n15304), .B1(n15270), .B2(n15298), .ZN(
        n15272) );
  AOI211_X1 U16856 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n15274), .A(n15273), .B(
        n15272), .ZN(n15283) );
  OAI21_X1 U16857 ( .B1(n15277), .B2(n15276), .A(n15275), .ZN(n15278) );
  AOI22_X1 U16858 ( .A1(n15281), .A2(n15280), .B1(n15279), .B2(n15278), .ZN(
        n15282) );
  NAND2_X1 U16859 ( .A1(n15283), .A2(n15282), .ZN(P3_U3189) );
  AOI21_X1 U16860 ( .B1(n15286), .B2(n15285), .A(n15284), .ZN(n15305) );
  OAI22_X1 U16861 ( .A1(n15290), .A2(n15289), .B1(n15288), .B2(n15287), .ZN(
        n15301) );
  AOI21_X1 U16862 ( .B1(n7841), .B2(n15292), .A(n15291), .ZN(n15299) );
  AOI21_X1 U16863 ( .B1(n15295), .B2(n15294), .A(n15293), .ZN(n15297) );
  OAI22_X1 U16864 ( .A1(n15299), .A2(n15298), .B1(n15297), .B2(n15296), .ZN(
        n15300) );
  NOR3_X1 U16865 ( .A1(n15302), .A2(n15301), .A3(n15300), .ZN(n15303) );
  OAI21_X1 U16866 ( .B1(n15305), .B2(n15304), .A(n15303), .ZN(P3_U3193) );
  XNOR2_X1 U16867 ( .A(n15306), .B(n8127), .ZN(n15313) );
  INV_X1 U16868 ( .A(n15313), .ZN(n15427) );
  OAI211_X1 U16869 ( .C1(n15308), .C2(n8127), .A(n15341), .B(n15307), .ZN(
        n15312) );
  AOI22_X1 U16870 ( .A1(n15326), .A2(n15310), .B1(n15324), .B2(n15309), .ZN(
        n15311) );
  OAI211_X1 U16871 ( .C1(n15345), .C2(n15313), .A(n15312), .B(n15311), .ZN(
        n15424) );
  AOI21_X1 U16872 ( .B1(n15390), .B2(n15427), .A(n15424), .ZN(n15317) );
  AND2_X1 U16873 ( .A1(n15314), .A2(n15410), .ZN(n15425) );
  AOI22_X1 U16874 ( .A1(n15349), .A2(n15425), .B1(n15395), .B2(n15315), .ZN(
        n15316) );
  OAI221_X1 U16875 ( .B1(n15398), .B2(n15317), .C1(n15396), .C2(n12041), .A(
        n15316), .ZN(P3_U3223) );
  XNOR2_X1 U16876 ( .A(n15318), .B(n15322), .ZN(n15422) );
  INV_X1 U16877 ( .A(n15319), .ZN(n15320) );
  AOI21_X1 U16878 ( .B1(n15322), .B2(n15321), .A(n15320), .ZN(n15329) );
  AOI22_X1 U16879 ( .A1(n15326), .A2(n15325), .B1(n15324), .B2(n15323), .ZN(
        n15328) );
  NAND2_X1 U16880 ( .A1(n15422), .A2(n15385), .ZN(n15327) );
  OAI211_X1 U16881 ( .C1(n15329), .C2(n15388), .A(n15328), .B(n15327), .ZN(
        n15420) );
  AOI21_X1 U16882 ( .B1(n15390), .B2(n15422), .A(n15420), .ZN(n15334) );
  AND2_X1 U16883 ( .A1(n15330), .A2(n15410), .ZN(n15421) );
  AOI22_X1 U16884 ( .A1(n15349), .A2(n15421), .B1(n15395), .B2(n15331), .ZN(
        n15332) );
  OAI221_X1 U16885 ( .B1(n15398), .B2(n15334), .C1(n15396), .C2(n15333), .A(
        n15332), .ZN(P3_U3224) );
  XNOR2_X1 U16886 ( .A(n15335), .B(n15336), .ZN(n15344) );
  INV_X1 U16887 ( .A(n15344), .ZN(n15418) );
  XOR2_X1 U16888 ( .A(n15337), .B(n15336), .Z(n15342) );
  OAI22_X1 U16889 ( .A1(n15339), .A2(n15382), .B1(n15338), .B2(n15381), .ZN(
        n15340) );
  AOI21_X1 U16890 ( .B1(n15342), .B2(n15341), .A(n15340), .ZN(n15343) );
  OAI21_X1 U16891 ( .B1(n15345), .B2(n15344), .A(n15343), .ZN(n15416) );
  AOI21_X1 U16892 ( .B1(n15390), .B2(n15418), .A(n15416), .ZN(n15352) );
  NOR2_X1 U16893 ( .A1(n15347), .A2(n15346), .ZN(n15417) );
  AOI22_X1 U16894 ( .A1(n15349), .A2(n15417), .B1(n15395), .B2(n15348), .ZN(
        n15350) );
  OAI221_X1 U16895 ( .B1(n15398), .B2(n15352), .C1(n15396), .C2(n15351), .A(
        n15350), .ZN(P3_U3225) );
  INV_X1 U16896 ( .A(n15353), .ZN(n15369) );
  OAI21_X1 U16897 ( .B1(n15369), .B2(n15355), .A(n15354), .ZN(n15356) );
  MUX2_X1 U16898 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n15356), .S(n15396), .Z(
        n15357) );
  AOI21_X1 U16899 ( .B1(n15374), .B2(n15358), .A(n15357), .ZN(n15359) );
  OAI21_X1 U16900 ( .B1(n15360), .B2(n15376), .A(n15359), .ZN(P3_U3228) );
  OAI21_X1 U16901 ( .B1(n15362), .B2(n15369), .A(n15361), .ZN(n15363) );
  MUX2_X1 U16902 ( .A(n15363), .B(P3_REG2_REG_4__SCAN_IN), .S(n15398), .Z(
        n15364) );
  AOI21_X1 U16903 ( .B1(n15374), .B2(n15365), .A(n15364), .ZN(n15366) );
  OAI21_X1 U16904 ( .B1(n15367), .B2(n15376), .A(n15366), .ZN(P3_U3229) );
  OAI21_X1 U16905 ( .B1(n15370), .B2(n15369), .A(n15368), .ZN(n15371) );
  MUX2_X1 U16906 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n15371), .S(n15396), .Z(
        n15372) );
  AOI21_X1 U16907 ( .B1(n15374), .B2(n15373), .A(n15372), .ZN(n15375) );
  OAI21_X1 U16908 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(n15376), .A(n15375), .ZN(
        P3_U3230) );
  XNOR2_X1 U16909 ( .A(n15379), .B(n15377), .ZN(n15387) );
  OAI21_X1 U16910 ( .B1(n15380), .B2(n15379), .A(n15378), .ZN(n15389) );
  OAI22_X1 U16911 ( .A1(n15383), .A2(n15382), .B1(n8111), .B2(n15381), .ZN(
        n15384) );
  AOI21_X1 U16912 ( .B1(n15389), .B2(n15385), .A(n15384), .ZN(n15386) );
  OAI21_X1 U16913 ( .B1(n15388), .B2(n15387), .A(n15386), .ZN(n15403) );
  INV_X1 U16914 ( .A(n15389), .ZN(n15407) );
  INV_X1 U16915 ( .A(n15390), .ZN(n15393) );
  NAND2_X1 U16916 ( .A1(n15391), .A2(n15410), .ZN(n15404) );
  OAI22_X1 U16917 ( .A1(n15407), .A2(n15393), .B1(n15392), .B2(n15404), .ZN(
        n15394) );
  AOI211_X1 U16918 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15395), .A(n15403), .B(
        n15394), .ZN(n15397) );
  AOI22_X1 U16919 ( .A1(n15398), .A2(n11006), .B1(n15397), .B2(n15396), .ZN(
        P3_U3231) );
  AOI211_X1 U16920 ( .C1(n15411), .C2(n15401), .A(n15400), .B(n15399), .ZN(
        n15432) );
  INV_X1 U16921 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15402) );
  AOI22_X1 U16922 ( .A1(n15430), .A2(n15432), .B1(n15402), .B2(n15428), .ZN(
        P3_U3393) );
  INV_X1 U16923 ( .A(n15426), .ZN(n15406) );
  INV_X1 U16924 ( .A(n15403), .ZN(n15405) );
  OAI211_X1 U16925 ( .C1(n15407), .C2(n15406), .A(n15405), .B(n15404), .ZN(
        n15433) );
  OAI22_X1 U16926 ( .A1(n15428), .A2(n15433), .B1(P3_REG0_REG_2__SCAN_IN), 
        .B2(n15430), .ZN(n15408) );
  INV_X1 U16927 ( .A(n15408), .ZN(P3_U3396) );
  AOI22_X1 U16928 ( .A1(n15412), .A2(n15411), .B1(n15410), .B2(n15409), .ZN(
        n15413) );
  AND2_X1 U16929 ( .A1(n15414), .A2(n15413), .ZN(n15435) );
  INV_X1 U16930 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15415) );
  AOI22_X1 U16931 ( .A1(n15430), .A2(n15435), .B1(n15415), .B2(n15428), .ZN(
        P3_U3411) );
  AOI211_X1 U16932 ( .C1(n15426), .C2(n15418), .A(n15417), .B(n15416), .ZN(
        n15436) );
  INV_X1 U16933 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15419) );
  AOI22_X1 U16934 ( .A1(n15430), .A2(n15436), .B1(n15419), .B2(n15428), .ZN(
        P3_U3414) );
  AOI211_X1 U16935 ( .C1(n15422), .C2(n15426), .A(n15421), .B(n15420), .ZN(
        n15437) );
  INV_X1 U16936 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15423) );
  AOI22_X1 U16937 ( .A1(n15430), .A2(n15437), .B1(n15423), .B2(n15428), .ZN(
        P3_U3417) );
  AOI211_X1 U16938 ( .C1(n15427), .C2(n15426), .A(n15425), .B(n15424), .ZN(
        n15440) );
  INV_X1 U16939 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15429) );
  AOI22_X1 U16940 ( .A1(n15430), .A2(n15440), .B1(n15429), .B2(n15428), .ZN(
        P3_U3420) );
  AOI22_X1 U16941 ( .A1(n15438), .A2(n15432), .B1(n15431), .B2(n15439), .ZN(
        P3_U3460) );
  OAI22_X1 U16942 ( .A1(n15439), .A2(n15433), .B1(P3_REG1_REG_2__SCAN_IN), 
        .B2(n15438), .ZN(n15434) );
  INV_X1 U16943 ( .A(n15434), .ZN(P3_U3461) );
  AOI22_X1 U16944 ( .A1(n15438), .A2(n15435), .B1(n7771), .B2(n15439), .ZN(
        P3_U3466) );
  AOI22_X1 U16945 ( .A1(n15438), .A2(n15436), .B1(n7788), .B2(n15439), .ZN(
        P3_U3467) );
  AOI22_X1 U16946 ( .A1(n15438), .A2(n15437), .B1(n7805), .B2(n15439), .ZN(
        P3_U3468) );
  AOI22_X1 U16947 ( .A1(n15438), .A2(n15440), .B1(n12028), .B2(n15439), .ZN(
        P3_U3469) );
  XNOR2_X1 U16948 ( .A(n15441), .B(n15442), .ZN(SUB_1596_U59) );
  XNOR2_X1 U16949 ( .A(n15443), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16950 ( .B1(n15445), .B2(n15444), .A(n15453), .ZN(SUB_1596_U53) );
  XOR2_X1 U16951 ( .A(n15447), .B(n15446), .Z(SUB_1596_U56) );
  OAI21_X1 U16952 ( .B1(n15450), .B2(n15449), .A(n15448), .ZN(n15451) );
  XNOR2_X1 U16953 ( .A(n15451), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16954 ( .A(n15453), .B(n15452), .Z(SUB_1596_U5) );
  INV_X1 U7255 ( .A(n13700), .ZN(n13607) );
  CLKBUF_X1 U7274 ( .A(n7721), .Z(n9570) );
  CLKBUF_X1 U7623 ( .A(n10182), .Z(n10413) );
endmodule

