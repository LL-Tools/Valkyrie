

module b21_C_AntiSAT_k_256_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479;

  AND2_X1 U4980 ( .A1(n4627), .A2(n4509), .ZN(n9630) );
  NAND2_X1 U4981 ( .A1(n4756), .A2(n4757), .ZN(n9750) );
  INV_X1 U4982 ( .A(n6865), .ZN(n10338) );
  CLKBUF_X2 U4985 ( .A(n5279), .Z(n4475) );
  CLKBUF_X2 U4986 ( .A(n6434), .Z(n4478) );
  NAND2_X1 U4987 ( .A1(n6217), .A2(n6216), .ZN(n9564) );
  AND3_X2 U4988 ( .A1(n6422), .A2(n6421), .A3(n6420), .ZN(n10171) );
  CLKBUF_X2 U4989 ( .A(n5055), .Z(n4951) );
  CLKBUF_X2 U4990 ( .A(n5598), .Z(n4481) );
  NAND2_X2 U4991 ( .A1(n5873), .A2(n5910), .ZN(n6522) );
  INV_X4 U4992 ( .A(n6557), .ZN(n6431) );
  INV_X1 U4993 ( .A(n6527), .ZN(n6213) );
  INV_X2 U4994 ( .A(n5247), .ZN(n5512) );
  CLKBUF_X2 U4995 ( .A(n5598), .Z(n4482) );
  INV_X1 U4996 ( .A(n6589), .ZN(n9035) );
  NOR2_X1 U4997 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5045) );
  INV_X1 U4998 ( .A(n5788), .ZN(n5782) );
  NOR2_X1 U4999 ( .A1(n7436), .A2(n5009), .ZN(n5008) );
  INV_X1 U5000 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5324) );
  INV_X1 U5001 ( .A(n8044), .ZN(n7946) );
  OR2_X1 U5002 ( .A1(n9472), .A2(n9527), .ZN(n6412) );
  INV_X1 U5003 ( .A(n9126), .ZN(n5222) );
  AOI21_X1 U5004 ( .B1(n8421), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8428), .ZN(
        n8067) );
  INV_X1 U5005 ( .A(n6506), .ZN(n7803) );
  NOR3_X1 U5006 ( .A1(n8515), .A2(n4740), .A3(n9037), .ZN(n8452) );
  INV_X1 U5007 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5479) );
  NAND2_X2 U5008 ( .A1(n6522), .A2(n6684), .ZN(n7945) );
  INV_X1 U5009 ( .A(n7947), .ZN(n8047) );
  NAND2_X1 U5010 ( .A1(n7767), .A2(n7766), .ZN(n9242) );
  XNOR2_X1 U5011 ( .A(n5217), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9122) );
  INV_X1 U5012 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U5013 ( .A1(n7696), .A2(n7695), .ZN(n9919) );
  CLKBUF_X2 U5014 ( .A(n6434), .Z(n4479) );
  NAND4_X1 U5015 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n10138)
         );
  NAND2_X1 U5016 ( .A1(n5867), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U5017 ( .A1(n5291), .A2(n5290), .ZN(n5293) );
  NAND4_X1 U5018 ( .A1(n5259), .A2(n5258), .A3(n5257), .A4(n5256), .ZN(n8382)
         );
  INV_X1 U5019 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U5020 ( .A1(n4711), .A2(n5195), .ZN(n9133) );
  INV_X1 U5021 ( .A(n6542), .ZN(n7802) );
  BUF_X1 U5022 ( .A(n6433), .Z(n4477) );
  NAND2_X2 U5023 ( .A1(n4861), .A2(n4860), .ZN(n8177) );
  AND2_X1 U5024 ( .A1(n5223), .A2(n5222), .ZN(n5608) );
  INV_X1 U5025 ( .A(n5608), .ZN(n4484) );
  NAND2_X1 U5026 ( .A1(n5942), .A2(n9964), .ZN(n6433) );
  AOI21_X2 U5027 ( .B1(n9618), .B2(n10135), .A(n9617), .ZN(n9852) );
  XNOR2_X2 U5028 ( .A(n5823), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6589) );
  OAI211_X2 U5029 ( .C1(n5329), .C2(n6416), .A(n5252), .B(n5251), .ZN(n6613)
         );
  XNOR2_X2 U5030 ( .A(n5868), .B(n4950), .ZN(n7613) );
  NAND2_X1 U5031 ( .A1(n8107), .A2(n5943), .ZN(n6434) );
  NOR2_X4 U5032 ( .A1(n5464), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5480) );
  OR2_X2 U5033 ( .A1(n5421), .A2(n4849), .ZN(n5464) );
  INV_X1 U5034 ( .A(n7945), .ZN(n4480) );
  NAND2_X1 U5035 ( .A1(n5223), .A2(n9126), .ZN(n5598) );
  OAI21_X1 U5036 ( .B1(n9532), .B2(n9531), .A(n9530), .ZN(n9542) );
  NOR2_X1 U5037 ( .A1(n8042), .A2(n4552), .ZN(n8065) );
  AND2_X1 U5038 ( .A1(n9040), .A2(n9039), .ZN(n4981) );
  OR2_X1 U5039 ( .A1(n8153), .A2(n8152), .ZN(n8154) );
  NAND2_X1 U5040 ( .A1(n9635), .A2(n9629), .ZN(n9640) );
  NAND2_X1 U5041 ( .A1(n8205), .A2(n8140), .ZN(n8307) );
  NAND2_X1 U5042 ( .A1(n9165), .A2(n9164), .ZN(n4908) );
  NAND2_X1 U5043 ( .A1(n4703), .A2(n4528), .ZN(n9165) );
  NAND2_X1 U5044 ( .A1(n9770), .A2(n9404), .ZN(n9758) );
  NAND2_X1 U5045 ( .A1(n7987), .A2(n9387), .ZN(n9806) );
  NAND2_X1 U5046 ( .A1(n7566), .A2(n4517), .ZN(n7724) );
  NAND2_X1 U5047 ( .A1(n7845), .A2(n7844), .ZN(n9889) );
  NAND2_X1 U5048 ( .A1(n5440), .A2(n5439), .ZN(n7581) );
  NAND2_X1 U5049 ( .A1(n7556), .A2(n7555), .ZN(n9928) );
  NAND2_X1 U5050 ( .A1(n5375), .A2(n5041), .ZN(n5102) );
  AND2_X1 U5051 ( .A1(n6780), .A2(n6779), .ZN(n7192) );
  INV_X1 U5052 ( .A(n10355), .ZN(n8289) );
  AND2_X2 U5053 ( .A1(n7025), .A2(n10150), .ZN(n10157) );
  AND2_X1 U5054 ( .A1(n6795), .A2(n6794), .ZN(n10190) );
  AND3_X1 U5055 ( .A1(n5313), .A2(n5312), .A3(n5311), .ZN(n10355) );
  AND3_X2 U5056 ( .A1(n6350), .A2(n6349), .A3(n6348), .ZN(n10223) );
  NAND4_X1 U5057 ( .A1(n6565), .A2(n6564), .A3(n6563), .A4(n6562), .ZN(n9559)
         );
  NAND2_X1 U5058 ( .A1(n5292), .A2(n5293), .ZN(n6540) );
  INV_X4 U5059 ( .A(n7945), .ZN(n7347) );
  NAND4_X1 U5060 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n8381)
         );
  NAND2_X4 U5061 ( .A1(n8107), .A2(n9964), .ZN(n6557) );
  INV_X1 U5062 ( .A(n5943), .ZN(n9964) );
  INV_X2 U5063 ( .A(n5329), .ZN(n4990) );
  OR2_X1 U5064 ( .A1(n6573), .A2(n6597), .ZN(n6115) );
  NAND2_X1 U5065 ( .A1(n5884), .A2(n5883), .ZN(n9472) );
  NAND2_X2 U5066 ( .A1(n5662), .A2(n8086), .ZN(n6576) );
  CLKBUF_X1 U5067 ( .A(n8505), .Z(n4573) );
  CLKBUF_X3 U5068 ( .A(n5611), .Z(n4483) );
  INV_X1 U5069 ( .A(n6600), .ZN(n5662) );
  NAND2_X1 U5070 ( .A1(n4872), .A2(n4871), .ZN(n5661) );
  NAND2_X1 U5071 ( .A1(n5221), .A2(n5220), .ZN(n9126) );
  MUX2_X1 U5072 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5219), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5221) );
  NAND2_X1 U5073 ( .A1(n5220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U5074 ( .A1(n5195), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4646) );
  OR2_X1 U5075 ( .A1(n5639), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5830) );
  INV_X2 U5076 ( .A(n9961), .ZN(n9971) );
  INV_X1 U5077 ( .A(n4948), .ZN(n4755) );
  AND2_X1 U5078 ( .A1(n4580), .A2(n5180), .ZN(n4579) );
  INV_X1 U5079 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5180) );
  INV_X1 U5080 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5831) );
  INV_X1 U5081 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5827) );
  INV_X1 U5082 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6479) );
  INV_X1 U5083 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4580) );
  NOR2_X1 U5084 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5892) );
  INV_X1 U5085 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5181) );
  INV_X2 U5086 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5087 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5856) );
  NOR2_X1 U5088 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5857) );
  NOR2_X1 U5089 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5858) );
  INV_X4 U5090 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OAI21_X2 U5091 ( .B1(n7512), .B2(n4841), .A(n4838), .ZN(n7664) );
  NAND2_X1 U5092 ( .A1(n9122), .A2(n9126), .ZN(n5611) );
  INV_X2 U5093 ( .A(n4484), .ZN(n4485) );
  XNOR2_X2 U5094 ( .A(n5888), .B(n5887), .ZN(n5956) );
  OR2_X1 U5095 ( .A1(n6576), .A2(n10326), .ZN(n4486) );
  NAND2_X2 U5096 ( .A1(n5565), .A2(n5564), .ZN(n9071) );
  AOI21_X1 U5097 ( .B1(n8351), .B2(n8168), .A(n4889), .ZN(n4888) );
  INV_X1 U5098 ( .A(n8209), .ZN(n4889) );
  NAND2_X1 U5099 ( .A1(n4845), .A2(n4844), .ZN(n8153) );
  AOI21_X1 U5100 ( .B1(n4846), .B2(n4848), .A(n4515), .ZN(n4844) );
  NAND2_X1 U5101 ( .A1(n8156), .A2(n6578), .ZN(n6117) );
  AND2_X1 U5102 ( .A1(n4955), .A2(n8537), .ZN(n4954) );
  OR2_X1 U5103 ( .A1(n9854), .A2(n9654), .ZN(n9444) );
  NAND2_X1 U5104 ( .A1(n4803), .A2(n4801), .ZN(n5593) );
  AOI21_X1 U5105 ( .B1(n4550), .B2(n4808), .A(n4802), .ZN(n4801) );
  INV_X1 U5106 ( .A(n5167), .ZN(n4802) );
  NAND2_X1 U5107 ( .A1(n5420), .A2(n5042), .ZN(n4727) );
  NAND2_X1 U5108 ( .A1(n8177), .A2(n8157), .ZN(n4869) );
  NAND2_X1 U5109 ( .A1(n4584), .A2(n4586), .ZN(n4581) );
  NAND2_X1 U5110 ( .A1(n4584), .A2(n10266), .ZN(n4582) );
  NAND2_X1 U5111 ( .A1(n9664), .A2(n4779), .ZN(n9645) );
  OR2_X1 U5112 ( .A1(n9667), .A2(n9547), .ZN(n4779) );
  NAND2_X1 U5113 ( .A1(n9958), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5939) );
  OR2_X1 U5114 ( .A1(n5940), .A2(n6035), .ZN(n5941) );
  NAND2_X1 U5115 ( .A1(n5019), .A2(n4496), .ZN(n5018) );
  INV_X1 U5116 ( .A(n5021), .ZN(n5019) );
  AOI21_X1 U5117 ( .B1(n4490), .B2(n5022), .A(n4566), .ZN(n5021) );
  NAND2_X1 U5118 ( .A1(n8381), .A2(n10344), .ZN(n5686) );
  NOR2_X1 U5119 ( .A1(n5162), .A2(n4810), .ZN(n4809) );
  INV_X1 U5120 ( .A(n5153), .ZN(n4642) );
  AOI21_X1 U5121 ( .B1(n4888), .B2(n4886), .A(n4536), .ZN(n4885) );
  INV_X1 U5122 ( .A(n8168), .ZN(n4886) );
  INV_X1 U5123 ( .A(n9122), .ZN(n5223) );
  NOR2_X1 U5124 ( .A1(n8458), .A2(n4523), .ZN(n8124) );
  NOR2_X1 U5125 ( .A1(n9049), .A2(n9056), .ZN(n4741) );
  NOR2_X1 U5126 ( .A1(n8482), .A2(n5032), .ZN(n5031) );
  INV_X1 U5127 ( .A(n5776), .ZN(n5032) );
  OR2_X1 U5128 ( .A1(n9066), .A2(n8297), .ZN(n5767) );
  OR2_X1 U5129 ( .A1(n9088), .A2(n8243), .ZN(n5748) );
  OR2_X1 U5130 ( .A1(n7607), .A2(n8278), .ZN(n5729) );
  INV_X1 U5131 ( .A(n5723), .ZN(n5009) );
  AOI21_X1 U5132 ( .B1(n10310), .B2(n10323), .A(n10324), .ZN(n9028) );
  NOR2_X1 U5133 ( .A1(n5189), .A2(n5188), .ZN(n5190) );
  INV_X1 U5134 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5187) );
  INV_X1 U5135 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U5136 ( .A1(n5824), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5825) );
  NOR2_X1 U5137 ( .A1(n5027), .A2(n5026), .ZN(n5025) );
  INV_X1 U5138 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5048) );
  INV_X1 U5139 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4830) );
  AND2_X1 U5140 ( .A1(n5376), .A2(n5044), .ZN(n5047) );
  INV_X1 U5141 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U5142 ( .A1(n9293), .A2(n9292), .ZN(n9463) );
  INV_X1 U5143 ( .A(n4760), .ZN(n4759) );
  OAI21_X1 U5144 ( .B1(n9781), .B2(n4761), .A(n7973), .ZN(n4760) );
  OR2_X1 U5145 ( .A1(n7319), .A2(n4794), .ZN(n4793) );
  INV_X1 U5146 ( .A(n7288), .ZN(n4794) );
  NAND2_X1 U5147 ( .A1(n9473), .A2(n9690), .ZN(n4909) );
  OR2_X1 U5148 ( .A1(n9844), .A2(n9616), .ZN(n9454) );
  NAND2_X1 U5149 ( .A1(n4812), .A2(n4811), .ZN(n5633) );
  AOI21_X1 U5150 ( .B1(n4814), .B2(n4816), .A(n4568), .ZN(n4811) );
  NAND2_X1 U5151 ( .A1(n4639), .A2(n5153), .ZN(n5563) );
  NAND2_X1 U5152 ( .A1(n5146), .A2(n5145), .ZN(n5537) );
  OAI21_X1 U5153 ( .B1(n5511), .B2(n5510), .A(n5141), .ZN(n5525) );
  AND2_X1 U5154 ( .A1(n5129), .A2(n5128), .ZN(n5462) );
  INV_X1 U5155 ( .A(n4632), .ZN(n4631) );
  OAI21_X1 U5156 ( .B1(n4635), .B2(n4503), .A(n5124), .ZN(n4632) );
  INV_X1 U5157 ( .A(n4617), .ZN(n4616) );
  OAI21_X1 U5158 ( .B1(n4618), .B2(n4505), .A(n5110), .ZN(n4617) );
  NAND2_X1 U5159 ( .A1(n5097), .A2(n5096), .ZN(n5375) );
  OAI21_X1 U5160 ( .B1(n6417), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n5052), .ZN(
        n5053) );
  NAND2_X1 U5161 ( .A1(n6417), .A2(n5051), .ZN(n5052) );
  INV_X1 U5162 ( .A(n4888), .ZN(n4887) );
  INV_X1 U5163 ( .A(n4885), .ZN(n4882) );
  NAND2_X1 U5164 ( .A1(n6118), .A2(n4837), .ZN(n4832) );
  INV_X1 U5165 ( .A(n8586), .ZN(n8243) );
  NAND2_X1 U5166 ( .A1(n4868), .A2(n4554), .ZN(n4867) );
  INV_X1 U5167 ( .A(n8293), .ZN(n4868) );
  NAND2_X1 U5168 ( .A1(n5830), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5823) );
  AND2_X1 U5169 ( .A1(n8397), .A2(n6340), .ZN(n6342) );
  OR2_X1 U5170 ( .A1(n8222), .A2(n5622), .ZN(n5229) );
  NAND2_X1 U5171 ( .A1(n4593), .A2(n4592), .ZN(n8511) );
  AOI21_X1 U5172 ( .B1(n4594), .B2(n4495), .A(n8524), .ZN(n4592) );
  NOR2_X1 U5173 ( .A1(n9066), .A2(n8549), .ZN(n8531) );
  XNOR2_X1 U5174 ( .A(n9071), .B(n8572), .ZN(n8556) );
  AND2_X1 U5175 ( .A1(n4595), .A2(n4597), .ZN(n8562) );
  NAND2_X1 U5176 ( .A1(n8579), .A2(n8113), .ZN(n4595) );
  AND2_X1 U5177 ( .A1(n8596), .A2(n5748), .ZN(n8585) );
  OR2_X1 U5178 ( .A1(n9098), .A2(n8111), .ZN(n5743) );
  NOR2_X1 U5179 ( .A1(n4603), .A2(n8112), .ZN(n4602) );
  INV_X1 U5180 ( .A(n4605), .ZN(n4603) );
  OR2_X1 U5181 ( .A1(n8110), .A2(n8647), .ZN(n4605) );
  NAND2_X1 U5182 ( .A1(n5409), .A2(n5408), .ZN(n7393) );
  NAND2_X1 U5183 ( .A1(n10239), .A2(n4971), .ZN(n6995) );
  AND2_X1 U5184 ( .A1(n6944), .A2(n6943), .ZN(n4971) );
  AND2_X1 U5185 ( .A1(n5247), .A2(n5055), .ZN(n5279) );
  NAND2_X1 U5186 ( .A1(n6937), .A2(n6936), .ZN(n10266) );
  NAND2_X1 U5187 ( .A1(n8382), .A2(n10261), .ZN(n4675) );
  NAND2_X2 U5188 ( .A1(n9133), .A2(n5844), .ZN(n5247) );
  NAND4_X1 U5189 ( .A1(n5185), .A2(n5025), .A3(n5190), .A4(n5047), .ZN(n5191)
         );
  XNOR2_X1 U5190 ( .A(n5660), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U5191 ( .A1(n4873), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5660) );
  AND2_X2 U5192 ( .A1(n5025), .A2(n5047), .ZN(n5394) );
  NAND2_X1 U5193 ( .A1(n5263), .A2(n5324), .ZN(n5024) );
  AND2_X1 U5194 ( .A1(n9192), .A2(n9179), .ZN(n4702) );
  NAND2_X1 U5195 ( .A1(n4533), .A2(n4902), .ZN(n9157) );
  NAND3_X1 U5196 ( .A1(n4902), .A2(n4704), .A3(n9230), .ZN(n4703) );
  AND2_X1 U5197 ( .A1(n4901), .A2(n9210), .ZN(n4704) );
  OR2_X1 U5198 ( .A1(n7921), .A2(n8938), .ZN(n7951) );
  NAND2_X1 U5199 ( .A1(n4539), .A2(n4489), .ZN(n4624) );
  NAND2_X1 U5200 ( .A1(n4489), .A2(n4626), .ZN(n4625) );
  INV_X1 U5201 ( .A(n4563), .ZN(n4626) );
  NOR2_X1 U5203 ( .A1(n7983), .A2(n7982), .ZN(n9664) );
  NOR2_X1 U5204 ( .A1(n9662), .A2(n9668), .ZN(n7982) );
  AND2_X1 U5205 ( .A1(n4511), .A2(n7693), .ZN(n4776) );
  NAND2_X1 U5206 ( .A1(n4775), .A2(n4511), .ZN(n4774) );
  INV_X1 U5207 ( .A(n4777), .ZN(n4775) );
  AOI21_X1 U5208 ( .B1(n4494), .B2(n7693), .A(n4524), .ZN(n4777) );
  NAND2_X1 U5209 ( .A1(n4764), .A2(n4762), .ZN(n7094) );
  AOI21_X1 U5210 ( .B1(n9304), .B2(n7009), .A(n4763), .ZN(n4762) );
  INV_X1 U5211 ( .A(n9306), .ZN(n4763) );
  NAND2_X1 U5212 ( .A1(n6542), .A2(n5055), .ZN(n6792) );
  NOR2_X1 U5213 ( .A1(n7674), .A2(n7613), .ZN(n5873) );
  AND2_X1 U5214 ( .A1(n5864), .A2(n4911), .ZN(n4910) );
  INV_X1 U5215 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5876) );
  XNOR2_X1 U5216 ( .A(n5563), .B(n5562), .ZN(n7880) );
  XNOR2_X1 U5217 ( .A(n6184), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U5218 ( .A1(n5865), .A2(n5864), .ZN(n6183) );
  INV_X1 U5219 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U5220 ( .A1(n5246), .A2(n5059), .ZN(n5060) );
  AND2_X1 U5221 ( .A1(n8154), .A2(n4564), .ZN(n4865) );
  AND2_X1 U5222 ( .A1(n8318), .A2(n8382), .ZN(n4676) );
  OAI21_X1 U5223 ( .B1(n7635), .B2(n7634), .A(n7640), .ZN(n7760) );
  INV_X1 U5224 ( .A(n9649), .ZN(n9859) );
  NAND2_X1 U5225 ( .A1(n5685), .A2(n5689), .ZN(n4664) );
  AND2_X1 U5226 ( .A1(n7439), .A2(n5724), .ZN(n4650) );
  NAND2_X1 U5227 ( .A1(n7583), .A2(n5728), .ZN(n4649) );
  AOI21_X1 U5228 ( .B1(n4656), .B2(n4493), .A(n4654), .ZN(n4653) );
  NAND2_X1 U5229 ( .A1(n5030), .A2(n5780), .ZN(n4654) );
  INV_X1 U5230 ( .A(n5774), .ZN(n4657) );
  NAND2_X1 U5231 ( .A1(n4493), .A2(n4529), .ZN(n4655) );
  INV_X1 U5232 ( .A(n4916), .ZN(n4914) );
  INV_X1 U5233 ( .A(n5583), .ZN(n4804) );
  AOI21_X1 U5234 ( .B1(n4535), .B2(n5018), .A(n4500), .ZN(n5015) );
  NOR2_X1 U5235 ( .A1(n5018), .A2(n4491), .ZN(n5017) );
  NOR2_X1 U5236 ( .A1(n9076), .A2(n4730), .ZN(n4729) );
  INV_X1 U5237 ( .A(n4731), .ZN(n4730) );
  INV_X1 U5238 ( .A(n4504), .ZN(n4600) );
  OR3_X1 U5239 ( .A1(n5454), .A2(n5453), .A3(n5452), .ZN(n5468) );
  NAND2_X1 U5240 ( .A1(n10021), .A2(n8278), .ZN(n4968) );
  NOR2_X1 U5241 ( .A1(n5012), .A2(n4985), .ZN(n4984) );
  INV_X1 U5242 ( .A(n7394), .ZN(n4985) );
  INV_X1 U5243 ( .A(n7081), .ZN(n4997) );
  INV_X1 U5244 ( .A(n5798), .ZN(n4998) );
  INV_X1 U5245 ( .A(n5693), .ZN(n5003) );
  OAI21_X1 U5246 ( .B1(n5800), .B2(n5003), .A(n5695), .ZN(n5002) );
  INV_X1 U5247 ( .A(SI_13_), .ZN(n8915) );
  NAND2_X1 U5248 ( .A1(n10255), .A2(n10256), .ZN(n5332) );
  AND2_X1 U5249 ( .A1(n5693), .A2(n5689), .ZN(n5800) );
  NAND2_X1 U5250 ( .A1(n6578), .A2(n10333), .ZN(n5795) );
  OR2_X1 U5251 ( .A1(n9063), .A2(n8539), .ZN(n5773) );
  AND2_X1 U5252 ( .A1(n5775), .A2(n5776), .ZN(n8495) );
  NAND2_X1 U5253 ( .A1(n5279), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4666) );
  AOI21_X1 U5254 ( .B1(n4875), .B2(P2_IR_REG_31__SCAN_IN), .A(
        P2_IR_REG_19__SCAN_IN), .ZN(n4874) );
  INV_X1 U5255 ( .A(n4512), .ZN(n4875) );
  NAND2_X1 U5256 ( .A1(n4537), .A2(n4850), .ZN(n4849) );
  AND2_X1 U5257 ( .A1(n5360), .A2(n5043), .ZN(n5376) );
  INV_X1 U5258 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5043) );
  INV_X1 U5259 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5851) );
  OR2_X1 U5260 ( .A1(n9849), .A2(n9638), .ZN(n9450) );
  OR2_X1 U5261 ( .A1(n9859), .A2(n9671), .ZN(n9440) );
  OR2_X1 U5262 ( .A1(n9667), .A2(n9687), .ZN(n9434) );
  AOI21_X1 U5263 ( .B1(n9511), .B2(n4917), .A(n9427), .ZN(n4916) );
  NAND2_X1 U5264 ( .A1(n4615), .A2(n4518), .ZN(n9424) );
  INV_X1 U5265 ( .A(n7900), .ZN(n4614) );
  AOI21_X1 U5266 ( .B1(n4942), .B2(n9757), .A(n4941), .ZN(n4940) );
  INV_X1 U5267 ( .A(n4768), .ZN(n4767) );
  OAI21_X1 U5268 ( .B1(n7975), .B2(n4769), .A(n7978), .ZN(n4768) );
  INV_X1 U5269 ( .A(n7977), .ZN(n4769) );
  AND2_X1 U5270 ( .A1(n9751), .A2(n9736), .ZN(n9718) );
  OR2_X1 U5271 ( .A1(n9883), .A2(n9709), .ZN(n9418) );
  OR2_X1 U5272 ( .A1(n9928), .A2(n9819), .ZN(n9375) );
  NOR2_X1 U5273 ( .A1(n4747), .A2(n7092), .ZN(n4745) );
  NAND2_X1 U5274 ( .A1(n10196), .A2(n7192), .ZN(n4747) );
  NOR2_X1 U5275 ( .A1(n4927), .A2(n4925), .ZN(n4924) );
  INV_X1 U5276 ( .A(n9491), .ZN(n4925) );
  OR2_X1 U5277 ( .A1(n9896), .A2(n9159), .ZN(n9415) );
  AND2_X1 U5278 ( .A1(n7427), .A2(n10053), .ZN(n7497) );
  OAI21_X1 U5279 ( .B1(n5633), .B2(n5632), .A(n5631), .ZN(n5649) );
  AND2_X1 U5280 ( .A1(n5178), .A2(n5177), .ZN(n5603) );
  AND2_X1 U5281 ( .A1(n5172), .A2(n5171), .ZN(n5592) );
  NOR2_X1 U5282 ( .A1(n4642), .A2(n4810), .ZN(n4638) );
  INV_X1 U5283 ( .A(n4641), .ZN(n4640) );
  OAI21_X1 U5284 ( .B1(n4643), .B2(n4642), .A(n5562), .ZN(n4641) );
  OR2_X1 U5285 ( .A1(n5537), .A2(n4828), .ZN(n4645) );
  INV_X1 U5286 ( .A(n6185), .ZN(n5865) );
  AND2_X1 U5287 ( .A1(n5145), .A2(n5144), .ZN(n5524) );
  AOI21_X1 U5288 ( .B1(n4716), .B2(n4718), .A(n4559), .ZN(n4714) );
  NOR2_X1 U5289 ( .A1(n5134), .A2(n4720), .ZN(n4719) );
  INV_X1 U5290 ( .A(n5129), .ZN(n4720) );
  NAND2_X1 U5291 ( .A1(n4630), .A2(n4628), .ZN(n4827) );
  AOI21_X1 U5292 ( .B1(n4631), .B2(n4503), .A(n4629), .ZN(n4628) );
  NAND2_X1 U5293 ( .A1(n4727), .A2(n4631), .ZN(n4630) );
  INV_X1 U5294 ( .A(n5462), .ZN(n4629) );
  AOI21_X1 U5295 ( .B1(n4820), .B2(n4987), .A(n4819), .ZN(n4818) );
  INV_X1 U5296 ( .A(n5082), .ZN(n4819) );
  AND2_X1 U5297 ( .A1(n5082), .A2(n5081), .ZN(n5328) );
  AND2_X1 U5298 ( .A1(n5077), .A2(n5076), .ZN(n5304) );
  AOI21_X1 U5299 ( .B1(n4885), .B2(n4887), .A(n8221), .ZN(n4884) );
  AND2_X1 U5300 ( .A1(n8241), .A2(n4847), .ZN(n4846) );
  NAND2_X1 U5301 ( .A1(n8308), .A2(n8147), .ZN(n4847) );
  INV_X1 U5302 ( .A(n8147), .ZN(n4848) );
  NAND2_X1 U5303 ( .A1(n4853), .A2(n4851), .ZN(n6743) );
  NOR2_X1 U5304 ( .A1(n6740), .A2(n4852), .ZN(n4851) );
  INV_X1 U5305 ( .A(n6304), .ZN(n4852) );
  NAND2_X1 U5306 ( .A1(n5207), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5529) );
  OR2_X1 U5307 ( .A1(n5529), .A2(n5528), .ZN(n5541) );
  NAND2_X1 U5308 ( .A1(n8146), .A2(n8145), .ZN(n8305) );
  INV_X1 U5309 ( .A(n6120), .ZN(n4831) );
  OR2_X1 U5310 ( .A1(n6144), .A2(n10309), .ZN(n6143) );
  AND3_X1 U5311 ( .A1(n5581), .A2(n5580), .A3(n5579), .ZN(n8297) );
  AND2_X1 U5312 ( .A1(n6488), .A2(n6487), .ZN(n8415) );
  AND2_X1 U5313 ( .A1(n5628), .A2(n5627), .ZN(n8460) );
  NAND2_X1 U5314 ( .A1(n8494), .A2(n5031), .ZN(n5033) );
  OAI21_X1 U5315 ( .B1(n8523), .B2(n4679), .A(n4532), .ZN(n8458) );
  INV_X1 U5316 ( .A(n5029), .ZN(n4679) );
  OR2_X1 U5317 ( .A1(n8464), .A2(n5778), .ZN(n5028) );
  OR2_X1 U5318 ( .A1(n9056), .A2(n8368), .ZN(n8115) );
  NAND2_X1 U5319 ( .A1(n5778), .A2(n5779), .ZN(n8482) );
  AND2_X1 U5320 ( .A1(n5607), .A2(n5597), .ZN(n8502) );
  AOI21_X1 U5321 ( .B1(n4954), .B2(n4590), .A(n4589), .ZN(n4594) );
  NOR2_X1 U5322 ( .A1(n4596), .A2(n8113), .ZN(n4590) );
  NAND2_X1 U5323 ( .A1(n4953), .A2(n4959), .ZN(n4589) );
  AOI21_X1 U5324 ( .B1(n4956), .B2(n8569), .A(n4534), .ZN(n4955) );
  INV_X1 U5325 ( .A(n8556), .ZN(n8547) );
  NAND2_X1 U5326 ( .A1(n8568), .A2(n5037), .ZN(n8555) );
  AND2_X1 U5327 ( .A1(n8556), .A2(n5757), .ZN(n5037) );
  OR2_X1 U5328 ( .A1(n9076), .A2(n8179), .ZN(n5757) );
  NAND2_X1 U5329 ( .A1(n8584), .A2(n5038), .ZN(n8568) );
  AND2_X1 U5330 ( .A1(n8569), .A2(n5750), .ZN(n5038) );
  NAND2_X1 U5331 ( .A1(n8585), .A2(n5549), .ZN(n8584) );
  NAND2_X1 U5332 ( .A1(n9086), .A2(n4551), .ZN(n8579) );
  INV_X1 U5333 ( .A(n8571), .ZN(n8593) );
  INV_X1 U5334 ( .A(n4690), .ZN(n4689) );
  AND2_X1 U5335 ( .A1(n4687), .A2(n5023), .ZN(n4686) );
  NOR2_X1 U5336 ( .A1(n8598), .A2(n4742), .ZN(n5023) );
  NAND2_X1 U5337 ( .A1(n5748), .A2(n5751), .ZN(n8598) );
  NAND2_X1 U5338 ( .A1(n8629), .A2(n4690), .ZN(n8615) );
  NAND2_X1 U5339 ( .A1(n8631), .A2(n8630), .ZN(n8629) );
  NAND2_X1 U5340 ( .A1(n5485), .A2(n5484), .ZN(n8110) );
  OAI21_X1 U5341 ( .B1(n7580), .B2(n4961), .A(n4960), .ZN(n7679) );
  NAND2_X1 U5342 ( .A1(n4965), .A2(n4967), .ZN(n4961) );
  NAND2_X1 U5343 ( .A1(n4538), .A2(n4967), .ZN(n4960) );
  NAND2_X1 U5344 ( .A1(n10015), .A2(n8370), .ZN(n4967) );
  NAND2_X1 U5345 ( .A1(n7679), .A2(n7678), .ZN(n8109) );
  AND2_X1 U5346 ( .A1(n4968), .A2(n4969), .ZN(n4966) );
  OAI21_X1 U5347 ( .B1(n7398), .B2(n7399), .A(n5008), .ZN(n5007) );
  NAND2_X1 U5348 ( .A1(n5012), .A2(n5726), .ZN(n5006) );
  NAND2_X1 U5349 ( .A1(n5005), .A2(n5726), .ZN(n5004) );
  INV_X1 U5350 ( .A(n5008), .ZN(n5005) );
  NAND2_X1 U5351 ( .A1(n5011), .A2(n5012), .ZN(n5010) );
  INV_X1 U5352 ( .A(n7398), .ZN(n5011) );
  OAI21_X1 U5353 ( .B1(n7079), .B2(n4611), .A(n4609), .ZN(n7437) );
  NAND2_X1 U5354 ( .A1(n4983), .A2(n7222), .ZN(n4611) );
  AND2_X1 U5355 ( .A1(n4610), .A2(n4982), .ZN(n4609) );
  NAND2_X1 U5356 ( .A1(n4983), .A2(n4519), .ZN(n4610) );
  NOR2_X2 U5357 ( .A1(n4726), .A2(n7435), .ZN(n7587) );
  NOR2_X1 U5358 ( .A1(n7227), .A2(n8189), .ZN(n4725) );
  OR2_X1 U5359 ( .A1(n5366), .A2(n5201), .ZN(n5384) );
  NAND2_X1 U5360 ( .A1(n6942), .A2(n6941), .ZN(n10239) );
  INV_X1 U5361 ( .A(n10236), .ZN(n6941) );
  INV_X1 U5362 ( .A(n10367), .ZN(n9012) );
  NAND2_X1 U5363 ( .A1(n5332), .A2(n5800), .ZN(n10258) );
  NAND2_X1 U5364 ( .A1(n6852), .A2(n6851), .ZN(n6935) );
  INV_X1 U5365 ( .A(n8381), .ZN(n10287) );
  NAND2_X1 U5366 ( .A1(n10351), .A2(n8380), .ZN(n10282) );
  NAND2_X1 U5367 ( .A1(n6586), .A2(n6865), .ZN(n6588) );
  INV_X1 U5368 ( .A(n10284), .ZN(n10261) );
  INV_X1 U5369 ( .A(n10286), .ZN(n10259) );
  NAND2_X1 U5370 ( .A1(n5621), .A2(n5620), .ZN(n9037) );
  NAND2_X1 U5371 ( .A1(n5197), .A2(n5196), .ZN(n9043) );
  NAND2_X1 U5372 ( .A1(n5575), .A2(n5574), .ZN(n9066) );
  NAND2_X1 U5373 ( .A1(n5501), .A2(n5500), .ZN(n9098) );
  NAND2_X1 U5374 ( .A1(n5279), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U5375 ( .A1(n5512), .A2(n6064), .ZN(n4606) );
  OR2_X1 U5376 ( .A1(n6505), .A2(n5329), .ZN(n4607) );
  AND2_X1 U5377 ( .A1(n6125), .A2(n6123), .ZN(n10310) );
  OR2_X1 U5378 ( .A1(n5825), .A2(n5828), .ZN(n5826) );
  AND2_X1 U5379 ( .A1(n5394), .A2(n4541), .ZN(n4691) );
  AND2_X1 U5380 ( .A1(n5185), .A2(n5190), .ZN(n4692) );
  NAND2_X1 U5381 ( .A1(n5825), .A2(n5828), .ZN(n5839) );
  NAND2_X1 U5382 ( .A1(n5480), .A2(n5181), .ZN(n5498) );
  INV_X1 U5383 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5348) );
  NOR2_X1 U5384 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5263) );
  NAND2_X1 U5385 ( .A1(n7935), .A2(n7936), .ZN(n4898) );
  INV_X1 U5386 ( .A(n4906), .ZN(n4905) );
  OAI21_X1 U5387 ( .B1(n7031), .B2(n4907), .A(n6904), .ZN(n4906) );
  AND2_X1 U5388 ( .A1(n6415), .A2(n6414), .ZN(n6426) );
  OR2_X1 U5389 ( .A1(n6413), .A2(n8047), .ZN(n6415) );
  NAND2_X1 U5390 ( .A1(n9192), .A2(n4701), .ZN(n4700) );
  INV_X1 U5391 ( .A(n7768), .ZN(n4701) );
  NAND2_X1 U5392 ( .A1(n9210), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U5393 ( .A1(n6625), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U5394 ( .A1(n7800), .A2(n7799), .ZN(n9230) );
  NOR2_X1 U5395 ( .A1(n8040), .A2(n4896), .ZN(n4895) );
  INV_X1 U5396 ( .A(n4900), .ZN(n4896) );
  OR2_X1 U5397 ( .A1(n9171), .A2(n9172), .ZN(n4897) );
  NAND2_X1 U5398 ( .A1(n9328), .A2(n9472), .ZN(n9468) );
  OR3_X1 U5399 ( .A1(n9474), .A2(n9524), .A3(n9327), .ZN(n9328) );
  NAND2_X1 U5400 ( .A1(n8093), .A2(n5039), .ZN(n9293) );
  INV_X1 U5401 ( .A(n4921), .ZN(n4920) );
  NOR2_X1 U5402 ( .A1(n9613), .A2(n4922), .ZN(n4921) );
  INV_X1 U5403 ( .A(n9444), .ZN(n4922) );
  AND2_X1 U5404 ( .A1(n7951), .A2(n7732), .ZN(n9647) );
  NAND2_X1 U5405 ( .A1(n4620), .A2(n4619), .ZN(n9662) );
  INV_X1 U5406 ( .A(n7981), .ZN(n4619) );
  INV_X1 U5407 ( .A(n9692), .ZN(n4620) );
  OR2_X1 U5408 ( .A1(n9878), .A2(n9688), .ZN(n9684) );
  NAND2_X1 U5409 ( .A1(n7899), .A2(n6907), .ZN(n4615) );
  NOR2_X1 U5410 ( .A1(n9896), .A2(n9764), .ZN(n9751) );
  AOI21_X1 U5411 ( .B1(n4759), .B2(n4761), .A(n4556), .ZN(n4757) );
  OR2_X1 U5412 ( .A1(n9900), .A2(n9785), .ZN(n9764) );
  AND2_X1 U5413 ( .A1(n9400), .A2(n9404), .ZN(n9772) );
  INV_X1 U5414 ( .A(n9260), .ZN(n4935) );
  NAND2_X1 U5415 ( .A1(n4938), .A2(n4937), .ZN(n4936) );
  INV_X1 U5416 ( .A(n9806), .ZN(n4938) );
  OR2_X1 U5417 ( .A1(n7570), .A2(n7569), .ZN(n7702) );
  NOR2_X1 U5418 ( .A1(n9916), .A2(n4750), .ZN(n4749) );
  OAI21_X1 U5419 ( .B1(n7692), .B2(n4773), .A(n4497), .ZN(n7968) );
  INV_X1 U5420 ( .A(n4774), .ZN(n4773) );
  NAND2_X1 U5421 ( .A1(n4772), .A2(n4774), .ZN(n4771) );
  OR2_X1 U5422 ( .A1(n6922), .A2(n7270), .ZN(n7272) );
  INV_X1 U5423 ( .A(n4792), .ZN(n4791) );
  OAI22_X1 U5424 ( .A1(n7095), .A2(n4793), .B1(n9556), .B2(n10203), .ZN(n4792)
         );
  INV_X1 U5425 ( .A(n7096), .ZN(n4795) );
  OR2_X1 U5426 ( .A1(n7287), .A2(n7291), .ZN(n9351) );
  AND2_X1 U5427 ( .A1(n6969), .A2(n6883), .ZN(n4796) );
  OR2_X1 U5428 ( .A1(n6973), .A2(n9304), .ZN(n7010) );
  AND2_X1 U5429 ( .A1(n7015), .A2(n7016), .ZN(n9303) );
  NAND2_X1 U5430 ( .A1(n6703), .A2(n9298), .ZN(n6884) );
  INV_X1 U5431 ( .A(n10140), .ZN(n9816) );
  INV_X1 U5432 ( .A(n10135), .ZN(n9807) );
  AND2_X1 U5433 ( .A1(n6671), .A2(n9467), .ZN(n10137) );
  NAND2_X1 U5434 ( .A1(n4623), .A2(n4622), .ZN(n9611) );
  AOI21_X1 U5435 ( .B1(n4624), .B2(n4625), .A(n9325), .ZN(n4622) );
  NAND2_X1 U5436 ( .A1(n7985), .A2(n7984), .ZN(n9844) );
  AND3_X1 U5437 ( .A1(n6545), .A2(n6544), .A3(n6543), .ZN(n10182) );
  AND2_X1 U5438 ( .A1(n4948), .A2(n4800), .ZN(n4799) );
  NOR2_X1 U5439 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4800) );
  XNOR2_X1 U5440 ( .A(n5649), .B(n5648), .ZN(n5647) );
  AND2_X1 U5441 ( .A1(n4513), .A2(n4949), .ZN(n4948) );
  AND2_X1 U5442 ( .A1(n5866), .A2(n5886), .ZN(n4949) );
  NOR2_X1 U5443 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5886) );
  XNOR2_X1 U5444 ( .A(n5872), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U5445 ( .A1(n4805), .A2(n4806), .ZN(n5584) );
  OR2_X1 U5446 ( .A1(n5563), .A2(n4808), .ZN(n4805) );
  XNOR2_X1 U5447 ( .A(n5877), .B(n5876), .ZN(n7451) );
  XNOR2_X1 U5448 ( .A(n5880), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9473) );
  OAI21_X1 U5449 ( .B1(n4727), .B2(n4503), .A(n4631), .ZN(n5463) );
  NAND2_X1 U5450 ( .A1(n4634), .A2(n5118), .ZN(n5447) );
  NAND2_X1 U5451 ( .A1(n5102), .A2(n4618), .ZN(n5404) );
  NAND2_X1 U5452 ( .A1(n5102), .A2(n5101), .ZN(n5392) );
  INV_X1 U5453 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5931) );
  NOR2_X1 U5454 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5848) );
  INV_X1 U5455 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U5456 ( .A1(n5061), .A2(n5060), .ZN(n5261) );
  INV_X1 U5457 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5049) );
  NAND2_X1 U5458 ( .A1(n5606), .A2(n5605), .ZN(n9049) );
  NAND2_X1 U5459 ( .A1(n4859), .A2(n4858), .ZN(n4857) );
  INV_X1 U5460 ( .A(n6284), .ZN(n4859) );
  INV_X1 U5461 ( .A(n6283), .ZN(n4858) );
  NAND2_X1 U5462 ( .A1(n8327), .A2(n4572), .ZN(n8205) );
  AND2_X1 U5463 ( .A1(n8196), .A2(n8136), .ZN(n4572) );
  NOR2_X1 U5464 ( .A1(n4882), .A2(n4890), .ZN(n4878) );
  NAND2_X1 U5465 ( .A1(n4832), .A2(n6148), .ZN(n6121) );
  NAND2_X1 U5466 ( .A1(n5539), .A2(n5538), .ZN(n9081) );
  INV_X1 U5467 ( .A(n4842), .ZN(n4841) );
  AOI21_X1 U5468 ( .B1(n4842), .B2(n4840), .A(n4839), .ZN(n4838) );
  NOR2_X1 U5469 ( .A1(n7657), .A2(n4843), .ZN(n4842) );
  INV_X1 U5470 ( .A(n8318), .ZN(n8357) );
  AND2_X1 U5471 ( .A1(n8287), .A2(n10259), .ZN(n8346) );
  NAND2_X1 U5472 ( .A1(n4672), .A2(n4670), .ZN(n4669) );
  NAND2_X1 U5473 ( .A1(n5822), .A2(n5821), .ZN(n4672) );
  NAND2_X1 U5474 ( .A1(n5819), .A2(n6576), .ZN(n4671) );
  XNOR2_X1 U5475 ( .A(n4824), .B(n4573), .ZN(n5816) );
  INV_X1 U5476 ( .A(n8297), .ZN(n8558) );
  OR2_X1 U5477 ( .A1(n4483), .A2(n5254), .ZN(n5259) );
  INV_X1 U5478 ( .A(n4508), .ZN(n4677) );
  NAND2_X1 U5479 ( .A1(n5655), .A2(n5654), .ZN(n9022) );
  AND2_X1 U5480 ( .A1(n4685), .A2(n4683), .ZN(n9040) );
  AOI21_X1 U5481 ( .B1(n8366), .B2(n10259), .A(n4684), .ZN(n4683) );
  NAND2_X1 U5482 ( .A1(n8127), .A2(n10264), .ZN(n4685) );
  AND2_X1 U5483 ( .A1(n8364), .A2(n8448), .ZN(n4684) );
  OR2_X1 U5484 ( .A1(n10309), .A2(n9025), .ZN(n10297) );
  NAND2_X1 U5485 ( .A1(n4576), .A2(n4973), .ZN(n9041) );
  NOR2_X1 U5486 ( .A1(n8123), .A2(n4492), .ZN(n4974) );
  AND2_X1 U5487 ( .A1(n4541), .A2(n5216), .ZN(n5034) );
  INV_X1 U5488 ( .A(n5191), .ZN(n5035) );
  INV_X1 U5489 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U5490 ( .A1(n5194), .A2(n5193), .ZN(n4711) );
  NAND2_X1 U5491 ( .A1(n5192), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5194) );
  INV_X1 U5492 ( .A(n8505), .ZN(n8086) );
  NAND2_X1 U5493 ( .A1(n7521), .A2(n7520), .ZN(n7635) );
  NAND2_X1 U5494 ( .A1(n7784), .A2(n7783), .ZN(n9906) );
  NAND2_X1 U5495 ( .A1(n6440), .A2(n6212), .ZN(n9234) );
  NAND2_X1 U5496 ( .A1(n8039), .A2(n8040), .ZN(n4709) );
  NAND2_X1 U5497 ( .A1(n4897), .A2(n4900), .ZN(n8039) );
  NAND2_X1 U5498 ( .A1(n4897), .A2(n4895), .ZN(n4899) );
  NAND2_X1 U5499 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  INV_X1 U5500 ( .A(n9687), .ZN(n9547) );
  OR3_X1 U5501 ( .A1(n7723), .A2(n7722), .A3(n7721), .ZN(n9550) );
  OR3_X1 U5502 ( .A1(n7539), .A2(n7538), .A3(n7537), .ZN(n9553) );
  AND2_X1 U5503 ( .A1(n7731), .A2(n7730), .ZN(n9649) );
  OR2_X2 U5504 ( .A1(n9956), .A2(n6319), .ZN(n10150) );
  INV_X1 U5505 ( .A(n9690), .ZN(n10148) );
  OAI21_X1 U5506 ( .B1(n9848), .B2(n9930), .A(n9847), .ZN(n4753) );
  INV_X1 U5507 ( .A(n4663), .ZN(n4662) );
  AOI21_X1 U5508 ( .B1(n5681), .B2(n5680), .A(n4664), .ZN(n4660) );
  INV_X1 U5509 ( .A(n5692), .ZN(n4661) );
  OAI21_X1 U5510 ( .B1(n4648), .B2(n4647), .A(n5733), .ZN(n5734) );
  NAND2_X1 U5511 ( .A1(n8644), .A2(n5731), .ZN(n4647) );
  AOI21_X1 U5512 ( .B1(n5725), .B2(n4650), .A(n4649), .ZN(n4648) );
  INV_X1 U5513 ( .A(n4499), .ZN(n5022) );
  INV_X1 U5514 ( .A(n5775), .ZN(n4659) );
  NAND2_X1 U5515 ( .A1(n4496), .A2(n4490), .ZN(n5020) );
  AND2_X1 U5516 ( .A1(n7435), .A2(n8372), .ZN(n4986) );
  AND2_X1 U5517 ( .A1(n4850), .A2(n5179), .ZN(n4578) );
  INV_X1 U5518 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5179) );
  INV_X1 U5519 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U5520 ( .A1(n5394), .A2(n5180), .ZN(n5421) );
  INV_X1 U5521 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4829) );
  INV_X1 U5522 ( .A(n9421), .ZN(n4941) );
  INV_X1 U5523 ( .A(n5178), .ZN(n4816) );
  INV_X1 U5524 ( .A(n4815), .ZN(n4814) );
  OAI21_X1 U5525 ( .B1(n5603), .B2(n4816), .A(n5615), .ZN(n4815) );
  NOR2_X1 U5526 ( .A1(n5550), .A2(n4644), .ZN(n4643) );
  INV_X1 U5527 ( .A(n5149), .ZN(n4644) );
  INV_X1 U5528 ( .A(n4717), .ZN(n4716) );
  OAI21_X1 U5529 ( .B1(n4719), .B2(n4718), .A(n5135), .ZN(n4717) );
  INV_X1 U5530 ( .A(n5133), .ZN(n4718) );
  INV_X1 U5531 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5130) );
  INV_X1 U5532 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5119) );
  INV_X1 U5533 ( .A(n4821), .ZN(n4820) );
  INV_X1 U5534 ( .A(n5077), .ZN(n4989) );
  AOI21_X1 U5535 ( .B1(n4653), .B2(n4655), .A(n4658), .ZN(n4651) );
  NAND2_X1 U5536 ( .A1(n8123), .A2(n4525), .ZN(n4658) );
  NAND2_X1 U5537 ( .A1(n4496), .A2(n4490), .ZN(n5814) );
  NAND2_X1 U5538 ( .A1(n8471), .A2(n4741), .ZN(n4740) );
  AND2_X1 U5539 ( .A1(n5030), .A2(n5031), .ZN(n5029) );
  NAND2_X1 U5540 ( .A1(n5029), .A2(n4681), .ZN(n4678) );
  NOR2_X1 U5541 ( .A1(n9081), .A2(n9088), .ZN(n4731) );
  INV_X1 U5542 ( .A(n5746), .ZN(n4742) );
  NAND2_X1 U5543 ( .A1(n4690), .A2(n4688), .ZN(n4687) );
  OR2_X1 U5544 ( .A1(n8110), .A2(n8330), .ZN(n5666) );
  NAND2_X1 U5545 ( .A1(n4965), .A2(n4964), .ZN(n4963) );
  INV_X1 U5546 ( .A(n4966), .ZN(n4964) );
  NOR2_X1 U5547 ( .A1(n7224), .A2(n4986), .ZN(n4983) );
  OR2_X1 U5548 ( .A1(n4984), .A2(n4986), .ZN(n4982) );
  OR2_X1 U5549 ( .A1(n7393), .A2(n7374), .ZN(n5804) );
  NAND2_X1 U5550 ( .A1(n5374), .A2(n5798), .ZN(n6996) );
  INV_X1 U5551 ( .A(n4585), .ZN(n4584) );
  OAI21_X1 U5552 ( .B1(n10265), .B2(n4586), .A(n9005), .ZN(n4585) );
  INV_X1 U5553 ( .A(n6939), .ZN(n4586) );
  AND2_X1 U5554 ( .A1(n10278), .A2(n5686), .ZN(n6585) );
  INV_X1 U5555 ( .A(n7336), .ZN(n6597) );
  NAND2_X1 U5556 ( .A1(n10267), .A2(n10361), .ZN(n9006) );
  NAND2_X1 U5557 ( .A1(n7879), .A2(n9219), .ZN(n7898) );
  INV_X1 U5558 ( .A(n9155), .ZN(n4901) );
  NAND2_X1 U5559 ( .A1(n4699), .A2(n4527), .ZN(n7797) );
  NOR2_X1 U5560 ( .A1(n6034), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6156) );
  OR2_X1 U5561 ( .A1(n6477), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6770) );
  NOR2_X1 U5562 ( .A1(n4914), .A2(n7989), .ZN(n4913) );
  OR2_X1 U5563 ( .A1(n7901), .A2(n9201), .ZN(n7919) );
  INV_X1 U5564 ( .A(n9415), .ZN(n4943) );
  INV_X1 U5565 ( .A(n7972), .ZN(n4761) );
  INV_X1 U5566 ( .A(n4776), .ZN(n4772) );
  OR2_X1 U5567 ( .A1(n9919), .A2(n9928), .ZN(n4750) );
  AND2_X1 U5568 ( .A1(n9275), .A2(n9367), .ZN(n9313) );
  INV_X1 U5569 ( .A(n4793), .ZN(n4790) );
  NAND2_X1 U5570 ( .A1(n6675), .A2(n4923), .ZN(n4926) );
  NOR2_X1 U5571 ( .A1(n6704), .A2(n4928), .ZN(n4923) );
  INV_X1 U5572 ( .A(n9482), .ZN(n4928) );
  NAND2_X1 U5573 ( .A1(n4946), .A2(n4945), .ZN(n4944) );
  NAND2_X1 U5574 ( .A1(n4746), .A2(n4745), .ZN(n7296) );
  INV_X1 U5575 ( .A(n4746), .ZN(n6979) );
  NAND2_X1 U5576 ( .A1(n9536), .A2(n10148), .ZN(n9460) );
  AOI21_X1 U5577 ( .B1(n4807), .B2(n4809), .A(n4561), .ZN(n4806) );
  INV_X1 U5578 ( .A(n5562), .ZN(n4807) );
  INV_X1 U5579 ( .A(n4809), .ZN(n4808) );
  INV_X1 U5580 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5853) );
  INV_X1 U5581 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5852) );
  INV_X1 U5582 ( .A(SI_16_), .ZN(n5125) );
  INV_X1 U5583 ( .A(n5118), .ZN(n4633) );
  NOR2_X1 U5584 ( .A1(n5115), .A2(n4636), .ZN(n4635) );
  INV_X1 U5585 ( .A(n5114), .ZN(n4636) );
  AND2_X1 U5586 ( .A1(n6770), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6478) );
  OR2_X1 U5587 ( .A1(n6374), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6477) );
  AND2_X1 U5588 ( .A1(n5391), .A2(n5101), .ZN(n4618) );
  NOR2_X1 U5589 ( .A1(n4822), .A2(n4989), .ZN(n4821) );
  INV_X1 U5590 ( .A(n5072), .ZN(n4822) );
  INV_X1 U5591 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4736) );
  INV_X1 U5592 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4738) );
  NAND2_X1 U5593 ( .A1(n7512), .A2(n7511), .ZN(n7600) );
  NAND2_X1 U5594 ( .A1(n4677), .A2(n6661), .ZN(n6610) );
  INV_X1 U5595 ( .A(n7599), .ZN(n4843) );
  INV_X1 U5596 ( .A(n7663), .ZN(n4839) );
  INV_X1 U5597 ( .A(n7511), .ZN(n4840) );
  NOR2_X1 U5598 ( .A1(n4864), .A2(n4564), .ZN(n4863) );
  NAND2_X1 U5599 ( .A1(n4856), .A2(n4854), .ZN(n4853) );
  INV_X1 U5600 ( .A(n6299), .ZN(n4855) );
  NAND2_X1 U5601 ( .A1(n7153), .A2(n7154), .ZN(n8186) );
  NAND2_X1 U5602 ( .A1(n5204), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U5603 ( .A1(n5208), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U5604 ( .A1(n8186), .A2(n8187), .ZN(n8185) );
  INV_X1 U5605 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U5606 ( .A1(n7600), .A2(n7599), .ZN(n8270) );
  AOI21_X1 U5607 ( .B1(n5015), .B2(n5017), .A(n4498), .ZN(n5014) );
  INV_X1 U5608 ( .A(n5814), .ZN(n4826) );
  NOR2_X1 U5609 ( .A1(n5813), .A2(n8464), .ZN(n4825) );
  AND2_X1 U5610 ( .A1(n8413), .A2(n6490), .ZN(n6493) );
  NAND2_X1 U5611 ( .A1(n6691), .A2(n4569), .ZN(n6693) );
  OR2_X1 U5612 ( .A1(n6692), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4569) );
  NAND2_X1 U5613 ( .A1(n6693), .A2(n6694), .ZN(n6956) );
  INV_X1 U5614 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5436) );
  NOR2_X1 U5615 ( .A1(n7246), .A2(n7247), .ZN(n8066) );
  AOI21_X1 U5616 ( .B1(n8071), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8066), .ZN(
        n8430) );
  NOR2_X1 U5617 ( .A1(n8515), .A2(n4739), .ZN(n8485) );
  INV_X1 U5618 ( .A(n4741), .ZN(n4739) );
  OR2_X1 U5619 ( .A1(n8515), .A2(n4740), .ZN(n8466) );
  INV_X1 U5620 ( .A(n8495), .ZN(n8492) );
  AND3_X1 U5621 ( .A1(n5591), .A2(n5590), .A3(n5589), .ZN(n8539) );
  NAND2_X1 U5622 ( .A1(n4710), .A2(n5582), .ZN(n8541) );
  OR2_X1 U5623 ( .A1(n5566), .A2(n8178), .ZN(n5577) );
  NAND2_X1 U5624 ( .A1(n8611), .A2(n4516), .ZN(n8549) );
  NAND2_X1 U5625 ( .A1(n8611), .A2(n4729), .ZN(n8563) );
  NAND2_X1 U5626 ( .A1(n4733), .A2(n8614), .ZN(n8602) );
  NAND2_X1 U5627 ( .A1(n8611), .A2(n8605), .ZN(n8600) );
  NOR2_X1 U5628 ( .A1(n4600), .A2(n4553), .ZN(n4599) );
  NAND2_X1 U5629 ( .A1(n8654), .A2(n10011), .ZN(n8624) );
  AND2_X1 U5630 ( .A1(n7395), .A2(n4984), .ZN(n7434) );
  NAND2_X1 U5631 ( .A1(n7395), .A2(n7394), .ZN(n7396) );
  NOR2_X1 U5632 ( .A1(n4724), .A2(n7393), .ZN(n4723) );
  INV_X1 U5633 ( .A(n4725), .ZN(n4724) );
  AND2_X1 U5634 ( .A1(n7223), .A2(n7222), .ZN(n7226) );
  NAND2_X1 U5635 ( .A1(n7226), .A2(n7225), .ZN(n7395) );
  NAND2_X1 U5636 ( .A1(n7079), .A2(n7082), .ZN(n7223) );
  NAND2_X1 U5637 ( .A1(n4996), .A2(n4994), .ZN(n4993) );
  NAND2_X1 U5638 ( .A1(n5374), .A2(n4996), .ZN(n4995) );
  AOI21_X1 U5639 ( .B1(n7076), .B2(n4998), .A(n4997), .ZN(n4996) );
  NAND2_X1 U5640 ( .A1(n6996), .A2(n7076), .ZN(n7083) );
  NAND2_X1 U5641 ( .A1(n7003), .A2(n10387), .ZN(n7228) );
  NAND2_X1 U5642 ( .A1(n5202), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U5643 ( .A1(n5001), .A2(n5003), .ZN(n4999) );
  INV_X1 U5644 ( .A(n5002), .ZN(n5001) );
  OR2_X1 U5645 ( .A1(n9006), .A2(n9012), .ZN(n10246) );
  NOR2_X1 U5646 ( .A1(n10294), .A2(n8289), .ZN(n10267) );
  INV_X1 U5647 ( .A(n10344), .ZN(n10292) );
  OR2_X1 U5648 ( .A1(n10293), .A2(n4722), .ZN(n10294) );
  OR2_X1 U5649 ( .A1(n10301), .A2(n10292), .ZN(n4722) );
  NOR2_X1 U5650 ( .A1(n6613), .A2(n6661), .ZN(n6864) );
  NAND2_X1 U5651 ( .A1(n4677), .A2(n4834), .ZN(n6368) );
  AND2_X1 U5652 ( .A1(n5781), .A2(n4499), .ZN(n8123) );
  OAI21_X1 U5653 ( .B1(n8463), .B2(n4976), .A(n4975), .ZN(n4577) );
  NAND2_X1 U5654 ( .A1(n8123), .A2(n4492), .ZN(n4975) );
  INV_X1 U5655 ( .A(n8123), .ZN(n4976) );
  NAND2_X1 U5656 ( .A1(n5586), .A2(n5585), .ZN(n9063) );
  INV_X1 U5657 ( .A(n10402), .ZN(n10295) );
  NAND2_X1 U5658 ( .A1(n10258), .A2(n5693), .ZN(n9015) );
  NAND2_X1 U5659 ( .A1(n5295), .A2(n4666), .ZN(n4665) );
  NOR2_X1 U5660 ( .A1(n6540), .A2(n5329), .ZN(n4667) );
  INV_X1 U5661 ( .A(n6613), .ZN(n10333) );
  INV_X1 U5662 ( .A(n10376), .ZN(n10400) );
  NOR2_X1 U5663 ( .A1(n9029), .A2(n9028), .ZN(n9105) );
  INV_X1 U5664 ( .A(n7672), .ZN(n6126) );
  NAND2_X1 U5665 ( .A1(n5191), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U5666 ( .A1(n4587), .A2(n5394), .ZN(n5195) );
  AND2_X1 U5667 ( .A1(n5185), .A2(n4588), .ZN(n4587) );
  AND2_X1 U5668 ( .A1(n5190), .A2(n5036), .ZN(n4588) );
  AND2_X1 U5669 ( .A1(n5834), .A2(n5191), .ZN(n6125) );
  OR2_X1 U5670 ( .A1(n5830), .A2(n5829), .ZN(n5835) );
  NAND2_X1 U5671 ( .A1(n5832), .A2(n5831), .ZN(n5837) );
  INV_X1 U5672 ( .A(n5835), .ZN(n5832) );
  AOI21_X1 U5673 ( .B1(n4874), .B2(n5479), .A(n5479), .ZN(n4871) );
  AND2_X1 U5674 ( .A1(n7031), .A2(n4907), .ZN(n4904) );
  XNOR2_X1 U5675 ( .A(n6548), .B(n7947), .ZN(n6775) );
  NOR2_X1 U5676 ( .A1(n7471), .A2(n4698), .ZN(n4697) );
  INV_X1 U5677 ( .A(n7467), .ZN(n4698) );
  NAND2_X1 U5678 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  OR2_X1 U5679 ( .A1(n7934), .A2(n7933), .ZN(n4900) );
  INV_X1 U5680 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7569) );
  AND2_X1 U5681 ( .A1(n9526), .A2(n9525), .ZN(n9533) );
  AND4_X1 U5682 ( .A1(n6827), .A2(n6826), .A3(n6825), .A4(n6824), .ZN(n7011)
         );
  NAND2_X1 U5683 ( .A1(n9640), .A2(n9444), .ZN(n9614) );
  NAND2_X1 U5684 ( .A1(n9444), .A2(n9442), .ZN(n9636) );
  INV_X1 U5685 ( .A(n9636), .ZN(n9629) );
  NAND2_X1 U5686 ( .A1(n9650), .A2(n9651), .ZN(n9656) );
  AND2_X1 U5687 ( .A1(n9440), .A2(n9441), .ZN(n9651) );
  NAND2_X1 U5688 ( .A1(n4915), .A2(n4916), .ZN(n9669) );
  AND2_X1 U5689 ( .A1(n7980), .A2(n9693), .ZN(n9692) );
  AND2_X1 U5690 ( .A1(n9426), .A2(n9424), .ZN(n9695) );
  INV_X1 U5691 ( .A(n9729), .ZN(n9688) );
  NAND2_X1 U5692 ( .A1(n9707), .A2(n9708), .ZN(n9712) );
  AOI21_X1 U5693 ( .B1(n4767), .B2(n4769), .A(n4526), .ZN(n4765) );
  NAND2_X1 U5694 ( .A1(n4944), .A2(n4942), .ZN(n9737) );
  NAND2_X1 U5695 ( .A1(n9718), .A2(n9724), .ZN(n9719) );
  AND2_X1 U5696 ( .A1(n9416), .A2(n9725), .ZN(n9744) );
  NAND2_X1 U5697 ( .A1(n6626), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7827) );
  OR2_X1 U5698 ( .A1(n7827), .A2(n9213), .ZN(n7847) );
  NAND2_X1 U5699 ( .A1(n4931), .A2(n4932), .ZN(n9771) );
  AOI21_X1 U5700 ( .B1(n9805), .B2(n4934), .A(n4933), .ZN(n4932) );
  NOR2_X2 U5701 ( .A1(n4751), .A2(n9911), .ZN(n9798) );
  NAND2_X1 U5702 ( .A1(n6624), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7719) );
  INV_X1 U5703 ( .A(n7702), .ZN(n6624) );
  NOR2_X1 U5704 ( .A1(n9814), .A2(n4930), .ZN(n4929) );
  INV_X1 U5705 ( .A(n9375), .ZN(n4930) );
  NOR2_X1 U5706 ( .A1(n7626), .A2(n4750), .ZN(n9825) );
  NAND2_X1 U5707 ( .A1(n7724), .A2(n9375), .ZN(n9815) );
  INV_X1 U5708 ( .A(n7532), .ZN(n6623) );
  INV_X1 U5709 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7472) );
  OR2_X1 U5710 ( .A1(n7473), .A2(n7472), .ZN(n7532) );
  INV_X1 U5711 ( .A(n4571), .ZN(n7626) );
  NOR2_X1 U5712 ( .A1(n4744), .A2(n10203), .ZN(n4743) );
  INV_X1 U5713 ( .A(n4745), .ZN(n4744) );
  INV_X1 U5714 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6919) );
  NOR2_X1 U5715 ( .A1(n6979), .A2(n7043), .ZN(n7023) );
  NOR3_X1 U5716 ( .A1(n6979), .A2(n7043), .A3(n7092), .ZN(n7109) );
  AND2_X1 U5717 ( .A1(n4926), .A2(n9490), .ZN(n6878) );
  NAND2_X1 U5718 ( .A1(n9488), .A2(n9490), .ZN(n9299) );
  NAND2_X1 U5719 ( .A1(n6675), .A2(n9482), .ZN(n6705) );
  AND3_X1 U5720 ( .A1(n6511), .A2(n6510), .A3(n6509), .ZN(n6681) );
  NAND2_X1 U5721 ( .A1(n8096), .A2(n8095), .ZN(n9840) );
  NAND2_X1 U5722 ( .A1(n7826), .A2(n7825), .ZN(n9896) );
  NAND2_X1 U5723 ( .A1(n7805), .A2(n7804), .ZN(n9900) );
  INV_X1 U5724 ( .A(n6681), .ZN(n6731) );
  AND2_X1 U5725 ( .A1(n6321), .A2(n9534), .ZN(n10000) );
  OR2_X1 U5726 ( .A1(n6654), .A2(n9527), .ZN(n10205) );
  INV_X1 U5727 ( .A(n10000), .ZN(n10204) );
  NAND2_X1 U5728 ( .A1(n9536), .A2(n9472), .ZN(n6654) );
  AND2_X1 U5729 ( .A1(n6318), .A2(n6348), .ZN(n6653) );
  INV_X1 U5730 ( .A(SI_30_), .ZN(n4823) );
  XNOR2_X1 U5731 ( .A(n5647), .B(SI_30_), .ZN(n8106) );
  XNOR2_X1 U5732 ( .A(n5633), .B(n5619), .ZN(n9125) );
  AND2_X1 U5733 ( .A1(n4948), .A2(n5889), .ZN(n4798) );
  XNOR2_X1 U5734 ( .A(n5616), .B(n5615), .ZN(n8004) );
  NAND2_X1 U5735 ( .A1(n4813), .A2(n5178), .ZN(n5616) );
  INV_X1 U5736 ( .A(n5878), .ZN(n5879) );
  NAND2_X1 U5737 ( .A1(n4507), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  AND2_X1 U5738 ( .A1(n4513), .A2(n5866), .ZN(n4947) );
  INV_X1 U5739 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5869) );
  INV_X1 U5740 ( .A(n4637), .ZN(n5573) );
  OAI21_X1 U5741 ( .B1(n5537), .B2(n4562), .A(n4502), .ZN(n4637) );
  NAND2_X1 U5742 ( .A1(n4645), .A2(n5149), .ZN(n5551) );
  INV_X1 U5743 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U5744 ( .A1(n4715), .A2(n5133), .ZN(n5497) );
  NAND2_X1 U5745 ( .A1(n4827), .A2(n4719), .ZN(n4715) );
  XNOR2_X1 U5746 ( .A(n5433), .B(n5432), .ZN(n7553) );
  OR2_X1 U5747 ( .A1(n5934), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6034) );
  INV_X1 U5748 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5922) );
  INV_X1 U5749 ( .A(n5328), .ZN(n4992) );
  NAND2_X1 U5750 ( .A1(n4817), .A2(n4987), .ZN(n5327) );
  NAND2_X1 U5751 ( .A1(n5293), .A2(n4821), .ZN(n4817) );
  OR2_X1 U5753 ( .A1(n5054), .A2(SI_1_), .ZN(n4712) );
  NAND2_X1 U5754 ( .A1(n5058), .A2(n5057), .ZN(n5242) );
  NAND2_X1 U5755 ( .A1(n6417), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U5756 ( .A1(n5055), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5057) );
  AND2_X1 U5757 ( .A1(n5338), .A2(n5337), .ZN(n10367) );
  NAND2_X1 U5758 ( .A1(n6761), .A2(n6760), .ZN(n8228) );
  AOI21_X1 U5759 ( .B1(n4884), .B2(n4882), .A(n4880), .ZN(n4879) );
  OAI21_X1 U5760 ( .B1(n4882), .B2(n4881), .A(n8220), .ZN(n4880) );
  NAND2_X1 U5761 ( .A1(n4887), .A2(n8219), .ZN(n4881) );
  INV_X1 U5762 ( .A(n4884), .ZN(n4883) );
  OAI21_X1 U5763 ( .B1(n8146), .B2(n4848), .A(n4846), .ZN(n8245) );
  NAND2_X1 U5764 ( .A1(n5467), .A2(n5466), .ZN(n10015) );
  NAND2_X1 U5765 ( .A1(n6749), .A2(n6748), .ZN(n8335) );
  INV_X1 U5766 ( .A(n8284), .ZN(n6749) );
  NAND2_X1 U5767 ( .A1(n4853), .A2(n6304), .ZN(n6741) );
  INV_X1 U5768 ( .A(n8375), .ZN(n7185) );
  INV_X1 U5769 ( .A(n8373), .ZN(n7374) );
  INV_X1 U5770 ( .A(n8346), .ZN(n8356) );
  NAND2_X1 U5771 ( .A1(n8135), .A2(n8323), .ZN(n8327) );
  AND2_X1 U5772 ( .A1(n6293), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8342) );
  INV_X1 U5773 ( .A(n8160), .ZN(n4866) );
  INV_X1 U5774 ( .A(n8362), .ZN(n8336) );
  NAND2_X1 U5775 ( .A1(n5451), .A2(n5450), .ZN(n7607) );
  OR2_X1 U5776 ( .A1(n4483), .A2(n5269), .ZN(n5272) );
  INV_X1 U5777 ( .A(P2_U3966), .ZN(n8383) );
  OR2_X1 U5778 ( .A1(n4483), .A2(n6617), .ZN(n5240) );
  INV_X1 U5779 ( .A(n10229), .ZN(n10224) );
  XNOR2_X1 U5780 ( .A(n8067), .B(n8078), .ZN(n8436) );
  NAND2_X1 U5781 ( .A1(n8436), .A2(n5505), .ZN(n8435) );
  AND2_X1 U5782 ( .A1(n5778), .A2(n5033), .ZN(n8459) );
  NAND2_X1 U5783 ( .A1(n8494), .A2(n5776), .ZN(n8476) );
  NAND2_X1 U5784 ( .A1(n5595), .A2(n5594), .ZN(n9056) );
  NAND2_X1 U5785 ( .A1(n4591), .A2(n4594), .ZN(n8513) );
  OR2_X1 U5786 ( .A1(n4495), .A2(n8579), .ZN(n4591) );
  OAI21_X1 U5787 ( .B1(n8562), .B2(n4957), .A(n4955), .ZN(n8530) );
  NAND2_X1 U5788 ( .A1(n4956), .A2(n4958), .ZN(n8546) );
  AND2_X1 U5789 ( .A1(n4958), .A2(n4510), .ZN(n8548) );
  NAND2_X1 U5790 ( .A1(n8562), .A2(n8114), .ZN(n4958) );
  AND2_X1 U5791 ( .A1(n8568), .A2(n5757), .ZN(n8557) );
  AND2_X1 U5792 ( .A1(n8584), .A2(n5750), .ZN(n8570) );
  NAND2_X1 U5793 ( .A1(n8599), .A2(n8598), .ZN(n9086) );
  NAND2_X1 U5794 ( .A1(n8615), .A2(n5746), .ZN(n8592) );
  AND2_X1 U5795 ( .A1(n8629), .A2(n5743), .ZN(n8616) );
  NAND2_X1 U5796 ( .A1(n4601), .A2(n4504), .ZN(n8610) );
  NAND2_X1 U5797 ( .A1(n8109), .A2(n4602), .ZN(n4601) );
  NAND2_X1 U5798 ( .A1(n8109), .A2(n4605), .ZN(n8622) );
  NAND2_X1 U5799 ( .A1(n4962), .A2(n4965), .ZN(n8645) );
  NAND2_X1 U5800 ( .A1(n7580), .A2(n4966), .ZN(n4962) );
  NAND2_X1 U5801 ( .A1(n7580), .A2(n4969), .ZN(n7677) );
  NAND2_X1 U5802 ( .A1(n5007), .A2(n5726), .ZN(n7584) );
  NAND2_X1 U5803 ( .A1(n5010), .A2(n5008), .ZN(n7438) );
  NAND2_X1 U5804 ( .A1(n5397), .A2(n5396), .ZN(n7227) );
  NAND2_X1 U5805 ( .A1(n6995), .A2(n6994), .ZN(n7075) );
  AND2_X1 U5806 ( .A1(n10239), .A2(n6943), .ZN(n6945) );
  NAND2_X1 U5807 ( .A1(n5352), .A2(n5351), .ZN(n10375) );
  NAND2_X1 U5808 ( .A1(n10266), .A2(n10265), .ZN(n4583) );
  INV_X1 U5809 ( .A(n10351), .ZN(n10301) );
  OR2_X1 U5810 ( .A1(n10304), .A2(n10402), .ZN(n10273) );
  AOI21_X1 U5811 ( .B1(n6608), .B2(n10264), .A(n4673), .ZN(n10334) );
  NAND2_X1 U5812 ( .A1(n4675), .A2(n4674), .ZN(n4673) );
  NAND2_X1 U5813 ( .A1(n4677), .A2(n10259), .ZN(n4674) );
  NAND2_X1 U5814 ( .A1(n6602), .A2(n10297), .ZN(n10299) );
  INV_X1 U5815 ( .A(n8627), .ZN(n10302) );
  INV_X1 U5816 ( .A(n10273), .ZN(n8637) );
  INV_X1 U5817 ( .A(n8639), .ZN(n10306) );
  INV_X1 U5818 ( .A(n10297), .ZN(n10245) );
  AND2_X2 U5819 ( .A1(n9105), .A2(n9103), .ZN(n10430) );
  INV_X1 U5820 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n4980) );
  AND2_X1 U5821 ( .A1(n6287), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10325) );
  INV_X1 U5822 ( .A(n10319), .ZN(n10322) );
  XNOR2_X1 U5823 ( .A(n5841), .B(n5840), .ZN(n7611) );
  INV_X1 U5824 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8899) );
  INV_X1 U5825 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8865) );
  INV_X1 U5826 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7284) );
  INV_X1 U5827 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7047) );
  NOR2_X1 U5828 ( .A1(n5483), .A2(n5482), .ZN(n8421) );
  INV_X1 U5829 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6640) );
  INV_X1 U5830 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6476) );
  INV_X1 U5831 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6378) );
  INV_X1 U5832 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6113) );
  AND2_X1 U5833 ( .A1(n5381), .A2(n5380), .ZN(n8396) );
  NAND2_X1 U5834 ( .A1(n5250), .A2(n5249), .ZN(n6062) );
  MUX2_X1 U5835 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5248), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5250) );
  OR2_X1 U5836 ( .A1(n6522), .A2(n6519), .ZN(n5957) );
  NAND2_X1 U5837 ( .A1(n6813), .A2(n7031), .ZN(n6906) );
  AND2_X1 U5838 ( .A1(n4694), .A2(n6808), .ZN(n6813) );
  OR2_X1 U5839 ( .A1(n9172), .A2(n4894), .ZN(n4893) );
  NAND2_X1 U5840 ( .A1(n4892), .A2(n4898), .ZN(n4891) );
  INV_X1 U5841 ( .A(n4898), .ZN(n4894) );
  NAND2_X1 U5842 ( .A1(n7883), .A2(n7882), .ZN(n9878) );
  NAND2_X1 U5843 ( .A1(n9230), .A2(n4902), .ZN(n9154) );
  NAND2_X1 U5844 ( .A1(n7468), .A2(n7467), .ZN(n7470) );
  AND2_X1 U5845 ( .A1(n7738), .A2(n7737), .ZN(n9671) );
  AND4_X1 U5846 ( .A1(n7791), .A2(n7790), .A3(n7789), .A4(n7788), .ZN(n9809)
         );
  AND2_X1 U5847 ( .A1(n4699), .A2(n4700), .ZN(n9190) );
  NAND2_X1 U5848 ( .A1(n9178), .A2(n7768), .ZN(n9191) );
  AND2_X1 U5849 ( .A1(n7927), .A2(n7926), .ZN(n9687) );
  AND2_X1 U5850 ( .A1(n4703), .A2(n4705), .ZN(n9208) );
  NAND2_X1 U5851 ( .A1(n9157), .A2(n9153), .ZN(n9209) );
  NAND2_X1 U5852 ( .A1(n7525), .A2(n7524), .ZN(n9932) );
  NAND2_X1 U5853 ( .A1(n7346), .A2(n7345), .ZN(n7352) );
  INV_X1 U5854 ( .A(n9203), .ZN(n9249) );
  MUX2_X1 U5855 ( .A(n9471), .B(n9470), .S(n10148), .Z(n9532) );
  INV_X1 U5856 ( .A(n9468), .ZN(n9329) );
  NAND2_X1 U5857 ( .A1(n9477), .A2(n9527), .ZN(n9531) );
  INV_X1 U5858 ( .A(n9671), .ZN(n9546) );
  OR3_X1 U5859 ( .A1(n7479), .A2(n7478), .A3(n7477), .ZN(n9554) );
  INV_X1 U5860 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6396) );
  AND4_X1 U5861 ( .A1(n6395), .A2(n6394), .A3(n6393), .A4(n6392), .ZN(n7619)
         );
  INV_X1 U5862 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5952) );
  AND4_X1 U5863 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n7422)
         );
  OR3_X1 U5864 ( .A1(n6926), .A2(n6925), .A3(n6924), .ZN(n9556) );
  AND4_X1 U5865 ( .A1(n6385), .A2(n6384), .A3(n6383), .A4(n6382), .ZN(n7291)
         );
  INV_X1 U5866 ( .A(n7011), .ZN(n9557) );
  NAND4_X1 U5867 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n9561)
         );
  INV_X1 U5868 ( .A(P1_U4006), .ZN(n9563) );
  INV_X1 U5869 ( .A(n9293), .ZN(n9839) );
  INV_X1 U5870 ( .A(n9840), .ZN(n9607) );
  AOI222_X1 U5871 ( .A1(n10135), .A2(n7997), .B1(n9544), .B2(n8103), .C1(n9545), .C2(n10137), .ZN(n9847) );
  NAND2_X1 U5872 ( .A1(n4920), .A2(n9451), .ZN(n4919) );
  NAND2_X1 U5873 ( .A1(n4621), .A2(n4624), .ZN(n9612) );
  OR2_X1 U5874 ( .A1(n9645), .A2(n4625), .ZN(n4621) );
  NAND2_X1 U5875 ( .A1(n7917), .A2(n7916), .ZN(n9667) );
  NAND2_X1 U5876 ( .A1(n4615), .A2(n7900), .ZN(n9875) );
  NAND2_X1 U5877 ( .A1(n9743), .A2(n7977), .ZN(n9717) );
  NAND2_X1 U5878 ( .A1(n4758), .A2(n7972), .ZN(n9763) );
  NAND2_X1 U5879 ( .A1(n9779), .A2(n9781), .ZN(n4758) );
  NAND2_X1 U5880 ( .A1(n4936), .A2(n9260), .ZN(n9780) );
  NAND2_X1 U5881 ( .A1(n4770), .A2(n4774), .ZN(n7710) );
  NAND2_X1 U5882 ( .A1(n7692), .A2(n4776), .ZN(n4770) );
  OAI21_X1 U5883 ( .B1(n7692), .B2(n4494), .A(n7693), .ZN(n9821) );
  NAND2_X1 U5884 ( .A1(n7458), .A2(n7457), .ZN(n7547) );
  NAND2_X1 U5885 ( .A1(n7342), .A2(n7341), .ZN(n7489) );
  NAND2_X1 U5886 ( .A1(n7259), .A2(n7258), .ZN(n10001) );
  NAND2_X1 U5887 ( .A1(n7289), .A2(n7288), .ZN(n7320) );
  NAND2_X1 U5888 ( .A1(n7010), .A2(n7009), .ZN(n7012) );
  INV_X1 U5889 ( .A(n9830), .ZN(n9799) );
  NAND2_X1 U5890 ( .A1(n6884), .A2(n6883), .ZN(n6968) );
  AND2_X1 U5891 ( .A1(n9810), .A2(n10149), .ZN(n9830) );
  INV_X1 U5892 ( .A(n9832), .ZN(n9733) );
  OAI211_X1 U5893 ( .C1(n9611), .C2(n9326), .A(n4785), .B(n4783), .ZN(n9848)
         );
  NAND2_X1 U5894 ( .A1(n4488), .A2(n9456), .ZN(n4785) );
  NOR2_X1 U5895 ( .A1(n4488), .A2(n9456), .ZN(n4784) );
  OR2_X1 U5896 ( .A1(n9847), .A2(n10211), .ZN(n4782) );
  INV_X1 U5897 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4788) );
  AOI21_X1 U5898 ( .B1(n9845), .B2(n10146), .A(n4754), .ZN(n9846) );
  AND2_X1 U5899 ( .A1(n9844), .A2(n10000), .ZN(n4754) );
  NAND2_X1 U5900 ( .A1(n6522), .A2(n5908), .ZN(n9956) );
  AND2_X1 U5901 ( .A1(n4799), .A2(n5938), .ZN(n4797) );
  INV_X1 U5902 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5938) );
  OAI21_X1 U5903 ( .B1(n5647), .B2(n4823), .A(n5650), .ZN(n5653) );
  INV_X1 U5904 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8783) );
  NAND2_X1 U5905 ( .A1(n5874), .A2(n5876), .ZN(n5867) );
  INV_X1 U5906 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7861) );
  INV_X1 U5907 ( .A(n9473), .ZN(n9536) );
  INV_X1 U5908 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7824) );
  INV_X1 U5909 ( .A(n9527), .ZN(n9528) );
  INV_X1 U5910 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8817) );
  XNOR2_X1 U5911 ( .A(n6187), .B(n5864), .ZN(n9690) );
  CLKBUF_X1 U5912 ( .A(n6185), .Z(n6186) );
  INV_X1 U5913 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6875) );
  INV_X1 U5914 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8891) );
  INV_X1 U5915 ( .A(n7554), .ZN(n7056) );
  INV_X1 U5916 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6376) );
  INV_X1 U5917 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6281) );
  INV_X1 U5918 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6037) );
  INV_X1 U5919 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U5920 ( .A1(n4991), .A2(n5327), .ZN(n6778) );
  NAND2_X1 U5921 ( .A1(n4952), .A2(n5260), .ZN(n5262) );
  INV_X1 U5922 ( .A(n5060), .ZN(n4952) );
  NOR2_X1 U5923 ( .A1(n8030), .A2(n10471), .ZN(n10460) );
  AOI21_X1 U5924 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10458), .ZN(n10457) );
  NOR2_X1 U5925 ( .A1(n10457), .A2(n10456), .ZN(n10455) );
  AOI21_X1 U5926 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10455), .ZN(n10454) );
  OAI21_X1 U5927 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10452), .ZN(n10450) );
  OAI21_X1 U5928 ( .B1(n6286), .B2(n6285), .A(n4857), .ZN(n6300) );
  AOI21_X1 U5929 ( .B1(n8346), .B2(n4677), .A(n4676), .ZN(n6146) );
  NAND2_X1 U5930 ( .A1(n4668), .A2(n5847), .ZN(P2_U3244) );
  OAI21_X1 U5931 ( .B1(n4669), .B2(n5820), .A(n7449), .ZN(n4668) );
  NAND2_X1 U5932 ( .A1(P2_U3966), .A2(n4677), .ZN(n5921) );
  MUX2_X1 U5933 ( .A(n8088), .B(n8087), .S(n8086), .Z(n8090) );
  OR2_X1 U5934 ( .A1(n10430), .A2(n5625), .ZN(n4682) );
  NAND2_X1 U5935 ( .A1(n4575), .A2(n10430), .ZN(n4574) );
  OAI21_X1 U5936 ( .B1(n9041), .B2(n10327), .A(n4981), .ZN(n4575) );
  NAND2_X1 U5937 ( .A1(n10409), .A2(n10407), .ZN(n4978) );
  NAND2_X1 U5938 ( .A1(n4708), .A2(n4707), .ZN(P1_U3238) );
  AOI21_X1 U5939 ( .B1(n9859), .B2(n9251), .A(n8041), .ZN(n4707) );
  NAND2_X1 U5940 ( .A1(n4612), .A2(n4752), .ZN(P1_U3552) );
  OR2_X1 U5941 ( .A1(n10223), .A2(n6634), .ZN(n4752) );
  OAI21_X1 U5942 ( .B1(n4753), .B2(n4613), .A(n10223), .ZN(n4612) );
  INV_X1 U5943 ( .A(n9846), .ZN(n4613) );
  OAI211_X1 U5944 ( .C1(n9848), .C2(n4786), .A(n4781), .B(n4780), .ZN(P1_U3520) );
  NAND2_X1 U5945 ( .A1(n10212), .A2(n10194), .ZN(n4786) );
  OR2_X1 U5946 ( .A1(n9846), .A2(n10211), .ZN(n4780) );
  AND2_X1 U5947 ( .A1(n4782), .A2(n4787), .ZN(n4781) );
  AND2_X1 U5948 ( .A1(n9849), .A2(n9545), .ZN(n4488) );
  OR2_X1 U5949 ( .A1(n9854), .A2(n4778), .ZN(n4489) );
  NAND2_X1 U5950 ( .A1(n9034), .A2(n8364), .ZN(n4490) );
  AND2_X1 U5951 ( .A1(n9034), .A2(n4499), .ZN(n4491) );
  AND2_X1 U5952 ( .A1(n8471), .A2(n8478), .ZN(n4492) );
  NOR2_X1 U5953 ( .A1(n8482), .A2(n5777), .ZN(n4493) );
  NAND2_X1 U5954 ( .A1(n9081), .A2(n8571), .ZN(n4597) );
  AND2_X1 U5955 ( .A1(n9928), .A2(n9553), .ZN(n4494) );
  NAND2_X1 U5956 ( .A1(n4954), .A2(n4597), .ZN(n4495) );
  INV_X1 U5957 ( .A(n4957), .ZN(n4956) );
  NAND2_X1 U5958 ( .A1(n8547), .A2(n4510), .ZN(n4957) );
  NAND2_X1 U5959 ( .A1(n8523), .A2(n4680), .ZN(n8494) );
  NAND2_X1 U5960 ( .A1(n6588), .A2(n5683), .ZN(n6582) );
  NAND2_X1 U5961 ( .A1(n7938), .A2(n7937), .ZN(n9854) );
  AND2_X1 U5962 ( .A1(n5757), .A2(n5758), .ZN(n8569) );
  NAND2_X1 U5963 ( .A1(n9022), .A2(n5657), .ZN(n4496) );
  INV_X1 U5964 ( .A(n9805), .ZN(n4937) );
  AND2_X1 U5965 ( .A1(n7709), .A2(n4771), .ZN(n4497) );
  AND2_X1 U5966 ( .A1(n5815), .A2(n4496), .ZN(n4498) );
  NAND2_X1 U5967 ( .A1(n9037), .A2(n8460), .ZN(n4499) );
  AND2_X1 U5968 ( .A1(n4491), .A2(n5016), .ZN(n4500) );
  NOR2_X1 U5969 ( .A1(n5027), .A2(n5024), .ZN(n4501) );
  INV_X1 U5970 ( .A(n9043), .ZN(n8471) );
  AND2_X1 U5971 ( .A1(n7958), .A2(n7957), .ZN(n9638) );
  INV_X1 U5972 ( .A(n9638), .ZN(n9545) );
  NAND2_X1 U5973 ( .A1(n7003), .A2(n4723), .ZN(n4726) );
  OR2_X1 U5974 ( .A1(n4640), .A2(n4810), .ZN(n4502) );
  OR2_X1 U5975 ( .A1(n5446), .A2(n4633), .ZN(n4503) );
  NAND2_X1 U5976 ( .A1(n5185), .A2(n5394), .ZN(n5639) );
  OR2_X1 U5977 ( .A1(n9049), .A2(n8498), .ZN(n5778) );
  AND2_X1 U5978 ( .A1(n5523), .A2(n5743), .ZN(n4690) );
  XNOR2_X1 U5979 ( .A(n5939), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5942) );
  OR2_X1 U5980 ( .A1(n7581), .A2(n7603), .ZN(n5726) );
  OR2_X1 U5981 ( .A1(n8628), .A2(n8111), .ZN(n4504) );
  INV_X1 U5982 ( .A(n8307), .ZN(n8146) );
  XNOR2_X1 U5983 ( .A(n9043), .B(n8478), .ZN(n8464) );
  INV_X1 U5984 ( .A(n8464), .ZN(n5030) );
  NAND2_X1 U5985 ( .A1(n5109), .A2(n5403), .ZN(n4505) );
  NAND2_X1 U5986 ( .A1(n7772), .A2(n7771), .ZN(n9911) );
  NAND2_X1 U5987 ( .A1(n5423), .A2(n5422), .ZN(n7435) );
  OR2_X1 U5988 ( .A1(n8515), .A2(n9056), .ZN(n4506) );
  NAND2_X1 U5989 ( .A1(n5878), .A2(n4947), .ZN(n4507) );
  AND4_X1 U5990 ( .A1(n5233), .A2(n5232), .A3(n5234), .A4(n5231), .ZN(n4508)
         );
  INV_X1 U5991 ( .A(n6661), .ZN(n4834) );
  NAND2_X1 U5992 ( .A1(n9859), .A2(n9546), .ZN(n4509) );
  NAND2_X1 U5993 ( .A1(n8567), .A2(n8179), .ZN(n4510) );
  OR2_X1 U5994 ( .A1(n9919), .A2(n9552), .ZN(n4511) );
  AND2_X1 U5995 ( .A1(n5181), .A2(n4876), .ZN(n4512) );
  NAND2_X1 U5996 ( .A1(n5527), .A2(n5526), .ZN(n9088) );
  INV_X1 U5997 ( .A(n9071), .ZN(n4728) );
  AND2_X1 U5998 ( .A1(n5715), .A2(n7217), .ZN(n5805) );
  INV_X1 U5999 ( .A(n8537), .ZN(n5582) );
  NAND2_X1 U6000 ( .A1(n8555), .A2(n5763), .ZN(n8536) );
  AND2_X1 U6001 ( .A1(n5876), .A2(n4950), .ZN(n4513) );
  OR2_X1 U6002 ( .A1(n6456), .A2(n6455), .ZN(n4514) );
  INV_X1 U6003 ( .A(n9757), .ZN(n4945) );
  INV_X1 U6004 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4850) );
  AND2_X1 U6005 ( .A1(n8150), .A2(n8149), .ZN(n4515) );
  NAND2_X1 U6006 ( .A1(n5553), .A2(n5552), .ZN(n9076) );
  AND2_X1 U6007 ( .A1(n4729), .A2(n4728), .ZN(n4516) );
  AND2_X1 U6008 ( .A1(n5708), .A2(n7081), .ZN(n7076) );
  INV_X1 U6009 ( .A(n7076), .ZN(n4994) );
  AND2_X1 U6010 ( .A1(n7567), .A2(n9367), .ZN(n4517) );
  NAND2_X1 U6011 ( .A1(n7700), .A2(n7699), .ZN(n9916) );
  INV_X1 U6012 ( .A(n7192), .ZN(n7043) );
  OR2_X1 U6013 ( .A1(n9037), .A2(n8460), .ZN(n5781) );
  INV_X1 U6014 ( .A(n5781), .ZN(n5016) );
  NOR2_X1 U6015 ( .A1(n9710), .A2(n4614), .ZN(n4518) );
  AND2_X1 U6016 ( .A1(n5743), .A2(n5741), .ZN(n8630) );
  INV_X1 U6017 ( .A(n8630), .ZN(n4688) );
  AND2_X1 U6018 ( .A1(n5805), .A2(n7222), .ZN(n4519) );
  NAND2_X1 U6019 ( .A1(n8611), .A2(n4731), .ZN(n4732) );
  AND2_X1 U6020 ( .A1(n4944), .A2(n9415), .ZN(n4520) );
  AND2_X1 U6021 ( .A1(n4936), .A2(n4934), .ZN(n4521) );
  NOR2_X1 U6022 ( .A1(n4905), .A2(n4904), .ZN(n4522) );
  AND2_X1 U6023 ( .A1(n8471), .A2(n8366), .ZN(n4523) );
  AND2_X1 U6024 ( .A1(n9919), .A2(n9552), .ZN(n4524) );
  AND2_X1 U6025 ( .A1(n5784), .A2(n5783), .ZN(n4525) );
  AND2_X1 U6026 ( .A1(n9883), .A2(n9738), .ZN(n4526) );
  AND2_X1 U6027 ( .A1(n4700), .A2(n7780), .ZN(n4527) );
  AND2_X1 U6028 ( .A1(n4705), .A2(n7841), .ZN(n4528) );
  INV_X1 U6029 ( .A(n4570), .ZN(n9646) );
  NOR2_X1 U6030 ( .A1(n9675), .A2(n9859), .ZN(n4570) );
  NOR2_X1 U6031 ( .A1(n5771), .A2(n4659), .ZN(n4529) );
  INV_X1 U6032 ( .A(n8219), .ZN(n4890) );
  INV_X1 U6033 ( .A(n4681), .ZN(n4680) );
  NAND2_X1 U6034 ( .A1(n8495), .A2(n5773), .ZN(n4681) );
  INV_X1 U6035 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4876) );
  INV_X1 U6036 ( .A(n4970), .ZN(n4604) );
  NOR2_X1 U6037 ( .A1(n8632), .A2(n9094), .ZN(n4970) );
  INV_X1 U6038 ( .A(n4597), .ZN(n4596) );
  NAND2_X1 U6039 ( .A1(n5878), .A2(n4798), .ZN(n4530) );
  OR2_X1 U6040 ( .A1(n5294), .A2(n5325), .ZN(n4531) );
  AND2_X1 U6041 ( .A1(n4678), .A2(n5028), .ZN(n4532) );
  OAI21_X1 U6042 ( .B1(n5770), .B2(n4659), .A(n4657), .ZN(n4656) );
  AND2_X1 U6043 ( .A1(n9230), .A2(n4901), .ZN(n4533) );
  AND2_X1 U6044 ( .A1(n5729), .A2(n5730), .ZN(n7583) );
  INV_X1 U6045 ( .A(n8524), .ZN(n8512) );
  AND2_X1 U6046 ( .A1(n5773), .A2(n5768), .ZN(n8524) );
  NOR2_X1 U6047 ( .A1(n4728), .A2(n8538), .ZN(n4534) );
  OR2_X1 U6048 ( .A1(n5020), .A2(n5016), .ZN(n4535) );
  INV_X1 U6049 ( .A(n9034), .ZN(n8454) );
  AND2_X1 U6050 ( .A1(n5635), .A2(n5634), .ZN(n9034) );
  AND2_X1 U6051 ( .A1(n8208), .A2(n8207), .ZN(n4536) );
  INV_X1 U6052 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U6053 ( .A1(n7583), .A2(n4968), .ZN(n4965) );
  AND2_X1 U6054 ( .A1(n5436), .A2(n4580), .ZN(n4537) );
  INV_X1 U6055 ( .A(n5815), .ZN(n5663) );
  NAND2_X1 U6056 ( .A1(n5789), .A2(n5787), .ZN(n5815) );
  NAND2_X1 U6057 ( .A1(n7976), .A2(n7975), .ZN(n9743) );
  NAND2_X1 U6058 ( .A1(n4963), .A2(n8643), .ZN(n4538) );
  NAND2_X1 U6059 ( .A1(n9636), .A2(n4509), .ZN(n4539) );
  NAND2_X1 U6060 ( .A1(n5247), .A2(n6417), .ZN(n5329) );
  INV_X1 U6061 ( .A(n6905), .ZN(n4907) );
  AND2_X1 U6062 ( .A1(n8523), .A2(n5773), .ZN(n4540) );
  AND2_X1 U6063 ( .A1(n5215), .A2(n5036), .ZN(n4541) );
  AND2_X1 U6064 ( .A1(n9640), .A2(n4921), .ZN(n4542) );
  NOR2_X1 U6065 ( .A1(n9781), .A2(n4935), .ZN(n4934) );
  NOR2_X1 U6066 ( .A1(n7975), .A2(n4943), .ZN(n4942) );
  AND2_X1 U6067 ( .A1(n7859), .A2(n7873), .ZN(n4543) );
  AND2_X1 U6068 ( .A1(n4992), .A2(n5077), .ZN(n4544) );
  AND2_X1 U6069 ( .A1(n7354), .A2(n7345), .ZN(n4545) );
  AND2_X1 U6070 ( .A1(n4604), .A2(n4602), .ZN(n4546) );
  AND2_X1 U6071 ( .A1(n4994), .A2(n6994), .ZN(n4547) );
  AND2_X1 U6072 ( .A1(n9451), .A2(n9629), .ZN(n4548) );
  OR2_X1 U6073 ( .A1(n4599), .A2(n4970), .ZN(n4549) );
  INV_X1 U6074 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5889) );
  INV_X1 U6075 ( .A(n4988), .ZN(n4987) );
  OAI21_X1 U6076 ( .B1(n5304), .B2(n4989), .A(n5328), .ZN(n4988) );
  INV_X1 U6077 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5036) );
  AND2_X1 U6078 ( .A1(n9332), .A2(n9334), .ZN(n9304) );
  AOI21_X1 U6079 ( .B1(n9632), .B2(n6213), .A(n7942), .ZN(n9654) );
  INV_X1 U6080 ( .A(n9654), .ZN(n4778) );
  AND2_X1 U6081 ( .A1(n5047), .A2(n4501), .ZN(n5379) );
  INV_X1 U6082 ( .A(n9153), .ZN(n4706) );
  INV_X1 U6083 ( .A(n5536), .ZN(n4828) );
  AND2_X1 U6084 ( .A1(n4806), .A2(n4804), .ZN(n4550) );
  NAND2_X1 U6085 ( .A1(n5514), .A2(n5513), .ZN(n9094) );
  INV_X1 U6086 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4950) );
  INV_X1 U6087 ( .A(n8632), .ZN(n8594) );
  NOR2_X1 U6088 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5360) );
  NAND2_X1 U6089 ( .A1(n9454), .A2(n9521), .ZN(n9456) );
  INV_X1 U6090 ( .A(n9397), .ZN(n4933) );
  AND2_X1 U6091 ( .A1(n5229), .A2(n5228), .ZN(n8478) );
  INV_X1 U6092 ( .A(n5159), .ZN(n4810) );
  AND2_X1 U6093 ( .A1(n9684), .A2(n9507), .ZN(n9708) );
  INV_X1 U6094 ( .A(n9708), .ZN(n4917) );
  OR2_X1 U6095 ( .A1(n8605), .A2(n8243), .ZN(n4551) );
  AND2_X1 U6096 ( .A1(n8043), .A2(n8051), .ZN(n4552) );
  INV_X1 U6097 ( .A(n4751), .ZN(n9797) );
  NAND2_X1 U6098 ( .A1(n4749), .A2(n4571), .ZN(n4751) );
  AND2_X1 U6099 ( .A1(n9094), .A2(n8632), .ZN(n4553) );
  NAND2_X1 U6100 ( .A1(n8158), .A2(n8299), .ZN(n4554) );
  AND2_X1 U6101 ( .A1(n7566), .A2(n9367), .ZN(n4555) );
  INV_X1 U6102 ( .A(n4733), .ZN(n8623) );
  NOR2_X1 U6103 ( .A1(n8624), .A2(n9098), .ZN(n4733) );
  AND2_X1 U6104 ( .A1(n9900), .A2(n9549), .ZN(n4556) );
  AND2_X1 U6105 ( .A1(n7913), .A2(n7912), .ZN(n4557) );
  AND2_X1 U6106 ( .A1(n5010), .A2(n5723), .ZN(n4558) );
  NAND2_X1 U6107 ( .A1(n7966), .A2(n7965), .ZN(n9849) );
  AND2_X1 U6108 ( .A1(n5136), .A2(SI_18_), .ZN(n4559) );
  OR2_X1 U6109 ( .A1(n7626), .A2(n9928), .ZN(n4560) );
  AND2_X1 U6110 ( .A1(n5161), .A2(SI_24_), .ZN(n4561) );
  NAND2_X1 U6111 ( .A1(n5536), .A2(n4638), .ZN(n4562) );
  AND2_X1 U6112 ( .A1(n9649), .A2(n9671), .ZN(n4563) );
  XOR2_X1 U6113 ( .A(n9071), .B(n8165), .Z(n4564) );
  INV_X1 U6114 ( .A(n4564), .ZN(n4870) );
  NOR2_X1 U6115 ( .A1(n8253), .A2(n4866), .ZN(n4565) );
  AND2_X2 U6116 ( .A1(n9105), .A2(n9104), .ZN(n10409) );
  INV_X1 U6117 ( .A(n10409), .ZN(n10408) );
  NOR2_X1 U6118 ( .A1(n8449), .A2(n7336), .ZN(n4566) );
  NAND2_X1 U6119 ( .A1(n4583), .A2(n6939), .ZN(n9004) );
  NAND2_X1 U6120 ( .A1(n4795), .A2(n7095), .ZN(n7289) );
  NAND2_X1 U6121 ( .A1(n10276), .A2(n5687), .ZN(n10255) );
  AND2_X1 U6122 ( .A1(n7003), .A2(n4725), .ZN(n4567) );
  INV_X1 U6123 ( .A(n7399), .ZN(n5012) );
  AND2_X1 U6124 ( .A1(n9388), .A2(n9387), .ZN(n9385) );
  INV_X1 U6125 ( .A(n9385), .ZN(n7709) );
  AND2_X1 U6126 ( .A1(n5618), .A2(n8951), .ZN(n4568) );
  AND2_X1 U6127 ( .A1(n5878), .A2(n5866), .ZN(n5874) );
  INV_X1 U6128 ( .A(n6808), .ZN(n4696) );
  INV_X1 U6129 ( .A(n9253), .ZN(n9211) );
  AND2_X2 U6130 ( .A1(n6653), .A2(n6349), .ZN(n10212) );
  AND2_X1 U6131 ( .A1(n10143), .A2(n9999), .ZN(n9930) );
  NAND2_X1 U6132 ( .A1(n7118), .A2(n7117), .ZN(n10203) );
  INV_X1 U6133 ( .A(n10203), .ZN(n4748) );
  INV_X1 U6134 ( .A(n9490), .ZN(n4927) );
  INV_X1 U6135 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4911) );
  AND2_X1 U6136 ( .A1(n9035), .A2(n7336), .ZN(n6141) );
  INV_X1 U6137 ( .A(n6141), .ZN(n10326) );
  NAND2_X1 U6138 ( .A1(n5278), .A2(n5067), .ZN(n5291) );
  NAND2_X1 U6139 ( .A1(n4721), .A2(n4818), .ZN(n5335) );
  NOR2_X1 U6140 ( .A1(n5053), .A2(n6189), .ZN(n5054) );
  NAND2_X1 U6141 ( .A1(n4645), .A2(n4643), .ZN(n4639) );
  AOI21_X1 U6142 ( .B1(n6064), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6232), .ZN(
        n6270) );
  AOI21_X1 U6143 ( .B1(n6066), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6268), .ZN(
        n6246) );
  AOI21_X1 U6144 ( .B1(n6070), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6257), .ZN(
        n6222) );
  AOI21_X1 U6145 ( .B1(n9979), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9975), .ZN(
        n9989) );
  INV_X1 U6146 ( .A(n6610), .ZN(n4836) );
  NAND2_X1 U6147 ( .A1(n4835), .A2(n4833), .ZN(n6120) );
  NOR2_X2 U6148 ( .A1(n9854), .A2(n9646), .ZN(n9631) );
  NOR2_X2 U6149 ( .A1(n6723), .A2(n6731), .ZN(n6711) );
  NOR2_X2 U6150 ( .A1(n7327), .A2(n10001), .ZN(n7427) );
  NOR2_X2 U6151 ( .A1(n6876), .A2(n6970), .ZN(n4746) );
  NOR2_X2 U6152 ( .A1(n7624), .A2(n9932), .ZN(n4571) );
  XNOR2_X2 U6153 ( .A(n8153), .B(n8151), .ZN(n8315) );
  NAND2_X2 U6154 ( .A1(n8315), .A2(n8314), .ZN(n8155) );
  NAND2_X1 U6155 ( .A1(n4574), .A2(n4682), .ZN(P2_U3549) );
  INV_X1 U6156 ( .A(n4577), .ZN(n4576) );
  NAND3_X1 U6157 ( .A1(n4579), .A2(n4578), .A3(n5436), .ZN(n5184) );
  NAND3_X1 U6158 ( .A1(n4582), .A2(n4581), .A3(n6940), .ZN(n10237) );
  NAND2_X1 U6159 ( .A1(n6995), .A2(n4547), .ZN(n7078) );
  NAND2_X1 U6160 ( .A1(n8579), .A2(n4594), .ZN(n4593) );
  NAND2_X1 U6161 ( .A1(n8109), .A2(n4546), .ZN(n4598) );
  NAND2_X1 U6162 ( .A1(n4598), .A2(n4549), .ZN(n8599) );
  AND3_X2 U6163 ( .A1(n4608), .A2(n4607), .A3(n4606), .ZN(n10344) );
  OAI21_X2 U6164 ( .B1(n5102), .B2(n4505), .A(n4616), .ZN(n5420) );
  NAND2_X1 U6165 ( .A1(n9645), .A2(n4624), .ZN(n4623) );
  OR2_X2 U6166 ( .A1(n9645), .A2(n4563), .ZN(n4627) );
  NAND2_X1 U6167 ( .A1(n4727), .A2(n4635), .ZN(n4634) );
  NAND2_X1 U6168 ( .A1(n4727), .A2(n5114), .ZN(n5433) );
  XNOR2_X2 U6169 ( .A(n4646), .B(n5215), .ZN(n5844) );
  NAND2_X1 U6170 ( .A1(n5772), .A2(n4653), .ZN(n4652) );
  NAND2_X1 U6171 ( .A1(n4652), .A2(n4651), .ZN(n5785) );
  OAI21_X1 U6172 ( .B1(n4661), .B2(n4660), .A(n4662), .ZN(n5697) );
  OAI21_X1 U6173 ( .B1(n5693), .B2(n5788), .A(n9014), .ZN(n4663) );
  NOR2_X2 U6174 ( .A1(n4667), .A2(n4665), .ZN(n10351) );
  NAND3_X1 U6175 ( .A1(n5818), .A2(n10326), .A3(n4671), .ZN(n4670) );
  NAND2_X1 U6176 ( .A1(n10279), .A2(n5672), .ZN(n10276) );
  NAND2_X1 U6177 ( .A1(n5282), .A2(n6585), .ZN(n10279) );
  OAI21_X2 U6178 ( .B1(n8631), .B2(n4689), .A(n4686), .ZN(n8596) );
  NAND2_X1 U6179 ( .A1(n4692), .A2(n4691), .ZN(n5218) );
  AND2_X2 U6180 ( .A1(n5865), .A2(n4910), .ZN(n5878) );
  AOI21_X2 U6181 ( .B1(n9199), .B2(n9200), .A(n4557), .ZN(n9171) );
  OAI21_X2 U6182 ( .B1(n9145), .B2(n9146), .A(n9143), .ZN(n9199) );
  NOR2_X2 U6183 ( .A1(n7898), .A2(n7897), .ZN(n9145) );
  NAND2_X1 U6184 ( .A1(n4695), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U6185 ( .A1(n6892), .A2(n6803), .ZN(n4694) );
  NAND2_X1 U6186 ( .A1(n4693), .A2(n4903), .ZN(n7130) );
  NOR2_X1 U6187 ( .A1(n4696), .A2(n4522), .ZN(n4695) );
  NAND2_X1 U6188 ( .A1(n7468), .A2(n4697), .ZN(n7521) );
  NAND3_X1 U6189 ( .A1(n9180), .A2(n4702), .A3(n9242), .ZN(n4699) );
  NAND3_X1 U6190 ( .A1(n9180), .A2(n9179), .A3(n9242), .ZN(n9178) );
  NAND2_X1 U6191 ( .A1(n10138), .A2(n7347), .ZN(n6204) );
  NAND3_X1 U6192 ( .A1(n4709), .A2(n4899), .A3(n9211), .ZN(n4708) );
  INV_X1 U6193 ( .A(n8536), .ZN(n4710) );
  NAND2_X1 U6194 ( .A1(n5241), .A2(n5242), .ZN(n5246) );
  AND2_X1 U6195 ( .A1(n5059), .A2(n4712), .ZN(n5241) );
  NAND2_X1 U6196 ( .A1(n4827), .A2(n4716), .ZN(n4713) );
  NAND2_X1 U6197 ( .A1(n4713), .A2(n4714), .ZN(n5511) );
  NAND2_X1 U6198 ( .A1(n4827), .A2(n5129), .ZN(n5478) );
  NAND3_X1 U6199 ( .A1(n5291), .A2(n5290), .A3(n4987), .ZN(n4721) );
  OAI21_X1 U6200 ( .B1(n5335), .B2(SI_7_), .A(n5333), .ZN(n5084) );
  INV_X1 U6201 ( .A(n4726), .ZN(n7405) );
  INV_X1 U6202 ( .A(n4732), .ZN(n8580) );
  NOR2_X2 U6203 ( .A1(n8652), .A2(n10015), .ZN(n8654) );
  AND2_X4 U6204 ( .A1(n4735), .A2(n4734), .ZN(n6417) );
  NAND3_X1 U6205 ( .A1(n5049), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4734) );
  NAND3_X1 U6206 ( .A1(n4738), .A2(n4737), .A3(n4736), .ZN(n4735) );
  NOR2_X2 U6207 ( .A1(n9701), .A2(n9875), .ZN(n9681) );
  OR2_X2 U6208 ( .A1(n9719), .A2(n9878), .ZN(n9701) );
  NAND2_X1 U6209 ( .A1(n4746), .A2(n4743), .ZN(n7327) );
  OAI21_X2 U6210 ( .B1(n5879), .B2(n4755), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5890) );
  NAND2_X1 U6211 ( .A1(n9779), .A2(n4759), .ZN(n4756) );
  NAND2_X1 U6212 ( .A1(n6973), .A2(n7009), .ZN(n4764) );
  NAND2_X1 U6213 ( .A1(n7976), .A2(n4767), .ZN(n4766) );
  NAND2_X2 U6214 ( .A1(n4766), .A2(n4765), .ZN(n9700) );
  NAND2_X1 U6215 ( .A1(n9611), .A2(n4784), .ZN(n4783) );
  OR2_X1 U6216 ( .A1(n10212), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U6217 ( .A1(n7096), .A2(n4790), .ZN(n4789) );
  NAND2_X1 U6218 ( .A1(n4789), .A2(n4791), .ZN(n7412) );
  NAND2_X1 U6219 ( .A1(n6884), .A2(n4796), .ZN(n6972) );
  AND2_X1 U6220 ( .A1(n5878), .A2(n4799), .ZN(n5940) );
  NAND2_X1 U6221 ( .A1(n5878), .A2(n4797), .ZN(n9958) );
  NOR2_X1 U6222 ( .A1(n4477), .A2(n10156), .ZN(n6215) );
  NOR2_X2 U6223 ( .A1(n10246), .A2(n10375), .ZN(n10249) );
  NAND2_X1 U6224 ( .A1(n5563), .A2(n4550), .ZN(n4803) );
  INV_X4 U6225 ( .A(n6417), .ZN(n5055) );
  NAND2_X1 U6226 ( .A1(n5604), .A2(n4814), .ZN(n4812) );
  NAND2_X1 U6227 ( .A1(n5604), .A2(n5603), .ZN(n4813) );
  NAND2_X1 U6228 ( .A1(n5293), .A2(n5072), .ZN(n5305) );
  NAND3_X1 U6229 ( .A1(n4826), .A2(n5663), .A3(n4825), .ZN(n4824) );
  NAND4_X1 U6230 ( .A1(n5048), .A2(n5324), .A3(n4830), .A4(n4829), .ZN(n5026)
         );
  NAND3_X1 U6231 ( .A1(n4832), .A2(n6148), .A3(n4831), .ZN(n6149) );
  NAND2_X1 U6232 ( .A1(n6116), .A2(n6117), .ZN(n6148) );
  INV_X1 U6233 ( .A(n8212), .ZN(n8165) );
  INV_X1 U6234 ( .A(n8156), .ZN(n8211) );
  NAND2_X1 U6235 ( .A1(n8212), .A2(n4834), .ZN(n4833) );
  NAND2_X4 U6236 ( .A1(n6115), .A2(n6591), .ZN(n8212) );
  NAND2_X1 U6237 ( .A1(n8156), .A2(n4836), .ZN(n4835) );
  INV_X1 U6238 ( .A(n6116), .ZN(n4837) );
  NAND2_X1 U6239 ( .A1(n8146), .A2(n4846), .ZN(n4845) );
  NAND2_X1 U6240 ( .A1(n6286), .A2(n4857), .ZN(n4856) );
  AOI21_X1 U6241 ( .B1(n6285), .B2(n4857), .A(n4855), .ZN(n4854) );
  NAND2_X1 U6242 ( .A1(n4865), .A2(n8155), .ZN(n4860) );
  NAND2_X1 U6243 ( .A1(n4862), .A2(n4870), .ZN(n4861) );
  NAND2_X1 U6244 ( .A1(n8155), .A2(n8154), .ZN(n4862) );
  NAND2_X1 U6245 ( .A1(n8155), .A2(n4863), .ZN(n8293) );
  INV_X1 U6246 ( .A(n8154), .ZN(n4864) );
  NAND3_X1 U6247 ( .A1(n4869), .A2(n4867), .A3(n8160), .ZN(n8257) );
  NAND3_X1 U6248 ( .A1(n4869), .A2(n4867), .A3(n4565), .ZN(n8164) );
  NAND2_X1 U6249 ( .A1(n5480), .A2(n4874), .ZN(n4872) );
  NAND2_X1 U6250 ( .A1(n5480), .A2(n4512), .ZN(n4873) );
  NAND2_X1 U6251 ( .A1(n8352), .A2(n4878), .ZN(n4877) );
  OAI211_X1 U6252 ( .C1(n8352), .C2(n4883), .A(n4879), .B(n4877), .ZN(n8225)
         );
  OAI21_X1 U6253 ( .B1(n8352), .B2(n8351), .A(n8168), .ZN(n8210) );
  OAI21_X1 U6254 ( .B1(n9171), .B2(n4893), .A(n4891), .ZN(n8042) );
  INV_X1 U6255 ( .A(n4895), .ZN(n4892) );
  NAND2_X1 U6256 ( .A1(n7346), .A2(n4545), .ZN(n7468) );
  NAND2_X2 U6257 ( .A1(n9229), .A2(n9232), .ZN(n4902) );
  NAND2_X1 U6258 ( .A1(n4905), .A2(n4907), .ZN(n4903) );
  NAND2_X1 U6259 ( .A1(n4908), .A2(n7859), .ZN(n7878) );
  NAND2_X1 U6260 ( .A1(n4908), .A2(n4543), .ZN(n9220) );
  NAND2_X2 U6261 ( .A1(n6412), .A2(n4909), .ZN(n7947) );
  NAND3_X1 U6262 ( .A1(n7132), .A2(n7133), .A3(n7131), .ZN(n7256) );
  NAND2_X1 U6263 ( .A1(n7256), .A2(n7255), .ZN(n7344) );
  NAND2_X1 U6264 ( .A1(n7132), .A2(n7131), .ZN(n7135) );
  INV_X1 U6265 ( .A(n9707), .ZN(n4912) );
  NAND2_X1 U6266 ( .A1(n4912), .A2(n9511), .ZN(n4915) );
  NAND2_X1 U6267 ( .A1(n4915), .A2(n4913), .ZN(n7990) );
  NAND2_X1 U6268 ( .A1(n4918), .A2(n4919), .ZN(n7991) );
  NAND2_X1 U6269 ( .A1(n9635), .A2(n4548), .ZN(n4918) );
  NAND2_X1 U6270 ( .A1(n4926), .A2(n4924), .ZN(n7018) );
  NAND2_X1 U6271 ( .A1(n7724), .A2(n4929), .ZN(n7725) );
  NAND2_X1 U6272 ( .A1(n9806), .A2(n4934), .ZN(n4931) );
  INV_X1 U6273 ( .A(n9758), .ZN(n4946) );
  NAND2_X1 U6274 ( .A1(n4939), .A2(n4940), .ZN(n7988) );
  NAND2_X1 U6275 ( .A1(n9758), .A2(n4942), .ZN(n4939) );
  MUX2_X1 U6276 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5055), .Z(n5063) );
  MUX2_X1 U6277 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5055), .Z(n5068) );
  MUX2_X1 U6278 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5055), .Z(n5073) );
  MUX2_X1 U6279 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5055), .Z(n5078) );
  MUX2_X1 U6280 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4951), .Z(n5333) );
  MUX2_X1 U6281 ( .A(n6386), .B(n5085), .S(n5055), .Z(n5087) );
  MUX2_X1 U6282 ( .A(n5091), .B(n6012), .S(n4951), .Z(n5093) );
  MUX2_X1 U6283 ( .A(n5952), .B(n6037), .S(n4951), .Z(n5098) );
  MUX2_X1 U6284 ( .A(n6113), .B(n6112), .S(n4951), .Z(n5107) );
  MUX2_X1 U6285 ( .A(n6396), .B(n6281), .S(n4951), .Z(n5104) );
  MUX2_X1 U6286 ( .A(n6378), .B(n6376), .S(n4951), .Z(n5111) );
  MUX2_X1 U6287 ( .A(n6476), .B(n8891), .S(n4951), .Z(n5116) );
  MUX2_X1 U6288 ( .A(n6640), .B(n5119), .S(n4951), .Z(n5121) );
  MUX2_X1 U6289 ( .A(n6774), .B(n6772), .S(n4951), .Z(n5126) );
  MUX2_X1 U6290 ( .A(n5130), .B(n6875), .S(n4951), .Z(n5131) );
  MUX2_X1 U6291 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4951), .Z(n5136) );
  MUX2_X1 U6292 ( .A(n7047), .B(n8817), .S(n4951), .Z(n5138) );
  MUX2_X1 U6293 ( .A(n7284), .B(n7824), .S(n4951), .Z(n5142) );
  MUX2_X1 U6294 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4951), .Z(n5148) );
  MUX2_X1 U6295 ( .A(n8865), .B(n7861), .S(n4951), .Z(n5150) );
  MUX2_X1 U6296 ( .A(n5154), .B(n7881), .S(n4951), .Z(n5156) );
  MUX2_X1 U6297 ( .A(n8899), .B(n8783), .S(n4951), .Z(n5160) );
  MUX2_X1 U6298 ( .A(n7673), .B(n7915), .S(n4951), .Z(n5164) );
  MUX2_X1 U6299 ( .A(n9138), .B(n9969), .S(n4951), .Z(n5169) );
  MUX2_X1 U6300 ( .A(n9135), .B(n9967), .S(n4951), .Z(n5175) );
  MUX2_X1 U6301 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4951), .Z(n5617) );
  MUX2_X1 U6302 ( .A(n9127), .B(n9965), .S(n4951), .Z(n5629) );
  MUX2_X1 U6303 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4951), .Z(n5648) );
  MUX2_X1 U6304 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4951), .Z(n5651) );
  NAND3_X1 U6305 ( .A1(n4955), .A2(n4957), .A3(n8537), .ZN(n4953) );
  OR2_X1 U6306 ( .A1(n9066), .A2(n8558), .ZN(n4959) );
  OR2_X1 U6307 ( .A1(n7581), .A2(n8371), .ZN(n4969) );
  NAND2_X1 U6308 ( .A1(n8463), .A2(n4974), .ZN(n4973) );
  OAI21_X1 U6309 ( .B1(n9041), .B2(n4978), .A(n4972), .ZN(P2_U3517) );
  AND2_X2 U6310 ( .A1(n4977), .A2(n4979), .ZN(n4972) );
  OR2_X2 U6311 ( .A1(n4981), .A2(n10408), .ZN(n4977) );
  OR2_X1 U6312 ( .A1(n10409), .A2(n4980), .ZN(n4979) );
  NAND2_X1 U6313 ( .A1(n5305), .A2(n5304), .ZN(n5307) );
  NAND2_X1 U6314 ( .A1(n5307), .A2(n4544), .ZN(n4991) );
  NAND3_X1 U6315 ( .A1(n4991), .A2(n5327), .A3(n4990), .ZN(n5331) );
  NAND3_X1 U6316 ( .A1(n4995), .A2(n5805), .A3(n4993), .ZN(n7080) );
  NAND3_X1 U6317 ( .A1(n5000), .A2(n4999), .A3(n5694), .ZN(n10235) );
  NAND2_X1 U6318 ( .A1(n5332), .A2(n5001), .ZN(n5000) );
  OAI211_X2 U6319 ( .C1(n7398), .C2(n5006), .A(n7583), .B(n5004), .ZN(n7582)
         );
  NAND2_X1 U6320 ( .A1(n5013), .A2(n5014), .ZN(n5658) );
  NAND2_X1 U6321 ( .A1(n8124), .A2(n5015), .ZN(n5013) );
  NAND2_X1 U6322 ( .A1(n5046), .A2(n5045), .ZN(n5027) );
  NAND2_X1 U6323 ( .A1(n5045), .A2(n5263), .ZN(n5294) );
  INV_X1 U6324 ( .A(n5033), .ZN(n8475) );
  NAND2_X1 U6325 ( .A1(n5035), .A2(n5034), .ZN(n5220) );
  AND2_X1 U6326 ( .A1(n6576), .A2(n6141), .ZN(n10376) );
  NAND2_X1 U6327 ( .A1(n6149), .A2(n6148), .ZN(n6286) );
  NAND2_X1 U6328 ( .A1(n5850), .A2(n5849), .ZN(n5903) );
  INV_X1 U6329 ( .A(n5900), .ZN(n5850) );
  INV_X1 U6330 ( .A(n5903), .ZN(n5863) );
  INV_X1 U6331 ( .A(n7797), .ZN(n7800) );
  INV_X1 U6332 ( .A(n5942), .ZN(n8107) );
  INV_X1 U6333 ( .A(n6585), .ZN(n6846) );
  NAND2_X1 U6334 ( .A1(n6584), .A2(n6583), .ZN(n6847) );
  OR2_X1 U6335 ( .A1(n4482), .A2(n5236), .ZN(n5239) );
  INV_X1 U6336 ( .A(n4481), .ZN(n5643) );
  AOI21_X1 U6337 ( .B1(n8502), .B2(n5614), .A(n5602), .ZN(n8477) );
  NAND2_X1 U6338 ( .A1(n5614), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5238) );
  INV_X1 U6339 ( .A(n5614), .ZN(n5622) );
  INV_X1 U6340 ( .A(n8578), .ZN(n5549) );
  INV_X1 U6341 ( .A(n7100), .ZN(n7095) );
  OR2_X1 U6342 ( .A1(n8094), .A2(n5927), .ZN(n5039) );
  AND2_X1 U6343 ( .A1(n5096), .A2(n5095), .ZN(n5040) );
  AND2_X1 U6344 ( .A1(n5101), .A2(n5100), .ZN(n5041) );
  INV_X1 U6345 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5452) );
  INV_X1 U6346 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5056) );
  INV_X1 U6347 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5887) );
  AND2_X1 U6348 ( .A1(n5114), .A2(n5113), .ZN(n5042) );
  AOI21_X1 U6349 ( .B1(n8486), .B2(n5614), .A(n5613), .ZN(n8498) );
  INV_X1 U6350 ( .A(n9049), .ZN(n8116) );
  INV_X1 U6351 ( .A(n8609), .ZN(n5523) );
  INV_X1 U6352 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5186) );
  INV_X1 U6353 ( .A(n5516), .ZN(n5207) );
  INV_X1 U6354 ( .A(n7136), .ZN(n7133) );
  INV_X1 U6355 ( .A(n7786), .ZN(n6625) );
  INV_X1 U6356 ( .A(n7864), .ZN(n6627) );
  INV_X1 U6357 ( .A(n9665), .ZN(n9668) );
  INV_X1 U6358 ( .A(n7272), .ZN(n6388) );
  NOR2_X1 U6359 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5866) );
  INV_X1 U6360 ( .A(SI_22_), .ZN(n8867) );
  INV_X1 U6361 ( .A(SI_19_), .ZN(n5137) );
  INV_X1 U6362 ( .A(SI_15_), .ZN(n5120) );
  INV_X1 U6363 ( .A(SI_10_), .ZN(n8947) );
  INV_X1 U6364 ( .A(n5541), .ZN(n5208) );
  INV_X1 U6365 ( .A(n8308), .ZN(n8145) );
  AND2_X1 U6366 ( .A1(n6576), .A2(n6575), .ZN(n6289) );
  OR2_X1 U6367 ( .A1(n5596), .A2(n8353), .ZN(n5607) );
  INV_X1 U6368 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6369 ( .A1(n8116), .A2(n8498), .ZN(n8117) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7881) );
  AND2_X1 U6371 ( .A1(n6350), .A2(n6652), .ZN(n6440) );
  NAND2_X1 U6372 ( .A1(n6627), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7885) );
  INV_X1 U6373 ( .A(n9744), .ZN(n7975) );
  OR2_X1 U6374 ( .A1(n7719), .A2(n7718), .ZN(n7786) );
  NAND2_X1 U6375 ( .A1(n6623), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7570) );
  NAND2_X1 U6376 ( .A1(n6388), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7274) );
  OR2_X1 U6377 ( .A1(n6920), .A2(n6919), .ZN(n6922) );
  INV_X1 U6378 ( .A(n6412), .ZN(n6684) );
  NAND2_X1 U6379 ( .A1(n6719), .A2(n9301), .ZN(n6718) );
  INV_X1 U6380 ( .A(SI_28_), .ZN(n8951) );
  AND2_X1 U6381 ( .A1(n5923), .A2(n5922), .ZN(n5932) );
  OR2_X1 U6382 ( .A1(n8218), .A2(n8217), .ZN(n8219) );
  OR2_X1 U6383 ( .A1(n5412), .A2(n5203), .ZN(n5424) );
  INV_X1 U6384 ( .A(n8648), .ZN(n8278) );
  OR2_X1 U6385 ( .A1(n5555), .A2(n5554), .ZN(n5566) );
  NOR2_X1 U6386 ( .A1(n10309), .A2(n6289), .ZN(n9026) );
  OR2_X1 U6387 ( .A1(n5502), .A2(n8825), .ZN(n5516) );
  INV_X1 U6388 ( .A(n6038), .ZN(n6575) );
  INV_X1 U6389 ( .A(n8342), .ZN(n8355) );
  INV_X1 U6390 ( .A(n4483), .ZN(n5642) );
  AND2_X1 U6391 ( .A1(n6125), .A2(n6126), .ZN(n5843) );
  OR2_X1 U6392 ( .A1(n4483), .A2(n10225), .ZN(n5234) );
  INV_X1 U6393 ( .A(n7583), .ZN(n7676) );
  INV_X1 U6394 ( .A(n5800), .ZN(n10265) );
  INV_X1 U6395 ( .A(n10264), .ZN(n10281) );
  NAND2_X1 U6396 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5036), .ZN(n5193) );
  XNOR2_X1 U6397 ( .A(n6832), .B(n7947), .ZN(n6904) );
  INV_X1 U6398 ( .A(n7928), .ZN(n7943) );
  INV_X1 U6399 ( .A(n7353), .ZN(n7354) );
  INV_X1 U6400 ( .A(n4479), .ZN(n7887) );
  INV_X1 U6401 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7270) );
  OR2_X1 U6402 ( .A1(n7847), .A2(n7846), .ZN(n7864) );
  INV_X1 U6403 ( .A(n9549), .ZN(n9783) );
  INV_X1 U6404 ( .A(n9550), .ZN(n9784) );
  AND2_X1 U6405 ( .A1(n9473), .A2(n9480), .ZN(n9467) );
  INV_X1 U6406 ( .A(n10205), .ZN(n10146) );
  INV_X1 U6407 ( .A(n10137), .ZN(n9818) );
  OR2_X1 U6408 ( .A1(n6885), .A2(n10148), .ZN(n10143) );
  AND2_X1 U6409 ( .A1(n5159), .A2(n5158), .ZN(n5562) );
  INV_X1 U6410 ( .A(n9088), .ZN(n8605) );
  NOR2_X1 U6411 ( .A1(n8263), .A2(n10284), .ZN(n8318) );
  AND2_X1 U6412 ( .A1(n5843), .A2(n5842), .ZN(n6040) );
  INV_X1 U6413 ( .A(n10226), .ZN(n9986) );
  AND2_X1 U6414 ( .A1(n6075), .A2(n6074), .ZN(n10226) );
  INV_X1 U6415 ( .A(n5805), .ZN(n7082) );
  AND2_X1 U6416 ( .A1(n10299), .A2(n6598), .ZN(n10251) );
  NAND2_X1 U6417 ( .A1(n6591), .A2(n6590), .ZN(n10264) );
  NOR2_X1 U6418 ( .A1(n6124), .A2(n10320), .ZN(n9103) );
  OR2_X1 U6419 ( .A1(n6600), .A2(n10326), .ZN(n10402) );
  AND2_X1 U6420 ( .A1(n10241), .A2(n10380), .ZN(n10327) );
  INV_X1 U6421 ( .A(n10327), .ZN(n10407) );
  NAND2_X1 U6422 ( .A1(n6288), .A2(n10325), .ZN(n10309) );
  AND2_X1 U6423 ( .A1(n5448), .A2(n5438), .ZN(n6957) );
  INV_X1 U6424 ( .A(n9245), .ZN(n9236) );
  NAND2_X1 U6425 ( .A1(n6188), .A2(n10150), .ZN(n9251) );
  AND3_X1 U6426 ( .A1(n7851), .A2(n7850), .A3(n7849), .ZN(n9760) );
  AND4_X1 U6427 ( .A1(n7708), .A2(n7707), .A3(n7706), .A4(n7705), .ZN(n9817)
         );
  INV_X1 U6428 ( .A(n10106), .ZN(n10120) );
  INV_X1 U6429 ( .A(n9590), .ZN(n10124) );
  NAND2_X1 U6430 ( .A1(n9450), .A2(n9451), .ZN(n9613) );
  AND2_X1 U6431 ( .A1(n9418), .A2(n9296), .ZN(n9726) );
  NAND2_X1 U6432 ( .A1(n6677), .A2(n6676), .ZN(n10135) );
  INV_X1 U6433 ( .A(n10143), .ZN(n7615) );
  NOR2_X1 U6434 ( .A1(n10157), .A2(n10144), .ZN(n9834) );
  AND2_X1 U6435 ( .A1(n5956), .A2(n9467), .ZN(n10140) );
  NOR2_X1 U6436 ( .A1(n9956), .A2(n6520), .ZN(n6348) );
  OR2_X1 U6437 ( .A1(n9460), .A2(n9527), .ZN(n9999) );
  INV_X1 U6438 ( .A(n9999), .ZN(n10210) );
  OAI211_X1 U6439 ( .C1(P1_B_REG_SCAN_IN), .C2(n7613), .A(n5910), .B(n5909), 
        .ZN(n10158) );
  AND2_X1 U6440 ( .A1(n6481), .A2(n6483), .ZN(n7554) );
  INV_X1 U6441 ( .A(n8091), .ZN(n10231) );
  INV_X1 U6442 ( .A(n8110), .ZN(n10011) );
  INV_X1 U6443 ( .A(n8360), .ZN(n8338) );
  NAND2_X1 U6444 ( .A1(n6140), .A2(n6138), .ZN(n8362) );
  INV_X1 U6445 ( .A(n8478), .ZN(n8366) );
  NAND2_X1 U6446 ( .A1(n6040), .A2(n10325), .ZN(n8379) );
  NAND2_X1 U6447 ( .A1(n10299), .A2(n6599), .ZN(n8627) );
  NAND2_X1 U6448 ( .A1(n10299), .A2(n6612), .ZN(n8639) );
  INV_X1 U6449 ( .A(n10430), .ZN(n10427) );
  AND2_X1 U6450 ( .A1(n10393), .A2(n10392), .ZN(n10424) );
  AND3_X1 U6451 ( .A1(n10360), .A2(n10359), .A3(n10358), .ZN(n10418) );
  NOR2_X1 U6452 ( .A1(n10310), .A2(n10309), .ZN(n10319) );
  AND2_X1 U6453 ( .A1(n9141), .A2(n7611), .ZN(n10320) );
  NAND2_X1 U6454 ( .A1(n5838), .A2(n5837), .ZN(n7672) );
  INV_X1 U6455 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6774) );
  INV_X1 U6456 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6386) );
  CLKBUF_X1 U6457 ( .A(n9139), .Z(n9134) );
  INV_X1 U6458 ( .A(n6666), .ZN(n10147) );
  INV_X1 U6459 ( .A(n7489), .ZN(n10053) );
  NAND2_X1 U6460 ( .A1(n6207), .A2(n6206), .ZN(n9253) );
  AND2_X1 U6461 ( .A1(n6637), .A2(n6636), .ZN(n9616) );
  INV_X1 U6462 ( .A(n9760), .ZN(n9728) );
  OR2_X1 U6463 ( .A1(n9592), .A2(n6671), .ZN(n9595) );
  OR2_X1 U6464 ( .A1(P1_U3083), .A2(n5958), .ZN(n10063) );
  NAND2_X1 U6465 ( .A1(n5960), .A2(n5959), .ZN(n10106) );
  NAND2_X1 U6466 ( .A1(n9810), .A2(n6886), .ZN(n9813) );
  OR2_X1 U6467 ( .A1(n9937), .A2(n9936), .ZN(n9955) );
  INV_X1 U6468 ( .A(n10212), .ZN(n10211) );
  INV_X1 U6469 ( .A(n10168), .ZN(n10165) );
  AND2_X1 U6470 ( .A1(n6171), .A2(n6170), .ZN(n9957) );
  XNOR2_X1 U6471 ( .A(n5870), .B(n5869), .ZN(n7674) );
  INV_X1 U6472 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6772) );
  INV_X1 U6473 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6112) );
  NOR2_X1 U6474 ( .A1(n10460), .A2(n10459), .ZN(n10458) );
  OAI21_X1 U6475 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10449), .ZN(n10447) );
  INV_X1 U6476 ( .A(n8379), .ZN(P2_U3966) );
  NOR2_X1 U6477 ( .A1(n5957), .A2(P1_U3084), .ZN(P1_U4006) );
  NOR2_X1 U6478 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5046) );
  MUX2_X1 U6479 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5055), .Z(n5050) );
  NAND2_X1 U6480 ( .A1(n5050), .A2(SI_2_), .ZN(n5062) );
  OAI21_X1 U6481 ( .B1(n5050), .B2(SI_2_), .A(n5062), .ZN(n5260) );
  INV_X1 U6482 ( .A(n5260), .ZN(n5061) );
  INV_X1 U6483 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6190) );
  INV_X1 U6484 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5051) );
  INV_X1 U6485 ( .A(SI_0_), .ZN(n6189) );
  NAND2_X1 U6486 ( .A1(n5054), .A2(SI_1_), .ZN(n5059) );
  NAND2_X1 U6487 ( .A1(n5261), .A2(n5062), .ZN(n5276) );
  NAND2_X1 U6488 ( .A1(n5063), .A2(SI_3_), .ZN(n5067) );
  INV_X1 U6489 ( .A(n5063), .ZN(n5065) );
  INV_X1 U6490 ( .A(SI_3_), .ZN(n5064) );
  NAND2_X1 U6491 ( .A1(n5065), .A2(n5064), .ZN(n5066) );
  AND2_X1 U6492 ( .A1(n5067), .A2(n5066), .ZN(n5275) );
  NAND2_X1 U6493 ( .A1(n5276), .A2(n5275), .ZN(n5278) );
  NAND2_X1 U6494 ( .A1(n5068), .A2(SI_4_), .ZN(n5072) );
  INV_X1 U6495 ( .A(n5068), .ZN(n5070) );
  INV_X1 U6496 ( .A(SI_4_), .ZN(n5069) );
  NAND2_X1 U6497 ( .A1(n5070), .A2(n5069), .ZN(n5071) );
  AND2_X1 U6498 ( .A1(n5072), .A2(n5071), .ZN(n5290) );
  NAND2_X1 U6499 ( .A1(n5073), .A2(SI_5_), .ZN(n5077) );
  INV_X1 U6500 ( .A(n5073), .ZN(n5075) );
  INV_X1 U6501 ( .A(SI_5_), .ZN(n5074) );
  NAND2_X1 U6502 ( .A1(n5075), .A2(n5074), .ZN(n5076) );
  NAND2_X1 U6503 ( .A1(n5078), .A2(SI_6_), .ZN(n5082) );
  INV_X1 U6504 ( .A(n5078), .ZN(n5080) );
  INV_X1 U6505 ( .A(SI_6_), .ZN(n5079) );
  NAND2_X1 U6506 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  NAND2_X1 U6507 ( .A1(n5335), .A2(SI_7_), .ZN(n5083) );
  NAND2_X1 U6508 ( .A1(n5084), .A2(n5083), .ZN(n5347) );
  INV_X1 U6509 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5085) );
  INV_X1 U6510 ( .A(SI_8_), .ZN(n5086) );
  NAND2_X1 U6511 ( .A1(n5087), .A2(n5086), .ZN(n5090) );
  INV_X1 U6512 ( .A(n5087), .ZN(n5088) );
  NAND2_X1 U6513 ( .A1(n5088), .A2(SI_8_), .ZN(n5089) );
  NAND2_X1 U6514 ( .A1(n5090), .A2(n5089), .ZN(n5346) );
  OAI21_X2 U6515 ( .B1(n5347), .B2(n5346), .A(n5090), .ZN(n5359) );
  INV_X1 U6516 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5091) );
  INV_X1 U6517 ( .A(SI_9_), .ZN(n5092) );
  NAND2_X1 U6518 ( .A1(n5093), .A2(n5092), .ZN(n5096) );
  INV_X1 U6519 ( .A(n5093), .ZN(n5094) );
  NAND2_X1 U6520 ( .A1(n5094), .A2(SI_9_), .ZN(n5095) );
  NAND2_X1 U6521 ( .A1(n5359), .A2(n5040), .ZN(n5097) );
  NAND2_X1 U6522 ( .A1(n5098), .A2(n8947), .ZN(n5101) );
  INV_X1 U6523 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6524 ( .A1(n5099), .A2(SI_10_), .ZN(n5100) );
  XNOR2_X1 U6525 ( .A(n5107), .B(SI_11_), .ZN(n5391) );
  INV_X1 U6526 ( .A(SI_12_), .ZN(n5103) );
  NAND2_X1 U6527 ( .A1(n5104), .A2(n5103), .ZN(n5110) );
  INV_X1 U6528 ( .A(n5104), .ZN(n5105) );
  NAND2_X1 U6529 ( .A1(n5105), .A2(SI_12_), .ZN(n5106) );
  NAND2_X1 U6530 ( .A1(n5110), .A2(n5106), .ZN(n5405) );
  INV_X1 U6531 ( .A(n5405), .ZN(n5109) );
  INV_X1 U6532 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6533 ( .A1(n5108), .A2(SI_11_), .ZN(n5403) );
  NAND2_X1 U6534 ( .A1(n5111), .A2(n8915), .ZN(n5114) );
  INV_X1 U6535 ( .A(n5111), .ZN(n5112) );
  NAND2_X1 U6536 ( .A1(n5112), .A2(SI_13_), .ZN(n5113) );
  XNOR2_X1 U6537 ( .A(n5116), .B(SI_14_), .ZN(n5432) );
  INV_X1 U6538 ( .A(n5432), .ZN(n5115) );
  INV_X1 U6539 ( .A(n5116), .ZN(n5117) );
  NAND2_X1 U6540 ( .A1(n5117), .A2(SI_14_), .ZN(n5118) );
  NAND2_X1 U6541 ( .A1(n5121), .A2(n5120), .ZN(n5124) );
  INV_X1 U6542 ( .A(n5121), .ZN(n5122) );
  NAND2_X1 U6543 ( .A1(n5122), .A2(SI_15_), .ZN(n5123) );
  NAND2_X1 U6544 ( .A1(n5124), .A2(n5123), .ZN(n5446) );
  NAND2_X1 U6545 ( .A1(n5126), .A2(n5125), .ZN(n5129) );
  INV_X1 U6546 ( .A(n5126), .ZN(n5127) );
  NAND2_X1 U6547 ( .A1(n5127), .A2(SI_16_), .ZN(n5128) );
  XNOR2_X1 U6548 ( .A(n5131), .B(SI_17_), .ZN(n5477) );
  INV_X1 U6549 ( .A(n5477), .ZN(n5134) );
  INV_X1 U6550 ( .A(n5131), .ZN(n5132) );
  NAND2_X1 U6551 ( .A1(n5132), .A2(SI_17_), .ZN(n5133) );
  XNOR2_X1 U6552 ( .A(n5136), .B(SI_18_), .ZN(n5496) );
  INV_X1 U6553 ( .A(n5496), .ZN(n5135) );
  NAND2_X1 U6554 ( .A1(n5138), .A2(n5137), .ZN(n5141) );
  INV_X1 U6555 ( .A(n5138), .ZN(n5139) );
  NAND2_X1 U6556 ( .A1(n5139), .A2(SI_19_), .ZN(n5140) );
  NAND2_X1 U6557 ( .A1(n5141), .A2(n5140), .ZN(n5510) );
  INV_X1 U6558 ( .A(SI_20_), .ZN(n8828) );
  NAND2_X1 U6559 ( .A1(n5142), .A2(n8828), .ZN(n5145) );
  INV_X1 U6560 ( .A(n5142), .ZN(n5143) );
  NAND2_X1 U6561 ( .A1(n5143), .A2(SI_20_), .ZN(n5144) );
  NAND2_X1 U6562 ( .A1(n5525), .A2(n5524), .ZN(n5146) );
  INV_X1 U6563 ( .A(SI_21_), .ZN(n5147) );
  XNOR2_X1 U6564 ( .A(n5148), .B(n5147), .ZN(n5536) );
  NAND2_X1 U6565 ( .A1(n5148), .A2(SI_21_), .ZN(n5149) );
  NAND2_X1 U6566 ( .A1(n5150), .A2(n8867), .ZN(n5153) );
  INV_X1 U6567 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6568 ( .A1(n5151), .A2(SI_22_), .ZN(n5152) );
  NAND2_X1 U6569 ( .A1(n5153), .A2(n5152), .ZN(n5550) );
  INV_X1 U6570 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5154) );
  INV_X1 U6571 ( .A(SI_23_), .ZN(n5155) );
  NAND2_X1 U6572 ( .A1(n5156), .A2(n5155), .ZN(n5159) );
  INV_X1 U6573 ( .A(n5156), .ZN(n5157) );
  NAND2_X1 U6574 ( .A1(n5157), .A2(SI_23_), .ZN(n5158) );
  XNOR2_X1 U6575 ( .A(n5160), .B(SI_24_), .ZN(n5572) );
  INV_X1 U6576 ( .A(n5572), .ZN(n5162) );
  INV_X1 U6577 ( .A(n5160), .ZN(n5161) );
  INV_X1 U6578 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7673) );
  INV_X1 U6579 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7915) );
  INV_X1 U6580 ( .A(SI_25_), .ZN(n5163) );
  NAND2_X1 U6581 ( .A1(n5164), .A2(n5163), .ZN(n5167) );
  INV_X1 U6582 ( .A(n5164), .ZN(n5165) );
  NAND2_X1 U6583 ( .A1(n5165), .A2(SI_25_), .ZN(n5166) );
  NAND2_X1 U6584 ( .A1(n5167), .A2(n5166), .ZN(n5583) );
  INV_X1 U6585 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9138) );
  INV_X1 U6586 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9969) );
  INV_X1 U6587 ( .A(SI_26_), .ZN(n5168) );
  NAND2_X1 U6588 ( .A1(n5169), .A2(n5168), .ZN(n5172) );
  INV_X1 U6589 ( .A(n5169), .ZN(n5170) );
  NAND2_X1 U6590 ( .A1(n5170), .A2(SI_26_), .ZN(n5171) );
  NAND2_X1 U6591 ( .A1(n5593), .A2(n5592), .ZN(n5173) );
  NAND2_X1 U6592 ( .A1(n5173), .A2(n5172), .ZN(n5604) );
  INV_X1 U6593 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9135) );
  INV_X1 U6594 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9967) );
  INV_X1 U6595 ( .A(SI_27_), .ZN(n5174) );
  NAND2_X1 U6596 ( .A1(n5175), .A2(n5174), .ZN(n5178) );
  INV_X1 U6597 ( .A(n5175), .ZN(n5176) );
  NAND2_X1 U6598 ( .A1(n5176), .A2(SI_27_), .ZN(n5177) );
  XNOR2_X1 U6599 ( .A(n5617), .B(n8951), .ZN(n5615) );
  NAND4_X1 U6600 ( .A1(n5659), .A2(n5182), .A3(n4876), .A4(n5181), .ZN(n5183)
         );
  NOR2_X2 U6601 ( .A1(n5184), .A2(n5183), .ZN(n5185) );
  NAND4_X1 U6602 ( .A1(n5187), .A2(n5840), .A3(n5831), .A4(n5186), .ZN(n5189)
         );
  NAND2_X1 U6603 ( .A1(n5828), .A2(n5827), .ZN(n5188) );
  NAND2_X1 U6604 ( .A1(n8004), .A2(n4990), .ZN(n5197) );
  NAND2_X1 U6605 ( .A1(n4475), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6606 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5296) );
  INV_X1 U6607 ( .A(n5296), .ZN(n5198) );
  NAND2_X1 U6608 ( .A1(n5198), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5315) );
  INV_X1 U6609 ( .A(n5315), .ZN(n5199) );
  NAND2_X1 U6610 ( .A1(n5199), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5339) );
  INV_X1 U6611 ( .A(n5339), .ZN(n5200) );
  NAND2_X1 U6612 ( .A1(n5200), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6613 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5201) );
  INV_X1 U6614 ( .A(n5384), .ZN(n5202) );
  NAND2_X1 U6615 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5203) );
  INV_X1 U6616 ( .A(n5424), .ZN(n5204) );
  INV_X1 U6617 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5453) );
  INV_X1 U6618 ( .A(n5468), .ZN(n5205) );
  NAND2_X1 U6619 ( .A1(n5205), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5486) );
  INV_X1 U6620 ( .A(n5486), .ZN(n5206) );
  NAND2_X1 U6621 ( .A1(n5206), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5502) );
  INV_X1 U6622 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5528) );
  INV_X1 U6623 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5554) );
  INV_X1 U6624 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8178) );
  INV_X1 U6625 ( .A(n5577), .ZN(n5209) );
  NAND2_X1 U6626 ( .A1(n5209), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5587) );
  INV_X1 U6627 ( .A(n5587), .ZN(n5210) );
  NAND2_X1 U6628 ( .A1(n5210), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5596) );
  INV_X1 U6629 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8353) );
  INV_X1 U6630 ( .A(n5607), .ZN(n5212) );
  AND2_X1 U6631 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5211) );
  NAND2_X1 U6632 ( .A1(n5212), .A2(n5211), .ZN(n8118) );
  INV_X1 U6633 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8169) );
  INV_X1 U6634 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5213) );
  OAI21_X1 U6635 ( .B1(n5607), .B2(n8169), .A(n5213), .ZN(n5214) );
  NAND2_X1 U6636 ( .A1(n8118), .A2(n5214), .ZN(n8222) );
  NAND2_X1 U6637 ( .A1(n5218), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5219) );
  AND2_X4 U6638 ( .A1(n9122), .A2(n5222), .ZN(n5614) );
  INV_X1 U6639 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6640 ( .A1(n5643), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6641 ( .A1(n5642), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5224) );
  OAI211_X1 U6642 ( .C1(n4484), .C2(n5226), .A(n5225), .B(n5224), .ZN(n5227)
         );
  INV_X1 U6643 ( .A(n5227), .ZN(n5228) );
  INV_X1 U6644 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10225) );
  NAND2_X1 U6645 ( .A1(n5608), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6646 ( .A1(n5614), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5232) );
  INV_X1 U6647 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5230) );
  OR2_X1 U6648 ( .A1(n5598), .A2(n5230), .ZN(n5231) );
  NAND2_X1 U6649 ( .A1(n6417), .A2(SI_0_), .ZN(n5235) );
  XNOR2_X1 U6650 ( .A(n5235), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9142) );
  MUX2_X1 U6651 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9142), .S(n5247), .Z(n6661) );
  NAND2_X1 U6652 ( .A1(n4508), .A2(n6661), .ZN(n6607) );
  INV_X1 U6653 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6617) );
  INV_X1 U6654 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6655 ( .A1(n5608), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5237) );
  NAND4_X2 U6656 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n6578)
         );
  INV_X1 U6657 ( .A(n6578), .ZN(n6659) );
  INV_X1 U6658 ( .A(n5241), .ZN(n5244) );
  INV_X1 U6659 ( .A(n5242), .ZN(n5243) );
  NAND2_X1 U6660 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  NAND2_X1 U6661 ( .A1(n5246), .A2(n5245), .ZN(n6416) );
  NAND2_X1 U6662 ( .A1(n5279), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6663 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5248) );
  INV_X1 U6664 ( .A(n5263), .ZN(n5249) );
  INV_X1 U6665 ( .A(n6062), .ZN(n9979) );
  NAND2_X1 U6666 ( .A1(n5512), .A2(n9979), .ZN(n5251) );
  NAND2_X1 U6667 ( .A1(n6659), .A2(n6613), .ZN(n5796) );
  NAND2_X1 U6668 ( .A1(n6607), .A2(n5796), .ZN(n5253) );
  NAND2_X1 U6669 ( .A1(n5253), .A2(n5795), .ZN(n5674) );
  INV_X1 U6670 ( .A(n5674), .ZN(n5268) );
  INV_X1 U6671 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5254) );
  INV_X1 U6672 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5255) );
  OR2_X1 U6673 ( .A1(n4481), .A2(n5255), .ZN(n5258) );
  NAND2_X1 U6674 ( .A1(n5608), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6675 ( .A1(n5614), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5256) );
  INV_X1 U6676 ( .A(n8382), .ZN(n6586) );
  NAND2_X1 U6677 ( .A1(n5262), .A2(n5261), .ZN(n6446) );
  NAND2_X1 U6678 ( .A1(n5279), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6679 ( .A1(n5263), .A2(n5479), .ZN(n5264) );
  XNOR2_X1 U6680 ( .A(n5264), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U6681 ( .A1(n5512), .A2(n9991), .ZN(n5265) );
  OAI211_X1 U6682 ( .C1(n5329), .C2(n6446), .A(n5266), .B(n5265), .ZN(n6865)
         );
  NAND2_X1 U6683 ( .A1(n8382), .A2(n10338), .ZN(n5683) );
  INV_X1 U6684 ( .A(n6582), .ZN(n5267) );
  NAND2_X1 U6685 ( .A1(n5268), .A2(n5267), .ZN(n6587) );
  NAND2_X1 U6686 ( .A1(n6587), .A2(n6588), .ZN(n5282) );
  NAND2_X1 U6687 ( .A1(n5614), .A2(n6294), .ZN(n5274) );
  NAND2_X1 U6688 ( .A1(n5608), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5273) );
  INV_X1 U6689 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5269) );
  INV_X1 U6690 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5270) );
  OR2_X1 U6691 ( .A1(n4481), .A2(n5270), .ZN(n5271) );
  OR2_X1 U6692 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  NAND2_X1 U6693 ( .A1(n5278), .A2(n5277), .ZN(n6505) );
  OR3_X1 U6694 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_IR_REG_1__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6695 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5280), .ZN(n5281) );
  XNOR2_X1 U6696 ( .A(n5281), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U6697 ( .A1(n10287), .A2(n10292), .ZN(n10278) );
  NAND2_X1 U6698 ( .A1(n4485), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5289) );
  OAI21_X1 U6699 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5296), .ZN(n10298) );
  INV_X1 U6700 ( .A(n10298), .ZN(n5283) );
  NAND2_X1 U6701 ( .A1(n5614), .A2(n5283), .ZN(n5288) );
  INV_X1 U6702 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5284) );
  OR2_X1 U6703 ( .A1(n4481), .A2(n5284), .ZN(n5287) );
  INV_X1 U6704 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5285) );
  OR2_X1 U6705 ( .A1(n4483), .A2(n5285), .ZN(n5286) );
  NAND4_X1 U6706 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n8380)
         );
  INV_X1 U6707 ( .A(n8380), .ZN(n6850) );
  OR2_X1 U6708 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  NAND2_X1 U6709 ( .A1(n5294), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5308) );
  XNOR2_X1 U6710 ( .A(n5308), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U6711 ( .A1(n5512), .A2(n6066), .ZN(n5295) );
  NAND2_X1 U6712 ( .A1(n6850), .A2(n10301), .ZN(n5794) );
  AND2_X1 U6713 ( .A1(n10278), .A2(n5794), .ZN(n5672) );
  NAND2_X1 U6714 ( .A1(n4485), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5303) );
  INV_X1 U6715 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U6716 ( .A1(n5296), .A2(n6247), .ZN(n5297) );
  AND2_X1 U6717 ( .A1(n5315), .A2(n5297), .ZN(n8288) );
  NAND2_X1 U6718 ( .A1(n5614), .A2(n8288), .ZN(n5302) );
  INV_X1 U6719 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5298) );
  OR2_X1 U6720 ( .A1(n4481), .A2(n5298), .ZN(n5301) );
  INV_X1 U6721 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5299) );
  OR2_X1 U6722 ( .A1(n4483), .A2(n5299), .ZN(n5300) );
  NAND4_X1 U6723 ( .A1(n5303), .A2(n5302), .A3(n5301), .A4(n5300), .ZN(n10260)
         );
  OR2_X1 U6724 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  AND2_X1 U6725 ( .A1(n5307), .A2(n5306), .ZN(n6793) );
  NAND2_X1 U6726 ( .A1(n4990), .A2(n6793), .ZN(n5313) );
  NAND2_X1 U6727 ( .A1(n4475), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6728 ( .A1(n5308), .A2(n5324), .ZN(n5309) );
  NAND2_X1 U6729 ( .A1(n5309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5310) );
  XNOR2_X1 U6730 ( .A(n5310), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U6731 ( .A1(n5512), .A2(n6068), .ZN(n5311) );
  NAND2_X1 U6732 ( .A1(n10260), .A2(n10355), .ZN(n5793) );
  AND2_X1 U6733 ( .A1(n10282), .A2(n5793), .ZN(n5687) );
  INV_X1 U6734 ( .A(n10260), .ZN(n10285) );
  NAND2_X1 U6735 ( .A1(n10285), .A2(n8289), .ZN(n10256) );
  NAND2_X1 U6736 ( .A1(n4485), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5322) );
  INV_X1 U6737 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6738 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  AND2_X1 U6739 ( .A1(n5339), .A2(n5316), .ZN(n10268) );
  NAND2_X1 U6740 ( .A1(n5614), .A2(n10268), .ZN(n5321) );
  INV_X1 U6741 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5317) );
  OR2_X1 U6742 ( .A1(n4482), .A2(n5317), .ZN(n5320) );
  INV_X1 U6743 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5318) );
  OR2_X1 U6744 ( .A1(n4483), .A2(n5318), .ZN(n5319) );
  NAND4_X1 U6745 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n8378)
         );
  INV_X1 U6746 ( .A(n8378), .ZN(n6938) );
  INV_X1 U6747 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6748 ( .A1(n5324), .A2(n5323), .ZN(n5325) );
  NAND2_X1 U6749 ( .A1(n4531), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5326) );
  XNOR2_X1 U6750 ( .A(n5326), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6070) );
  INV_X1 U6751 ( .A(n6070), .ZN(n6265) );
  NAND2_X1 U6752 ( .A1(n4475), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5330) );
  OAI211_X1 U6753 ( .C1(n5247), .C2(n6265), .A(n5331), .B(n5330), .ZN(n10271)
         );
  NAND2_X1 U6754 ( .A1(n6938), .A2(n10271), .ZN(n5693) );
  INV_X1 U6755 ( .A(n10271), .ZN(n10361) );
  NAND2_X1 U6756 ( .A1(n8378), .A2(n10361), .ZN(n5689) );
  XNOR2_X1 U6757 ( .A(n5333), .B(SI_7_), .ZN(n5334) );
  XNOR2_X1 U6758 ( .A(n5335), .B(n5334), .ZN(n6814) );
  NAND2_X1 U6759 ( .A1(n6814), .A2(n4990), .ZN(n5338) );
  OR2_X1 U6760 ( .A1(n4501), .A2(n5479), .ZN(n5336) );
  XNOR2_X1 U6761 ( .A(n5336), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6071) );
  AOI22_X1 U6762 ( .A1(n4475), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5512), .B2(
        n6071), .ZN(n5337) );
  NAND2_X1 U6763 ( .A1(n4485), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5345) );
  INV_X1 U6764 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U6765 ( .A1(n5339), .A2(n6764), .ZN(n5340) );
  AND2_X1 U6766 ( .A1(n5366), .A2(n5340), .ZN(n9008) );
  NAND2_X1 U6767 ( .A1(n5614), .A2(n9008), .ZN(n5344) );
  INV_X1 U6768 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5341) );
  OR2_X1 U6769 ( .A1(n4482), .A2(n5341), .ZN(n5343) );
  INV_X1 U6770 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9010) );
  OR2_X1 U6771 ( .A1(n4483), .A2(n9010), .ZN(n5342) );
  NAND4_X1 U6772 ( .A1(n5345), .A2(n5344), .A3(n5343), .A4(n5342), .ZN(n10262)
         );
  NAND2_X1 U6773 ( .A1(n10367), .A2(n10262), .ZN(n5695) );
  INV_X1 U6774 ( .A(n10262), .ZN(n8339) );
  NAND2_X1 U6775 ( .A1(n8339), .A2(n9012), .ZN(n5694) );
  XNOR2_X1 U6776 ( .A(n5346), .B(n5347), .ZN(n5930) );
  NAND2_X1 U6777 ( .A1(n5930), .A2(n4990), .ZN(n5352) );
  AND2_X1 U6778 ( .A1(n5348), .A2(n4501), .ZN(n5349) );
  OR2_X1 U6779 ( .A1(n5349), .A2(n5479), .ZN(n5350) );
  XNOR2_X1 U6780 ( .A(n5350), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6334) );
  AOI22_X1 U6781 ( .A1(n4475), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5512), .B2(
        n6334), .ZN(n5351) );
  NAND2_X1 U6782 ( .A1(n4485), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5357) );
  XNOR2_X1 U6783 ( .A(n5366), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n10244) );
  NAND2_X1 U6784 ( .A1(n5614), .A2(n10244), .ZN(n5356) );
  INV_X1 U6785 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5353) );
  OR2_X1 U6786 ( .A1(n4481), .A2(n5353), .ZN(n5355) );
  INV_X1 U6787 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6061) );
  OR2_X1 U6788 ( .A1(n4483), .A2(n6061), .ZN(n5354) );
  NAND4_X1 U6789 ( .A1(n5357), .A2(n5356), .A3(n5355), .A4(n5354), .ZN(n8377)
         );
  XNOR2_X1 U6790 ( .A(n10375), .B(n8377), .ZN(n10236) );
  NAND2_X1 U6791 ( .A1(n10235), .A2(n10236), .ZN(n5358) );
  INV_X1 U6792 ( .A(n8377), .ZN(n5699) );
  NAND2_X1 U6793 ( .A1(n10375), .A2(n5699), .ZN(n5698) );
  NAND2_X1 U6794 ( .A1(n5358), .A2(n5698), .ZN(n6933) );
  XNOR2_X1 U6795 ( .A(n5359), .B(n5040), .ZN(n7115) );
  NAND2_X1 U6796 ( .A1(n7115), .A2(n4990), .ZN(n5364) );
  NAND2_X1 U6797 ( .A1(n4501), .A2(n5360), .ZN(n5361) );
  NAND2_X1 U6798 ( .A1(n5361), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5362) );
  XNOR2_X1 U6799 ( .A(n5362), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8384) );
  AOI22_X1 U6800 ( .A1(n4475), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5512), .B2(
        n8384), .ZN(n5363) );
  NAND2_X1 U6801 ( .A1(n5364), .A2(n5363), .ZN(n7167) );
  NAND2_X1 U6802 ( .A1(n4485), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5373) );
  INV_X1 U6803 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8235) );
  INV_X1 U6804 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5365) );
  OAI21_X1 U6805 ( .B1(n5366), .B2(n8235), .A(n5365), .ZN(n5367) );
  AND2_X1 U6806 ( .A1(n5367), .A2(n5384), .ZN(n7160) );
  NAND2_X1 U6807 ( .A1(n5614), .A2(n7160), .ZN(n5372) );
  INV_X1 U6808 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5368) );
  OR2_X1 U6809 ( .A1(n4482), .A2(n5368), .ZN(n5371) );
  INV_X1 U6810 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5369) );
  OR2_X1 U6811 ( .A1(n4483), .A2(n5369), .ZN(n5370) );
  NAND4_X1 U6812 ( .A1(n5373), .A2(n5372), .A3(n5371), .A4(n5370), .ZN(n8376)
         );
  INV_X1 U6813 ( .A(n8376), .ZN(n7164) );
  OR2_X1 U6814 ( .A1(n7167), .A2(n7164), .ZN(n5799) );
  NAND2_X1 U6815 ( .A1(n6933), .A2(n5799), .ZN(n5374) );
  NAND2_X1 U6816 ( .A1(n7167), .A2(n7164), .ZN(n5798) );
  XNOR2_X1 U6817 ( .A(n5375), .B(n5041), .ZN(n7257) );
  NAND2_X1 U6818 ( .A1(n7257), .A2(n4990), .ZN(n5383) );
  NAND2_X1 U6819 ( .A1(n4501), .A2(n5376), .ZN(n5377) );
  NAND2_X1 U6820 ( .A1(n5377), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5378) );
  MUX2_X1 U6821 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5378), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5381) );
  INV_X1 U6822 ( .A(n5379), .ZN(n5380) );
  AOI22_X1 U6823 ( .A1(n4475), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5512), .B2(
        n8396), .ZN(n5382) );
  NAND2_X1 U6824 ( .A1(n5383), .A2(n5382), .ZN(n8189) );
  NAND2_X1 U6825 ( .A1(n4485), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5390) );
  INV_X1 U6826 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U6827 ( .A1(n5384), .A2(n8830), .ZN(n5385) );
  AND2_X1 U6828 ( .A1(n5412), .A2(n5385), .ZN(n8188) );
  NAND2_X1 U6829 ( .A1(n5614), .A2(n8188), .ZN(n5389) );
  INV_X1 U6830 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5386) );
  OR2_X1 U6831 ( .A1(n4482), .A2(n5386), .ZN(n5388) );
  INV_X1 U6832 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6339) );
  OR2_X1 U6833 ( .A1(n4483), .A2(n6339), .ZN(n5387) );
  NAND4_X1 U6834 ( .A1(n5390), .A2(n5389), .A3(n5388), .A4(n5387), .ZN(n8375)
         );
  OR2_X1 U6835 ( .A1(n8189), .A2(n7185), .ZN(n5708) );
  NAND2_X1 U6836 ( .A1(n8189), .A2(n7185), .ZN(n7081) );
  XNOR2_X1 U6837 ( .A(n5392), .B(n5391), .ZN(n7339) );
  NAND2_X1 U6838 ( .A1(n7339), .A2(n4990), .ZN(n5397) );
  NOR2_X1 U6839 ( .A1(n5379), .A2(n5479), .ZN(n5393) );
  MUX2_X1 U6840 ( .A(n5479), .B(n5393), .S(P2_IR_REG_11__SCAN_IN), .Z(n5395)
         );
  OR2_X1 U6841 ( .A1(n5395), .A2(n5394), .ZN(n6486) );
  INV_X1 U6842 ( .A(n6486), .ZN(n6496) );
  AOI22_X1 U6843 ( .A1(n4475), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5512), .B2(
        n6496), .ZN(n5396) );
  NAND2_X1 U6844 ( .A1(n4485), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5402) );
  XNOR2_X1 U6845 ( .A(n5412), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n7188) );
  NAND2_X1 U6846 ( .A1(n5614), .A2(n7188), .ZN(n5401) );
  INV_X1 U6847 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5398) );
  OR2_X1 U6848 ( .A1(n4481), .A2(n5398), .ZN(n5400) );
  INV_X1 U6849 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7087) );
  OR2_X1 U6850 ( .A1(n4483), .A2(n7087), .ZN(n5399) );
  NAND4_X1 U6851 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n8374)
         );
  INV_X1 U6852 ( .A(n8374), .ZN(n7314) );
  OR2_X1 U6853 ( .A1(n7227), .A2(n7314), .ZN(n5715) );
  NAND2_X1 U6854 ( .A1(n7227), .A2(n7314), .ZN(n7217) );
  NAND2_X1 U6855 ( .A1(n5404), .A2(n5403), .ZN(n5406) );
  XNOR2_X1 U6856 ( .A(n5406), .B(n5405), .ZN(n7455) );
  NAND2_X1 U6857 ( .A1(n7455), .A2(n4990), .ZN(n5409) );
  OR2_X1 U6858 ( .A1(n5394), .A2(n5479), .ZN(n5407) );
  XNOR2_X1 U6859 ( .A(n5407), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6497) );
  AOI22_X1 U6860 ( .A1(n4475), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5512), .B2(
        n6497), .ZN(n5408) );
  NAND2_X1 U6861 ( .A1(n4485), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5418) );
  INV_X1 U6862 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5411) );
  INV_X1 U6863 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5410) );
  OAI21_X1 U6864 ( .B1(n5412), .B2(n5411), .A(n5410), .ZN(n5413) );
  AND2_X1 U6865 ( .A1(n5413), .A2(n5424), .ZN(n7316) );
  NAND2_X1 U6866 ( .A1(n5614), .A2(n7316), .ZN(n5417) );
  INV_X1 U6867 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5414) );
  OR2_X1 U6868 ( .A1(n4482), .A2(n5414), .ZN(n5416) );
  INV_X1 U6869 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6489) );
  OR2_X1 U6870 ( .A1(n4483), .A2(n6489), .ZN(n5415) );
  NAND4_X1 U6871 ( .A1(n5418), .A2(n5417), .A3(n5416), .A4(n5415), .ZN(n8373)
         );
  NAND2_X1 U6872 ( .A1(n7393), .A2(n7374), .ZN(n5803) );
  AND2_X1 U6873 ( .A1(n5803), .A2(n7217), .ZN(n5714) );
  NAND2_X1 U6874 ( .A1(n7080), .A2(n5714), .ZN(n5419) );
  NAND2_X1 U6875 ( .A1(n5419), .A2(n5804), .ZN(n7398) );
  XNOR2_X1 U6876 ( .A(n5420), .B(n5042), .ZN(n7522) );
  NAND2_X1 U6877 ( .A1(n7522), .A2(n4990), .ZN(n5423) );
  NAND2_X1 U6878 ( .A1(n5421), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5434) );
  XNOR2_X1 U6879 ( .A(n5434), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6692) );
  AOI22_X1 U6880 ( .A1(n4475), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5512), .B2(
        n6692), .ZN(n5422) );
  NAND2_X1 U6881 ( .A1(n4485), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5431) );
  INV_X1 U6882 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U6883 ( .A1(n5424), .A2(n8917), .ZN(n5425) );
  AND2_X1 U6884 ( .A1(n5454), .A2(n5425), .ZN(n7406) );
  NAND2_X1 U6885 ( .A1(n5614), .A2(n7406), .ZN(n5430) );
  INV_X1 U6886 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n5426) );
  OR2_X1 U6887 ( .A1(n4481), .A2(n5426), .ZN(n5429) );
  INV_X1 U6888 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5427) );
  OR2_X1 U6889 ( .A1(n4483), .A2(n5427), .ZN(n5428) );
  NAND4_X1 U6890 ( .A1(n5431), .A2(n5430), .A3(n5429), .A4(n5428), .ZN(n8372)
         );
  INV_X1 U6891 ( .A(n8372), .ZN(n7503) );
  OR2_X1 U6892 ( .A1(n7435), .A2(n7503), .ZN(n5722) );
  NAND2_X1 U6893 ( .A1(n7435), .A2(n7503), .ZN(n5723) );
  NAND2_X1 U6894 ( .A1(n5722), .A2(n5723), .ZN(n7399) );
  NAND2_X1 U6895 ( .A1(n7553), .A2(n4990), .ZN(n5440) );
  NAND2_X1 U6896 ( .A1(n5434), .A2(n4850), .ZN(n5435) );
  NAND2_X1 U6897 ( .A1(n5435), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6898 ( .A1(n5437), .A2(n5436), .ZN(n5448) );
  OR2_X1 U6899 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  AOI22_X1 U6900 ( .A1(n4475), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5512), .B2(
        n6957), .ZN(n5439) );
  NAND2_X1 U6901 ( .A1(n4485), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5445) );
  XNOR2_X1 U6902 ( .A(n5454), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U6903 ( .A1(n5614), .A2(n7442), .ZN(n5444) );
  INV_X1 U6904 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5441) );
  OR2_X1 U6905 ( .A1(n4482), .A2(n5441), .ZN(n5443) );
  INV_X1 U6906 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7443) );
  OR2_X1 U6907 ( .A1(n4483), .A2(n7443), .ZN(n5442) );
  NAND4_X1 U6908 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n8371)
         );
  INV_X1 U6909 ( .A(n8371), .ZN(n7603) );
  NAND2_X1 U6910 ( .A1(n7581), .A2(n7603), .ZN(n5727) );
  NAND2_X1 U6911 ( .A1(n5726), .A2(n5727), .ZN(n7436) );
  XNOR2_X1 U6912 ( .A(n5447), .B(n5446), .ZN(n7694) );
  NAND2_X1 U6913 ( .A1(n7694), .A2(n4990), .ZN(n5451) );
  NAND2_X1 U6914 ( .A1(n5448), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5449) );
  XNOR2_X1 U6915 ( .A(n5449), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7235) );
  AOI22_X1 U6916 ( .A1(n4475), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5512), .B2(
        n7235), .ZN(n5450) );
  NAND2_X1 U6917 ( .A1(n4485), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5461) );
  OAI21_X1 U6918 ( .B1(n5454), .B2(n5453), .A(n5452), .ZN(n5455) );
  AND2_X1 U6919 ( .A1(n5455), .A2(n5468), .ZN(n7590) );
  NAND2_X1 U6920 ( .A1(n5614), .A2(n7590), .ZN(n5460) );
  INV_X1 U6921 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5456) );
  OR2_X1 U6922 ( .A1(n4481), .A2(n5456), .ZN(n5459) );
  INV_X1 U6923 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5457) );
  OR2_X1 U6924 ( .A1(n4483), .A2(n5457), .ZN(n5458) );
  NAND4_X1 U6925 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n8648)
         );
  NAND2_X1 U6926 ( .A1(n7607), .A2(n8278), .ZN(n5730) );
  NAND2_X1 U6927 ( .A1(n7582), .A2(n5729), .ZN(n8642) );
  INV_X1 U6928 ( .A(n8642), .ZN(n5476) );
  XNOR2_X1 U6929 ( .A(n5463), .B(n5462), .ZN(n7697) );
  NAND2_X1 U6930 ( .A1(n7697), .A2(n4990), .ZN(n5467) );
  NAND2_X1 U6931 ( .A1(n5464), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5465) );
  XNOR2_X1 U6932 ( .A(n5465), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8071) );
  AOI22_X1 U6933 ( .A1(n4475), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5512), .B2(
        n8071), .ZN(n5466) );
  NAND2_X1 U6934 ( .A1(n4485), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5475) );
  INV_X1 U6935 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U6936 ( .A1(n5468), .A2(n8276), .ZN(n5469) );
  AND2_X1 U6937 ( .A1(n5486), .A2(n5469), .ZN(n8655) );
  NAND2_X1 U6938 ( .A1(n5614), .A2(n8655), .ZN(n5474) );
  INV_X1 U6939 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5470) );
  OR2_X1 U6940 ( .A1(n4483), .A2(n5470), .ZN(n5473) );
  INV_X1 U6941 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5471) );
  OR2_X1 U6942 ( .A1(n4482), .A2(n5471), .ZN(n5472) );
  NAND4_X1 U6943 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n8370)
         );
  INV_X1 U6944 ( .A(n8370), .ZN(n7604) );
  OR2_X1 U6945 ( .A1(n10015), .A2(n7604), .ZN(n5732) );
  NAND2_X1 U6946 ( .A1(n10015), .A2(n7604), .ZN(n7682) );
  NAND2_X1 U6947 ( .A1(n5732), .A2(n7682), .ZN(n8643) );
  NAND2_X1 U6948 ( .A1(n5476), .A2(n8644), .ZN(n8640) );
  XNOR2_X1 U6949 ( .A(n5478), .B(n5477), .ZN(n7769) );
  NAND2_X1 U6950 ( .A1(n7769), .A2(n4990), .ZN(n5485) );
  NOR2_X1 U6951 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  MUX2_X1 U6952 ( .A(n5479), .B(n5481), .S(P2_IR_REG_17__SCAN_IN), .Z(n5483)
         );
  INV_X1 U6953 ( .A(n5498), .ZN(n5482) );
  AOI22_X1 U6954 ( .A1(n4475), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8421), .B2(
        n5512), .ZN(n5484) );
  NAND2_X1 U6955 ( .A1(n4485), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5493) );
  INV_X1 U6956 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7668) );
  NAND2_X1 U6957 ( .A1(n5486), .A2(n7668), .ZN(n5487) );
  AND2_X1 U6958 ( .A1(n5502), .A2(n5487), .ZN(n7686) );
  NAND2_X1 U6959 ( .A1(n5614), .A2(n7686), .ZN(n5492) );
  INV_X1 U6960 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5488) );
  OR2_X1 U6961 ( .A1(n4481), .A2(n5488), .ZN(n5491) );
  INV_X1 U6962 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n5489) );
  OR2_X1 U6963 ( .A1(n4483), .A2(n5489), .ZN(n5490) );
  NAND4_X1 U6964 ( .A1(n5493), .A2(n5492), .A3(n5491), .A4(n5490), .ZN(n8647)
         );
  INV_X1 U6965 ( .A(n8647), .ZN(n8330) );
  NAND2_X1 U6966 ( .A1(n8110), .A2(n8330), .ZN(n5665) );
  NAND2_X1 U6967 ( .A1(n5666), .A2(n5665), .ZN(n7678) );
  INV_X1 U6968 ( .A(n7682), .ZN(n5494) );
  NOR2_X1 U6969 ( .A1(n7678), .A2(n5494), .ZN(n5495) );
  NAND2_X1 U6970 ( .A1(n8640), .A2(n5495), .ZN(n7680) );
  NAND2_X1 U6971 ( .A1(n7680), .A2(n5666), .ZN(n8631) );
  XNOR2_X1 U6972 ( .A(n5497), .B(n5496), .ZN(n7781) );
  NAND2_X1 U6973 ( .A1(n7781), .A2(n4990), .ZN(n5501) );
  NAND2_X1 U6974 ( .A1(n5498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5499) );
  XNOR2_X1 U6975 ( .A(n5499), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8078) );
  AOI22_X1 U6976 ( .A1(n4475), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5512), .B2(
        n8078), .ZN(n5500) );
  NAND2_X1 U6977 ( .A1(n4485), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U6978 ( .A1(n5502), .A2(n8825), .ZN(n5503) );
  AND2_X1 U6979 ( .A1(n5516), .A2(n5503), .ZN(n8625) );
  NAND2_X1 U6980 ( .A1(n5614), .A2(n8625), .ZN(n5508) );
  INV_X1 U6981 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5504) );
  OR2_X1 U6982 ( .A1(n4481), .A2(n5504), .ZN(n5507) );
  INV_X1 U6983 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5505) );
  OR2_X1 U6984 ( .A1(n4483), .A2(n5505), .ZN(n5506) );
  NAND4_X1 U6985 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), .ZN(n8369)
         );
  INV_X1 U6986 ( .A(n8369), .ZN(n8111) );
  NAND2_X1 U6987 ( .A1(n9098), .A2(n8111), .ZN(n5741) );
  XNOR2_X1 U6988 ( .A(n5511), .B(n5510), .ZN(n7801) );
  NAND2_X1 U6989 ( .A1(n7801), .A2(n4990), .ZN(n5514) );
  AOI22_X1 U6990 ( .A1(n4475), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4573), .B2(
        n5512), .ZN(n5513) );
  NAND2_X1 U6991 ( .A1(n4485), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5522) );
  INV_X1 U6992 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U6993 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  AND2_X1 U6994 ( .A1(n5529), .A2(n5517), .ZN(n8612) );
  NAND2_X1 U6995 ( .A1(n5614), .A2(n8612), .ZN(n5521) );
  INV_X1 U6996 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8878) );
  OR2_X1 U6997 ( .A1(n4482), .A2(n8878), .ZN(n5520) );
  INV_X1 U6998 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5518) );
  OR2_X1 U6999 ( .A1(n4483), .A2(n5518), .ZN(n5519) );
  NAND4_X1 U7000 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), .ZN(n8632)
         );
  XNOR2_X1 U7001 ( .A(n9094), .B(n8594), .ZN(n8609) );
  NAND2_X1 U7002 ( .A1(n9094), .A2(n8594), .ZN(n5746) );
  XNOR2_X1 U7003 ( .A(n5525), .B(n5524), .ZN(n7823) );
  NAND2_X1 U7004 ( .A1(n7823), .A2(n4990), .ZN(n5527) );
  NAND2_X1 U7005 ( .A1(n4475), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7006 ( .A1(n4485), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7007 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  AND2_X1 U7008 ( .A1(n5541), .A2(n5530), .ZN(n8603) );
  NAND2_X1 U7009 ( .A1(n5614), .A2(n8603), .ZN(n5534) );
  INV_X1 U7010 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8905) );
  OR2_X1 U7011 ( .A1(n4482), .A2(n8905), .ZN(n5533) );
  INV_X1 U7012 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5531) );
  OR2_X1 U7013 ( .A1(n4483), .A2(n5531), .ZN(n5532) );
  NAND4_X1 U7014 ( .A1(n5535), .A2(n5534), .A3(n5533), .A4(n5532), .ZN(n8586)
         );
  NAND2_X1 U7015 ( .A1(n9088), .A2(n8243), .ZN(n5751) );
  XNOR2_X1 U7016 ( .A(n5537), .B(n5536), .ZN(n7842) );
  NAND2_X1 U7017 ( .A1(n7842), .A2(n4990), .ZN(n5539) );
  NAND2_X1 U7018 ( .A1(n4475), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7019 ( .A1(n4485), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5548) );
  INV_X1 U7020 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7021 ( .A1(n5541), .A2(n5540), .ZN(n5542) );
  AND2_X1 U7022 ( .A1(n5555), .A2(n5542), .ZN(n8581) );
  NAND2_X1 U7023 ( .A1(n5614), .A2(n8581), .ZN(n5547) );
  INV_X1 U7024 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5543) );
  OR2_X1 U7025 ( .A1(n4482), .A2(n5543), .ZN(n5546) );
  INV_X1 U7026 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5544) );
  OR2_X1 U7027 ( .A1(n4483), .A2(n5544), .ZN(n5545) );
  NAND4_X1 U7028 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), .ZN(n8571)
         );
  XNOR2_X1 U7029 ( .A(n9081), .B(n8593), .ZN(n8578) );
  NAND2_X1 U7030 ( .A1(n9081), .A2(n8593), .ZN(n5750) );
  XNOR2_X1 U7031 ( .A(n5551), .B(n5550), .ZN(n7860) );
  NAND2_X1 U7032 ( .A1(n7860), .A2(n4990), .ZN(n5553) );
  NAND2_X1 U7033 ( .A1(n4475), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7034 ( .A1(n4485), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7035 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  AND2_X1 U7036 ( .A1(n5566), .A2(n5556), .ZN(n8565) );
  NAND2_X1 U7037 ( .A1(n5614), .A2(n8565), .ZN(n5560) );
  INV_X1 U7038 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8919) );
  OR2_X1 U7039 ( .A1(n4482), .A2(n8919), .ZN(n5559) );
  INV_X1 U7040 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5557) );
  OR2_X1 U7041 ( .A1(n4483), .A2(n5557), .ZN(n5558) );
  NAND4_X1 U7042 ( .A1(n5561), .A2(n5560), .A3(n5559), .A4(n5558), .ZN(n8587)
         );
  INV_X1 U7043 ( .A(n8587), .ZN(n8179) );
  NAND2_X1 U7044 ( .A1(n9076), .A2(n8179), .ZN(n5758) );
  NAND2_X1 U7045 ( .A1(n7880), .A2(n4990), .ZN(n5565) );
  NAND2_X1 U7046 ( .A1(n4475), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7047 ( .A1(n5566), .A2(n8178), .ZN(n5567) );
  NAND2_X1 U7048 ( .A1(n5577), .A2(n5567), .ZN(n8551) );
  NAND2_X1 U7049 ( .A1(n4485), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5569) );
  INV_X1 U7050 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8953) );
  OR2_X1 U7051 ( .A1(n4481), .A2(n8953), .ZN(n5568) );
  AND2_X1 U7052 ( .A1(n5569), .A2(n5568), .ZN(n5571) );
  NAND2_X1 U7053 ( .A1(n5642), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5570) );
  OAI211_X1 U7054 ( .C1(n5622), .C2(n8551), .A(n5571), .B(n5570), .ZN(n8572)
         );
  INV_X1 U7055 ( .A(n8572), .ZN(n8538) );
  NAND2_X1 U7056 ( .A1(n9071), .A2(n8538), .ZN(n5763) );
  XNOR2_X1 U7057 ( .A(n5573), .B(n5572), .ZN(n7899) );
  NAND2_X1 U7058 ( .A1(n7899), .A2(n4990), .ZN(n5575) );
  NAND2_X1 U7059 ( .A1(n4475), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5574) );
  INV_X1 U7060 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7061 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  NAND2_X1 U7062 ( .A1(n5587), .A2(n5578), .ZN(n8532) );
  OR2_X1 U7063 ( .A1(n8532), .A2(n5622), .ZN(n5581) );
  AOI22_X1 U7064 ( .A1(n4485), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n5643), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7065 ( .A1(n5642), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7066 ( .A1(n9066), .A2(n8297), .ZN(n5765) );
  NAND2_X1 U7067 ( .A1(n5767), .A2(n5765), .ZN(n8537) );
  NAND2_X1 U7068 ( .A1(n8541), .A2(n5767), .ZN(n8525) );
  XNOR2_X1 U7069 ( .A(n5584), .B(n5583), .ZN(n7914) );
  NAND2_X1 U7070 ( .A1(n7914), .A2(n4990), .ZN(n5586) );
  NAND2_X1 U7071 ( .A1(n4475), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5585) );
  INV_X1 U7072 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U7073 ( .A1(n5587), .A2(n8262), .ZN(n5588) );
  NAND2_X1 U7074 ( .A1(n5596), .A2(n5588), .ZN(n8519) );
  OR2_X1 U7075 ( .A1(n8519), .A2(n5622), .ZN(n5591) );
  AOI22_X1 U7076 ( .A1(n4485), .A2(P2_REG1_REG_25__SCAN_IN), .B1(n5642), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n5590) );
  INV_X1 U7077 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8929) );
  OR2_X1 U7078 ( .A1(n4481), .A2(n8929), .ZN(n5589) );
  NAND2_X1 U7079 ( .A1(n9063), .A2(n8539), .ZN(n5768) );
  NAND2_X1 U7080 ( .A1(n8525), .A2(n8524), .ZN(n8523) );
  XNOR2_X1 U7081 ( .A(n5593), .B(n5592), .ZN(n9136) );
  NAND2_X1 U7082 ( .A1(n9136), .A2(n4990), .ZN(n5595) );
  NAND2_X1 U7083 ( .A1(n4475), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7084 ( .A1(n5596), .A2(n8353), .ZN(n5597) );
  INV_X1 U7085 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7086 ( .A1(n4485), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5600) );
  INV_X1 U7087 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8941) );
  OR2_X1 U7088 ( .A1(n4482), .A2(n8941), .ZN(n5599) );
  OAI211_X1 U7089 ( .C1(n5601), .C2(n4483), .A(n5600), .B(n5599), .ZN(n5602)
         );
  OR2_X1 U7090 ( .A1(n9056), .A2(n8477), .ZN(n5775) );
  NAND2_X1 U7091 ( .A1(n9056), .A2(n8477), .ZN(n5776) );
  XNOR2_X1 U7092 ( .A(n5604), .B(n5603), .ZN(n9132) );
  NAND2_X1 U7093 ( .A1(n9132), .A2(n4990), .ZN(n5606) );
  NAND2_X1 U7094 ( .A1(n4475), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5605) );
  XNOR2_X1 U7095 ( .A(n5607), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8486) );
  INV_X1 U7096 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7097 ( .A1(n5643), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7098 ( .A1(n4485), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5609) );
  OAI211_X1 U7099 ( .C1(n5612), .C2(n4483), .A(n5610), .B(n5609), .ZN(n5613)
         );
  NAND2_X1 U7100 ( .A1(n9049), .A2(n8498), .ZN(n5779) );
  INV_X1 U7101 ( .A(n5617), .ZN(n5618) );
  INV_X1 U7102 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9127) );
  INV_X1 U7103 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9965) );
  XNOR2_X1 U7104 ( .A(n5629), .B(SI_29_), .ZN(n5619) );
  NAND2_X1 U7105 ( .A1(n9125), .A2(n4990), .ZN(n5621) );
  NAND2_X1 U7106 ( .A1(n4475), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5620) );
  OR2_X1 U7107 ( .A1(n8118), .A2(n5622), .ZN(n5628) );
  INV_X1 U7108 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7109 ( .A1(n5642), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U7110 ( .A1(n5643), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5623) );
  OAI211_X1 U7111 ( .C1(n4484), .C2(n5625), .A(n5624), .B(n5623), .ZN(n5626)
         );
  INV_X1 U7112 ( .A(n5626), .ZN(n5627) );
  INV_X1 U7113 ( .A(n5629), .ZN(n5630) );
  NOR2_X1 U7114 ( .A1(n5630), .A2(SI_29_), .ZN(n5632) );
  NAND2_X1 U7115 ( .A1(n5630), .A2(SI_29_), .ZN(n5631) );
  NAND2_X1 U7116 ( .A1(n8106), .A2(n4990), .ZN(n5635) );
  NAND2_X1 U7117 ( .A1(n5279), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5634) );
  INV_X1 U7118 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7119 ( .A1(n5643), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7120 ( .A1(n5642), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5636) );
  OAI211_X1 U7121 ( .C1(n4484), .C2(n5638), .A(n5637), .B(n5636), .ZN(n8364)
         );
  NAND2_X1 U7122 ( .A1(n5639), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5640) );
  MUX2_X1 U7123 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5640), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5641) );
  NAND2_X1 U7124 ( .A1(n5641), .A2(n5830), .ZN(n7336) );
  INV_X1 U7125 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7126 ( .A1(n5642), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7127 ( .A1(n5643), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5644) );
  OAI211_X1 U7128 ( .C1(n4484), .C2(n5646), .A(n5645), .B(n5644), .ZN(n8449)
         );
  NAND2_X1 U7129 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  XNOR2_X1 U7130 ( .A(n5651), .B(SI_31_), .ZN(n5652) );
  XNOR2_X1 U7131 ( .A(n5653), .B(n5652), .ZN(n8092) );
  NAND2_X1 U7132 ( .A1(n8092), .A2(n4990), .ZN(n5655) );
  NAND2_X1 U7133 ( .A1(n4475), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5654) );
  INV_X1 U7134 ( .A(n8449), .ZN(n5657) );
  OR2_X1 U7135 ( .A1(n9022), .A2(n5657), .ZN(n5789) );
  INV_X1 U7136 ( .A(n8364), .ZN(n5656) );
  NAND2_X1 U7137 ( .A1(n8454), .A2(n5656), .ZN(n5787) );
  XOR2_X1 U7138 ( .A(n4573), .B(n5658), .Z(n5822) );
  XNOR2_X2 U7139 ( .A(n5661), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6600) );
  OR2_X4 U7140 ( .A1(n6576), .A2(n10326), .ZN(n8156) );
  NAND2_X1 U7141 ( .A1(n6600), .A2(n6597), .ZN(n6591) );
  NAND2_X1 U7142 ( .A1(n4486), .A2(n6591), .ZN(n5821) );
  AND2_X1 U7143 ( .A1(n9035), .A2(n6597), .ZN(n5664) );
  NAND2_X1 U7144 ( .A1(n4573), .A2(n5664), .ZN(n5788) );
  MUX2_X1 U7145 ( .A(n5815), .B(n5814), .S(n5788), .Z(n5792) );
  MUX2_X1 U7146 ( .A(n4499), .B(n5781), .S(n5782), .Z(n5786) );
  INV_X1 U7147 ( .A(n5665), .ZN(n5668) );
  NAND2_X1 U7148 ( .A1(n5743), .A2(n5666), .ZN(n5667) );
  MUX2_X1 U7149 ( .A(n5668), .B(n5667), .S(n5788), .Z(n5669) );
  INV_X1 U7150 ( .A(n5669), .ZN(n5736) );
  INV_X1 U7151 ( .A(n7678), .ZN(n7681) );
  INV_X1 U7152 ( .A(n8643), .ZN(n8644) );
  NAND2_X1 U7153 ( .A1(n10256), .A2(n5794), .ZN(n5671) );
  INV_X1 U7154 ( .A(n5687), .ZN(n5670) );
  MUX2_X1 U7155 ( .A(n5671), .B(n5670), .S(n5788), .Z(n5688) );
  OAI211_X1 U7156 ( .C1(n5688), .C2(n5672), .A(n5693), .B(n10256), .ZN(n5673)
         );
  NAND2_X1 U7157 ( .A1(n5673), .A2(n5788), .ZN(n5681) );
  NAND3_X1 U7158 ( .A1(n5795), .A2(n6368), .A3(n6597), .ZN(n5676) );
  INV_X1 U7159 ( .A(n5683), .ZN(n5675) );
  AOI21_X1 U7160 ( .B1(n5674), .B2(n5676), .A(n5675), .ZN(n5679) );
  NAND2_X1 U7161 ( .A1(n6588), .A2(n5788), .ZN(n5678) );
  INV_X1 U7162 ( .A(n5688), .ZN(n5677) );
  OAI211_X1 U7163 ( .C1(n5679), .C2(n5678), .A(n5677), .B(n6585), .ZN(n5680)
         );
  NAND2_X1 U7164 ( .A1(n5795), .A2(n6368), .ZN(n5682) );
  NAND3_X1 U7165 ( .A1(n6588), .A2(n5796), .A3(n5682), .ZN(n5684) );
  NAND3_X1 U7166 ( .A1(n5684), .A2(n5782), .A3(n5683), .ZN(n5685) );
  AOI22_X1 U7167 ( .A1(n5688), .A2(n5793), .B1(n5687), .B2(n5686), .ZN(n5691)
         );
  INV_X1 U7168 ( .A(n5689), .ZN(n5690) );
  OAI21_X1 U7169 ( .B1(n5691), .B2(n5690), .A(n5782), .ZN(n5692) );
  NAND2_X1 U7170 ( .A1(n5695), .A2(n5694), .ZN(n9005) );
  INV_X1 U7171 ( .A(n9005), .ZN(n9014) );
  MUX2_X1 U7172 ( .A(n5695), .B(n5694), .S(n5788), .Z(n5696) );
  NAND3_X1 U7173 ( .A1(n5697), .A2(n10236), .A3(n5696), .ZN(n5704) );
  INV_X1 U7174 ( .A(n5698), .ZN(n5701) );
  OAI21_X1 U7175 ( .B1(n5699), .B2(n10375), .A(n5799), .ZN(n5700) );
  MUX2_X1 U7176 ( .A(n5701), .B(n5700), .S(n5788), .Z(n5702) );
  INV_X1 U7177 ( .A(n5702), .ZN(n5703) );
  NAND3_X1 U7178 ( .A1(n5704), .A2(n5798), .A3(n5703), .ZN(n5707) );
  AND2_X1 U7179 ( .A1(n7081), .A2(n5798), .ZN(n5705) );
  MUX2_X1 U7180 ( .A(n5799), .B(n5705), .S(n5788), .Z(n5706) );
  NAND3_X1 U7181 ( .A1(n5707), .A2(n5708), .A3(n5706), .ZN(n5712) );
  AND2_X1 U7182 ( .A1(n7217), .A2(n7081), .ZN(n5710) );
  AND2_X1 U7183 ( .A1(n5715), .A2(n5708), .ZN(n5709) );
  MUX2_X1 U7184 ( .A(n5710), .B(n5709), .S(n5788), .Z(n5711) );
  NAND2_X1 U7185 ( .A1(n5712), .A2(n5711), .ZN(n5718) );
  INV_X1 U7186 ( .A(n5804), .ZN(n5713) );
  AOI21_X1 U7187 ( .B1(n5718), .B2(n5714), .A(n5713), .ZN(n5720) );
  AND2_X1 U7188 ( .A1(n5804), .A2(n5715), .ZN(n5717) );
  INV_X1 U7189 ( .A(n5803), .ZN(n5716) );
  AOI21_X1 U7190 ( .B1(n5718), .B2(n5717), .A(n5716), .ZN(n5719) );
  MUX2_X1 U7191 ( .A(n5720), .B(n5719), .S(n5782), .Z(n5721) );
  NAND2_X1 U7192 ( .A1(n5721), .A2(n5012), .ZN(n5725) );
  INV_X1 U7193 ( .A(n7436), .ZN(n7439) );
  MUX2_X1 U7194 ( .A(n5723), .B(n5722), .S(n5782), .Z(n5724) );
  MUX2_X1 U7195 ( .A(n5727), .B(n5726), .S(n5788), .Z(n5728) );
  MUX2_X1 U7196 ( .A(n5730), .B(n5729), .S(n5782), .Z(n5731) );
  MUX2_X1 U7197 ( .A(n5732), .B(n7682), .S(n5782), .Z(n5733) );
  NAND2_X1 U7198 ( .A1(n7681), .A2(n5734), .ZN(n5735) );
  NAND2_X1 U7199 ( .A1(n5736), .A2(n5735), .ZN(n5745) );
  OR2_X1 U7200 ( .A1(n9094), .A2(n8594), .ZN(n5742) );
  INV_X1 U7201 ( .A(n5742), .ZN(n5737) );
  AOI21_X1 U7202 ( .B1(n5745), .B2(n5741), .A(n5737), .ZN(n5739) );
  NAND2_X1 U7203 ( .A1(n5751), .A2(n5746), .ZN(n5738) );
  OR2_X1 U7204 ( .A1(n9081), .A2(n8593), .ZN(n5753) );
  OAI211_X1 U7205 ( .C1(n5739), .C2(n5738), .A(n5748), .B(n5753), .ZN(n5740)
         );
  NAND3_X1 U7206 ( .A1(n5740), .A2(n5758), .A3(n5750), .ZN(n5756) );
  INV_X1 U7207 ( .A(n5741), .ZN(n5744) );
  OAI211_X1 U7208 ( .C1(n5745), .C2(n5744), .A(n5743), .B(n5742), .ZN(n5747)
         );
  NAND2_X1 U7209 ( .A1(n5747), .A2(n5746), .ZN(n5749) );
  NAND2_X1 U7210 ( .A1(n5749), .A2(n5748), .ZN(n5752) );
  NAND3_X1 U7211 ( .A1(n5752), .A2(n5751), .A3(n5750), .ZN(n5754) );
  NAND3_X1 U7212 ( .A1(n5754), .A2(n5757), .A3(n5753), .ZN(n5755) );
  MUX2_X1 U7213 ( .A(n5756), .B(n5755), .S(n5782), .Z(n5759) );
  AND3_X1 U7214 ( .A1(n5759), .A2(n8556), .A3(n5757), .ZN(n5762) );
  NAND3_X1 U7215 ( .A1(n5759), .A2(n8556), .A3(n5758), .ZN(n5760) );
  OAI211_X1 U7216 ( .C1(n8538), .C2(n9071), .A(n5582), .B(n5760), .ZN(n5761)
         );
  MUX2_X1 U7217 ( .A(n5762), .B(n5761), .S(n5782), .Z(n5766) );
  NAND2_X1 U7218 ( .A1(n5765), .A2(n5763), .ZN(n5764) );
  AOI22_X1 U7219 ( .A1(n5766), .A2(n5765), .B1(n5788), .B2(n5764), .ZN(n5772)
         );
  OAI21_X1 U7220 ( .B1(n5782), .B2(n5767), .A(n8524), .ZN(n5771) );
  INV_X1 U7221 ( .A(n5768), .ZN(n5769) );
  OAI21_X1 U7222 ( .B1(n8492), .B2(n5769), .A(n5788), .ZN(n5770) );
  AOI21_X1 U7223 ( .B1(n5775), .B2(n5773), .A(n5788), .ZN(n5774) );
  NOR2_X1 U7224 ( .A1(n5776), .A2(n5788), .ZN(n5777) );
  MUX2_X1 U7225 ( .A(n5779), .B(n5778), .S(n5782), .Z(n5780) );
  OR3_X1 U7226 ( .A1(n9043), .A2(n8478), .A3(n5782), .ZN(n5784) );
  NAND3_X1 U7227 ( .A1(n9043), .A2(n8478), .A3(n5782), .ZN(n5783) );
  AND4_X1 U7228 ( .A1(n4490), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n5791)
         );
  MUX2_X1 U7229 ( .A(n4496), .B(n5789), .S(n5788), .Z(n5790) );
  OAI21_X1 U7230 ( .B1(n5792), .B2(n5791), .A(n5790), .ZN(n5818) );
  INV_X1 U7231 ( .A(n8482), .ZN(n5812) );
  AND2_X1 U7232 ( .A1(n10256), .A2(n5793), .ZN(n6841) );
  NAND2_X1 U7233 ( .A1(n6607), .A2(n6368), .ZN(n6660) );
  NAND2_X1 U7234 ( .A1(n5794), .A2(n10282), .ZN(n10291) );
  NAND2_X1 U7235 ( .A1(n5796), .A2(n5795), .ZN(n6609) );
  NOR4_X1 U7236 ( .A1(n6582), .A2(n6660), .A3(n10291), .A4(n6609), .ZN(n5797)
         );
  NAND4_X1 U7237 ( .A1(n6841), .A2(n6585), .A3(n6600), .A4(n5797), .ZN(n5801)
         );
  NAND2_X1 U7238 ( .A1(n5799), .A2(n5798), .ZN(n6944) );
  NOR4_X1 U7239 ( .A1(n5801), .A2(n6944), .A3(n9005), .A4(n10265), .ZN(n5802)
         );
  NAND3_X1 U7240 ( .A1(n7076), .A2(n5802), .A3(n10236), .ZN(n5806) );
  NAND2_X1 U7241 ( .A1(n5804), .A2(n5803), .ZN(n7225) );
  NOR4_X1 U7242 ( .A1(n7399), .A2(n5806), .A3(n7225), .A4(n7082), .ZN(n5807)
         );
  NAND4_X1 U7243 ( .A1(n8644), .A2(n7583), .A3(n7439), .A4(n5807), .ZN(n5808)
         );
  NOR4_X1 U7244 ( .A1(n8598), .A2(n4688), .A3(n7678), .A4(n5808), .ZN(n5809)
         );
  NAND4_X1 U7245 ( .A1(n8569), .A2(n5809), .A3(n5549), .A4(n5523), .ZN(n5810)
         );
  NOR4_X1 U7246 ( .A1(n8512), .A2(n8537), .A3(n8547), .A4(n5810), .ZN(n5811)
         );
  NAND4_X1 U7247 ( .A1(n8123), .A2(n5812), .A3(n8495), .A4(n5811), .ZN(n5813)
         );
  AND2_X1 U7248 ( .A1(n5662), .A2(n4573), .ZN(n9036) );
  AOI22_X1 U7249 ( .A1(n5816), .A2(n7336), .B1(n9036), .B2(n6589), .ZN(n5817)
         );
  AOI21_X1 U7250 ( .B1(n5662), .B2(n5818), .A(n5817), .ZN(n5820) );
  NAND2_X1 U7251 ( .A1(n5662), .A2(n9035), .ZN(n5819) );
  NAND2_X1 U7252 ( .A1(n5823), .A2(n5827), .ZN(n5824) );
  NAND2_X1 U7253 ( .A1(n5839), .A2(n5826), .ZN(n6287) );
  OR2_X1 U7254 ( .A1(n6287), .A2(P2_U3152), .ZN(n6039) );
  NAND3_X1 U7255 ( .A1(n5828), .A2(n5827), .A3(n5840), .ZN(n5829) );
  NAND2_X1 U7256 ( .A1(n5837), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5833) );
  MUX2_X1 U7257 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5833), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5834) );
  NAND2_X1 U7258 ( .A1(n5835), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5836) );
  MUX2_X1 U7259 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5836), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5838) );
  NAND2_X1 U7260 ( .A1(n5839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5841) );
  INV_X1 U7261 ( .A(n7611), .ZN(n5842) );
  INV_X1 U7262 ( .A(n6040), .ZN(n6288) );
  NAND2_X1 U7263 ( .A1(n6589), .A2(n6597), .ZN(n6038) );
  OR2_X1 U7264 ( .A1(n5844), .A2(n6038), .ZN(n10286) );
  NOR4_X1 U7265 ( .A1(n10309), .A2(n9133), .A3(n6576), .A4(n10286), .ZN(n5846)
         );
  OAI21_X1 U7266 ( .B1(n6039), .B2(n6589), .A(P2_B_REG_SCAN_IN), .ZN(n5845) );
  OR2_X1 U7267 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  NAND2_X1 U7268 ( .A1(n5892), .A2(n5848), .ZN(n5900) );
  NAND2_X1 U7269 ( .A1(n6479), .A2(n5851), .ZN(n6769) );
  INV_X1 U7270 ( .A(n6769), .ZN(n5855) );
  NOR2_X1 U7271 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5854) );
  NAND4_X1 U7272 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n5861)
         );
  NOR2_X1 U7273 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5859) );
  NAND4_X1 U7274 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n5860)
         );
  NOR2_X1 U7275 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  NAND2_X1 U7276 ( .A1(n5863), .A2(n5862), .ZN(n6185) );
  NAND2_X1 U7277 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U7278 ( .A1(n5871), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5872) );
  INV_X1 U7279 ( .A(n5874), .ZN(n5875) );
  NAND2_X1 U7280 ( .A1(n5875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5877) );
  INV_X1 U7281 ( .A(n7451), .ZN(n6519) );
  NAND2_X1 U7282 ( .A1(n5879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7283 ( .A1(n5882), .A2(n5881), .ZN(n5884) );
  NAND2_X1 U7284 ( .A1(n5884), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5880) );
  OR2_X1 U7285 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  INV_X1 U7286 ( .A(n9472), .ZN(n9480) );
  NAND2_X1 U7287 ( .A1(n9467), .A2(n7451), .ZN(n5885) );
  NAND2_X1 U7288 ( .A1(n5957), .A2(n5885), .ZN(n5955) );
  NAND2_X1 U7289 ( .A1(n4530), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5888) );
  XNOR2_X2 U7290 ( .A(n5890), .B(n5889), .ZN(n10065) );
  NAND2_X2 U7291 ( .A1(n5956), .A2(n10065), .ZN(n6542) );
  OAI21_X1 U7292 ( .B1(n5955), .B2(n7802), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  NOR2_X1 U7293 ( .A1(n6417), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9129) );
  INV_X1 U7294 ( .A(n9129), .ZN(n9137) );
  NAND2_X1 U7295 ( .A1(n6417), .A2(P2_U3152), .ZN(n9139) );
  OAI222_X1 U7296 ( .A1(n9137), .A2(n5056), .B1(n9134), .B2(n6416), .C1(n6062), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  INV_X1 U7297 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5891) );
  INV_X1 U7298 ( .A(n9991), .ZN(n6049) );
  OAI222_X1 U7299 ( .A1(n9137), .A2(n5891), .B1(n9134), .B2(n6446), .C1(n6049), 
        .C2(P2_U3152), .ZN(P2_U3356) );
  OR2_X1 U7300 ( .A1(n5892), .A2(n6035), .ZN(n5894) );
  INV_X1 U7301 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7302 ( .A1(n5894), .A2(n5893), .ZN(n5897) );
  OAI21_X1 U7303 ( .B1(n5894), .B2(n5893), .A(n5897), .ZN(n6448) );
  NOR2_X1 U7304 ( .A1(n6417), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9961) );
  INV_X1 U7305 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6447) );
  AND2_X1 U7306 ( .A1(n6417), .A2(P1_U3084), .ZN(n7452) );
  INV_X1 U7307 ( .A(n7452), .ZN(n9968) );
  OAI222_X1 U7308 ( .A1(P1_U3084), .A2(n6448), .B1(n9971), .B2(n6446), .C1(
        n6447), .C2(n9968), .ZN(P1_U3351) );
  INV_X1 U7309 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7310 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5895) );
  XNOR2_X1 U7311 ( .A(n5896), .B(n5895), .ZN(n6419) );
  INV_X1 U7312 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6418) );
  OAI222_X1 U7313 ( .A1(P1_U3084), .A2(n6419), .B1(n9971), .B2(n6416), .C1(
        n6418), .C2(n9968), .ZN(P1_U3352) );
  NAND2_X1 U7314 ( .A1(n5897), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5899) );
  INV_X1 U7315 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5898) );
  XNOR2_X1 U7316 ( .A(n5899), .B(n5898), .ZN(n6508) );
  INV_X1 U7317 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6507) );
  OAI222_X1 U7318 ( .A1(P1_U3084), .A2(n6508), .B1(n9971), .B2(n6505), .C1(
        n6507), .C2(n9968), .ZN(P1_U3350) );
  INV_X1 U7319 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8876) );
  INV_X1 U7320 ( .A(n6064), .ZN(n6241) );
  OAI222_X1 U7321 ( .A1(n9137), .A2(n8876), .B1(n9134), .B2(n6505), .C1(n6241), 
        .C2(P2_U3152), .ZN(P2_U3355) );
  NAND2_X1 U7322 ( .A1(n5900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5901) );
  XNOR2_X1 U7323 ( .A(n5901), .B(n5849), .ZN(n6541) );
  INV_X1 U7324 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8864) );
  OAI222_X1 U7325 ( .A1(P1_U3084), .A2(n6541), .B1(n9971), .B2(n6540), .C1(
        n8864), .C2(n9968), .ZN(P1_U3349) );
  INV_X1 U7326 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5902) );
  INV_X1 U7327 ( .A(n6066), .ZN(n6277) );
  OAI222_X1 U7328 ( .A1(n9137), .A2(n5902), .B1(n9134), .B2(n6540), .C1(n6277), 
        .C2(P2_U3152), .ZN(P2_U3354) );
  INV_X1 U7329 ( .A(n6793), .ZN(n5906) );
  NAND2_X1 U7330 ( .A1(n5915), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5904) );
  XNOR2_X1 U7331 ( .A(n5904), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10080) );
  AOI22_X1 U7332 ( .A1(n10080), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n7452), .ZN(n5905) );
  OAI21_X1 U7333 ( .B1(n5906), .B2(n9971), .A(n5905), .ZN(P1_U3348) );
  INV_X1 U7334 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5907) );
  INV_X1 U7335 ( .A(n6068), .ZN(n6254) );
  OAI222_X1 U7336 ( .A1(n9137), .A2(n5907), .B1(n9134), .B2(n5906), .C1(n6254), 
        .C2(P2_U3152), .ZN(P2_U3353) );
  AND2_X1 U7337 ( .A1(n7451), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5908) );
  INV_X1 U7338 ( .A(n9956), .ZN(n10159) );
  INV_X1 U7339 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5914) );
  NAND3_X1 U7340 ( .A1(n7674), .A2(P1_B_REG_SCAN_IN), .A3(n7613), .ZN(n5909)
         );
  OR2_X1 U7341 ( .A1(n10158), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5912) );
  INV_X1 U7342 ( .A(n5910), .ZN(n9973) );
  NAND2_X1 U7343 ( .A1(n9973), .A2(n7674), .ZN(n5911) );
  NAND2_X1 U7344 ( .A1(n5912), .A2(n5911), .ZN(n6320) );
  INV_X1 U7345 ( .A(n6320), .ZN(n6652) );
  NAND2_X1 U7346 ( .A1(n6652), .A2(n10159), .ZN(n5913) );
  OAI21_X1 U7347 ( .B1(n10159), .B2(n5914), .A(n5913), .ZN(P1_U3441) );
  NOR2_X1 U7348 ( .A1(n5915), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5923) );
  INV_X1 U7349 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6035) );
  OR2_X1 U7350 ( .A1(n5923), .A2(n6035), .ZN(n5916) );
  XNOR2_X1 U7351 ( .A(n5916), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10098) );
  AOI22_X1 U7352 ( .A1(n10098), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7452), .ZN(n5917) );
  OAI21_X1 U7353 ( .B1(n6778), .B2(n9971), .A(n5917), .ZN(P1_U3347) );
  INV_X1 U7354 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5918) );
  OAI222_X1 U7355 ( .A1(n9137), .A2(n5918), .B1(n9134), .B2(n6778), .C1(n6265), 
        .C2(P2_U3152), .ZN(P2_U3352) );
  OAI21_X1 U7356 ( .B1(n10309), .B2(n6038), .A(n5247), .ZN(n5920) );
  NAND2_X1 U7357 ( .A1(n10309), .A2(n6039), .ZN(n5919) );
  NAND2_X1 U7358 ( .A1(n5920), .A2(n5919), .ZN(n8091) );
  NOR2_X1 U7359 ( .A1(n10231), .A2(P2_U3966), .ZN(P2_U3151) );
  OAI21_X1 U7360 ( .B1(n6190), .B2(P2_U3966), .A(n5921), .ZN(P2_U3552) );
  INV_X1 U7361 ( .A(n6814), .ZN(n5928) );
  OR2_X1 U7362 ( .A1(n5932), .A2(n6035), .ZN(n5924) );
  XNOR2_X1 U7363 ( .A(n5924), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U7364 ( .A1(n6815), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7452), .ZN(n5925) );
  OAI21_X1 U7365 ( .B1(n5928), .B2(n9971), .A(n5925), .ZN(P1_U3346) );
  INV_X1 U7366 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7367 ( .A1(n8449), .A2(P2_U3966), .ZN(n5926) );
  OAI21_X1 U7368 ( .B1(n5927), .B2(P2_U3966), .A(n5926), .ZN(P2_U3583) );
  INV_X1 U7369 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5929) );
  INV_X1 U7370 ( .A(n6071), .ZN(n6229) );
  OAI222_X1 U7371 ( .A1(n9137), .A2(n5929), .B1(n9139), .B2(n5928), .C1(
        P2_U3152), .C2(n6229), .ZN(P2_U3351) );
  INV_X1 U7372 ( .A(n5930), .ZN(n5937) );
  NAND2_X1 U7373 ( .A1(n5932), .A2(n5931), .ZN(n5934) );
  NAND2_X1 U7374 ( .A1(n5934), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5933) );
  MUX2_X1 U7375 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5933), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5935) );
  AND2_X1 U7376 ( .A1(n5935), .A2(n6034), .ZN(n6908) );
  AOI22_X1 U7377 ( .A1(n6908), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7452), .ZN(n5936) );
  OAI21_X1 U7378 ( .B1(n5937), .B2(n9971), .A(n5936), .ZN(P1_U3345) );
  INV_X1 U7379 ( .A(n6334), .ZN(n6328) );
  OAI222_X1 U7380 ( .A1(n9137), .A2(n6386), .B1(n9139), .B2(n5937), .C1(
        P2_U3152), .C2(n6328), .ZN(P2_U3350) );
  XNOR2_X2 U7381 ( .A(n5941), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7382 ( .A1(n6431), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5951) );
  INV_X1 U7383 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6091) );
  OR2_X1 U7384 ( .A1(n4478), .A2(n6091), .ZN(n5950) );
  NAND2_X2 U7385 ( .A1(n5943), .A2(n5942), .ZN(n6527) );
  NAND3_X1 U7386 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6782) );
  INV_X1 U7387 ( .A(n6782), .ZN(n5944) );
  NAND2_X1 U7388 ( .A1(n5944), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6821) );
  INV_X1 U7389 ( .A(n6821), .ZN(n5945) );
  NAND2_X1 U7390 ( .A1(n5945), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6823) );
  INV_X1 U7391 ( .A(n6823), .ZN(n5946) );
  NAND2_X1 U7392 ( .A1(n5946), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U7393 ( .A1(n6922), .A2(n7270), .ZN(n5947) );
  NAND2_X1 U7394 ( .A1(n7272), .A2(n5947), .ZN(n7330) );
  OR2_X1 U7395 ( .A1(n6527), .A2(n7330), .ZN(n5949) );
  INV_X1 U7396 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7331) );
  OR2_X1 U7397 ( .A1(n4477), .A2(n7331), .ZN(n5948) );
  MUX2_X1 U7398 ( .A(n5952), .B(n7422), .S(P1_U4006), .Z(n5953) );
  INV_X1 U7399 ( .A(n5953), .ZN(P1_U3565) );
  INV_X1 U7400 ( .A(n7115), .ZN(n6011) );
  AOI22_X1 U7401 ( .A1(n8384), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9129), .ZN(n5954) );
  OAI21_X1 U7402 ( .B1(n6011), .B2(n9134), .A(n5954), .ZN(P2_U3349) );
  NOR2_X1 U7403 ( .A1(n5955), .A2(P1_U3084), .ZN(n5960) );
  INV_X1 U7404 ( .A(n10065), .ZN(n7995) );
  NAND2_X1 U7405 ( .A1(n5960), .A2(n7995), .ZN(n9592) );
  INV_X1 U7406 ( .A(n5956), .ZN(n6671) );
  INV_X1 U7407 ( .A(n5957), .ZN(n5958) );
  INV_X1 U7408 ( .A(n10063), .ZN(n10122) );
  NOR2_X1 U7409 ( .A1(n5956), .A2(n7995), .ZN(n5959) );
  INV_X1 U7410 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10213) );
  MUX2_X1 U7411 ( .A(n10213), .B(P1_REG1_REG_1__SCAN_IN), .S(n6419), .Z(n5962)
         );
  AND2_X1 U7412 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n5961) );
  NAND2_X1 U7413 ( .A1(n5962), .A2(n5961), .ZN(n5976) );
  OAI21_X1 U7414 ( .B1(n5962), .B2(n5961), .A(n5976), .ZN(n5963) );
  INV_X1 U7415 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10151) );
  OAI22_X1 U7416 ( .A1(n10106), .A2(n5963), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10151), .ZN(n5964) );
  AOI21_X1 U7417 ( .B1(n10122), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n5964), .ZN(
        n5968) );
  INV_X1 U7418 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10156) );
  MUX2_X1 U7419 ( .A(n10156), .B(P1_REG2_REG_1__SCAN_IN), .S(n6419), .Z(n5966)
         );
  AND2_X1 U7420 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n5965) );
  OR2_X1 U7421 ( .A1(n9592), .A2(n5956), .ZN(n9590) );
  NAND2_X1 U7422 ( .A1(n5966), .A2(n5965), .ZN(n5970) );
  OAI211_X1 U7423 ( .C1(n5966), .C2(n5965), .A(n10124), .B(n5970), .ZN(n5967)
         );
  OAI211_X1 U7424 ( .C1(n9595), .C2(n6419), .A(n5968), .B(n5967), .ZN(P1_U3242) );
  XNOR2_X1 U7425 ( .A(n6508), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n5973) );
  INV_X1 U7426 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6725) );
  MUX2_X1 U7427 ( .A(n6725), .B(P1_REG2_REG_2__SCAN_IN), .S(n6448), .Z(n6363)
         );
  INV_X1 U7428 ( .A(n6419), .ZN(n5974) );
  NAND2_X1 U7429 ( .A1(n5974), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7430 ( .A1(n5970), .A2(n5969), .ZN(n6362) );
  NAND2_X1 U7431 ( .A1(n6363), .A2(n6362), .ZN(n6361) );
  INV_X1 U7432 ( .A(n6448), .ZN(n5977) );
  NAND2_X1 U7433 ( .A1(n5977), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7434 ( .A1(n6361), .A2(n5971), .ZN(n5972) );
  NAND2_X1 U7435 ( .A1(n5972), .A2(n5973), .ZN(n5989) );
  OAI211_X1 U7436 ( .C1(n5973), .C2(n5972), .A(n10124), .B(n5989), .ZN(n5987)
         );
  INV_X1 U7437 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n5984) );
  AND2_X1 U7438 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6533) );
  INV_X1 U7439 ( .A(n6533), .ZN(n5983) );
  INV_X1 U7440 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10215) );
  MUX2_X1 U7441 ( .A(n10215), .B(P1_REG1_REG_2__SCAN_IN), .S(n6448), .Z(n6359)
         );
  NAND2_X1 U7442 ( .A1(n5974), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7443 ( .A1(n5976), .A2(n5975), .ZN(n6358) );
  NAND2_X1 U7444 ( .A1(n6359), .A2(n6358), .ZN(n6357) );
  NAND2_X1 U7445 ( .A1(n5977), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7446 ( .A1(n6357), .A2(n5978), .ZN(n5980) );
  XNOR2_X1 U7447 ( .A(n6508), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n5979) );
  AND2_X1 U7448 ( .A1(n5980), .A2(n5979), .ZN(n6000) );
  NOR2_X1 U7449 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  OR3_X1 U7450 ( .A1(n10106), .A2(n6000), .A3(n5981), .ZN(n5982) );
  OAI211_X1 U7451 ( .C1(n10063), .C2(n5984), .A(n5983), .B(n5982), .ZN(n5985)
         );
  INV_X1 U7452 ( .A(n5985), .ZN(n5986) );
  OAI211_X1 U7453 ( .C1(n9595), .C2(n6508), .A(n5987), .B(n5986), .ZN(P1_U3244) );
  INV_X1 U7454 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6009) );
  INV_X1 U7455 ( .A(n9595), .ZN(n10118) );
  INV_X1 U7456 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6465) );
  OR2_X1 U7457 ( .A1(n6508), .A2(n6465), .ZN(n5988) );
  NAND2_X1 U7458 ( .A1(n5989), .A2(n5988), .ZN(n9572) );
  INV_X1 U7459 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6710) );
  XNOR2_X1 U7460 ( .A(n6541), .B(n6710), .ZN(n9573) );
  OR2_X1 U7461 ( .A1(n9572), .A2(n9573), .ZN(n9574) );
  NAND2_X1 U7462 ( .A1(n6541), .A2(n6710), .ZN(n5990) );
  NAND2_X1 U7463 ( .A1(n9574), .A2(n5990), .ZN(n10082) );
  NOR2_X1 U7464 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10080), .ZN(n5991) );
  AOI21_X1 U7465 ( .B1(n10080), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5991), .ZN(
        n10083) );
  NAND2_X1 U7466 ( .A1(n10082), .A2(n10083), .ZN(n10081) );
  OR2_X1 U7467 ( .A1(n10080), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5992) );
  AND2_X1 U7468 ( .A1(n10081), .A2(n5992), .ZN(n10092) );
  INV_X1 U7469 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8880) );
  MUX2_X1 U7470 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n8880), .S(n10098), .Z(n10093) );
  NAND2_X1 U7471 ( .A1(n10092), .A2(n10093), .ZN(n10091) );
  NAND2_X1 U7472 ( .A1(n10098), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5993) );
  AND2_X1 U7473 ( .A1(n10091), .A2(n5993), .ZN(n5996) );
  NOR2_X1 U7474 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6815), .ZN(n5994) );
  AOI21_X1 U7475 ( .B1(n6815), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5994), .ZN(
        n5995) );
  NAND2_X1 U7476 ( .A1(n5995), .A2(n5996), .ZN(n6013) );
  OAI21_X1 U7477 ( .B1(n5996), .B2(n5995), .A(n6013), .ZN(n5997) );
  AOI22_X1 U7478 ( .A1(n6815), .A2(n10118), .B1(n10124), .B2(n5997), .ZN(n6008) );
  NOR2_X1 U7479 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6815), .ZN(n5998) );
  AOI21_X1 U7480 ( .B1(n6815), .B2(P1_REG1_REG_7__SCAN_IN), .A(n5998), .ZN(
        n6005) );
  INV_X1 U7481 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5999) );
  MUX2_X1 U7482 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n5999), .S(n10098), .Z(n6003)
         );
  INV_X1 U7483 ( .A(n6541), .ZN(n9578) );
  INV_X1 U7484 ( .A(n6508), .ZN(n6001) );
  AOI21_X1 U7485 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6001), .A(n6000), .ZN(
        n9566) );
  XNOR2_X1 U7486 ( .A(n6541), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U7487 ( .A1(n9566), .A2(n9567), .ZN(n9565) );
  OAI21_X1 U7488 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9578), .A(n9565), .ZN(
        n10077) );
  NAND2_X1 U7489 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n10080), .ZN(n6002) );
  OAI21_X1 U7490 ( .B1(n10080), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6002), .ZN(
        n10076) );
  NOR2_X1 U7491 ( .A1(n10077), .A2(n10076), .ZN(n10075) );
  AOI21_X1 U7492 ( .B1(n10080), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10075), .ZN(
        n10089) );
  NAND2_X1 U7493 ( .A1(n6003), .A2(n10089), .ZN(n10088) );
  OAI21_X1 U7494 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10098), .A(n10088), .ZN(
        n6004) );
  NAND2_X1 U7495 ( .A1(n6005), .A2(n6004), .ZN(n6015) );
  OAI21_X1 U7496 ( .B1(n6005), .B2(n6004), .A(n6015), .ZN(n6006) );
  AND2_X1 U7497 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6835) );
  AOI21_X1 U7498 ( .B1(n10120), .B2(n6006), .A(n6835), .ZN(n6007) );
  OAI211_X1 U7499 ( .C1(n10063), .C2(n6009), .A(n6008), .B(n6007), .ZN(
        P1_U3248) );
  NAND2_X1 U7500 ( .A1(n6034), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7501 ( .A(n6010), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7116) );
  INV_X1 U7502 ( .A(n7116), .ZN(n6108) );
  OAI222_X1 U7503 ( .A1(n9968), .A2(n6012), .B1(n9971), .B2(n6011), .C1(n6108), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U7504 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7108) );
  OR2_X1 U7505 ( .A1(n6815), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7506 ( .A1(n6014), .A2(n6013), .ZN(n6022) );
  NOR3_X1 U7507 ( .A1(n9590), .A2(n7108), .A3(n6022), .ZN(n6018) );
  INV_X1 U7508 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6379) );
  OR2_X1 U7509 ( .A1(n6815), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7510 ( .A1(n6016), .A2(n6015), .ZN(n6024) );
  NOR3_X1 U7511 ( .A1(n10106), .A2(n6379), .A3(n6024), .ZN(n6017) );
  NOR3_X1 U7512 ( .A1(n6018), .A2(n10118), .A3(n6017), .ZN(n6032) );
  INV_X1 U7513 ( .A(n6908), .ZN(n6031) );
  OR2_X1 U7514 ( .A1(n6908), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6021) );
  INV_X1 U7515 ( .A(n6021), .ZN(n6023) );
  NAND2_X1 U7516 ( .A1(n6908), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7517 ( .A1(n6019), .A2(n6022), .ZN(n6020) );
  AND2_X1 U7518 ( .A1(n6021), .A2(n6020), .ZN(n6106) );
  AOI211_X1 U7519 ( .C1(n6023), .C2(n6022), .A(n6106), .B(n9590), .ZN(n6029)
         );
  NOR2_X1 U7520 ( .A1(n6908), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6025) );
  OAI22_X1 U7521 ( .A1(n6025), .A2(n6024), .B1(n6379), .B2(n6031), .ZN(n6103)
         );
  AOI211_X1 U7522 ( .C1(n6025), .C2(n6024), .A(n6103), .B(n10106), .ZN(n6028)
         );
  INV_X1 U7523 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6380) );
  NOR2_X1 U7524 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6380), .ZN(n6928) );
  INV_X1 U7525 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6026) );
  NOR2_X1 U7526 ( .A1(n10063), .A2(n6026), .ZN(n6027) );
  NOR4_X1 U7527 ( .A1(n6029), .A2(n6028), .A3(n6928), .A4(n6027), .ZN(n6030)
         );
  OAI21_X1 U7528 ( .B1(n6032), .B2(n6031), .A(n6030), .ZN(P1_U3249) );
  INV_X1 U7529 ( .A(n7257), .ZN(n6036) );
  AOI22_X1 U7530 ( .A1(n8396), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9129), .ZN(n6033) );
  OAI21_X1 U7531 ( .B1(n6036), .B2(n9134), .A(n6033), .ZN(P2_U3348) );
  OR2_X1 U7532 ( .A1(n6156), .A2(n6035), .ZN(n6081) );
  XNOR2_X1 U7533 ( .A(n6081), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10101) );
  INV_X1 U7534 ( .A(n10101), .ZN(n6092) );
  OAI222_X1 U7535 ( .A1(n9968), .A2(n6037), .B1(n9971), .B2(n6036), .C1(n6092), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  OR2_X1 U7536 ( .A1(n10309), .A2(n6575), .ZN(n6042) );
  NOR2_X1 U7537 ( .A1(n5844), .A2(P2_U3152), .ZN(n9128) );
  INV_X1 U7538 ( .A(n6039), .ZN(n7449) );
  AOI21_X1 U7539 ( .B1(n6040), .B2(n9128), .A(n7449), .ZN(n6041) );
  NAND2_X1 U7540 ( .A1(n6042), .A2(n6041), .ZN(n6056) );
  NAND2_X1 U7541 ( .A1(n6056), .A2(n5247), .ZN(n6043) );
  NAND2_X1 U7542 ( .A1(n6043), .A2(n8383), .ZN(n6075) );
  NAND2_X1 U7543 ( .A1(n6075), .A2(n5844), .ZN(n10227) );
  AND2_X1 U7544 ( .A1(P2_U3152), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7545 ( .A1(n6071), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6054) );
  INV_X1 U7546 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6044) );
  MUX2_X1 U7547 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6044), .S(n6071), .Z(n6225)
         );
  NAND2_X1 U7548 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n6070), .ZN(n6053) );
  INV_X1 U7549 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6045) );
  MUX2_X1 U7550 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6045), .S(n6070), .Z(n6261)
         );
  NAND2_X1 U7551 ( .A1(n6068), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6052) );
  INV_X1 U7552 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6046) );
  MUX2_X1 U7553 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6046), .S(n6068), .Z(n6250)
         );
  NAND2_X1 U7554 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n6066), .ZN(n6051) );
  INV_X1 U7555 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6047) );
  MUX2_X1 U7556 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6047), .S(n6066), .Z(n6273)
         );
  NAND2_X1 U7557 ( .A1(n6064), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6050) );
  INV_X1 U7558 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6048) );
  MUX2_X1 U7559 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6048), .S(n6064), .Z(n6238)
         );
  INV_X1 U7560 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10414) );
  MUX2_X1 U7561 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10414), .S(n9991), .Z(n9994)
         );
  INV_X1 U7562 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10412) );
  MUX2_X1 U7563 ( .A(n10412), .B(P2_REG1_REG_1__SCAN_IN), .S(n6062), .Z(n9981)
         );
  NAND3_X1 U7564 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9981), .ZN(n9980) );
  OAI21_X1 U7565 ( .B1(n6062), .B2(n10412), .A(n9980), .ZN(n9995) );
  NAND2_X1 U7566 ( .A1(n9994), .A2(n9995), .ZN(n9993) );
  OAI21_X1 U7567 ( .B1(n6049), .B2(n10414), .A(n9993), .ZN(n6237) );
  NAND2_X1 U7568 ( .A1(n6238), .A2(n6237), .ZN(n6236) );
  NAND2_X1 U7569 ( .A1(n6050), .A2(n6236), .ZN(n6274) );
  NAND2_X1 U7570 ( .A1(n6273), .A2(n6274), .ZN(n6272) );
  NAND2_X1 U7571 ( .A1(n6051), .A2(n6272), .ZN(n6251) );
  NAND2_X1 U7572 ( .A1(n6250), .A2(n6251), .ZN(n6249) );
  NAND2_X1 U7573 ( .A1(n6052), .A2(n6249), .ZN(n6262) );
  NAND2_X1 U7574 ( .A1(n6261), .A2(n6262), .ZN(n6260) );
  NAND2_X1 U7575 ( .A1(n6053), .A2(n6260), .ZN(n6226) );
  NAND2_X1 U7576 ( .A1(n6225), .A2(n6226), .ZN(n6224) );
  AND2_X1 U7577 ( .A1(n6054), .A2(n6224), .ZN(n6058) );
  INV_X1 U7578 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10421) );
  MUX2_X1 U7579 ( .A(n10421), .B(P2_REG1_REG_8__SCAN_IN), .S(n6334), .Z(n6057)
         );
  NOR2_X1 U7580 ( .A1(n6058), .A2(n6057), .ZN(n6326) );
  AND2_X1 U7581 ( .A1(n5247), .A2(n9133), .ZN(n6055) );
  NAND2_X1 U7582 ( .A1(n6056), .A2(n6055), .ZN(n10229) );
  AOI211_X1 U7583 ( .C1(n6058), .C2(n6057), .A(n6326), .B(n10229), .ZN(n6059)
         );
  AOI211_X1 U7584 ( .C1(n10231), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6060), .B(
        n6059), .ZN(n6079) );
  XNOR2_X1 U7585 ( .A(n6334), .B(n6061), .ZN(n6077) );
  NAND2_X1 U7586 ( .A1(n6071), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6073) );
  XNOR2_X1 U7587 ( .A(n6062), .B(n6617), .ZN(n9976) );
  NOR3_X1 U7588 ( .A1(n4830), .A2(n10225), .A3(n9976), .ZN(n9975) );
  XNOR2_X1 U7589 ( .A(n9991), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9988) );
  NOR2_X1 U7590 ( .A1(n9989), .A2(n9988), .ZN(n9987) );
  AOI21_X1 U7591 ( .B1(n9991), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9987), .ZN(
        n6234) );
  NAND2_X1 U7592 ( .A1(n6064), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6063) );
  OAI21_X1 U7593 ( .B1(n6064), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6063), .ZN(
        n6233) );
  NOR2_X1 U7594 ( .A1(n6234), .A2(n6233), .ZN(n6232) );
  NAND2_X1 U7595 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n6066), .ZN(n6065) );
  OAI21_X1 U7596 ( .B1(n6066), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6065), .ZN(
        n6269) );
  NOR2_X1 U7597 ( .A1(n6270), .A2(n6269), .ZN(n6268) );
  NAND2_X1 U7598 ( .A1(n6068), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6067) );
  OAI21_X1 U7599 ( .B1(n6068), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6067), .ZN(
        n6245) );
  NOR2_X1 U7600 ( .A1(n6246), .A2(n6245), .ZN(n6244) );
  AOI21_X1 U7601 ( .B1(n6068), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6244), .ZN(
        n6259) );
  NAND2_X1 U7602 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n6070), .ZN(n6069) );
  OAI21_X1 U7603 ( .B1(n6070), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6069), .ZN(
        n6258) );
  NOR2_X1 U7604 ( .A1(n6259), .A2(n6258), .ZN(n6257) );
  OAI21_X1 U7605 ( .B1(n6071), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6073), .ZN(
        n6221) );
  NOR2_X1 U7606 ( .A1(n6222), .A2(n6221), .ZN(n6220) );
  INV_X1 U7607 ( .A(n6220), .ZN(n6072) );
  NAND2_X1 U7608 ( .A1(n6073), .A2(n6072), .ZN(n6076) );
  NOR2_X1 U7609 ( .A1(n5844), .A2(n9133), .ZN(n6074) );
  NAND2_X1 U7610 ( .A1(n6077), .A2(n6076), .ZN(n6336) );
  OAI211_X1 U7611 ( .C1(n6077), .C2(n6076), .A(n10226), .B(n6336), .ZN(n6078)
         );
  OAI211_X1 U7612 ( .C1(n10227), .C2(n6328), .A(n6079), .B(n6078), .ZN(
        P2_U3253) );
  INV_X1 U7613 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7614 ( .A1(n6081), .A2(n6080), .ZN(n6082) );
  NAND2_X1 U7615 ( .A1(n6082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6083) );
  XNOR2_X1 U7616 ( .A(n6083), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7340) );
  INV_X1 U7617 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6084) );
  INV_X1 U7618 ( .A(n7340), .ZN(n6154) );
  AOI22_X1 U7619 ( .A1(n7340), .A2(n6084), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n6154), .ZN(n6089) );
  NAND2_X1 U7620 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10101), .ZN(n6087) );
  MUX2_X1 U7621 ( .A(n7331), .B(P1_REG2_REG_10__SCAN_IN), .S(n10101), .Z(n6085) );
  INV_X1 U7622 ( .A(n6085), .ZN(n10109) );
  NAND2_X1 U7623 ( .A1(n7116), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6086) );
  INV_X1 U7624 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6917) );
  MUX2_X1 U7625 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6917), .S(n7116), .Z(n6105)
         );
  NAND2_X1 U7626 ( .A1(n6106), .A2(n6105), .ZN(n6104) );
  NAND2_X1 U7627 ( .A1(n6086), .A2(n6104), .ZN(n10110) );
  NAND2_X1 U7628 ( .A1(n10109), .A2(n10110), .ZN(n10108) );
  NAND2_X1 U7629 ( .A1(n6087), .A2(n10108), .ZN(n6088) );
  NOR2_X1 U7630 ( .A1(n6089), .A2(n6088), .ZN(n6164) );
  AOI21_X1 U7631 ( .B1(n6089), .B2(n6088), .A(n6164), .ZN(n6100) );
  NOR2_X1 U7632 ( .A1(n7116), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6090) );
  INV_X1 U7633 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U7634 ( .A1(n7116), .A2(n10221), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6108), .ZN(n6102) );
  NOR2_X1 U7635 ( .A1(n6103), .A2(n6102), .ZN(n6101) );
  NOR2_X1 U7636 ( .A1(n6090), .A2(n6101), .ZN(n10105) );
  MUX2_X1 U7637 ( .A(n6091), .B(P1_REG1_REG_10__SCAN_IN), .S(n10101), .Z(
        n10104) );
  NOR2_X1 U7638 ( .A1(n10105), .A2(n10104), .ZN(n10103) );
  AOI21_X1 U7639 ( .B1(n6091), .B2(n6092), .A(n10103), .ZN(n6094) );
  INV_X1 U7640 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U7641 ( .A1(n7340), .A2(n10057), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n6154), .ZN(n6093) );
  NOR2_X1 U7642 ( .A1(n6094), .A2(n6093), .ZN(n6153) );
  AOI21_X1 U7643 ( .B1(n6094), .B2(n6093), .A(n6153), .ZN(n6095) );
  OR2_X1 U7644 ( .A1(n6095), .A2(n10106), .ZN(n6099) );
  AND2_X1 U7645 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7356) );
  INV_X1 U7646 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6096) );
  NOR2_X1 U7647 ( .A1(n10063), .A2(n6096), .ZN(n6097) );
  AOI211_X1 U7648 ( .C1(n10118), .C2(n7340), .A(n7356), .B(n6097), .ZN(n6098)
         );
  OAI211_X1 U7649 ( .C1(n6100), .C2(n9590), .A(n6099), .B(n6098), .ZN(P1_U3252) );
  AOI21_X1 U7650 ( .B1(n6103), .B2(n6102), .A(n6101), .ZN(n6111) );
  AND2_X1 U7651 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7138) );
  OAI211_X1 U7652 ( .C1(n6106), .C2(n6105), .A(n10124), .B(n6104), .ZN(n6107)
         );
  OAI21_X1 U7653 ( .B1(n9595), .B2(n6108), .A(n6107), .ZN(n6109) );
  AOI211_X1 U7654 ( .C1(n10122), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7138), .B(
        n6109), .ZN(n6110) );
  OAI21_X1 U7655 ( .B1(n6111), .B2(n10106), .A(n6110), .ZN(P1_U3250) );
  INV_X1 U7656 ( .A(n7339), .ZN(n6114) );
  OAI222_X1 U7657 ( .A1(n9968), .A2(n6112), .B1(n9971), .B2(n6114), .C1(n6154), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  OAI222_X1 U7658 ( .A1(P2_U3152), .A2(n6486), .B1(n9139), .B2(n6114), .C1(
        n6113), .C2(n9137), .ZN(P2_U3347) );
  NOR2_X1 U7659 ( .A1(n8505), .A2(n9035), .ZN(n6573) );
  XNOR2_X1 U7660 ( .A(n8212), .B(n6613), .ZN(n6116) );
  INV_X1 U7661 ( .A(n6117), .ZN(n6118) );
  INV_X1 U7662 ( .A(n6149), .ZN(n6119) );
  AOI21_X1 U7663 ( .B1(n6121), .B2(n6120), .A(n6119), .ZN(n6147) );
  XNOR2_X1 U7664 ( .A(n7611), .B(P2_B_REG_SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7665 ( .A1(n7672), .A2(n6122), .ZN(n6123) );
  INV_X1 U7666 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10321) );
  AND2_X1 U7667 ( .A1(n10310), .A2(n10321), .ZN(n6124) );
  INV_X1 U7668 ( .A(n6125), .ZN(n9141) );
  INV_X1 U7669 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10323) );
  NOR2_X1 U7670 ( .A1(n6126), .A2(n6125), .ZN(n10324) );
  NOR4_X1 U7671 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6130) );
  NOR4_X1 U7672 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6129) );
  NOR4_X1 U7673 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6128) );
  NOR4_X1 U7674 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6127) );
  NAND4_X1 U7675 ( .A1(n6130), .A2(n6129), .A3(n6128), .A4(n6127), .ZN(n6136)
         );
  NOR2_X1 U7676 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n6134) );
  NOR4_X1 U7677 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6133) );
  NOR4_X1 U7678 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6132) );
  NOR4_X1 U7679 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6131) );
  NAND4_X1 U7680 ( .A1(n6134), .A2(n6133), .A3(n6132), .A4(n6131), .ZN(n6135)
         );
  OAI21_X1 U7681 ( .B1(n6136), .B2(n6135), .A(n10310), .ZN(n9027) );
  NAND2_X1 U7682 ( .A1(n9028), .A2(n9027), .ZN(n6595) );
  INV_X1 U7683 ( .A(n6595), .ZN(n6137) );
  NAND2_X1 U7684 ( .A1(n9103), .A2(n6137), .ZN(n6144) );
  INV_X1 U7685 ( .A(n6143), .ZN(n6140) );
  NOR2_X1 U7686 ( .A1(n10376), .A2(n6575), .ZN(n6138) );
  INV_X1 U7687 ( .A(n6576), .ZN(n6139) );
  NAND2_X1 U7688 ( .A1(n6140), .A2(n6139), .ZN(n8263) );
  NAND2_X1 U7689 ( .A1(n6575), .A2(n5844), .ZN(n10284) );
  INV_X1 U7690 ( .A(n8263), .ZN(n8287) );
  AND2_X1 U7691 ( .A1(n6600), .A2(n6141), .ZN(n6599) );
  INV_X1 U7692 ( .A(n6599), .ZN(n6142) );
  NAND2_X1 U7693 ( .A1(n9036), .A2(n6141), .ZN(n9025) );
  OAI21_X2 U7694 ( .B1(n6143), .B2(n6142), .A(n10297), .ZN(n8360) );
  NAND2_X1 U7695 ( .A1(n6144), .A2(n9025), .ZN(n6292) );
  NAND2_X1 U7696 ( .A1(n9026), .A2(n6292), .ZN(n6370) );
  AOI22_X1 U7697 ( .A1(n8360), .A2(n6613), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n6370), .ZN(n6145) );
  OAI211_X1 U7698 ( .C1(n6147), .C2(n8362), .A(n6146), .B(n6145), .ZN(P2_U3224) );
  XNOR2_X1 U7699 ( .A(n8212), .B(n6865), .ZN(n6284) );
  NAND2_X1 U7700 ( .A1(n8382), .A2(n8156), .ZN(n6283) );
  XNOR2_X1 U7701 ( .A(n6283), .B(n6284), .ZN(n6285) );
  XNOR2_X1 U7702 ( .A(n6286), .B(n6285), .ZN(n6152) );
  AOI22_X1 U7703 ( .A1(n8318), .A2(n8381), .B1(n8346), .B2(n6578), .ZN(n6151)
         );
  AOI22_X1 U7704 ( .A1(n8360), .A2(n6865), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n6370), .ZN(n6150) );
  OAI211_X1 U7705 ( .C1(n8362), .C2(n6152), .A(n6151), .B(n6150), .ZN(P2_U3239) );
  AOI21_X1 U7706 ( .B1(n6154), .B2(n10057), .A(n6153), .ZN(n6159) );
  NOR2_X1 U7707 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6155) );
  NAND2_X1 U7708 ( .A1(n6156), .A2(n6155), .ZN(n6374) );
  NAND2_X1 U7709 ( .A1(n6374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6157) );
  XNOR2_X1 U7710 ( .A(n6157), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7456) );
  INV_X1 U7711 ( .A(n7456), .ZN(n6399) );
  INV_X1 U7712 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U7713 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6399), .B1(n7456), .B2(
        n10050), .ZN(n6158) );
  NOR2_X1 U7714 ( .A1(n6159), .A2(n6158), .ZN(n6398) );
  AOI21_X1 U7715 ( .B1(n6159), .B2(n6158), .A(n6398), .ZN(n6169) );
  INV_X1 U7716 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7717 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6160) );
  OAI21_X1 U7718 ( .B1(n10063), .B2(n6161), .A(n6160), .ZN(n6162) );
  AOI21_X1 U7719 ( .B1(n7456), .B2(n10118), .A(n6162), .ZN(n6168) );
  NOR2_X1 U7720 ( .A1(n7340), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6163) );
  NOR2_X1 U7721 ( .A1(n6164), .A2(n6163), .ZN(n6166) );
  INV_X1 U7722 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7496) );
  MUX2_X1 U7723 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n7496), .S(n7456), .Z(n6165)
         );
  NAND2_X1 U7724 ( .A1(n6165), .A2(n6166), .ZN(n6403) );
  OAI211_X1 U7725 ( .C1(n6166), .C2(n6165), .A(n10124), .B(n6403), .ZN(n6167)
         );
  OAI211_X1 U7726 ( .C1(n6169), .C2(n10106), .A(n6168), .B(n6167), .ZN(
        P1_U3253) );
  OR2_X1 U7727 ( .A1(n10158), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7728 ( .A1(n9973), .A2(n7613), .ZN(n6170) );
  NOR2_X1 U7729 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n6175) );
  NOR4_X1 U7730 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6174) );
  NOR4_X1 U7731 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6173) );
  NOR4_X1 U7732 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6172) );
  NAND4_X1 U7733 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n6181)
         );
  NOR4_X1 U7734 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6179) );
  NOR4_X1 U7735 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6178) );
  NOR4_X1 U7736 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6177) );
  NOR4_X1 U7737 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6176) );
  NAND4_X1 U7738 ( .A1(n6179), .A2(n6178), .A3(n6177), .A4(n6176), .ZN(n6180)
         );
  NOR2_X1 U7739 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  OR2_X1 U7740 ( .A1(n10158), .A2(n6182), .ZN(n6316) );
  AND2_X1 U7741 ( .A1(n9957), .A2(n6316), .ZN(n6350) );
  INV_X1 U7742 ( .A(n6440), .ZN(n6210) );
  NOR2_X1 U7743 ( .A1(n6210), .A2(n9956), .ZN(n6207) );
  NAND2_X1 U7744 ( .A1(n6183), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6184) );
  NOR2_X1 U7745 ( .A1(n6654), .A2(n9528), .ZN(n10149) );
  NAND2_X1 U7746 ( .A1(n6207), .A2(n10149), .ZN(n6188) );
  NAND2_X1 U7747 ( .A1(n6186), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6187) );
  OR2_X1 U7748 ( .A1(n10205), .A2(n9690), .ZN(n6319) );
  INV_X1 U7749 ( .A(n9251), .ZN(n9218) );
  NOR2_X1 U7750 ( .A1(n6417), .A2(n6189), .ZN(n6191) );
  XNOR2_X1 U7751 ( .A(n6191), .B(n6190), .ZN(n9974) );
  MUX2_X1 U7752 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9974), .S(n6542), .Z(n6666) );
  NAND2_X1 U7753 ( .A1(n7887), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6197) );
  INV_X1 U7754 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10062) );
  OR2_X1 U7755 ( .A1(n6527), .A2(n10062), .ZN(n6196) );
  INV_X1 U7756 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6192) );
  OR2_X1 U7757 ( .A1(n6557), .A2(n6192), .ZN(n6195) );
  INV_X1 U7758 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6193) );
  OR2_X1 U7759 ( .A1(n4477), .A2(n6193), .ZN(n6194) );
  AND2_X4 U7760 ( .A1(n6522), .A2(n6412), .ZN(n8044) );
  NAND2_X1 U7761 ( .A1(n9528), .A2(n9690), .ZN(n9534) );
  INV_X1 U7762 ( .A(n9534), .ZN(n6198) );
  NAND2_X1 U7763 ( .A1(n9536), .A2(n6198), .ZN(n6199) );
  AND2_X2 U7764 ( .A1(n8044), .A2(n6199), .ZN(n7928) );
  INV_X1 U7765 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U7766 ( .A1(n6666), .A2(n4480), .ZN(n6200) );
  OAI21_X1 U7767 ( .B1(n6522), .B2(n6355), .A(n6200), .ZN(n6201) );
  AOI21_X1 U7768 ( .B1(n10138), .B2(n7928), .A(n6201), .ZN(n6205) );
  INV_X1 U7769 ( .A(n6522), .ZN(n6202) );
  AOI22_X1 U7770 ( .A1(n6666), .A2(n8044), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n6202), .ZN(n6203) );
  NAND2_X1 U7771 ( .A1(n6204), .A2(n6203), .ZN(n6413) );
  NAND2_X1 U7772 ( .A1(n6205), .A2(n6413), .ZN(n6414) );
  OAI21_X1 U7773 ( .B1(n6205), .B2(n6413), .A(n6414), .ZN(n6353) );
  INV_X1 U7774 ( .A(n6654), .ZN(n6321) );
  NOR2_X1 U7775 ( .A1(n10000), .A2(n9467), .ZN(n6206) );
  NAND2_X1 U7776 ( .A1(n6353), .A2(n9211), .ZN(n6219) );
  INV_X1 U7777 ( .A(n10149), .ZN(n6208) );
  NOR2_X1 U7778 ( .A1(n9956), .A2(n6208), .ZN(n6209) );
  NAND2_X1 U7779 ( .A1(n6210), .A2(n6209), .ZN(n6525) );
  NAND2_X1 U7780 ( .A1(n6210), .A2(n10204), .ZN(n6523) );
  AND2_X1 U7781 ( .A1(n9467), .A2(n9534), .ZN(n6520) );
  NAND3_X1 U7782 ( .A1(n6525), .A2(n6523), .A3(n6348), .ZN(n6473) );
  NAND3_X1 U7783 ( .A1(n6684), .A2(n9473), .A3(n9690), .ZN(n6665) );
  INV_X1 U7784 ( .A(n6665), .ZN(n6322) );
  NAND2_X1 U7785 ( .A1(n5956), .A2(n6322), .ZN(n6211) );
  NOR2_X1 U7786 ( .A1(n9956), .A2(n6211), .ZN(n6212) );
  INV_X1 U7787 ( .A(n9234), .ZN(n9247) );
  AOI22_X1 U7788 ( .A1(n6431), .A2(P1_REG0_REG_1__SCAN_IN), .B1(n6213), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6217) );
  NOR2_X1 U7789 ( .A1(n6434), .A2(n10213), .ZN(n6214) );
  NOR2_X1 U7790 ( .A1(n6215), .A2(n6214), .ZN(n6216) );
  AOI22_X1 U7791 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n6473), .B1(n9247), .B2(
        n9564), .ZN(n6218) );
  OAI211_X1 U7792 ( .C1(n9218), .C2(n10147), .A(n6219), .B(n6218), .ZN(
        P1_U3230) );
  AOI211_X1 U7793 ( .C1(n6222), .C2(n6221), .A(n6220), .B(n9986), .ZN(n6231)
         );
  NOR2_X1 U7794 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6764), .ZN(n6223) );
  AOI21_X1 U7795 ( .B1(n10231), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6223), .ZN(
        n6228) );
  OAI211_X1 U7796 ( .C1(n6226), .C2(n6225), .A(n10224), .B(n6224), .ZN(n6227)
         );
  OAI211_X1 U7797 ( .C1(n10227), .C2(n6229), .A(n6228), .B(n6227), .ZN(n6230)
         );
  OR2_X1 U7798 ( .A1(n6231), .A2(n6230), .ZN(P2_U3252) );
  AOI211_X1 U7799 ( .C1(n6234), .C2(n6233), .A(n6232), .B(n9986), .ZN(n6243)
         );
  INV_X1 U7800 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6294) );
  NOR2_X1 U7801 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6294), .ZN(n6235) );
  AOI21_X1 U7802 ( .B1(n10231), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6235), .ZN(
        n6240) );
  OAI211_X1 U7803 ( .C1(n6238), .C2(n6237), .A(n10224), .B(n6236), .ZN(n6239)
         );
  OAI211_X1 U7804 ( .C1(n10227), .C2(n6241), .A(n6240), .B(n6239), .ZN(n6242)
         );
  OR2_X1 U7805 ( .A1(n6243), .A2(n6242), .ZN(P2_U3248) );
  AOI211_X1 U7806 ( .C1(n6246), .C2(n6245), .A(n6244), .B(n9986), .ZN(n6256)
         );
  NOR2_X1 U7807 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6247), .ZN(n6248) );
  AOI21_X1 U7808 ( .B1(n10231), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6248), .ZN(
        n6253) );
  OAI211_X1 U7809 ( .C1(n6251), .C2(n6250), .A(n10224), .B(n6249), .ZN(n6252)
         );
  OAI211_X1 U7810 ( .C1(n10227), .C2(n6254), .A(n6253), .B(n6252), .ZN(n6255)
         );
  OR2_X1 U7811 ( .A1(n6256), .A2(n6255), .ZN(P2_U3250) );
  AOI211_X1 U7812 ( .C1(n6259), .C2(n6258), .A(n6257), .B(n9986), .ZN(n6267)
         );
  AND2_X1 U7813 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8341) );
  AOI21_X1 U7814 ( .B1(n10231), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8341), .ZN(
        n6264) );
  OAI211_X1 U7815 ( .C1(n6262), .C2(n6261), .A(n10224), .B(n6260), .ZN(n6263)
         );
  OAI211_X1 U7816 ( .C1(n10227), .C2(n6265), .A(n6264), .B(n6263), .ZN(n6266)
         );
  OR2_X1 U7817 ( .A1(n6267), .A2(n6266), .ZN(P2_U3251) );
  AOI211_X1 U7818 ( .C1(n6270), .C2(n6269), .A(n6268), .B(n9986), .ZN(n6279)
         );
  NAND2_X1 U7819 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6311) );
  INV_X1 U7820 ( .A(n6311), .ZN(n6271) );
  AOI21_X1 U7821 ( .B1(n10231), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6271), .ZN(
        n6276) );
  OAI211_X1 U7822 ( .C1(n6274), .C2(n6273), .A(n10224), .B(n6272), .ZN(n6275)
         );
  OAI211_X1 U7823 ( .C1(n10227), .C2(n6277), .A(n6276), .B(n6275), .ZN(n6278)
         );
  OR2_X1 U7824 ( .A1(n6279), .A2(n6278), .ZN(P2_U3249) );
  INV_X1 U7825 ( .A(n7455), .ZN(n6280) );
  INV_X1 U7826 ( .A(n6497), .ZN(n8416) );
  OAI222_X1 U7827 ( .A1(n9137), .A2(n6396), .B1(n9139), .B2(n6280), .C1(
        P2_U3152), .C2(n8416), .ZN(P2_U3346) );
  OAI222_X1 U7828 ( .A1(n9968), .A2(n6281), .B1(n9971), .B2(n6280), .C1(
        P1_U3084), .C2(n6399), .ZN(P1_U3341) );
  INV_X1 U7829 ( .A(n9563), .ZN(n9562) );
  NAND2_X1 U7830 ( .A1(n10138), .A2(n9562), .ZN(n6282) );
  OAI21_X1 U7831 ( .B1(n9562), .B2(n5051), .A(n6282), .ZN(P1_U3555) );
  XNOR2_X1 U7832 ( .A(n8212), .B(n10344), .ZN(n6303) );
  NAND2_X1 U7833 ( .A1(n8381), .A2(n4486), .ZN(n6301) );
  XNOR2_X1 U7834 ( .A(n6303), .B(n6301), .ZN(n6299) );
  XNOR2_X1 U7835 ( .A(n6300), .B(n6299), .ZN(n6298) );
  NAND2_X1 U7836 ( .A1(n6288), .A2(n6287), .ZN(n6290) );
  NOR2_X1 U7837 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  NAND2_X1 U7838 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  OAI22_X1 U7839 ( .A1(n8355), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n6294), .ZN(n6296) );
  OAI22_X1 U7840 ( .A1(n8357), .A2(n6850), .B1(n10344), .B2(n8338), .ZN(n6295)
         );
  AOI211_X1 U7841 ( .C1(n8346), .C2(n8382), .A(n6296), .B(n6295), .ZN(n6297)
         );
  OAI21_X1 U7842 ( .B1(n6298), .B2(n8362), .A(n6297), .ZN(P2_U3220) );
  INV_X1 U7843 ( .A(n6301), .ZN(n6302) );
  NAND2_X1 U7844 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  XNOR2_X1 U7845 ( .A(n8212), .B(n10351), .ZN(n6308) );
  INV_X1 U7846 ( .A(n6308), .ZN(n6306) );
  AND2_X1 U7847 ( .A1(n8380), .A2(n8156), .ZN(n6307) );
  INV_X1 U7848 ( .A(n6307), .ZN(n6305) );
  NAND2_X1 U7849 ( .A1(n6306), .A2(n6305), .ZN(n6742) );
  INV_X1 U7850 ( .A(n6742), .ZN(n6309) );
  AND2_X1 U7851 ( .A1(n6308), .A2(n6307), .ZN(n6740) );
  NOR2_X1 U7852 ( .A1(n6309), .A2(n6740), .ZN(n6310) );
  XNOR2_X1 U7853 ( .A(n6741), .B(n6310), .ZN(n6315) );
  OAI21_X1 U7854 ( .B1(n8355), .B2(n10298), .A(n6311), .ZN(n6313) );
  OAI22_X1 U7855 ( .A1(n8357), .A2(n10285), .B1(n10351), .B2(n8338), .ZN(n6312) );
  AOI211_X1 U7856 ( .C1(n8346), .C2(n8381), .A(n6313), .B(n6312), .ZN(n6314)
         );
  OAI21_X1 U7857 ( .B1(n6315), .B2(n8362), .A(n6314), .ZN(P2_U3232) );
  INV_X1 U7858 ( .A(n6316), .ZN(n6317) );
  NOR2_X1 U7859 ( .A1(n9957), .A2(n6317), .ZN(n6318) );
  AND2_X1 U7860 ( .A1(n6320), .A2(n6319), .ZN(n6349) );
  NOR2_X1 U7861 ( .A1(n10138), .A2(n10147), .ZN(n10133) );
  AND2_X1 U7862 ( .A1(n10138), .A2(n10147), .ZN(n9478) );
  OR2_X1 U7863 ( .A1(n10133), .A2(n9478), .ZN(n9300) );
  NOR2_X1 U7864 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  AOI22_X1 U7865 ( .A1(n9300), .A2(n6323), .B1(n10140), .B2(n9564), .ZN(n6658)
         );
  OAI21_X1 U7866 ( .B1(n10147), .B2(n6654), .A(n6658), .ZN(n6351) );
  NAND2_X1 U7867 ( .A1(n6351), .A2(n10212), .ZN(n6324) );
  OAI21_X1 U7868 ( .B1(n10212), .B2(n6192), .A(n6324), .ZN(P1_U3454) );
  NAND2_X1 U7869 ( .A1(n8384), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6329) );
  INV_X1 U7870 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6325) );
  MUX2_X1 U7871 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6325), .S(n8384), .Z(n8391)
         );
  INV_X1 U7872 ( .A(n6326), .ZN(n6327) );
  OAI21_X1 U7873 ( .B1(n10421), .B2(n6328), .A(n6327), .ZN(n8390) );
  NAND2_X1 U7874 ( .A1(n8391), .A2(n8390), .ZN(n8389) );
  NAND2_X1 U7875 ( .A1(n6329), .A2(n8389), .ZN(n8403) );
  INV_X1 U7876 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6330) );
  MUX2_X1 U7877 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6330), .S(n8396), .Z(n8402)
         );
  NAND2_X1 U7878 ( .A1(n8403), .A2(n8402), .ZN(n8401) );
  NAND2_X1 U7879 ( .A1(n8396), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6332) );
  INV_X1 U7880 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10425) );
  MUX2_X1 U7881 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10425), .S(n6486), .Z(n6331) );
  AOI21_X1 U7882 ( .B1(n8401), .B2(n6332), .A(n6331), .ZN(n6495) );
  NAND3_X1 U7883 ( .A1(n8401), .A2(n6332), .A3(n6331), .ZN(n6333) );
  NAND2_X1 U7884 ( .A1(n10224), .A2(n6333), .ZN(n6347) );
  NAND2_X1 U7885 ( .A1(n6334), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7886 ( .A1(n6336), .A2(n6335), .ZN(n8386) );
  OR2_X1 U7887 ( .A1(n8384), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7888 ( .A1(n8384), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6338) );
  AND2_X1 U7889 ( .A1(n6337), .A2(n6338), .ZN(n8387) );
  NAND2_X1 U7890 ( .A1(n8386), .A2(n8387), .ZN(n8385) );
  NAND2_X1 U7891 ( .A1(n8385), .A2(n6338), .ZN(n8398) );
  XNOR2_X1 U7892 ( .A(n8396), .B(n6339), .ZN(n8399) );
  NAND2_X1 U7893 ( .A1(n8398), .A2(n8399), .ZN(n8397) );
  NAND2_X1 U7894 ( .A1(n8396), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6340) );
  MUX2_X1 U7895 ( .A(n7087), .B(P2_REG2_REG_11__SCAN_IN), .S(n6486), .Z(n6341)
         );
  NAND2_X1 U7896 ( .A1(n6342), .A2(n6341), .ZN(n6488) );
  OAI21_X1 U7897 ( .B1(n6342), .B2(n6341), .A(n6488), .ZN(n6345) );
  NOR2_X1 U7898 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5411), .ZN(n7187) );
  AOI21_X1 U7899 ( .B1(n10231), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7187), .ZN(
        n6343) );
  OAI21_X1 U7900 ( .B1(n10227), .B2(n6486), .A(n6343), .ZN(n6344) );
  AOI21_X1 U7901 ( .B1(n10226), .B2(n6345), .A(n6344), .ZN(n6346) );
  OAI21_X1 U7902 ( .B1(n6495), .B2(n6347), .A(n6346), .ZN(P2_U3256) );
  INV_X1 U7903 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U7904 ( .A1(n6351), .A2(n10223), .ZN(n6352) );
  OAI21_X1 U7905 ( .B1(n10223), .B2(n10071), .A(n6352), .ZN(P1_U3523) );
  MUX2_X1 U7906 ( .A(n6355), .B(n6353), .S(n10065), .Z(n6356) );
  NOR2_X1 U7907 ( .A1(n10065), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6354) );
  OR2_X1 U7908 ( .A1(n6354), .A2(n5956), .ZN(n10068) );
  NAND2_X1 U7909 ( .A1(n10068), .A2(n6355), .ZN(n10066) );
  OAI211_X1 U7910 ( .C1(n6356), .C2(n10068), .A(n9562), .B(n10066), .ZN(n9581)
         );
  OAI21_X1 U7911 ( .B1(n6359), .B2(n6358), .A(n6357), .ZN(n6360) );
  INV_X1 U7912 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6432) );
  OAI22_X1 U7913 ( .A1(n10106), .A2(n6360), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6432), .ZN(n6366) );
  OAI211_X1 U7914 ( .C1(n6363), .C2(n6362), .A(n10124), .B(n6361), .ZN(n6364)
         );
  OAI21_X1 U7915 ( .B1(n9595), .B2(n6448), .A(n6364), .ZN(n6365) );
  AOI211_X1 U7916 ( .C1(n10122), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n6366), .B(
        n6365), .ZN(n6367) );
  NAND2_X1 U7917 ( .A1(n9581), .A2(n6367), .ZN(P1_U3243) );
  OR2_X1 U7918 ( .A1(n8362), .A2(n8211), .ZN(n8345) );
  INV_X1 U7919 ( .A(n8345), .ZN(n8313) );
  INV_X1 U7920 ( .A(n6368), .ZN(n6369) );
  AOI22_X1 U7921 ( .A1(n8318), .A2(n6578), .B1(n8313), .B2(n6369), .ZN(n6373)
         );
  OAI21_X1 U7922 ( .B1(n4834), .B2(n8156), .A(n6607), .ZN(n6371) );
  AOI22_X1 U7923 ( .A1(n8336), .A2(n6371), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n6370), .ZN(n6372) );
  OAI211_X1 U7924 ( .C1(n8338), .C2(n4834), .A(n6373), .B(n6372), .ZN(P2_U3234) );
  INV_X1 U7925 ( .A(n7522), .ZN(n6377) );
  NAND2_X1 U7926 ( .A1(n6477), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6375) );
  XNOR2_X1 U7927 ( .A(n6375), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7523) );
  INV_X1 U7928 ( .A(n7523), .ZN(n6642) );
  OAI222_X1 U7929 ( .A1(n9968), .A2(n6376), .B1(n9971), .B2(n6377), .C1(n6642), 
        .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U7930 ( .A(n6692), .ZN(n6688) );
  OAI222_X1 U7931 ( .A1(n9137), .A2(n6378), .B1(n9139), .B2(n6377), .C1(n6688), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  NAND2_X1 U7932 ( .A1(n6431), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6385) );
  OR2_X1 U7933 ( .A1(n4479), .A2(n6379), .ZN(n6384) );
  NAND2_X1 U7934 ( .A1(n6823), .A2(n6380), .ZN(n6381) );
  NAND2_X1 U7935 ( .A1(n6920), .A2(n6381), .ZN(n7107) );
  OR2_X1 U7936 ( .A1(n6527), .A2(n7107), .ZN(n6383) );
  OR2_X1 U7937 ( .A1(n4476), .A2(n7108), .ZN(n6382) );
  MUX2_X1 U7938 ( .A(n6386), .B(n7291), .S(n9562), .Z(n6387) );
  INV_X1 U7939 ( .A(n6387), .ZN(P1_U3563) );
  NAND2_X1 U7940 ( .A1(n6431), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6395) );
  OR2_X1 U7941 ( .A1(n4478), .A2(n10050), .ZN(n6394) );
  INV_X1 U7942 ( .A(n7274), .ZN(n6389) );
  NAND2_X1 U7943 ( .A1(n6389), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7473) );
  INV_X1 U7944 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7945 ( .A1(n7274), .A2(n6390), .ZN(n6391) );
  NAND2_X1 U7946 ( .A1(n7473), .A2(n6391), .ZN(n7495) );
  OR2_X1 U7947 ( .A1(n6527), .A2(n7495), .ZN(n6393) );
  OR2_X1 U7948 ( .A1(n4476), .A2(n7496), .ZN(n6392) );
  MUX2_X1 U7949 ( .A(n6396), .B(n7619), .S(n9562), .Z(n6397) );
  INV_X1 U7950 ( .A(n6397), .ZN(P1_U3567) );
  AOI21_X1 U7951 ( .B1(n10050), .B2(n6399), .A(n6398), .ZN(n6401) );
  INV_X1 U7952 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7476) );
  AOI22_X1 U7953 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n6642), .B1(n7523), .B2(
        n7476), .ZN(n6400) );
  NOR2_X1 U7954 ( .A1(n6401), .A2(n6400), .ZN(n6641) );
  AOI21_X1 U7955 ( .B1(n6401), .B2(n6400), .A(n6641), .ZN(n6411) );
  AND2_X1 U7956 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7541) );
  NOR2_X1 U7957 ( .A1(n9595), .A2(n6642), .ZN(n6402) );
  AOI211_X1 U7958 ( .C1(n10122), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7541), .B(
        n6402), .ZN(n6410) );
  NAND2_X1 U7959 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7456), .ZN(n6404) );
  NAND2_X1 U7960 ( .A1(n6404), .A2(n6403), .ZN(n6408) );
  INV_X1 U7961 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6405) );
  MUX2_X1 U7962 ( .A(n6405), .B(P1_REG2_REG_13__SCAN_IN), .S(n7523), .Z(n6406)
         );
  INV_X1 U7963 ( .A(n6406), .ZN(n6407) );
  NAND2_X1 U7964 ( .A1(n6407), .A2(n6408), .ZN(n6646) );
  OAI211_X1 U7965 ( .C1(n6408), .C2(n6407), .A(n10124), .B(n6646), .ZN(n6409)
         );
  OAI211_X1 U7966 ( .C1(n6411), .C2(n10106), .A(n6410), .B(n6409), .ZN(
        P1_U3254) );
  NAND2_X1 U7967 ( .A1(n9564), .A2(n7347), .ZN(n6424) );
  OR2_X1 U7968 ( .A1(n6792), .A2(n6416), .ZN(n6422) );
  NAND2_X1 U7969 ( .A1(n6542), .A2(n6417), .ZN(n6506) );
  OR2_X1 U7970 ( .A1(n6506), .A2(n6418), .ZN(n6421) );
  OR2_X1 U7971 ( .A1(n6542), .A2(n6419), .ZN(n6420) );
  OR2_X1 U7972 ( .A1(n10171), .A2(n7946), .ZN(n6423) );
  NAND2_X1 U7973 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  XNOR2_X1 U7974 ( .A(n6425), .B(n7947), .ZN(n6427) );
  NAND2_X1 U7975 ( .A1(n6426), .A2(n6427), .ZN(n6458) );
  INV_X1 U7976 ( .A(n6426), .ZN(n6429) );
  INV_X1 U7977 ( .A(n6427), .ZN(n6428) );
  NAND2_X1 U7978 ( .A1(n6429), .A2(n6428), .ZN(n6459) );
  NAND2_X1 U7979 ( .A1(n6458), .A2(n6459), .ZN(n6430) );
  INV_X1 U7980 ( .A(n10171), .ZN(n6667) );
  AOI22_X1 U7981 ( .A1(n9564), .A2(n7928), .B1(n6667), .B2(n7347), .ZN(n6457)
         );
  XNOR2_X1 U7982 ( .A(n6430), .B(n6457), .ZN(n6445) );
  NAND2_X1 U7983 ( .A1(n6431), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6438) );
  OR2_X1 U7984 ( .A1(n6527), .A2(n6432), .ZN(n6437) );
  OR2_X1 U7985 ( .A1(n4477), .A2(n6725), .ZN(n6436) );
  OR2_X1 U7986 ( .A1(n4478), .A2(n10215), .ZN(n6435) );
  NAND4_X2 U7987 ( .A1(n6438), .A2(n6437), .A3(n6436), .A4(n6435), .ZN(n10139)
         );
  INV_X1 U7988 ( .A(n10139), .ZN(n9485) );
  INV_X1 U7989 ( .A(n10138), .ZN(n6441) );
  OR3_X1 U7990 ( .A1(n9956), .A2(n5956), .A3(n6665), .ZN(n9539) );
  INV_X1 U7991 ( .A(n9539), .ZN(n6439) );
  NAND2_X1 U7992 ( .A1(n6440), .A2(n6439), .ZN(n9245) );
  OAI22_X1 U7993 ( .A1(n9485), .A2(n9234), .B1(n6441), .B2(n9245), .ZN(n6443)
         );
  NOR2_X1 U7994 ( .A1(n9218), .A2(n10171), .ZN(n6442) );
  AOI211_X1 U7995 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n6473), .A(n6443), .B(
        n6442), .ZN(n6444) );
  OAI21_X1 U7996 ( .B1(n6445), .B2(n9253), .A(n6444), .ZN(P1_U3220) );
  OR2_X1 U7997 ( .A1(n6792), .A2(n6446), .ZN(n6451) );
  OR2_X1 U7998 ( .A1(n6506), .A2(n6447), .ZN(n6450) );
  OR2_X1 U7999 ( .A1(n6542), .A2(n6448), .ZN(n6449) );
  AND3_X2 U8000 ( .A1(n6451), .A2(n6450), .A3(n6449), .ZN(n10176) );
  NAND2_X1 U8001 ( .A1(n10139), .A2(n7347), .ZN(n6453) );
  OR2_X1 U8002 ( .A1(n10176), .A2(n7946), .ZN(n6452) );
  NAND2_X1 U8003 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  XNOR2_X1 U8004 ( .A(n6454), .B(n8047), .ZN(n6456) );
  INV_X1 U8005 ( .A(n10176), .ZN(n9484) );
  AOI22_X1 U8006 ( .A1(n10139), .A2(n7928), .B1(n9484), .B2(n7347), .ZN(n6455)
         );
  NAND2_X1 U8007 ( .A1(n6456), .A2(n6455), .ZN(n6515) );
  AND2_X1 U8008 ( .A1(n4514), .A2(n6515), .ZN(n6462) );
  NAND2_X1 U8009 ( .A1(n6458), .A2(n6457), .ZN(n6460) );
  NAND2_X1 U8010 ( .A1(n6461), .A2(n6462), .ZN(n6516) );
  OAI21_X1 U8011 ( .B1(n6462), .B2(n6461), .A(n6516), .ZN(n6463) );
  NAND2_X1 U8012 ( .A1(n6463), .A2(n9211), .ZN(n6475) );
  INV_X1 U8013 ( .A(n9564), .ZN(n6471) );
  NAND2_X1 U8014 ( .A1(n6431), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6469) );
  INV_X1 U8015 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6464) );
  OR2_X1 U8016 ( .A1(n4479), .A2(n6464), .ZN(n6468) );
  OR2_X1 U8017 ( .A1(n4476), .A2(n6465), .ZN(n6467) );
  OR2_X1 U8018 ( .A1(n6527), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6466) );
  INV_X1 U8019 ( .A(n9561), .ZN(n6470) );
  OAI22_X1 U8020 ( .A1(n6471), .A2(n9245), .B1(n6470), .B2(n9234), .ZN(n6472)
         );
  AOI21_X1 U8021 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6473), .A(n6472), .ZN(
        n6474) );
  OAI211_X1 U8022 ( .C1(n10176), .C2(n9218), .A(n6475), .B(n6474), .ZN(
        P1_U3235) );
  INV_X1 U8023 ( .A(n7553), .ZN(n6482) );
  INV_X1 U8024 ( .A(n6957), .ZN(n6960) );
  OAI222_X1 U8025 ( .A1(n9137), .A2(n6476), .B1(n9139), .B2(n6482), .C1(n6960), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U8026 ( .A1(n6478), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6481) );
  INV_X1 U8027 ( .A(n6478), .ZN(n6480) );
  NAND2_X1 U8028 ( .A1(n6480), .A2(n6479), .ZN(n6483) );
  OAI222_X1 U8029 ( .A1(n9968), .A2(n8891), .B1(n9971), .B2(n6482), .C1(n7056), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8030 ( .A(n7694), .ZN(n6639) );
  NAND2_X1 U8031 ( .A1(n6483), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6484) );
  XNOR2_X1 U8032 ( .A(n6484), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U8033 ( .A1(n10117), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n7452), .ZN(n6485) );
  OAI21_X1 U8034 ( .B1(n6639), .B2(n9971), .A(n6485), .ZN(P1_U3338) );
  NAND2_X1 U8035 ( .A1(n6486), .A2(n7087), .ZN(n6487) );
  XNOR2_X1 U8036 ( .A(n6497), .B(n6489), .ZN(n8414) );
  NAND2_X1 U8037 ( .A1(n8415), .A2(n8414), .ZN(n8413) );
  NAND2_X1 U8038 ( .A1(n6497), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6490) );
  NOR2_X1 U8039 ( .A1(n6692), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6491) );
  AOI21_X1 U8040 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n6692), .A(n6491), .ZN(
        n6492) );
  NAND2_X1 U8041 ( .A1(n6493), .A2(n6492), .ZN(n6691) );
  OAI21_X1 U8042 ( .B1(n6493), .B2(n6492), .A(n6691), .ZN(n6503) );
  AND2_X1 U8043 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7376) );
  AOI21_X1 U8044 ( .B1(n10231), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7376), .ZN(
        n6494) );
  OAI21_X1 U8045 ( .B1(n10227), .B2(n6688), .A(n6494), .ZN(n6502) );
  INV_X1 U8046 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10428) );
  AOI21_X1 U8047 ( .B1(n6496), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6495), .ZN(
        n8409) );
  MUX2_X1 U8048 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10428), .S(n6497), .Z(n8408) );
  AND2_X1 U8049 ( .A1(n8409), .A2(n8408), .ZN(n8410) );
  AOI21_X1 U8050 ( .B1(n10428), .B2(n8416), .A(n8410), .ZN(n6499) );
  INV_X1 U8051 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U8052 ( .A1(n6692), .A2(n10038), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n6688), .ZN(n6498) );
  NOR2_X1 U8053 ( .A1(n6499), .A2(n6498), .ZN(n6687) );
  AOI21_X1 U8054 ( .B1(n6499), .B2(n6498), .A(n6687), .ZN(n6500) );
  NOR2_X1 U8055 ( .A1(n6500), .A2(n10229), .ZN(n6501) );
  AOI211_X1 U8056 ( .C1(n10226), .C2(n6503), .A(n6502), .B(n6501), .ZN(n6504)
         );
  INV_X1 U8057 ( .A(n6504), .ZN(P2_U3258) );
  NAND2_X1 U8058 ( .A1(n9561), .A2(n7347), .ZN(n6513) );
  OR2_X1 U8059 ( .A1(n6792), .A2(n6505), .ZN(n6511) );
  OR2_X1 U8060 ( .A1(n6506), .A2(n6507), .ZN(n6510) );
  OR2_X1 U8061 ( .A1(n6542), .A2(n6508), .ZN(n6509) );
  OR2_X1 U8062 ( .A1(n6681), .A2(n7946), .ZN(n6512) );
  NAND2_X1 U8063 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  XNOR2_X1 U8064 ( .A(n6514), .B(n7947), .ZN(n6549) );
  AOI22_X1 U8065 ( .A1(n9561), .A2(n7928), .B1(n6731), .B2(n7347), .ZN(n6550)
         );
  XNOR2_X1 U8066 ( .A(n6549), .B(n6550), .ZN(n6518) );
  NAND2_X1 U8067 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  NAND2_X1 U8068 ( .A1(n6517), .A2(n6518), .ZN(n6552) );
  OAI21_X1 U8069 ( .B1(n6518), .B2(n6517), .A(n6552), .ZN(n6538) );
  NOR2_X1 U8070 ( .A1(n6520), .A2(n6519), .ZN(n6521) );
  NAND3_X1 U8071 ( .A1(n6523), .A2(n6522), .A3(n6521), .ZN(n6524) );
  NAND2_X1 U8072 ( .A1(n6524), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6526) );
  NAND2_X1 U8073 ( .A1(n6526), .A2(n6525), .ZN(n9203) );
  NOR2_X1 U8074 ( .A1(n9249), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8075 ( .A1(n6431), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6532) );
  OR2_X1 U8076 ( .A1(n4476), .A2(n6710), .ZN(n6531) );
  XNOR2_X1 U8077 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6709) );
  OR2_X1 U8078 ( .A1(n6527), .A2(n6709), .ZN(n6530) );
  INV_X1 U8079 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6528) );
  OR2_X1 U8080 ( .A1(n4479), .A2(n6528), .ZN(n6529) );
  NAND4_X1 U8081 ( .A1(n6532), .A2(n6531), .A3(n6530), .A4(n6529), .ZN(n9560)
         );
  INV_X1 U8082 ( .A(n9560), .ZN(n6898) );
  NAND2_X1 U8083 ( .A1(n9251), .A2(n6731), .ZN(n6535) );
  AOI21_X1 U8084 ( .B1(n9236), .B2(n10139), .A(n6533), .ZN(n6534) );
  OAI211_X1 U8085 ( .C1(n6898), .C2(n9234), .A(n6535), .B(n6534), .ZN(n6536)
         );
  AOI211_X1 U8086 ( .C1(n6538), .C2(n9211), .A(n6537), .B(n6536), .ZN(n6539)
         );
  INV_X1 U8087 ( .A(n6539), .ZN(P1_U3216) );
  NAND2_X1 U8088 ( .A1(n9560), .A2(n7347), .ZN(n6547) );
  OR2_X1 U8089 ( .A1(n6792), .A2(n6540), .ZN(n6545) );
  OR2_X1 U8090 ( .A1(n8094), .A2(n8864), .ZN(n6544) );
  OR2_X1 U8091 ( .A1(n6542), .A2(n6541), .ZN(n6543) );
  OR2_X1 U8092 ( .A1(n10182), .A2(n7946), .ZN(n6546) );
  NAND2_X1 U8093 ( .A1(n6547), .A2(n6546), .ZN(n6548) );
  INV_X1 U8094 ( .A(n10182), .ZN(n6882) );
  AOI22_X1 U8095 ( .A1(n9560), .A2(n7928), .B1(n6882), .B2(n7347), .ZN(n6776)
         );
  XNOR2_X1 U8096 ( .A(n6775), .B(n6776), .ZN(n6554) );
  INV_X1 U8097 ( .A(n6549), .ZN(n6551) );
  NAND2_X1 U8098 ( .A1(n6551), .A2(n6550), .ZN(n6555) );
  AND2_X1 U8099 ( .A1(n6554), .A2(n6555), .ZN(n6553) );
  NAND2_X1 U8100 ( .A1(n6553), .A2(n6552), .ZN(n6892) );
  NAND2_X1 U8101 ( .A1(n6892), .A2(n9211), .ZN(n6572) );
  AOI21_X1 U8102 ( .B1(n6552), .B2(n6555), .A(n6554), .ZN(n6571) );
  INV_X1 U8103 ( .A(n6709), .ZN(n6569) );
  NAND2_X1 U8104 ( .A1(n7992), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6565) );
  INV_X1 U8105 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6556) );
  OR2_X1 U8106 ( .A1(n4479), .A2(n6556), .ZN(n6564) );
  INV_X1 U8107 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6558) );
  OR2_X1 U8108 ( .A1(n6557), .A2(n6558), .ZN(n6563) );
  INV_X1 U8109 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U8110 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6559) );
  NAND2_X1 U8111 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  NAND2_X1 U8112 ( .A1(n6782), .A2(n6561), .ZN(n6899) );
  OR2_X1 U8113 ( .A1(n6527), .A2(n6899), .ZN(n6562) );
  INV_X1 U8114 ( .A(n9559), .ZN(n7040) );
  NAND2_X1 U8115 ( .A1(n9251), .A2(n6882), .ZN(n6567) );
  AND2_X1 U8116 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9570) );
  AOI21_X1 U8117 ( .B1(n9236), .B2(n9561), .A(n9570), .ZN(n6566) );
  OAI211_X1 U8118 ( .C1(n7040), .C2(n9234), .A(n6567), .B(n6566), .ZN(n6568)
         );
  AOI21_X1 U8119 ( .B1(n6569), .B2(n9203), .A(n6568), .ZN(n6570) );
  OAI21_X1 U8120 ( .B1(n6572), .B2(n6571), .A(n6570), .ZN(P1_U3228) );
  NAND2_X1 U8121 ( .A1(n6573), .A2(n6600), .ZN(n6574) );
  OAI21_X1 U8122 ( .B1(n6576), .B2(n6575), .A(n6574), .ZN(n6577) );
  NAND2_X1 U8123 ( .A1(n6577), .A2(n10326), .ZN(n10241) );
  INV_X1 U8124 ( .A(n10241), .ZN(n8646) );
  NAND2_X1 U8125 ( .A1(n6578), .A2(n6613), .ZN(n6579) );
  NAND2_X1 U8126 ( .A1(n6610), .A2(n6579), .ZN(n6581) );
  NAND2_X1 U8127 ( .A1(n6659), .A2(n10333), .ZN(n6580) );
  NAND2_X1 U8128 ( .A1(n6581), .A2(n6580), .ZN(n6859) );
  NAND2_X1 U8129 ( .A1(n6582), .A2(n6859), .ZN(n6584) );
  NAND2_X1 U8130 ( .A1(n6586), .A2(n10338), .ZN(n6583) );
  XNOR2_X1 U8131 ( .A(n6847), .B(n6846), .ZN(n10348) );
  OAI22_X1 U8132 ( .A1(n6850), .A2(n10284), .B1(n6586), .B2(n10286), .ZN(n6594) );
  NAND3_X1 U8133 ( .A1(n6587), .A2(n6846), .A3(n6588), .ZN(n6592) );
  NAND2_X1 U8134 ( .A1(n4573), .A2(n6589), .ZN(n6590) );
  AOI21_X1 U8135 ( .B1(n10279), .B2(n6592), .A(n10281), .ZN(n6593) );
  AOI211_X1 U8136 ( .C1(n8646), .C2(n10348), .A(n6594), .B(n6593), .ZN(n10345)
         );
  NOR2_X1 U8137 ( .A1(n9103), .A2(n6595), .ZN(n6596) );
  NAND2_X1 U8138 ( .A1(n9026), .A2(n6596), .ZN(n6602) );
  INV_X2 U8139 ( .A(n10299), .ZN(n10308) );
  NAND2_X1 U8140 ( .A1(n9036), .A2(n6597), .ZN(n6611) );
  INV_X1 U8141 ( .A(n6611), .ZN(n6598) );
  NAND2_X1 U8142 ( .A1(n6864), .A2(n10338), .ZN(n10293) );
  XNOR2_X1 U8143 ( .A(n10293), .B(n10344), .ZN(n6601) );
  NAND2_X1 U8144 ( .A1(n6601), .A2(n10295), .ZN(n10343) );
  OR2_X1 U8145 ( .A1(n6602), .A2(n4573), .ZN(n10304) );
  OAI22_X1 U8146 ( .A1(n8627), .A2(n10344), .B1(n10343), .B2(n10304), .ZN(
        n6603) );
  AOI21_X1 U8147 ( .B1(n10251), .B2(n10348), .A(n6603), .ZN(n6606) );
  OAI22_X1 U8148 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n10297), .B1(n5269), .B2(
        n10299), .ZN(n6604) );
  INV_X1 U8149 ( .A(n6604), .ZN(n6605) );
  OAI211_X1 U8150 ( .C1(n10345), .C2(n10308), .A(n6606), .B(n6605), .ZN(
        P2_U3293) );
  XNOR2_X1 U8151 ( .A(n6607), .B(n6609), .ZN(n6608) );
  XOR2_X1 U8152 ( .A(n6610), .B(n6609), .Z(n10331) );
  NAND2_X1 U8153 ( .A1(n10241), .A2(n6611), .ZN(n6612) );
  NOR2_X1 U8154 ( .A1(n10331), .A2(n8639), .ZN(n6621) );
  NOR2_X1 U8155 ( .A1(n8627), .A2(n10333), .ZN(n6620) );
  NAND2_X1 U8156 ( .A1(n6613), .A2(n6661), .ZN(n6614) );
  NAND2_X1 U8157 ( .A1(n10295), .A2(n6614), .ZN(n6615) );
  OR2_X1 U8158 ( .A1(n6615), .A2(n6864), .ZN(n10332) );
  INV_X1 U8159 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6616) );
  OAI22_X1 U8160 ( .A1(n10304), .A2(n10332), .B1(n6616), .B2(n10297), .ZN(
        n6619) );
  NOR2_X1 U8161 ( .A1(n10299), .A2(n6617), .ZN(n6618) );
  NOR4_X1 U8162 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n6622)
         );
  OAI21_X1 U8163 ( .B1(n10308), .B2(n10334), .A(n6622), .ZN(P2_U3295) );
  INV_X1 U8164 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7718) );
  INV_X1 U8165 ( .A(n7807), .ZN(n6626) );
  INV_X1 U8166 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9213) );
  INV_X1 U8167 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n7846) );
  INV_X1 U8168 ( .A(n7885), .ZN(n6628) );
  NAND2_X1 U8169 ( .A1(n6628), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7901) );
  INV_X1 U8170 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9201) );
  INV_X1 U8171 ( .A(n7919), .ZN(n6629) );
  NAND2_X1 U8172 ( .A1(n6629), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7921) );
  INV_X1 U8173 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8938) );
  INV_X1 U8174 ( .A(n7951), .ZN(n6631) );
  AND2_X1 U8175 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6630) );
  NAND2_X1 U8176 ( .A1(n6631), .A2(n6630), .ZN(n7998) );
  OR2_X1 U8177 ( .A1(n7998), .A2(n6527), .ZN(n6637) );
  INV_X1 U8178 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U8179 ( .A1(n7992), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U8180 ( .A1(n6431), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6632) );
  OAI211_X1 U8181 ( .C1(n4479), .C2(n6634), .A(n6633), .B(n6632), .ZN(n6635)
         );
  INV_X1 U8182 ( .A(n6635), .ZN(n6636) );
  NAND2_X1 U8183 ( .A1(n9563), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6638) );
  OAI21_X1 U8184 ( .B1(n9616), .B2(n9563), .A(n6638), .ZN(P1_U3584) );
  INV_X1 U8185 ( .A(n7235), .ZN(n7242) );
  OAI222_X1 U8186 ( .A1(n9137), .A2(n6640), .B1(n9139), .B2(n6639), .C1(
        P2_U3152), .C2(n7242), .ZN(P2_U3343) );
  AOI21_X1 U8187 ( .B1(n7476), .B2(n6642), .A(n6641), .ZN(n6644) );
  INV_X1 U8188 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7535) );
  AOI22_X1 U8189 ( .A1(n7554), .A2(n7535), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n7056), .ZN(n6643) );
  NOR2_X1 U8190 ( .A1(n6644), .A2(n6643), .ZN(n7055) );
  AOI21_X1 U8191 ( .B1(n6644), .B2(n6643), .A(n7055), .ZN(n6651) );
  INV_X1 U8192 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7531) );
  NOR2_X1 U8193 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7531), .ZN(n7647) );
  NOR2_X1 U8194 ( .A1(n9595), .A2(n7056), .ZN(n6645) );
  AOI211_X1 U8195 ( .C1(n10122), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7647), .B(
        n6645), .ZN(n6650) );
  NAND2_X1 U8196 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7523), .ZN(n6647) );
  NAND2_X1 U8197 ( .A1(n6647), .A2(n6646), .ZN(n7063) );
  XNOR2_X1 U8198 ( .A(n7063), .B(n7056), .ZN(n6648) );
  NAND2_X1 U8199 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n6648), .ZN(n7064) );
  OAI211_X1 U8200 ( .C1(n6648), .C2(P1_REG2_REG_14__SCAN_IN), .A(n10124), .B(
        n7064), .ZN(n6649) );
  OAI211_X1 U8201 ( .C1(n6651), .C2(n10106), .A(n6650), .B(n6649), .ZN(
        P1_U3255) );
  NAND2_X1 U8202 ( .A1(n6653), .A2(n6652), .ZN(n7025) );
  INV_X1 U8203 ( .A(n10150), .ZN(n9789) );
  AOI22_X1 U8204 ( .A1(n10157), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9789), .ZN(n6657) );
  NOR2_X1 U8205 ( .A1(n6654), .A2(n9534), .ZN(n6655) );
  NAND2_X1 U8206 ( .A1(n9810), .A2(n6655), .ZN(n9832) );
  INV_X2 U8207 ( .A(n10157), .ZN(n9810) );
  OAI21_X1 U8208 ( .B1(n9733), .B2(n9830), .A(n6666), .ZN(n6656) );
  OAI211_X1 U8209 ( .C1(n6658), .C2(n10157), .A(n6657), .B(n6656), .ZN(
        P1_U3291) );
  INV_X1 U8210 ( .A(n6660), .ZN(n10328) );
  OAI22_X1 U8211 ( .A1(n10328), .A2(n10281), .B1(n6659), .B2(n10284), .ZN(
        n10330) );
  AOI21_X1 U8212 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n10245), .A(n10330), .ZN(
        n6664) );
  AOI22_X1 U8213 ( .A1(n10306), .A2(n6660), .B1(n10308), .B2(
        P2_REG2_REG_0__SCAN_IN), .ZN(n6663) );
  OAI21_X1 U8214 ( .B1(n8637), .B2(n10302), .A(n6661), .ZN(n6662) );
  OAI211_X1 U8215 ( .C1(n6664), .C2(n10308), .A(n6663), .B(n6662), .ZN(
        P2_U3296) );
  NAND2_X1 U8216 ( .A1(n7947), .A2(n6665), .ZN(n6885) );
  XNOR2_X2 U8217 ( .A(n9564), .B(n10171), .ZN(n10132) );
  AND2_X1 U8218 ( .A1(n10138), .A2(n6666), .ZN(n10131) );
  NAND2_X1 U8219 ( .A1(n10132), .A2(n10131), .ZN(n10130) );
  NAND2_X1 U8220 ( .A1(n9564), .A2(n6667), .ZN(n6668) );
  AND2_X1 U8221 ( .A1(n10130), .A2(n6668), .ZN(n6719) );
  XNOR2_X1 U8222 ( .A(n10139), .B(n10176), .ZN(n9301) );
  OR2_X1 U8223 ( .A1(n10139), .A2(n9484), .ZN(n6669) );
  NAND2_X1 U8224 ( .A1(n6718), .A2(n6669), .ZN(n6670) );
  OR2_X1 U8225 ( .A1(n9561), .A2(n6681), .ZN(n9488) );
  NAND2_X1 U8226 ( .A1(n9561), .A2(n6681), .ZN(n9490) );
  NAND2_X1 U8227 ( .A1(n6670), .A2(n9299), .ZN(n6702) );
  OAI21_X1 U8228 ( .B1(n6670), .B2(n9299), .A(n6702), .ZN(n6730) );
  OAI22_X1 U8229 ( .A1(n9485), .A2(n9818), .B1(n6898), .B2(n9816), .ZN(n6680)
         );
  INV_X1 U8230 ( .A(n10132), .ZN(n10134) );
  NAND2_X1 U8231 ( .A1(n10134), .A2(n10133), .ZN(n6673) );
  OR2_X1 U8232 ( .A1(n9564), .A2(n10171), .ZN(n6672) );
  NAND2_X1 U8233 ( .A1(n6673), .A2(n6672), .ZN(n9487) );
  INV_X1 U8234 ( .A(n9301), .ZN(n6674) );
  NAND2_X1 U8235 ( .A1(n9487), .A2(n6674), .ZN(n6675) );
  OR2_X1 U8236 ( .A1(n10139), .A2(n10176), .ZN(n9482) );
  XNOR2_X1 U8237 ( .A(n6705), .B(n9299), .ZN(n6678) );
  NAND2_X1 U8238 ( .A1(n9473), .A2(n10148), .ZN(n6677) );
  NAND2_X1 U8239 ( .A1(n9480), .A2(n9527), .ZN(n6676) );
  NOR2_X1 U8240 ( .A1(n6678), .A2(n9807), .ZN(n6679) );
  AOI211_X1 U8241 ( .C1(n7615), .C2(n6730), .A(n6680), .B(n6679), .ZN(n6734)
         );
  NAND2_X1 U8242 ( .A1(n10171), .A2(n10147), .ZN(n10145) );
  OR2_X1 U8243 ( .A1(n10145), .A2(n9484), .ZN(n6723) );
  AOI21_X1 U8244 ( .B1(n6731), .B2(n6723), .A(n6711), .ZN(n6732) );
  OAI22_X1 U8245 ( .A1(n9810), .A2(n6465), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10150), .ZN(n6683) );
  NOR2_X1 U8246 ( .A1(n9799), .A2(n6681), .ZN(n6682) );
  AOI211_X1 U8247 ( .C1(n6732), .C2(n9733), .A(n6683), .B(n6682), .ZN(n6686)
         );
  NAND2_X1 U8248 ( .A1(n6684), .A2(n10148), .ZN(n10144) );
  NAND2_X1 U8249 ( .A1(n6730), .A2(n9834), .ZN(n6685) );
  OAI211_X1 U8250 ( .C1(n6734), .C2(n10157), .A(n6686), .B(n6685), .ZN(
        P1_U3288) );
  AOI21_X1 U8251 ( .B1(n6688), .B2(n10038), .A(n6687), .ZN(n6690) );
  INV_X1 U8252 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10032) );
  AOI22_X1 U8253 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6960), .B1(n6957), .B2(
        n10032), .ZN(n6689) );
  NOR2_X1 U8254 ( .A1(n6690), .A2(n6689), .ZN(n6959) );
  AOI21_X1 U8255 ( .B1(n6690), .B2(n6689), .A(n6959), .ZN(n6700) );
  AOI22_X1 U8256 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6957), .B1(n6960), .B2(
        n7443), .ZN(n6694) );
  OAI21_X1 U8257 ( .B1(n6694), .B2(n6693), .A(n6956), .ZN(n6695) );
  NAND2_X1 U8258 ( .A1(n6695), .A2(n10226), .ZN(n6699) );
  INV_X1 U8259 ( .A(n10227), .ZN(n9992) );
  INV_X1 U8260 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U8261 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7507) );
  OAI21_X1 U8262 ( .B1(n8091), .B2(n6696), .A(n7507), .ZN(n6697) );
  AOI21_X1 U8263 ( .B1(n9992), .B2(n6957), .A(n6697), .ZN(n6698) );
  OAI211_X1 U8264 ( .C1(n6700), .C2(n10229), .A(n6699), .B(n6698), .ZN(
        P2_U3259) );
  OR2_X1 U8265 ( .A1(n9561), .A2(n6731), .ZN(n6701) );
  NAND2_X1 U8266 ( .A1(n6702), .A2(n6701), .ZN(n6703) );
  OR2_X1 U8267 ( .A1(n9560), .A2(n10182), .ZN(n7014) );
  NAND2_X1 U8268 ( .A1(n9560), .A2(n10182), .ZN(n9491) );
  NAND2_X1 U8269 ( .A1(n7014), .A2(n9491), .ZN(n9298) );
  OAI21_X1 U8270 ( .B1(n6703), .B2(n9298), .A(n6884), .ZN(n10186) );
  INV_X1 U8271 ( .A(n10186), .ZN(n6717) );
  INV_X1 U8272 ( .A(n9834), .ZN(n7633) );
  INV_X1 U8273 ( .A(n9488), .ZN(n6704) );
  XNOR2_X1 U8274 ( .A(n6878), .B(n9298), .ZN(n6708) );
  NAND2_X1 U8275 ( .A1(n10186), .A2(n7615), .ZN(n6707) );
  AOI22_X1 U8276 ( .A1(n10137), .A2(n9561), .B1(n9559), .B2(n10140), .ZN(n6706) );
  OAI211_X1 U8277 ( .C1(n9807), .C2(n6708), .A(n6707), .B(n6706), .ZN(n10184)
         );
  NAND2_X1 U8278 ( .A1(n10184), .A2(n9810), .ZN(n6716) );
  OAI22_X1 U8279 ( .A1(n9810), .A2(n6710), .B1(n6709), .B2(n10150), .ZN(n6714)
         );
  NAND2_X1 U8280 ( .A1(n6711), .A2(n10182), .ZN(n6876) );
  OR2_X1 U8281 ( .A1(n6711), .A2(n10182), .ZN(n6712) );
  NAND2_X1 U8282 ( .A1(n6876), .A2(n6712), .ZN(n10183) );
  NOR2_X1 U8283 ( .A1(n10183), .A2(n9832), .ZN(n6713) );
  AOI211_X1 U8284 ( .C1(n9830), .C2(n6882), .A(n6714), .B(n6713), .ZN(n6715)
         );
  OAI211_X1 U8285 ( .C1(n6717), .C2(n7633), .A(n6716), .B(n6715), .ZN(P1_U3287) );
  XNOR2_X1 U8286 ( .A(n9487), .B(n9301), .ZN(n6722) );
  OAI21_X1 U8287 ( .B1(n6719), .B2(n9301), .A(n6718), .ZN(n10180) );
  NAND2_X1 U8288 ( .A1(n10180), .A2(n7615), .ZN(n6721) );
  AOI22_X1 U8289 ( .A1(n10137), .A2(n9564), .B1(n9561), .B2(n10140), .ZN(n6720) );
  OAI211_X1 U8290 ( .C1(n9807), .C2(n6722), .A(n6721), .B(n6720), .ZN(n10178)
         );
  INV_X1 U8291 ( .A(n10178), .ZN(n6729) );
  INV_X1 U8292 ( .A(n10145), .ZN(n6724) );
  OAI21_X1 U8293 ( .B1(n6724), .B2(n10176), .A(n6723), .ZN(n10177) );
  OAI22_X1 U8294 ( .A1(n9799), .A2(n10176), .B1(n10177), .B2(n9832), .ZN(n6727) );
  OAI22_X1 U8295 ( .A1(n10150), .A2(n6432), .B1(n6725), .B2(n9810), .ZN(n6726)
         );
  AOI211_X1 U8296 ( .C1(n9834), .C2(n10180), .A(n6727), .B(n6726), .ZN(n6728)
         );
  OAI21_X1 U8297 ( .B1(n10157), .B2(n6729), .A(n6728), .ZN(P1_U3289) );
  INV_X1 U8298 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6737) );
  INV_X1 U8299 ( .A(n6730), .ZN(n6735) );
  AOI22_X1 U8300 ( .A1(n6732), .A2(n10146), .B1(n10000), .B2(n6731), .ZN(n6733) );
  OAI211_X1 U8301 ( .C1(n6735), .C2(n9999), .A(n6734), .B(n6733), .ZN(n6738)
         );
  NAND2_X1 U8302 ( .A1(n6738), .A2(n10212), .ZN(n6736) );
  OAI21_X1 U8303 ( .B1(n10212), .B2(n6737), .A(n6736), .ZN(P1_U3463) );
  NAND2_X1 U8304 ( .A1(n6738), .A2(n10223), .ZN(n6739) );
  OAI21_X1 U8305 ( .B1(n10223), .B2(n6464), .A(n6739), .ZN(P1_U3526) );
  NAND2_X1 U8306 ( .A1(n6743), .A2(n6742), .ZN(n8284) );
  XNOR2_X1 U8307 ( .A(n8289), .B(n8212), .ZN(n8343) );
  NAND2_X1 U8308 ( .A1(n10260), .A2(n8156), .ZN(n6744) );
  NAND2_X1 U8309 ( .A1(n8343), .A2(n6744), .ZN(n6747) );
  INV_X1 U8310 ( .A(n8343), .ZN(n6746) );
  INV_X1 U8311 ( .A(n6744), .ZN(n6745) );
  NAND2_X1 U8312 ( .A1(n6746), .A2(n6745), .ZN(n6750) );
  NAND2_X1 U8313 ( .A1(n6747), .A2(n6750), .ZN(n8283) );
  INV_X1 U8314 ( .A(n8283), .ZN(n6748) );
  XNOR2_X1 U8315 ( .A(n8212), .B(n10271), .ZN(n6754) );
  AND2_X1 U8316 ( .A1(n8378), .A2(n8156), .ZN(n6752) );
  XNOR2_X1 U8317 ( .A(n6754), .B(n6752), .ZN(n8344) );
  AND2_X1 U8318 ( .A1(n8344), .A2(n6750), .ZN(n6751) );
  NAND2_X1 U8319 ( .A1(n8335), .A2(n6751), .ZN(n8334) );
  INV_X1 U8320 ( .A(n6752), .ZN(n6753) );
  NAND2_X1 U8321 ( .A1(n6754), .A2(n6753), .ZN(n6755) );
  AND2_X2 U8322 ( .A1(n8334), .A2(n6755), .ZN(n6761) );
  XNOR2_X1 U8323 ( .A(n10367), .B(n8212), .ZN(n6756) );
  AND2_X1 U8324 ( .A1(n10262), .A2(n8156), .ZN(n6757) );
  NAND2_X1 U8325 ( .A1(n6756), .A2(n6757), .ZN(n7143) );
  INV_X1 U8326 ( .A(n6756), .ZN(n8229) );
  INV_X1 U8327 ( .A(n6757), .ZN(n6758) );
  NAND2_X1 U8328 ( .A1(n8229), .A2(n6758), .ZN(n6759) );
  AND2_X1 U8329 ( .A1(n7143), .A2(n6759), .ZN(n6760) );
  OAI211_X1 U8330 ( .C1(n6761), .C2(n6760), .A(n8228), .B(n8336), .ZN(n6768)
         );
  NAND2_X1 U8331 ( .A1(n8377), .A2(n10261), .ZN(n6763) );
  NAND2_X1 U8332 ( .A1(n8378), .A2(n10259), .ZN(n6762) );
  NAND2_X1 U8333 ( .A1(n6763), .A2(n6762), .ZN(n9016) );
  INV_X1 U8334 ( .A(n9016), .ZN(n6765) );
  OAI22_X1 U8335 ( .A1(n8263), .A2(n6765), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6764), .ZN(n6766) );
  AOI21_X1 U8336 ( .B1(n9008), .B2(n8342), .A(n6766), .ZN(n6767) );
  OAI211_X1 U8337 ( .C1(n10367), .C2(n8338), .A(n6768), .B(n6767), .ZN(
        P2_U3215) );
  INV_X1 U8338 ( .A(n7697), .ZN(n6773) );
  NOR2_X1 U8339 ( .A1(n6770), .A2(n6769), .ZN(n6872) );
  OR2_X1 U8340 ( .A1(n6872), .A2(n6035), .ZN(n6771) );
  XNOR2_X1 U8341 ( .A(n6771), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7698) );
  INV_X1 U8342 ( .A(n7698), .ZN(n7203) );
  OAI222_X1 U8343 ( .A1(n9968), .A2(n6772), .B1(n9971), .B2(n6773), .C1(n7203), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8344 ( .A(n8071), .ZN(n7250) );
  OAI222_X1 U8345 ( .A1(n9137), .A2(n6774), .B1(n9139), .B2(n6773), .C1(n7250), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8346 ( .A(n6775), .ZN(n6777) );
  OR2_X1 U8347 ( .A1(n6777), .A2(n6776), .ZN(n6891) );
  OR2_X1 U8348 ( .A1(n6778), .A2(n6792), .ZN(n6780) );
  AOI22_X1 U8349 ( .A1(n7803), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7802), .B2(
        n10098), .ZN(n6779) );
  NAND2_X1 U8350 ( .A1(n7887), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6787) );
  INV_X1 U8351 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6781) );
  OR2_X1 U8352 ( .A1(n6557), .A2(n6781), .ZN(n6786) );
  INV_X1 U8353 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7038) );
  NAND2_X1 U8354 ( .A1(n6782), .A2(n7038), .ZN(n6783) );
  NAND2_X1 U8355 ( .A1(n6821), .A2(n6783), .ZN(n7191) );
  OR2_X1 U8356 ( .A1(n6527), .A2(n7191), .ZN(n6785) );
  OR2_X1 U8357 ( .A1(n4476), .A2(n8880), .ZN(n6784) );
  NAND4_X1 U8358 ( .A1(n6787), .A2(n6786), .A3(n6785), .A4(n6784), .ZN(n9558)
         );
  NAND2_X1 U8359 ( .A1(n9558), .A2(n7347), .ZN(n6788) );
  OAI21_X1 U8360 ( .B1(n7192), .B2(n7946), .A(n6788), .ZN(n6789) );
  XNOR2_X1 U8361 ( .A(n6789), .B(n7947), .ZN(n6809) );
  OR2_X1 U8362 ( .A1(n7192), .A2(n7945), .ZN(n6791) );
  NAND2_X1 U8363 ( .A1(n9558), .A2(n7928), .ZN(n6790) );
  NAND2_X1 U8364 ( .A1(n6791), .A2(n6790), .ZN(n6810) );
  NAND2_X1 U8365 ( .A1(n6809), .A2(n6810), .ZN(n7032) );
  NAND2_X1 U8366 ( .A1(n9559), .A2(n7347), .ZN(n6797) );
  AOI22_X1 U8367 ( .A1(n7803), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7802), .B2(
        n10080), .ZN(n6795) );
  INV_X2 U8368 ( .A(n6792), .ZN(n6907) );
  NAND2_X1 U8369 ( .A1(n6793), .A2(n6907), .ZN(n6794) );
  OR2_X1 U8370 ( .A1(n10190), .A2(n7946), .ZN(n6796) );
  NAND2_X1 U8371 ( .A1(n6797), .A2(n6796), .ZN(n6798) );
  XNOR2_X1 U8372 ( .A(n6798), .B(n8047), .ZN(n6893) );
  INV_X1 U8373 ( .A(n6893), .ZN(n6801) );
  NAND2_X1 U8374 ( .A1(n9559), .A2(n7928), .ZN(n6800) );
  OR2_X1 U8375 ( .A1(n10190), .A2(n7945), .ZN(n6799) );
  AND2_X1 U8376 ( .A1(n6800), .A2(n6799), .ZN(n6805) );
  INV_X1 U8377 ( .A(n6805), .ZN(n6896) );
  NAND2_X1 U8378 ( .A1(n6801), .A2(n6896), .ZN(n6802) );
  AND2_X1 U8379 ( .A1(n7032), .A2(n6802), .ZN(n6804) );
  AND2_X1 U8380 ( .A1(n6891), .A2(n6804), .ZN(n6803) );
  INV_X1 U8381 ( .A(n6804), .ZN(n6807) );
  NAND2_X1 U8382 ( .A1(n6893), .A2(n6805), .ZN(n6806) );
  OR2_X1 U8383 ( .A1(n6807), .A2(n6806), .ZN(n6808) );
  INV_X1 U8384 ( .A(n6809), .ZN(n6812) );
  INV_X1 U8385 ( .A(n6810), .ZN(n6811) );
  NAND2_X1 U8386 ( .A1(n6812), .A2(n6811), .ZN(n7031) );
  NAND2_X1 U8387 ( .A1(n6814), .A2(n6907), .ZN(n6817) );
  AOI22_X1 U8388 ( .A1(n7803), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7802), .B2(
        n6815), .ZN(n6816) );
  NAND2_X1 U8389 ( .A1(n6817), .A2(n6816), .ZN(n7092) );
  NAND2_X1 U8390 ( .A1(n7092), .A2(n7347), .ZN(n6829) );
  INV_X1 U8391 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6818) );
  OR2_X1 U8392 ( .A1(n6557), .A2(n6818), .ZN(n6827) );
  INV_X1 U8393 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6819) );
  OR2_X1 U8394 ( .A1(n4479), .A2(n6819), .ZN(n6826) );
  INV_X1 U8395 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6820) );
  NAND2_X1 U8396 ( .A1(n6821), .A2(n6820), .ZN(n6822) );
  NAND2_X1 U8397 ( .A1(n6823), .A2(n6822), .ZN(n7021) );
  OR2_X1 U8398 ( .A1(n6527), .A2(n7021), .ZN(n6825) );
  INV_X1 U8399 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7026) );
  OR2_X1 U8400 ( .A1(n4477), .A2(n7026), .ZN(n6824) );
  OR2_X1 U8401 ( .A1(n7011), .A2(n7943), .ZN(n6828) );
  AND2_X1 U8402 ( .A1(n6829), .A2(n6828), .ZN(n6905) );
  NAND2_X1 U8403 ( .A1(n7092), .A2(n8044), .ZN(n6831) );
  OR2_X1 U8404 ( .A1(n7011), .A2(n7945), .ZN(n6830) );
  NAND2_X1 U8405 ( .A1(n6831), .A2(n6830), .ZN(n6832) );
  XOR2_X1 U8406 ( .A(n6905), .B(n6904), .Z(n6833) );
  XNOR2_X1 U8407 ( .A(n6906), .B(n6833), .ZN(n6839) );
  NOR2_X1 U8408 ( .A1(n7291), .A2(n9234), .ZN(n6834) );
  AOI211_X1 U8409 ( .C1(n9236), .C2(n9558), .A(n6835), .B(n6834), .ZN(n6836)
         );
  OAI21_X1 U8410 ( .B1(n9249), .B2(n7021), .A(n6836), .ZN(n6837) );
  AOI21_X1 U8411 ( .B1(n7092), .B2(n9251), .A(n6837), .ZN(n6838) );
  OAI21_X1 U8412 ( .B1(n6839), .B2(n9253), .A(n6838), .ZN(P1_U3211) );
  INV_X1 U8413 ( .A(n7769), .ZN(n6874) );
  AOI22_X1 U8414 ( .A1(n8421), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9129), .ZN(n6840) );
  OAI21_X1 U8415 ( .B1(n6874), .B2(n9134), .A(n6840), .ZN(P2_U3341) );
  NAND2_X1 U8416 ( .A1(n10276), .A2(n10282), .ZN(n6842) );
  INV_X1 U8417 ( .A(n6841), .ZN(n6934) );
  XNOR2_X1 U8418 ( .A(n6842), .B(n6934), .ZN(n6845) );
  NAND2_X1 U8419 ( .A1(n8378), .A2(n10261), .ZN(n6844) );
  NAND2_X1 U8420 ( .A1(n8380), .A2(n10259), .ZN(n6843) );
  NAND2_X1 U8421 ( .A1(n6844), .A2(n6843), .ZN(n8286) );
  AOI21_X1 U8422 ( .B1(n6845), .B2(n10264), .A(n8286), .ZN(n10360) );
  NAND2_X1 U8423 ( .A1(n6847), .A2(n6846), .ZN(n6849) );
  NAND2_X1 U8424 ( .A1(n10287), .A2(n10344), .ZN(n6848) );
  NAND2_X1 U8425 ( .A1(n6849), .A2(n6848), .ZN(n10290) );
  NAND2_X1 U8426 ( .A1(n10290), .A2(n10291), .ZN(n6852) );
  NAND2_X1 U8427 ( .A1(n6850), .A2(n10351), .ZN(n6851) );
  XNOR2_X1 U8428 ( .A(n6935), .B(n6934), .ZN(n10357) );
  NAND2_X1 U8429 ( .A1(n10294), .A2(n8289), .ZN(n6853) );
  NAND2_X1 U8430 ( .A1(n6853), .A2(n10295), .ZN(n6854) );
  OR2_X1 U8431 ( .A1(n6854), .A2(n10267), .ZN(n10354) );
  AOI22_X1 U8432 ( .A1(n10308), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n8288), .B2(
        n10245), .ZN(n6856) );
  NAND2_X1 U8433 ( .A1(n10302), .A2(n8289), .ZN(n6855) );
  OAI211_X1 U8434 ( .C1(n10304), .C2(n10354), .A(n6856), .B(n6855), .ZN(n6857)
         );
  AOI21_X1 U8435 ( .B1(n10357), .B2(n10306), .A(n6857), .ZN(n6858) );
  OAI21_X1 U8436 ( .B1(n10360), .B2(n10308), .A(n6858), .ZN(P2_U3291) );
  XNOR2_X1 U8437 ( .A(n6859), .B(n6582), .ZN(n10342) );
  INV_X1 U8438 ( .A(n10342), .ZN(n6870) );
  NAND2_X1 U8439 ( .A1(n5674), .A2(n6582), .ZN(n6860) );
  NAND2_X1 U8440 ( .A1(n6587), .A2(n6860), .ZN(n6861) );
  NAND2_X1 U8441 ( .A1(n6861), .A2(n10264), .ZN(n6863) );
  AOI22_X1 U8442 ( .A1(n10259), .A2(n6578), .B1(n8381), .B2(n10261), .ZN(n6862) );
  NAND2_X1 U8443 ( .A1(n6863), .A2(n6862), .ZN(n10340) );
  OAI21_X1 U8444 ( .B1(n6864), .B2(n10338), .A(n10293), .ZN(n10339) );
  AOI22_X1 U8445 ( .A1(n10308), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n10245), .ZN(n6867) );
  NAND2_X1 U8446 ( .A1(n10302), .A2(n6865), .ZN(n6866) );
  OAI211_X1 U8447 ( .C1(n10273), .C2(n10339), .A(n6867), .B(n6866), .ZN(n6868)
         );
  AOI21_X1 U8448 ( .B1(n10299), .B2(n10340), .A(n6868), .ZN(n6869) );
  OAI21_X1 U8449 ( .B1(n6870), .B2(n8639), .A(n6869), .ZN(P2_U3294) );
  INV_X1 U8450 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6871) );
  NAND2_X1 U8451 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  NAND2_X1 U8452 ( .A1(n6873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6988) );
  XNOR2_X1 U8453 ( .A(n6988), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7770) );
  INV_X1 U8454 ( .A(n7770), .ZN(n7380) );
  OAI222_X1 U8455 ( .A1(n9968), .A2(n6875), .B1(n9971), .B2(n6874), .C1(n7380), 
        .C2(P1_U3084), .ZN(P1_U3336) );
  INV_X1 U8456 ( .A(n6876), .ZN(n6877) );
  INV_X1 U8457 ( .A(n10190), .ZN(n6970) );
  OAI211_X1 U8458 ( .C1(n6877), .C2(n10190), .A(n10146), .B(n6979), .ZN(n10189) );
  INV_X1 U8459 ( .A(n10189), .ZN(n6881) );
  NAND2_X1 U8460 ( .A1(n9558), .A2(n10140), .ZN(n10188) );
  OAI21_X1 U8461 ( .B1(n10150), .B2(n6899), .A(n10188), .ZN(n6880) );
  AND2_X1 U8462 ( .A1(n7018), .A2(n7014), .ZN(n6975) );
  OR2_X1 U8463 ( .A1(n9559), .A2(n10190), .ZN(n7015) );
  NAND2_X1 U8464 ( .A1(n9559), .A2(n10190), .ZN(n7016) );
  XNOR2_X1 U8465 ( .A(n6975), .B(n9303), .ZN(n6879) );
  OAI22_X1 U8466 ( .A1(n6879), .A2(n9807), .B1(n6898), .B2(n9818), .ZN(n10191)
         );
  AOI211_X1 U8467 ( .C1(n6881), .C2(n9690), .A(n6880), .B(n10191), .ZN(n6890)
         );
  OR2_X1 U8468 ( .A1(n9560), .A2(n6882), .ZN(n6883) );
  XOR2_X1 U8469 ( .A(n9303), .B(n6968), .Z(n10193) );
  INV_X1 U8470 ( .A(n6885), .ZN(n6886) );
  INV_X1 U8471 ( .A(n9813), .ZN(n9746) );
  INV_X1 U8472 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6887) );
  OAI22_X1 U8473 ( .A1(n9799), .A2(n10190), .B1(n6887), .B2(n9810), .ZN(n6888)
         );
  AOI21_X1 U8474 ( .B1(n10193), .B2(n9746), .A(n6888), .ZN(n6889) );
  OAI21_X1 U8475 ( .B1(n6890), .B2(n10157), .A(n6889), .ZN(P1_U3286) );
  AND2_X1 U8476 ( .A1(n6892), .A2(n6891), .ZN(n6894) );
  NAND2_X1 U8477 ( .A1(n6894), .A2(n6893), .ZN(n7033) );
  OAI21_X1 U8478 ( .B1(n6894), .B2(n6893), .A(n7033), .ZN(n6895) );
  NOR2_X1 U8479 ( .A1(n6895), .A2(n6896), .ZN(n7035) );
  AOI21_X1 U8480 ( .B1(n6896), .B2(n6895), .A(n7035), .ZN(n6903) );
  AND2_X1 U8481 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10079) );
  AOI21_X1 U8482 ( .B1(n9247), .B2(n9558), .A(n10079), .ZN(n6897) );
  OAI21_X1 U8483 ( .B1(n6898), .B2(n9245), .A(n6897), .ZN(n6901) );
  NOR2_X1 U8484 ( .A1(n9249), .A2(n6899), .ZN(n6900) );
  AOI211_X1 U8485 ( .C1(n6970), .C2(n9251), .A(n6901), .B(n6900), .ZN(n6902)
         );
  OAI21_X1 U8486 ( .B1(n6903), .B2(n9253), .A(n6902), .ZN(P1_U3225) );
  NAND2_X1 U8487 ( .A1(n5930), .A2(n6907), .ZN(n6910) );
  AOI22_X1 U8488 ( .A1(n7803), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7802), .B2(
        n6908), .ZN(n6909) );
  NAND2_X1 U8489 ( .A1(n6910), .A2(n6909), .ZN(n7287) );
  NAND2_X1 U8490 ( .A1(n7287), .A2(n7347), .ZN(n6912) );
  OR2_X1 U8491 ( .A1(n7291), .A2(n7943), .ZN(n6911) );
  NAND2_X1 U8492 ( .A1(n6912), .A2(n6911), .ZN(n7129) );
  NAND2_X1 U8493 ( .A1(n7287), .A2(n8044), .ZN(n6914) );
  OR2_X1 U8494 ( .A1(n7291), .A2(n7945), .ZN(n6913) );
  NAND2_X1 U8495 ( .A1(n6914), .A2(n6913), .ZN(n6915) );
  XNOR2_X1 U8496 ( .A(n6915), .B(n7947), .ZN(n7128) );
  XOR2_X1 U8497 ( .A(n7129), .B(n7128), .Z(n6916) );
  XNOR2_X1 U8498 ( .A(n7130), .B(n6916), .ZN(n6932) );
  OR2_X1 U8499 ( .A1(n4477), .A2(n6917), .ZN(n6918) );
  OAI21_X1 U8500 ( .B1(n4478), .B2(n10221), .A(n6918), .ZN(n6926) );
  NAND2_X1 U8501 ( .A1(n6920), .A2(n6919), .ZN(n6921) );
  NAND2_X1 U8502 ( .A1(n6922), .A2(n6921), .ZN(n7295) );
  NOR2_X1 U8503 ( .A1(n6527), .A2(n7295), .ZN(n6925) );
  INV_X1 U8504 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6923) );
  NOR2_X1 U8505 ( .A1(n6557), .A2(n6923), .ZN(n6924) );
  NOR2_X1 U8506 ( .A1(n7011), .A2(n9245), .ZN(n6927) );
  AOI211_X1 U8507 ( .C1(n9247), .C2(n9556), .A(n6928), .B(n6927), .ZN(n6929)
         );
  OAI21_X1 U8508 ( .B1(n9249), .B2(n7107), .A(n6929), .ZN(n6930) );
  AOI21_X1 U8509 ( .B1(n7287), .B2(n9251), .A(n6930), .ZN(n6931) );
  OAI21_X1 U8510 ( .B1(n6932), .B2(n9253), .A(n6931), .ZN(P1_U3219) );
  XNOR2_X1 U8511 ( .A(n6933), .B(n6944), .ZN(n6949) );
  NAND2_X1 U8512 ( .A1(n6935), .A2(n6934), .ZN(n6937) );
  NAND2_X1 U8513 ( .A1(n10285), .A2(n10355), .ZN(n6936) );
  NAND2_X1 U8514 ( .A1(n6938), .A2(n10361), .ZN(n6939) );
  NAND2_X1 U8515 ( .A1(n10367), .A2(n8339), .ZN(n6940) );
  INV_X1 U8516 ( .A(n10237), .ZN(n6942) );
  NAND2_X1 U8517 ( .A1(n10375), .A2(n8377), .ZN(n6943) );
  OAI21_X1 U8518 ( .B1(n6945), .B2(n6944), .A(n6995), .ZN(n10386) );
  NAND2_X1 U8519 ( .A1(n8375), .A2(n10261), .ZN(n6947) );
  NAND2_X1 U8520 ( .A1(n8377), .A2(n10259), .ZN(n6946) );
  NAND2_X1 U8521 ( .A1(n6947), .A2(n6946), .ZN(n7161) );
  AOI21_X1 U8522 ( .B1(n10386), .B2(n8646), .A(n7161), .ZN(n6948) );
  OAI21_X1 U8523 ( .B1(n10281), .B2(n6949), .A(n6948), .ZN(n10384) );
  INV_X1 U8524 ( .A(n10384), .ZN(n6955) );
  INV_X1 U8525 ( .A(n7167), .ZN(n10383) );
  AND2_X1 U8526 ( .A1(n10249), .A2(n10383), .ZN(n7003) );
  INV_X1 U8527 ( .A(n7003), .ZN(n6950) );
  OAI211_X1 U8528 ( .C1(n10383), .C2(n10249), .A(n6950), .B(n10295), .ZN(
        n10382) );
  AOI22_X1 U8529 ( .A1(n10308), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7160), .B2(
        n10245), .ZN(n6952) );
  NAND2_X1 U8530 ( .A1(n10302), .A2(n7167), .ZN(n6951) );
  OAI211_X1 U8531 ( .C1(n10382), .C2(n10304), .A(n6952), .B(n6951), .ZN(n6953)
         );
  AOI21_X1 U8532 ( .B1(n10386), .B2(n10251), .A(n6953), .ZN(n6954) );
  OAI21_X1 U8533 ( .B1(n6955), .B2(n10308), .A(n6954), .ZN(P2_U3287) );
  OAI21_X1 U8534 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6957), .A(n6956), .ZN(
        n7241) );
  XNOR2_X1 U8535 ( .A(n7241), .B(n7235), .ZN(n6958) );
  NAND2_X1 U8536 ( .A1(n6958), .A2(n5457), .ZN(n7243) );
  OAI21_X1 U8537 ( .B1(n6958), .B2(n5457), .A(n7243), .ZN(n6966) );
  AOI21_X1 U8538 ( .B1(n10032), .B2(n6960), .A(n6959), .ZN(n7234) );
  XNOR2_X1 U8539 ( .A(n7234), .B(n7242), .ZN(n6961) );
  NAND2_X1 U8540 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n6961), .ZN(n7236) );
  OAI211_X1 U8541 ( .C1(n6961), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10224), .B(
        n7236), .ZN(n6964) );
  NOR2_X1 U8542 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5452), .ZN(n6962) );
  AOI21_X1 U8543 ( .B1(n10231), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n6962), .ZN(
        n6963) );
  OAI211_X1 U8544 ( .C1(n10227), .C2(n7242), .A(n6964), .B(n6963), .ZN(n6965)
         );
  AOI21_X1 U8545 ( .B1(n10226), .B2(n6966), .A(n6965), .ZN(n6967) );
  INV_X1 U8546 ( .A(n6967), .ZN(P2_U3260) );
  INV_X1 U8547 ( .A(n9303), .ZN(n6969) );
  NAND2_X1 U8548 ( .A1(n9559), .A2(n6970), .ZN(n6971) );
  NAND2_X1 U8549 ( .A1(n6972), .A2(n6971), .ZN(n6973) );
  OR2_X1 U8550 ( .A1(n7192), .A2(n9558), .ZN(n9332) );
  NAND2_X1 U8551 ( .A1(n7192), .A2(n9558), .ZN(n9334) );
  NAND2_X1 U8552 ( .A1(n6973), .A2(n9304), .ZN(n6974) );
  NAND2_X1 U8553 ( .A1(n7010), .A2(n6974), .ZN(n7200) );
  INV_X1 U8554 ( .A(n7200), .ZN(n6983) );
  NAND2_X1 U8555 ( .A1(n6975), .A2(n7015), .ZN(n6976) );
  NAND2_X1 U8556 ( .A1(n6976), .A2(n7016), .ZN(n9333) );
  NAND2_X1 U8557 ( .A1(n9333), .A2(n9304), .ZN(n9341) );
  OAI211_X1 U8558 ( .C1(n9333), .C2(n9304), .A(n9341), .B(n10135), .ZN(n6978)
         );
  AOI22_X1 U8559 ( .A1(n9557), .A2(n10140), .B1(n10137), .B2(n9559), .ZN(n6977) );
  AND2_X1 U8560 ( .A1(n6978), .A2(n6977), .ZN(n7196) );
  NAND2_X1 U8561 ( .A1(n6979), .A2(n7043), .ZN(n6980) );
  NAND2_X1 U8562 ( .A1(n6980), .A2(n10146), .ZN(n6981) );
  NOR2_X1 U8563 ( .A1(n7023), .A2(n6981), .ZN(n7193) );
  AOI21_X1 U8564 ( .B1(n10000), .B2(n7043), .A(n7193), .ZN(n6982) );
  OAI211_X1 U8565 ( .C1(n6983), .C2(n9930), .A(n7196), .B(n6982), .ZN(n6985)
         );
  NAND2_X1 U8566 ( .A1(n6985), .A2(n10212), .ZN(n6984) );
  OAI21_X1 U8567 ( .B1(n10212), .B2(n6781), .A(n6984), .ZN(P1_U3472) );
  NAND2_X1 U8568 ( .A1(n6985), .A2(n10223), .ZN(n6986) );
  OAI21_X1 U8569 ( .B1(n10223), .B2(n5999), .A(n6986), .ZN(P1_U3529) );
  INV_X1 U8570 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6991) );
  INV_X1 U8571 ( .A(n7781), .ZN(n6992) );
  INV_X1 U8572 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6987) );
  NAND2_X1 U8573 ( .A1(n6988), .A2(n6987), .ZN(n6989) );
  NAND2_X1 U8574 ( .A1(n6989), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6990) );
  XNOR2_X1 U8575 ( .A(n6990), .B(P1_IR_REG_18__SCAN_IN), .ZN(n7782) );
  INV_X1 U8576 ( .A(n7782), .ZN(n9587) );
  OAI222_X1 U8577 ( .A1(n9968), .A2(n6991), .B1(n9971), .B2(n6992), .C1(
        P1_U3084), .C2(n9587), .ZN(P1_U3335) );
  INV_X1 U8578 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6993) );
  INV_X1 U8579 ( .A(n8078), .ZN(n8444) );
  OAI222_X1 U8580 ( .A1(n9137), .A2(n6993), .B1(n9139), .B2(n6992), .C1(
        P2_U3152), .C2(n8444), .ZN(P2_U3340) );
  OR2_X1 U8581 ( .A1(n7167), .A2(n8376), .ZN(n6994) );
  XNOR2_X1 U8582 ( .A(n7075), .B(n4994), .ZN(n10391) );
  NAND2_X1 U8583 ( .A1(n10391), .A2(n8646), .ZN(n7002) );
  OAI21_X1 U8584 ( .B1(n7076), .B2(n6996), .A(n7083), .ZN(n7000) );
  NAND2_X1 U8585 ( .A1(n8374), .A2(n10261), .ZN(n6998) );
  NAND2_X1 U8586 ( .A1(n8376), .A2(n10259), .ZN(n6997) );
  NAND2_X1 U8587 ( .A1(n6998), .A2(n6997), .ZN(n6999) );
  AOI21_X1 U8588 ( .B1(n7000), .B2(n10264), .A(n6999), .ZN(n7001) );
  AND2_X1 U8589 ( .A1(n7002), .A2(n7001), .ZN(n10393) );
  INV_X1 U8590 ( .A(n8189), .ZN(n10387) );
  OR2_X1 U8591 ( .A1(n7003), .A2(n10387), .ZN(n7004) );
  NAND2_X1 U8592 ( .A1(n7228), .A2(n7004), .ZN(n10388) );
  AOI22_X1 U8593 ( .A1(n10308), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8188), .B2(
        n10245), .ZN(n7006) );
  NAND2_X1 U8594 ( .A1(n10302), .A2(n8189), .ZN(n7005) );
  OAI211_X1 U8595 ( .C1(n10388), .C2(n10273), .A(n7006), .B(n7005), .ZN(n7007)
         );
  AOI21_X1 U8596 ( .B1(n10391), .B2(n10251), .A(n7007), .ZN(n7008) );
  OAI21_X1 U8597 ( .B1(n10393), .B2(n10308), .A(n7008), .ZN(P2_U3286) );
  OR2_X1 U8598 ( .A1(n9558), .A2(n7043), .ZN(n7009) );
  OR2_X1 U8599 ( .A1(n7092), .A2(n7011), .ZN(n9338) );
  NAND2_X1 U8600 ( .A1(n7092), .A2(n7011), .ZN(n9336) );
  NAND2_X1 U8601 ( .A1(n9338), .A2(n9336), .ZN(n9306) );
  OAI21_X1 U8602 ( .B1(n7012), .B2(n9306), .A(n7094), .ZN(n7013) );
  INV_X1 U8603 ( .A(n7013), .ZN(n7051) );
  AND3_X1 U8604 ( .A1(n9332), .A2(n7015), .A3(n7014), .ZN(n9493) );
  INV_X1 U8605 ( .A(n7016), .ZN(n7017) );
  AND2_X1 U8606 ( .A1(n9332), .A2(n7017), .ZN(n9495) );
  AOI21_X1 U8607 ( .B1(n7018), .B2(n9493), .A(n9495), .ZN(n7098) );
  NAND2_X1 U8608 ( .A1(n7098), .A2(n9334), .ZN(n7019) );
  XNOR2_X1 U8609 ( .A(n7019), .B(n9306), .ZN(n7020) );
  INV_X1 U8610 ( .A(n7291), .ZN(n7286) );
  AOI222_X1 U8611 ( .A1(n10135), .A2(n7020), .B1(n7286), .B2(n10140), .C1(
        n9558), .C2(n10137), .ZN(n7050) );
  OAI21_X1 U8612 ( .B1(n7021), .B2(n10150), .A(n7050), .ZN(n7022) );
  NAND2_X1 U8613 ( .A1(n7022), .A2(n9810), .ZN(n7030) );
  INV_X1 U8614 ( .A(n7092), .ZN(n7027) );
  OAI21_X1 U8615 ( .B1(n7023), .B2(n7027), .A(n10146), .ZN(n7024) );
  NOR2_X1 U8616 ( .A1(n7024), .A2(n7109), .ZN(n7048) );
  NOR2_X1 U8617 ( .A1(n7025), .A2(n10148), .ZN(n7714) );
  OAI22_X1 U8618 ( .A1(n9799), .A2(n7027), .B1(n7026), .B2(n9810), .ZN(n7028)
         );
  AOI21_X1 U8619 ( .B1(n7048), .B2(n7714), .A(n7028), .ZN(n7029) );
  OAI211_X1 U8620 ( .C1(n7051), .C2(n9813), .A(n7030), .B(n7029), .ZN(P1_U3284) );
  NAND2_X1 U8621 ( .A1(n7032), .A2(n7031), .ZN(n7037) );
  INV_X1 U8622 ( .A(n7033), .ZN(n7034) );
  NOR2_X1 U8623 ( .A1(n7035), .A2(n7034), .ZN(n7036) );
  XOR2_X1 U8624 ( .A(n7037), .B(n7036), .Z(n7045) );
  NOR2_X1 U8625 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7038), .ZN(n10096) );
  AOI21_X1 U8626 ( .B1(n9557), .B2(n9247), .A(n10096), .ZN(n7039) );
  OAI21_X1 U8627 ( .B1(n7040), .B2(n9245), .A(n7039), .ZN(n7042) );
  NOR2_X1 U8628 ( .A1(n9249), .A2(n7191), .ZN(n7041) );
  AOI211_X1 U8629 ( .C1(n7043), .C2(n9251), .A(n7042), .B(n7041), .ZN(n7044)
         );
  OAI21_X1 U8630 ( .B1(n7045), .B2(n9253), .A(n7044), .ZN(P1_U3237) );
  INV_X1 U8631 ( .A(n7801), .ZN(n7046) );
  OAI222_X1 U8632 ( .A1(n9968), .A2(n8817), .B1(n9971), .B2(n7046), .C1(n9690), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8633 ( .A1(n9137), .A2(n7047), .B1(n9139), .B2(n7046), .C1(
        P2_U3152), .C2(n8086), .ZN(P2_U3339) );
  AOI21_X1 U8634 ( .B1(n10000), .B2(n7092), .A(n7048), .ZN(n7049) );
  OAI211_X1 U8635 ( .C1(n7051), .C2(n9930), .A(n7050), .B(n7049), .ZN(n7053)
         );
  NAND2_X1 U8636 ( .A1(n7053), .A2(n10212), .ZN(n7052) );
  OAI21_X1 U8637 ( .B1(n10212), .B2(n6818), .A(n7052), .ZN(P1_U3475) );
  NAND2_X1 U8638 ( .A1(n7053), .A2(n10223), .ZN(n7054) );
  OAI21_X1 U8639 ( .B1(n10223), .B2(n6819), .A(n7054), .ZN(P1_U3530) );
  INV_X1 U8640 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7704) );
  AOI22_X1 U8641 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(n7698), .B1(n7203), .B2(
        n7704), .ZN(n7060) );
  AOI21_X1 U8642 ( .B1(n7056), .B2(n7535), .A(n7055), .ZN(n7057) );
  NAND2_X1 U8643 ( .A1(n10117), .A2(n7057), .ZN(n7058) );
  XOR2_X1 U8644 ( .A(n10117), .B(n7057), .Z(n10121) );
  NAND2_X1 U8645 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10121), .ZN(n10119) );
  NAND2_X1 U8646 ( .A1(n7058), .A2(n10119), .ZN(n7059) );
  NAND2_X1 U8647 ( .A1(n7060), .A2(n7059), .ZN(n7202) );
  OAI21_X1 U8648 ( .B1(n7060), .B2(n7059), .A(n7202), .ZN(n7074) );
  INV_X1 U8649 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U8650 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9183) );
  OAI21_X1 U8651 ( .B1(n10063), .B2(n7061), .A(n9183), .ZN(n7062) );
  AOI21_X1 U8652 ( .B1(n7698), .B2(n10118), .A(n7062), .ZN(n7073) );
  NAND2_X1 U8653 ( .A1(n7554), .A2(n7063), .ZN(n7065) );
  NAND2_X1 U8654 ( .A1(n7065), .A2(n7064), .ZN(n7066) );
  NAND2_X1 U8655 ( .A1(n10117), .A2(n7066), .ZN(n7067) );
  XOR2_X1 U8656 ( .A(n10117), .B(n7066), .Z(n10125) );
  NAND2_X1 U8657 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n10125), .ZN(n10123) );
  NAND2_X1 U8658 ( .A1(n7067), .A2(n10123), .ZN(n7071) );
  INV_X1 U8659 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7068) );
  MUX2_X1 U8660 ( .A(n7068), .B(P1_REG2_REG_16__SCAN_IN), .S(n7698), .Z(n7069)
         );
  INV_X1 U8661 ( .A(n7069), .ZN(n7070) );
  NAND2_X1 U8662 ( .A1(n7070), .A2(n7071), .ZN(n7208) );
  OAI211_X1 U8663 ( .C1(n7071), .C2(n7070), .A(n10124), .B(n7208), .ZN(n7072)
         );
  OAI211_X1 U8664 ( .C1(n7074), .C2(n10106), .A(n7073), .B(n7072), .ZN(
        P1_U3257) );
  NAND2_X1 U8665 ( .A1(n8189), .A2(n8375), .ZN(n7077) );
  NAND2_X1 U8666 ( .A1(n7078), .A2(n7077), .ZN(n7079) );
  OAI21_X1 U8667 ( .B1(n7079), .B2(n7082), .A(n7223), .ZN(n10394) );
  NAND3_X1 U8668 ( .A1(n7083), .A2(n7082), .A3(n7081), .ZN(n7084) );
  AND2_X1 U8669 ( .A1(n7080), .A2(n7084), .ZN(n7085) );
  OAI222_X1 U8670 ( .A1(n10284), .A2(n7374), .B1(n10286), .B2(n7185), .C1(
        n10281), .C2(n7085), .ZN(n10397) );
  NAND2_X1 U8671 ( .A1(n10397), .A2(n10299), .ZN(n7091) );
  INV_X1 U8672 ( .A(n7188), .ZN(n7086) );
  OAI22_X1 U8673 ( .A1(n10299), .A2(n7087), .B1(n7086), .B2(n10297), .ZN(n7089) );
  XNOR2_X1 U8674 ( .A(n7228), .B(n7227), .ZN(n10396) );
  NOR2_X1 U8675 ( .A1(n10396), .A2(n10273), .ZN(n7088) );
  AOI211_X1 U8676 ( .C1(n10302), .C2(n7227), .A(n7089), .B(n7088), .ZN(n7090)
         );
  OAI211_X1 U8677 ( .C1(n10394), .C2(n8639), .A(n7091), .B(n7090), .ZN(
        P2_U3285) );
  OR2_X1 U8678 ( .A1(n7092), .A2(n9557), .ZN(n7093) );
  NAND2_X1 U8679 ( .A1(n7094), .A2(n7093), .ZN(n7096) );
  NAND2_X1 U8680 ( .A1(n7287), .A2(n7291), .ZN(n9353) );
  AND2_X1 U8681 ( .A1(n9351), .A2(n9353), .ZN(n7100) );
  NAND2_X1 U8682 ( .A1(n7096), .A2(n7100), .ZN(n7097) );
  NAND2_X1 U8683 ( .A1(n7289), .A2(n7097), .ZN(n10195) );
  AOI22_X1 U8684 ( .A1(n9557), .A2(n10137), .B1(n10140), .B2(n9556), .ZN(n7106) );
  INV_X1 U8685 ( .A(n9351), .ZN(n7104) );
  AND2_X1 U8686 ( .A1(n9338), .A2(n9334), .ZN(n9497) );
  NAND2_X1 U8687 ( .A1(n7098), .A2(n9497), .ZN(n7099) );
  AND2_X1 U8688 ( .A1(n9353), .A2(n9336), .ZN(n9499) );
  NAND2_X1 U8689 ( .A1(n7099), .A2(n9499), .ZN(n9280) );
  INV_X1 U8690 ( .A(n7099), .ZN(n7102) );
  INV_X1 U8691 ( .A(n9336), .ZN(n7101) );
  OAI21_X1 U8692 ( .B1(n7102), .B2(n7101), .A(n7095), .ZN(n7103) );
  OAI211_X1 U8693 ( .C1(n7104), .C2(n9280), .A(n7103), .B(n10135), .ZN(n7105)
         );
  OAI211_X1 U8694 ( .C1(n10195), .C2(n10143), .A(n7106), .B(n7105), .ZN(n10198) );
  NAND2_X1 U8695 ( .A1(n10198), .A2(n9810), .ZN(n7114) );
  OAI22_X1 U8696 ( .A1(n9810), .A2(n7108), .B1(n7107), .B2(n10150), .ZN(n7112)
         );
  INV_X1 U8697 ( .A(n7287), .ZN(n10196) );
  OR2_X1 U8698 ( .A1(n7109), .A2(n10196), .ZN(n7110) );
  NAND2_X1 U8699 ( .A1(n7296), .A2(n7110), .ZN(n10197) );
  NOR2_X1 U8700 ( .A1(n10197), .A2(n9832), .ZN(n7111) );
  AOI211_X1 U8701 ( .C1(n9830), .C2(n7287), .A(n7112), .B(n7111), .ZN(n7113)
         );
  OAI211_X1 U8702 ( .C1(n10195), .C2(n7633), .A(n7114), .B(n7113), .ZN(
        P1_U3283) );
  NAND2_X1 U8703 ( .A1(n7115), .A2(n6907), .ZN(n7118) );
  AOI22_X1 U8704 ( .A1(n7803), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7802), .B2(
        n7116), .ZN(n7117) );
  NAND2_X1 U8705 ( .A1(n10203), .A2(n8044), .ZN(n7120) );
  NAND2_X1 U8706 ( .A1(n9556), .A2(n7347), .ZN(n7119) );
  NAND2_X1 U8707 ( .A1(n7120), .A2(n7119), .ZN(n7121) );
  XNOR2_X1 U8708 ( .A(n7121), .B(n8047), .ZN(n7123) );
  AND2_X1 U8709 ( .A1(n9556), .A2(n7928), .ZN(n7122) );
  AOI21_X1 U8710 ( .B1(n10203), .B2(n7347), .A(n7122), .ZN(n7124) );
  NAND2_X1 U8711 ( .A1(n7123), .A2(n7124), .ZN(n7255) );
  INV_X1 U8712 ( .A(n7123), .ZN(n7126) );
  INV_X1 U8713 ( .A(n7124), .ZN(n7125) );
  NAND2_X1 U8714 ( .A1(n7126), .A2(n7125), .ZN(n7127) );
  NAND2_X1 U8715 ( .A1(n7255), .A2(n7127), .ZN(n7136) );
  OAI21_X1 U8716 ( .B1(n7130), .B2(n7129), .A(n7128), .ZN(n7132) );
  NAND2_X1 U8717 ( .A1(n7130), .A2(n7129), .ZN(n7131) );
  INV_X1 U8718 ( .A(n7256), .ZN(n7134) );
  AOI21_X1 U8719 ( .B1(n7136), .B2(n7135), .A(n7134), .ZN(n7142) );
  INV_X1 U8720 ( .A(n7422), .ZN(n7413) );
  NOR2_X1 U8721 ( .A1(n7291), .A2(n9245), .ZN(n7137) );
  AOI211_X1 U8722 ( .C1(n9247), .C2(n7413), .A(n7138), .B(n7137), .ZN(n7139)
         );
  OAI21_X1 U8723 ( .B1(n9249), .B2(n7295), .A(n7139), .ZN(n7140) );
  AOI21_X1 U8724 ( .B1(n10203), .B2(n9251), .A(n7140), .ZN(n7141) );
  OAI21_X1 U8725 ( .B1(n7142), .B2(n9253), .A(n7141), .ZN(P1_U3229) );
  NAND2_X1 U8726 ( .A1(n8228), .A2(n7143), .ZN(n7144) );
  XNOR2_X1 U8727 ( .A(n10375), .B(n8165), .ZN(n7147) );
  NAND2_X1 U8728 ( .A1(n8377), .A2(n8156), .ZN(n7145) );
  XNOR2_X1 U8729 ( .A(n7147), .B(n7145), .ZN(n8226) );
  NAND2_X1 U8730 ( .A1(n7144), .A2(n8226), .ZN(n8230) );
  INV_X1 U8731 ( .A(n7145), .ZN(n7146) );
  NAND2_X1 U8732 ( .A1(n7147), .A2(n7146), .ZN(n7148) );
  NAND2_X1 U8733 ( .A1(n8230), .A2(n7148), .ZN(n7156) );
  XNOR2_X1 U8734 ( .A(n7167), .B(n8212), .ZN(n7150) );
  NAND2_X1 U8735 ( .A1(n8376), .A2(n8156), .ZN(n7151) );
  NAND2_X1 U8736 ( .A1(n7150), .A2(n7151), .ZN(n7149) );
  NAND2_X1 U8737 ( .A1(n7156), .A2(n7149), .ZN(n7153) );
  INV_X1 U8738 ( .A(n7150), .ZN(n7158) );
  INV_X1 U8739 ( .A(n7151), .ZN(n7152) );
  NAND2_X1 U8740 ( .A1(n7158), .A2(n7152), .ZN(n7154) );
  INV_X1 U8741 ( .A(n8186), .ZN(n7159) );
  INV_X1 U8742 ( .A(n7153), .ZN(n7155) );
  NAND2_X1 U8743 ( .A1(n7155), .A2(n7154), .ZN(n7157) );
  AOI22_X1 U8744 ( .A1(n7159), .A2(n7158), .B1(n7157), .B2(n7156), .ZN(n7169)
         );
  INV_X1 U8745 ( .A(n7160), .ZN(n7163) );
  AOI22_X1 U8746 ( .A1(n8287), .A2(n7161), .B1(P2_REG3_REG_9__SCAN_IN), .B2(
        P2_U3152), .ZN(n7162) );
  OAI21_X1 U8747 ( .B1(n7163), .B2(n8355), .A(n7162), .ZN(n7166) );
  NOR3_X1 U8748 ( .A1(n8186), .A2(n7164), .A3(n8345), .ZN(n7165) );
  AOI211_X1 U8749 ( .C1(n7167), .C2(n8360), .A(n7166), .B(n7165), .ZN(n7168)
         );
  OAI21_X1 U8750 ( .B1(n7169), .B2(n8362), .A(n7168), .ZN(P2_U3233) );
  INV_X1 U8751 ( .A(n7227), .ZN(n10395) );
  XNOR2_X1 U8752 ( .A(n8189), .B(n8165), .ZN(n7170) );
  AND2_X1 U8753 ( .A1(n8375), .A2(n8156), .ZN(n7171) );
  NAND2_X1 U8754 ( .A1(n7170), .A2(n7171), .ZN(n7180) );
  INV_X1 U8755 ( .A(n7170), .ZN(n7179) );
  INV_X1 U8756 ( .A(n7171), .ZN(n7172) );
  NAND2_X1 U8757 ( .A1(n7179), .A2(n7172), .ZN(n7173) );
  AND2_X1 U8758 ( .A1(n7180), .A2(n7173), .ZN(n8187) );
  XNOR2_X1 U8759 ( .A(n7227), .B(n8165), .ZN(n7174) );
  AND2_X1 U8760 ( .A1(n8374), .A2(n8156), .ZN(n7175) );
  NAND2_X1 U8761 ( .A1(n7174), .A2(n7175), .ZN(n7308) );
  INV_X1 U8762 ( .A(n7174), .ZN(n7307) );
  INV_X1 U8763 ( .A(n7175), .ZN(n7176) );
  NAND2_X1 U8764 ( .A1(n7307), .A2(n7176), .ZN(n7177) );
  AND2_X1 U8765 ( .A1(n7308), .A2(n7177), .ZN(n7181) );
  INV_X1 U8766 ( .A(n7181), .ZN(n7178) );
  AOI21_X1 U8767 ( .B1(n8185), .B2(n7178), .A(n8362), .ZN(n7184) );
  NOR3_X1 U8768 ( .A1(n7179), .A2(n7185), .A3(n8345), .ZN(n7183) );
  NAND2_X1 U8769 ( .A1(n8185), .A2(n7180), .ZN(n7182) );
  NAND2_X1 U8770 ( .A1(n7182), .A2(n7181), .ZN(n7309) );
  OAI21_X1 U8771 ( .B1(n7184), .B2(n7183), .A(n7309), .ZN(n7190) );
  OAI22_X1 U8772 ( .A1(n8357), .A2(n7374), .B1(n8356), .B2(n7185), .ZN(n7186)
         );
  AOI211_X1 U8773 ( .C1(n8342), .C2(n7188), .A(n7187), .B(n7186), .ZN(n7189)
         );
  OAI211_X1 U8774 ( .C1(n10395), .C2(n8338), .A(n7190), .B(n7189), .ZN(
        P2_U3238) );
  OAI22_X1 U8775 ( .A1(n9799), .A2(n7192), .B1(n7191), .B2(n10150), .ZN(n7199)
         );
  NAND2_X1 U8776 ( .A1(n7200), .A2(n7615), .ZN(n7195) );
  NAND2_X1 U8777 ( .A1(n7193), .A2(n9690), .ZN(n7194) );
  NAND3_X1 U8778 ( .A1(n7196), .A2(n7195), .A3(n7194), .ZN(n7197) );
  MUX2_X1 U8779 ( .A(n7197), .B(P1_REG2_REG_6__SCAN_IN), .S(n10157), .Z(n7198)
         );
  AOI211_X1 U8780 ( .C1(n9834), .C2(n7200), .A(n7199), .B(n7198), .ZN(n7201)
         );
  INV_X1 U8781 ( .A(n7201), .ZN(P1_U3285) );
  INV_X1 U8782 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7717) );
  AOI22_X1 U8783 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(n7770), .B1(n7380), .B2(
        n7717), .ZN(n7205) );
  OAI21_X1 U8784 ( .B1(n7203), .B2(n7704), .A(n7202), .ZN(n7204) );
  NAND2_X1 U8785 ( .A1(n7205), .A2(n7204), .ZN(n7379) );
  OAI21_X1 U8786 ( .B1(n7205), .B2(n7204), .A(n7379), .ZN(n7216) );
  INV_X1 U8787 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7206) );
  NAND2_X1 U8788 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9194) );
  OAI21_X1 U8789 ( .B1(n10063), .B2(n7206), .A(n9194), .ZN(n7207) );
  AOI21_X1 U8790 ( .B1(n7770), .B2(n10118), .A(n7207), .ZN(n7215) );
  NAND2_X1 U8791 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7698), .ZN(n7209) );
  NAND2_X1 U8792 ( .A1(n7209), .A2(n7208), .ZN(n7213) );
  INV_X1 U8793 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7211) );
  NAND2_X1 U8794 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n7770), .ZN(n7386) );
  INV_X1 U8795 ( .A(n7386), .ZN(n7210) );
  AOI21_X1 U8796 ( .B1(n7211), .B2(n7380), .A(n7210), .ZN(n7212) );
  NAND2_X1 U8797 ( .A1(n7212), .A2(n7213), .ZN(n7385) );
  OAI211_X1 U8798 ( .C1(n7213), .C2(n7212), .A(n10124), .B(n7385), .ZN(n7214)
         );
  OAI211_X1 U8799 ( .C1(n7216), .C2(n10106), .A(n7215), .B(n7214), .ZN(
        P1_U3258) );
  NAND2_X1 U8800 ( .A1(n7080), .A2(n7217), .ZN(n7218) );
  INV_X1 U8801 ( .A(n7225), .ZN(n7224) );
  XNOR2_X1 U8802 ( .A(n7218), .B(n7224), .ZN(n7219) );
  NAND2_X1 U8803 ( .A1(n7219), .A2(n10264), .ZN(n7221) );
  AOI22_X1 U8804 ( .A1(n10259), .A2(n8374), .B1(n8372), .B2(n10261), .ZN(n7220) );
  NAND2_X1 U8805 ( .A1(n7221), .A2(n7220), .ZN(n10404) );
  INV_X1 U8806 ( .A(n10404), .ZN(n7233) );
  NAND2_X1 U8807 ( .A1(n7227), .A2(n8374), .ZN(n7222) );
  OAI21_X1 U8808 ( .B1(n7226), .B2(n7225), .A(n7395), .ZN(n10406) );
  INV_X1 U8809 ( .A(n7393), .ZN(n10401) );
  OAI21_X1 U8810 ( .B1(n10401), .B2(n4567), .A(n4726), .ZN(n10403) );
  AOI22_X1 U8811 ( .A1(n10308), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7316), .B2(
        n10245), .ZN(n7230) );
  NAND2_X1 U8812 ( .A1(n7393), .A2(n10302), .ZN(n7229) );
  OAI211_X1 U8813 ( .C1(n10403), .C2(n10273), .A(n7230), .B(n7229), .ZN(n7231)
         );
  AOI21_X1 U8814 ( .B1(n10406), .B2(n10306), .A(n7231), .ZN(n7232) );
  OAI21_X1 U8815 ( .B1(n10308), .B2(n7233), .A(n7232), .ZN(P2_U3284) );
  NAND2_X1 U8816 ( .A1(n7235), .A2(n7234), .ZN(n7237) );
  NAND2_X1 U8817 ( .A1(n7237), .A2(n7236), .ZN(n7240) );
  INV_X1 U8818 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7238) );
  MUX2_X1 U8819 ( .A(n7238), .B(P2_REG1_REG_16__SCAN_IN), .S(n8071), .Z(n7239)
         );
  NOR2_X1 U8820 ( .A1(n7239), .A2(n7240), .ZN(n8072) );
  AOI21_X1 U8821 ( .B1(n7240), .B2(n7239), .A(n8072), .ZN(n7254) );
  NAND2_X1 U8822 ( .A1(n7242), .A2(n7241), .ZN(n7244) );
  NAND2_X1 U8823 ( .A1(n7244), .A2(n7243), .ZN(n7247) );
  NAND2_X1 U8824 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8071), .ZN(n7245) );
  OAI21_X1 U8825 ( .B1(n8071), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7245), .ZN(
        n7246) );
  AOI211_X1 U8826 ( .C1(n7247), .C2(n7246), .A(n8066), .B(n9986), .ZN(n7252)
         );
  NOR2_X1 U8827 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8276), .ZN(n7248) );
  AOI21_X1 U8828 ( .B1(n10231), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7248), .ZN(
        n7249) );
  OAI21_X1 U8829 ( .B1(n10227), .B2(n7250), .A(n7249), .ZN(n7251) );
  NOR2_X1 U8830 ( .A1(n7252), .A2(n7251), .ZN(n7253) );
  OAI21_X1 U8831 ( .B1(n7254), .B2(n10229), .A(n7253), .ZN(P2_U3261) );
  NAND2_X1 U8832 ( .A1(n7257), .A2(n6907), .ZN(n7259) );
  AOI22_X1 U8833 ( .A1(n7803), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7802), .B2(
        n10101), .ZN(n7258) );
  NAND2_X1 U8834 ( .A1(n10001), .A2(n8044), .ZN(n7261) );
  OR2_X1 U8835 ( .A1(n7422), .A2(n7945), .ZN(n7260) );
  NAND2_X1 U8836 ( .A1(n7261), .A2(n7260), .ZN(n7262) );
  XNOR2_X1 U8837 ( .A(n7262), .B(n7947), .ZN(n7265) );
  NAND2_X1 U8838 ( .A1(n10001), .A2(n7347), .ZN(n7264) );
  OR2_X1 U8839 ( .A1(n7422), .A2(n7943), .ZN(n7263) );
  NAND2_X1 U8840 ( .A1(n7264), .A2(n7263), .ZN(n7266) );
  NAND2_X1 U8841 ( .A1(n7265), .A2(n7266), .ZN(n7343) );
  INV_X1 U8842 ( .A(n7265), .ZN(n7268) );
  INV_X1 U8843 ( .A(n7266), .ZN(n7267) );
  NAND2_X1 U8844 ( .A1(n7268), .A2(n7267), .ZN(n7345) );
  NAND2_X1 U8845 ( .A1(n7343), .A2(n7345), .ZN(n7269) );
  XNOR2_X1 U8846 ( .A(n7344), .B(n7269), .ZN(n7283) );
  NOR2_X1 U8847 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7270), .ZN(n10102) );
  NAND2_X1 U8848 ( .A1(n6431), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7278) );
  OR2_X1 U8849 ( .A1(n4478), .A2(n10057), .ZN(n7277) );
  INV_X1 U8850 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7271) );
  NAND2_X1 U8851 ( .A1(n7272), .A2(n7271), .ZN(n7273) );
  NAND2_X1 U8852 ( .A1(n7274), .A2(n7273), .ZN(n7426) );
  OR2_X1 U8853 ( .A1(n6527), .A2(n7426), .ZN(n7276) );
  OR2_X1 U8854 ( .A1(n4476), .A2(n6084), .ZN(n7275) );
  NAND4_X1 U8855 ( .A1(n7278), .A2(n7277), .A3(n7276), .A4(n7275), .ZN(n9555)
         );
  INV_X1 U8856 ( .A(n9555), .ZN(n7491) );
  NOR2_X1 U8857 ( .A1(n7491), .A2(n9234), .ZN(n7279) );
  AOI211_X1 U8858 ( .C1(n9236), .C2(n9556), .A(n10102), .B(n7279), .ZN(n7280)
         );
  OAI21_X1 U8859 ( .B1(n9249), .B2(n7330), .A(n7280), .ZN(n7281) );
  AOI21_X1 U8860 ( .B1(n10001), .B2(n9251), .A(n7281), .ZN(n7282) );
  OAI21_X1 U8861 ( .B1(n7283), .B2(n9253), .A(n7282), .ZN(P1_U3215) );
  INV_X1 U8862 ( .A(n7823), .ZN(n7285) );
  OAI222_X1 U8863 ( .A1(P1_U3084), .A2(n9528), .B1(n9971), .B2(n7285), .C1(
        n7824), .C2(n9968), .ZN(P1_U3333) );
  OAI222_X1 U8864 ( .A1(P2_U3152), .A2(n5662), .B1(n9139), .B2(n7285), .C1(
        n7284), .C2(n9137), .ZN(P2_U3338) );
  NAND2_X1 U8865 ( .A1(n7287), .A2(n7286), .ZN(n7288) );
  INV_X1 U8866 ( .A(n9556), .ZN(n7290) );
  OR2_X1 U8867 ( .A1(n10203), .A2(n7290), .ZN(n9345) );
  NAND2_X1 U8868 ( .A1(n10203), .A2(n7290), .ZN(n9265) );
  NAND2_X1 U8869 ( .A1(n9345), .A2(n9265), .ZN(n9307) );
  XNOR2_X1 U8870 ( .A(n7320), .B(n9307), .ZN(n10202) );
  NAND2_X1 U8871 ( .A1(n9280), .A2(n9351), .ZN(n7321) );
  XNOR2_X1 U8872 ( .A(n7321), .B(n9307), .ZN(n7293) );
  OAI22_X1 U8873 ( .A1(n7291), .A2(n9818), .B1(n7422), .B2(n9816), .ZN(n7292)
         );
  AOI21_X1 U8874 ( .B1(n7293), .B2(n10135), .A(n7292), .ZN(n7294) );
  OAI21_X1 U8875 ( .B1(n10202), .B2(n10143), .A(n7294), .ZN(n10207) );
  NAND2_X1 U8876 ( .A1(n10207), .A2(n9810), .ZN(n7301) );
  OAI22_X1 U8877 ( .A1(n9810), .A2(n6917), .B1(n7295), .B2(n10150), .ZN(n7299)
         );
  NAND2_X1 U8878 ( .A1(n7296), .A2(n10203), .ZN(n7297) );
  NAND2_X1 U8879 ( .A1(n7327), .A2(n7297), .ZN(n10206) );
  NOR2_X1 U8880 ( .A1(n10206), .A2(n9832), .ZN(n7298) );
  AOI211_X1 U8881 ( .C1(n9830), .C2(n10203), .A(n7299), .B(n7298), .ZN(n7300)
         );
  OAI211_X1 U8882 ( .C1(n10202), .C2(n7633), .A(n7301), .B(n7300), .ZN(
        P1_U3282) );
  XNOR2_X1 U8883 ( .A(n7393), .B(n8165), .ZN(n7302) );
  AND2_X1 U8884 ( .A1(n8373), .A2(n8156), .ZN(n7303) );
  NAND2_X1 U8885 ( .A1(n7302), .A2(n7303), .ZN(n7368) );
  INV_X1 U8886 ( .A(n7302), .ZN(n7367) );
  INV_X1 U8887 ( .A(n7303), .ZN(n7304) );
  NAND2_X1 U8888 ( .A1(n7367), .A2(n7304), .ZN(n7305) );
  AND2_X1 U8889 ( .A1(n7368), .A2(n7305), .ZN(n7310) );
  INV_X1 U8890 ( .A(n7310), .ZN(n7306) );
  AOI21_X1 U8891 ( .B1(n7309), .B2(n7306), .A(n8362), .ZN(n7313) );
  NOR3_X1 U8892 ( .A1(n7307), .A2(n7314), .A3(n8345), .ZN(n7312) );
  NAND2_X1 U8893 ( .A1(n7309), .A2(n7308), .ZN(n7311) );
  NAND2_X1 U8894 ( .A1(n7311), .A2(n7310), .ZN(n7369) );
  OAI21_X1 U8895 ( .B1(n7313), .B2(n7312), .A(n7369), .ZN(n7318) );
  AND2_X1 U8896 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8412) );
  OAI22_X1 U8897 ( .A1(n8357), .A2(n7503), .B1(n8356), .B2(n7314), .ZN(n7315)
         );
  AOI211_X1 U8898 ( .C1(n7316), .C2(n8342), .A(n8412), .B(n7315), .ZN(n7317)
         );
  OAI211_X1 U8899 ( .C1(n10401), .C2(n8338), .A(n7318), .B(n7317), .ZN(
        P2_U3226) );
  AND2_X1 U8900 ( .A1(n10203), .A2(n9556), .ZN(n7319) );
  OR2_X1 U8901 ( .A1(n10001), .A2(n7422), .ZN(n9348) );
  NAND2_X1 U8902 ( .A1(n10001), .A2(n7422), .ZN(n9357) );
  NAND2_X1 U8903 ( .A1(n9348), .A2(n9357), .ZN(n9310) );
  XNOR2_X1 U8904 ( .A(n7412), .B(n9310), .ZN(n10005) );
  NAND2_X1 U8905 ( .A1(n7321), .A2(n9265), .ZN(n7420) );
  NAND2_X1 U8906 ( .A1(n7420), .A2(n9345), .ZN(n7323) );
  INV_X1 U8907 ( .A(n9310), .ZN(n7322) );
  XNOR2_X1 U8908 ( .A(n7323), .B(n7322), .ZN(n7325) );
  AOI22_X1 U8909 ( .A1(n10137), .A2(n9556), .B1(n9555), .B2(n10140), .ZN(n7324) );
  OAI21_X1 U8910 ( .B1(n7325), .B2(n9807), .A(n7324), .ZN(n7326) );
  AOI21_X1 U8911 ( .B1(n10005), .B2(n7615), .A(n7326), .ZN(n10007) );
  NAND2_X1 U8912 ( .A1(n7327), .A2(n10001), .ZN(n7328) );
  NAND2_X1 U8913 ( .A1(n7328), .A2(n10146), .ZN(n7329) );
  OR2_X1 U8914 ( .A1(n7427), .A2(n7329), .ZN(n10003) );
  INV_X1 U8915 ( .A(n7714), .ZN(n7498) );
  OAI22_X1 U8916 ( .A1(n9810), .A2(n7331), .B1(n7330), .B2(n10150), .ZN(n7332)
         );
  AOI21_X1 U8917 ( .B1(n10001), .B2(n9830), .A(n7332), .ZN(n7333) );
  OAI21_X1 U8918 ( .B1(n10003), .B2(n7498), .A(n7333), .ZN(n7334) );
  AOI21_X1 U8919 ( .B1(n10005), .B2(n9834), .A(n7334), .ZN(n7335) );
  OAI21_X1 U8920 ( .B1(n10007), .B2(n10157), .A(n7335), .ZN(P1_U3281) );
  INV_X1 U8921 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7337) );
  INV_X1 U8922 ( .A(n7842), .ZN(n7338) );
  OAI222_X1 U8923 ( .A1(n9137), .A2(n7337), .B1(n9139), .B2(n7338), .C1(n7336), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U8924 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7843) );
  OAI222_X1 U8925 ( .A1(n9968), .A2(n7843), .B1(P1_U3084), .B2(n9472), .C1(
        n9971), .C2(n7338), .ZN(P1_U3332) );
  NAND2_X1 U8926 ( .A1(n7339), .A2(n6907), .ZN(n7342) );
  AOI22_X1 U8927 ( .A1(n7803), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7802), .B2(
        n7340), .ZN(n7341) );
  NAND2_X1 U8928 ( .A1(n7344), .A2(n7343), .ZN(n7346) );
  NAND2_X1 U8929 ( .A1(n7489), .A2(n8044), .ZN(n7349) );
  NAND2_X1 U8930 ( .A1(n9555), .A2(n7347), .ZN(n7348) );
  NAND2_X1 U8931 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  XNOR2_X1 U8932 ( .A(n7350), .B(n8047), .ZN(n7463) );
  AND2_X1 U8933 ( .A1(n9555), .A2(n7928), .ZN(n7351) );
  AOI21_X1 U8934 ( .B1(n7489), .B2(n7347), .A(n7351), .ZN(n7464) );
  XNOR2_X1 U8935 ( .A(n7463), .B(n7464), .ZN(n7353) );
  AOI21_X1 U8936 ( .B1(n7352), .B2(n7353), .A(n9253), .ZN(n7355) );
  NAND2_X1 U8937 ( .A1(n7355), .A2(n7468), .ZN(n7361) );
  INV_X1 U8938 ( .A(n7426), .ZN(n7359) );
  AOI21_X1 U8939 ( .B1(n7413), .B2(n9236), .A(n7356), .ZN(n7357) );
  OAI21_X1 U8940 ( .B1(n7619), .B2(n9234), .A(n7357), .ZN(n7358) );
  AOI21_X1 U8941 ( .B1(n7359), .B2(n9203), .A(n7358), .ZN(n7360) );
  OAI211_X1 U8942 ( .C1(n10053), .C2(n9218), .A(n7361), .B(n7360), .ZN(
        P1_U3234) );
  INV_X1 U8943 ( .A(n7435), .ZN(n10033) );
  XNOR2_X1 U8944 ( .A(n7435), .B(n8165), .ZN(n7362) );
  AND2_X1 U8945 ( .A1(n8372), .A2(n8156), .ZN(n7363) );
  NAND2_X1 U8946 ( .A1(n7362), .A2(n7363), .ZN(n7510) );
  INV_X1 U8947 ( .A(n7362), .ZN(n7504) );
  INV_X1 U8948 ( .A(n7363), .ZN(n7364) );
  NAND2_X1 U8949 ( .A1(n7504), .A2(n7364), .ZN(n7365) );
  AND2_X1 U8950 ( .A1(n7510), .A2(n7365), .ZN(n7370) );
  INV_X1 U8951 ( .A(n7370), .ZN(n7366) );
  AOI21_X1 U8952 ( .B1(n7369), .B2(n7366), .A(n8362), .ZN(n7373) );
  NOR3_X1 U8953 ( .A1(n7367), .A2(n7374), .A3(n8345), .ZN(n7372) );
  NAND2_X1 U8954 ( .A1(n7369), .A2(n7368), .ZN(n7371) );
  NAND2_X1 U8955 ( .A1(n7371), .A2(n7370), .ZN(n7512) );
  OAI21_X1 U8956 ( .B1(n7373), .B2(n7372), .A(n7512), .ZN(n7378) );
  OAI22_X1 U8957 ( .A1(n8357), .A2(n7603), .B1(n8356), .B2(n7374), .ZN(n7375)
         );
  AOI211_X1 U8958 ( .C1(n8342), .C2(n7406), .A(n7376), .B(n7375), .ZN(n7377)
         );
  OAI211_X1 U8959 ( .C1(n10033), .C2(n8338), .A(n7378), .B(n7377), .ZN(
        P2_U3236) );
  INV_X1 U8960 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9583) );
  AOI22_X1 U8961 ( .A1(n7782), .A2(n9583), .B1(P1_REG1_REG_18__SCAN_IN), .B2(
        n9587), .ZN(n7382) );
  OAI21_X1 U8962 ( .B1(n7380), .B2(n7717), .A(n7379), .ZN(n7381) );
  NOR2_X1 U8963 ( .A1(n7382), .A2(n7381), .ZN(n9582) );
  AOI21_X1 U8964 ( .B1(n7382), .B2(n7381), .A(n9582), .ZN(n7391) );
  INV_X1 U8965 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n7383) );
  NAND2_X1 U8966 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9233) );
  OAI21_X1 U8967 ( .B1(n10063), .B2(n7383), .A(n9233), .ZN(n7384) );
  AOI21_X1 U8968 ( .B1(n7782), .B2(n10118), .A(n7384), .ZN(n7390) );
  NAND2_X1 U8969 ( .A1(n7386), .A2(n7385), .ZN(n7388) );
  XNOR2_X1 U8970 ( .A(n9587), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n7387) );
  NAND2_X1 U8971 ( .A1(n7387), .A2(n7388), .ZN(n9586) );
  OAI211_X1 U8972 ( .C1(n7388), .C2(n7387), .A(n10124), .B(n9586), .ZN(n7389)
         );
  OAI211_X1 U8973 ( .C1(n7391), .C2(n10106), .A(n7390), .B(n7389), .ZN(
        P1_U3259) );
  INV_X1 U8974 ( .A(n7860), .ZN(n7392) );
  OAI222_X1 U8975 ( .A1(n9968), .A2(n7861), .B1(n9971), .B2(n7392), .C1(
        P1_U3084), .C2(n9536), .ZN(P1_U3331) );
  OAI222_X1 U8976 ( .A1(n9137), .A2(n8865), .B1(n9134), .B2(n7392), .C1(
        P2_U3152), .C2(n9035), .ZN(P2_U3336) );
  OR2_X1 U8977 ( .A1(n7393), .A2(n8373), .ZN(n7394) );
  AND2_X1 U8978 ( .A1(n7396), .A2(n5012), .ZN(n7397) );
  OR2_X1 U8979 ( .A1(n7397), .A2(n7434), .ZN(n7403) );
  AOI22_X1 U8980 ( .A1(n10259), .A2(n8373), .B1(n8371), .B2(n10261), .ZN(n7402) );
  XNOR2_X1 U8981 ( .A(n7398), .B(n7399), .ZN(n7400) );
  NAND2_X1 U8982 ( .A1(n7400), .A2(n10264), .ZN(n7401) );
  OAI211_X1 U8983 ( .C1(n7403), .C2(n10241), .A(n7402), .B(n7401), .ZN(n10035)
         );
  INV_X1 U8984 ( .A(n10035), .ZN(n7411) );
  INV_X1 U8985 ( .A(n7403), .ZN(n10037) );
  INV_X1 U8986 ( .A(n7587), .ZN(n7404) );
  OAI21_X1 U8987 ( .B1(n10033), .B2(n7405), .A(n7404), .ZN(n10034) );
  AOI22_X1 U8988 ( .A1(n10308), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7406), .B2(
        n10245), .ZN(n7408) );
  NAND2_X1 U8989 ( .A1(n7435), .A2(n10302), .ZN(n7407) );
  OAI211_X1 U8990 ( .C1(n10034), .C2(n10273), .A(n7408), .B(n7407), .ZN(n7409)
         );
  AOI21_X1 U8991 ( .B1(n10037), .B2(n10251), .A(n7409), .ZN(n7410) );
  OAI21_X1 U8992 ( .B1(n7411), .B2(n10308), .A(n7410), .ZN(P2_U3283) );
  NAND2_X1 U8993 ( .A1(n7412), .A2(n9310), .ZN(n7415) );
  OR2_X1 U8994 ( .A1(n10001), .A2(n7413), .ZN(n7414) );
  NAND2_X1 U8995 ( .A1(n7415), .A2(n7414), .ZN(n7418) );
  INV_X1 U8996 ( .A(n7418), .ZN(n7417) );
  XNOR2_X1 U8997 ( .A(n7489), .B(n9555), .ZN(n9361) );
  INV_X1 U8998 ( .A(n9361), .ZN(n7416) );
  NAND2_X1 U8999 ( .A1(n7417), .A2(n7416), .ZN(n7486) );
  NAND2_X1 U9000 ( .A1(n7418), .A2(n9361), .ZN(n7419) );
  NAND2_X1 U9001 ( .A1(n7486), .A2(n7419), .ZN(n10051) );
  AND2_X1 U9002 ( .A1(n9348), .A2(n9345), .ZN(n9356) );
  NAND2_X1 U9003 ( .A1(n7420), .A2(n9356), .ZN(n7421) );
  NAND2_X1 U9004 ( .A1(n7421), .A2(n9357), .ZN(n7563) );
  XNOR2_X1 U9005 ( .A(n7563), .B(n9361), .ZN(n7424) );
  OAI22_X1 U9006 ( .A1(n7619), .A2(n9816), .B1(n7422), .B2(n9818), .ZN(n7423)
         );
  AOI21_X1 U9007 ( .B1(n7424), .B2(n10135), .A(n7423), .ZN(n7425) );
  OAI21_X1 U9008 ( .B1(n10051), .B2(n10143), .A(n7425), .ZN(n10054) );
  NAND2_X1 U9009 ( .A1(n10054), .A2(n9810), .ZN(n7433) );
  OAI22_X1 U9010 ( .A1(n9810), .A2(n6084), .B1(n7426), .B2(n10150), .ZN(n7431)
         );
  NOR2_X1 U9011 ( .A1(n7427), .A2(n10053), .ZN(n7428) );
  OR3_X1 U9012 ( .A1(n7497), .A2(n7428), .A3(n10205), .ZN(n10052) );
  NOR2_X1 U9013 ( .A1(n10157), .A2(n10148), .ZN(n9804) );
  INV_X1 U9014 ( .A(n9804), .ZN(n7429) );
  NOR2_X1 U9015 ( .A1(n10052), .A2(n7429), .ZN(n7430) );
  AOI211_X1 U9016 ( .C1(n9830), .C2(n7489), .A(n7431), .B(n7430), .ZN(n7432)
         );
  OAI211_X1 U9017 ( .C1(n10051), .C2(n7633), .A(n7433), .B(n7432), .ZN(
        P1_U3280) );
  NAND2_X1 U9018 ( .A1(n7437), .A2(n7436), .ZN(n7580) );
  OAI21_X1 U9019 ( .B1(n7437), .B2(n7436), .A(n7580), .ZN(n10031) );
  INV_X1 U9020 ( .A(n10031), .ZN(n7448) );
  OAI211_X1 U9021 ( .C1(n4558), .C2(n7439), .A(n10264), .B(n7438), .ZN(n7441)
         );
  AOI22_X1 U9022 ( .A1(n10259), .A2(n8372), .B1(n8648), .B2(n10261), .ZN(n7440) );
  NAND2_X1 U9023 ( .A1(n7441), .A2(n7440), .ZN(n10030) );
  INV_X1 U9024 ( .A(n7581), .ZN(n10027) );
  XNOR2_X1 U9025 ( .A(n7587), .B(n10027), .ZN(n10028) );
  INV_X1 U9026 ( .A(n7442), .ZN(n7509) );
  OAI22_X1 U9027 ( .A1(n10299), .A2(n7443), .B1(n7509), .B2(n10297), .ZN(n7444) );
  AOI21_X1 U9028 ( .B1(n7581), .B2(n10302), .A(n7444), .ZN(n7445) );
  OAI21_X1 U9029 ( .B1(n10028), .B2(n10273), .A(n7445), .ZN(n7446) );
  AOI21_X1 U9030 ( .B1(n10030), .B2(n10299), .A(n7446), .ZN(n7447) );
  OAI21_X1 U9031 ( .B1(n7448), .B2(n8639), .A(n7447), .ZN(P2_U3282) );
  INV_X1 U9032 ( .A(n7880), .ZN(n7454) );
  AOI21_X1 U9033 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9129), .A(n7449), .ZN(
        n7450) );
  OAI21_X1 U9034 ( .B1(n7454), .B2(n9134), .A(n7450), .ZN(P2_U3335) );
  NOR2_X1 U9035 ( .A1(n7451), .A2(P1_U3084), .ZN(n9537) );
  AOI21_X1 U9036 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n7452), .A(n9537), .ZN(
        n7453) );
  OAI21_X1 U9037 ( .B1(n7454), .B2(n9971), .A(n7453), .ZN(P1_U3330) );
  NAND2_X1 U9038 ( .A1(n7455), .A2(n6907), .ZN(n7458) );
  AOI22_X1 U9039 ( .A1(n7803), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7802), .B2(
        n7456), .ZN(n7457) );
  NAND2_X1 U9040 ( .A1(n7547), .A2(n8044), .ZN(n7460) );
  OR2_X1 U9041 ( .A1(n7619), .A2(n7945), .ZN(n7459) );
  NAND2_X1 U9042 ( .A1(n7460), .A2(n7459), .ZN(n7461) );
  XNOR2_X1 U9043 ( .A(n7461), .B(n8047), .ZN(n7519) );
  NOR2_X1 U9044 ( .A1(n7619), .A2(n7943), .ZN(n7462) );
  AOI21_X1 U9045 ( .B1(n7547), .B2(n7347), .A(n7462), .ZN(n7518) );
  XNOR2_X1 U9046 ( .A(n7519), .B(n7518), .ZN(n7471) );
  INV_X1 U9047 ( .A(n7463), .ZN(n7466) );
  INV_X1 U9048 ( .A(n7464), .ZN(n7465) );
  NAND2_X1 U9049 ( .A1(n7466), .A2(n7465), .ZN(n7467) );
  INV_X1 U9050 ( .A(n7521), .ZN(n7469) );
  AOI21_X1 U9051 ( .B1(n7471), .B2(n7470), .A(n7469), .ZN(n7484) );
  NAND2_X1 U9052 ( .A1(n7473), .A2(n7472), .ZN(n7474) );
  NAND2_X1 U9053 ( .A1(n7532), .A2(n7474), .ZN(n7627) );
  OR2_X1 U9054 ( .A1(n6527), .A2(n7627), .ZN(n7475) );
  OAI21_X1 U9055 ( .B1(n4476), .B2(n6405), .A(n7475), .ZN(n7479) );
  INV_X1 U9056 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8771) );
  NOR2_X1 U9057 ( .A1(n6557), .A2(n8771), .ZN(n7478) );
  NOR2_X1 U9058 ( .A1(n4478), .A2(n7476), .ZN(n7477) );
  AOI22_X1 U9059 ( .A1(n9247), .A2(n9554), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7481) );
  NAND2_X1 U9060 ( .A1(n9236), .A2(n9555), .ZN(n7480) );
  OAI211_X1 U9061 ( .C1(n9249), .C2(n7495), .A(n7481), .B(n7480), .ZN(n7482)
         );
  AOI21_X1 U9062 ( .B1(n7547), .B2(n9251), .A(n7482), .ZN(n7483) );
  OAI21_X1 U9063 ( .B1(n7484), .B2(n9253), .A(n7483), .ZN(P1_U3222) );
  NAND2_X1 U9064 ( .A1(n7489), .A2(n9555), .ZN(n7485) );
  NAND2_X1 U9065 ( .A1(n7486), .A2(n7485), .ZN(n7487) );
  OR2_X1 U9066 ( .A1(n7547), .A2(n7619), .ZN(n9369) );
  NAND2_X1 U9067 ( .A1(n7547), .A2(n7619), .ZN(n9363) );
  NAND2_X1 U9068 ( .A1(n9369), .A2(n9363), .ZN(n9297) );
  NAND2_X1 U9069 ( .A1(n7487), .A2(n9297), .ZN(n7549) );
  OR2_X1 U9070 ( .A1(n7487), .A2(n9297), .ZN(n7488) );
  NAND2_X1 U9071 ( .A1(n7549), .A2(n7488), .ZN(n10044) );
  OR2_X1 U9072 ( .A1(n7489), .A2(n7491), .ZN(n7562) );
  AND2_X1 U9073 ( .A1(n7489), .A2(n7491), .ZN(n9263) );
  AOI21_X1 U9074 ( .B1(n7563), .B2(n7562), .A(n9263), .ZN(n7490) );
  XNOR2_X1 U9075 ( .A(n7490), .B(n9297), .ZN(n7493) );
  INV_X1 U9076 ( .A(n9554), .ZN(n7565) );
  OAI22_X1 U9077 ( .A1(n7565), .A2(n9816), .B1(n7491), .B2(n9818), .ZN(n7492)
         );
  AOI21_X1 U9078 ( .B1(n7493), .B2(n10135), .A(n7492), .ZN(n7494) );
  OAI21_X1 U9079 ( .B1(n10044), .B2(n10143), .A(n7494), .ZN(n10047) );
  NAND2_X1 U9080 ( .A1(n10047), .A2(n9810), .ZN(n7502) );
  OAI22_X1 U9081 ( .A1(n9810), .A2(n7496), .B1(n7495), .B2(n10150), .ZN(n7500)
         );
  INV_X1 U9082 ( .A(n7547), .ZN(n10046) );
  NAND2_X1 U9083 ( .A1(n7497), .A2(n10046), .ZN(n7624) );
  OAI211_X1 U9084 ( .C1(n7497), .C2(n10046), .A(n10146), .B(n7624), .ZN(n10045) );
  NOR2_X1 U9085 ( .A1(n10045), .A2(n7498), .ZN(n7499) );
  AOI211_X1 U9086 ( .C1(n9830), .C2(n7547), .A(n7500), .B(n7499), .ZN(n7501)
         );
  OAI211_X1 U9087 ( .C1(n10044), .C2(n7633), .A(n7502), .B(n7501), .ZN(
        P1_U3279) );
  XNOR2_X1 U9088 ( .A(n7581), .B(n8165), .ZN(n7596) );
  NAND2_X1 U9089 ( .A1(n8371), .A2(n4486), .ZN(n7597) );
  XNOR2_X1 U9090 ( .A(n7596), .B(n7597), .ZN(n7517) );
  INV_X1 U9091 ( .A(n7512), .ZN(n7506) );
  NOR3_X1 U9092 ( .A1(n7504), .A2(n7503), .A3(n8345), .ZN(n7505) );
  AOI21_X1 U9093 ( .B1(n7506), .B2(n8336), .A(n7505), .ZN(n7516) );
  AOI22_X1 U9094 ( .A1(n8318), .A2(n8648), .B1(n8346), .B2(n8372), .ZN(n7508)
         );
  OAI211_X1 U9095 ( .C1(n8355), .C2(n7509), .A(n7508), .B(n7507), .ZN(n7514)
         );
  AND2_X1 U9096 ( .A1(n7517), .A2(n7510), .ZN(n7511) );
  NOR2_X1 U9097 ( .A1(n7600), .A2(n8362), .ZN(n7513) );
  AOI211_X1 U9098 ( .C1(n7581), .C2(n8360), .A(n7514), .B(n7513), .ZN(n7515)
         );
  OAI21_X1 U9099 ( .B1(n7517), .B2(n7516), .A(n7515), .ZN(P2_U3217) );
  NAND2_X1 U9100 ( .A1(n7519), .A2(n7518), .ZN(n7520) );
  NAND2_X1 U9101 ( .A1(n7522), .A2(n6907), .ZN(n7525) );
  AOI22_X1 U9102 ( .A1(n7803), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7802), .B2(
        n7523), .ZN(n7524) );
  NAND2_X1 U9103 ( .A1(n9932), .A2(n8044), .ZN(n7527) );
  NAND2_X1 U9104 ( .A1(n9554), .A2(n7347), .ZN(n7526) );
  NAND2_X1 U9105 ( .A1(n7527), .A2(n7526), .ZN(n7528) );
  XNOR2_X1 U9106 ( .A(n7528), .B(n8047), .ZN(n7636) );
  AND2_X1 U9107 ( .A1(n9554), .A2(n7928), .ZN(n7529) );
  AOI21_X1 U9108 ( .B1(n9932), .B2(n7347), .A(n7529), .ZN(n7637) );
  XNOR2_X1 U9109 ( .A(n7636), .B(n7637), .ZN(n7530) );
  XNOR2_X1 U9110 ( .A(n7635), .B(n7530), .ZN(n7545) );
  INV_X1 U9111 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U9112 ( .A1(n7532), .A2(n7531), .ZN(n7533) );
  NAND2_X1 U9113 ( .A1(n7570), .A2(n7533), .ZN(n7649) );
  OR2_X1 U9114 ( .A1(n6527), .A2(n7649), .ZN(n7534) );
  OAI21_X1 U9115 ( .B1(n4477), .B2(n7559), .A(n7534), .ZN(n7539) );
  NOR2_X1 U9116 ( .A1(n4479), .A2(n7535), .ZN(n7538) );
  INV_X1 U9117 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7536) );
  NOR2_X1 U9118 ( .A1(n6557), .A2(n7536), .ZN(n7537) );
  NOR2_X1 U9119 ( .A1(n7619), .A2(n9245), .ZN(n7540) );
  AOI211_X1 U9120 ( .C1(n9247), .C2(n9553), .A(n7541), .B(n7540), .ZN(n7542)
         );
  OAI21_X1 U9121 ( .B1(n9249), .B2(n7627), .A(n7542), .ZN(n7543) );
  AOI21_X1 U9122 ( .B1(n9932), .B2(n9251), .A(n7543), .ZN(n7544) );
  OAI21_X1 U9123 ( .B1(n7545), .B2(n9253), .A(n7544), .ZN(P1_U3232) );
  INV_X1 U9124 ( .A(n7619), .ZN(n7546) );
  NAND2_X1 U9125 ( .A1(n7547), .A2(n7546), .ZN(n7548) );
  NAND2_X1 U9126 ( .A1(n7549), .A2(n7548), .ZN(n7614) );
  OR2_X1 U9127 ( .A1(n9932), .A2(n9554), .ZN(n7550) );
  NAND2_X1 U9128 ( .A1(n7614), .A2(n7550), .ZN(n7552) );
  NAND2_X1 U9129 ( .A1(n9932), .A2(n9554), .ZN(n7551) );
  NAND2_X1 U9130 ( .A1(n7552), .A2(n7551), .ZN(n7692) );
  NAND2_X1 U9131 ( .A1(n7553), .A2(n6907), .ZN(n7556) );
  AOI22_X1 U9132 ( .A1(n7803), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7802), .B2(
        n7554), .ZN(n7555) );
  INV_X1 U9133 ( .A(n9553), .ZN(n9819) );
  NAND2_X1 U9134 ( .A1(n9928), .A2(n9819), .ZN(n9377) );
  NAND2_X1 U9135 ( .A1(n9375), .A2(n9377), .ZN(n9315) );
  XNOR2_X1 U9136 ( .A(n7692), .B(n9315), .ZN(n9931) );
  INV_X1 U9137 ( .A(n4560), .ZN(n7557) );
  AOI211_X1 U9138 ( .C1(n9928), .C2(n7626), .A(n10205), .B(n7557), .ZN(n9927)
         );
  INV_X1 U9139 ( .A(n9928), .ZN(n7558) );
  NOR2_X1 U9140 ( .A1(n7558), .A2(n9799), .ZN(n7561) );
  OAI22_X1 U9141 ( .A1(n9810), .A2(n7559), .B1(n7649), .B2(n10150), .ZN(n7560)
         );
  AOI211_X1 U9142 ( .C1(n9927), .C2(n7714), .A(n7561), .B(n7560), .ZN(n7579)
         );
  AND2_X1 U9143 ( .A1(n9369), .A2(n7562), .ZN(n9270) );
  OAI21_X1 U9144 ( .B1(n7563), .B2(n9263), .A(n9270), .ZN(n7564) );
  NAND2_X1 U9145 ( .A1(n7564), .A2(n9363), .ZN(n7617) );
  OR2_X1 U9146 ( .A1(n9932), .A2(n7565), .ZN(n9275) );
  NAND2_X1 U9147 ( .A1(n9932), .A2(n7565), .ZN(n9367) );
  NAND2_X1 U9148 ( .A1(n7617), .A2(n9313), .ZN(n7566) );
  INV_X1 U9149 ( .A(n9315), .ZN(n7567) );
  OAI211_X1 U9150 ( .C1(n4555), .C2(n7567), .A(n7724), .B(n10135), .ZN(n7577)
         );
  NAND2_X1 U9151 ( .A1(n6431), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7575) );
  INV_X1 U9152 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7568) );
  OR2_X1 U9153 ( .A1(n4478), .A2(n7568), .ZN(n7574) );
  NAND2_X1 U9154 ( .A1(n7570), .A2(n7569), .ZN(n7571) );
  NAND2_X1 U9155 ( .A1(n7702), .A2(n7571), .ZN(n9827) );
  OR2_X1 U9156 ( .A1(n6527), .A2(n9827), .ZN(n7573) );
  INV_X1 U9157 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9828) );
  OR2_X1 U9158 ( .A1(n4476), .A2(n9828), .ZN(n7572) );
  NAND4_X1 U9159 ( .A1(n7575), .A2(n7574), .A3(n7573), .A4(n7572), .ZN(n9552)
         );
  AOI22_X1 U9160 ( .A1(n10137), .A2(n9554), .B1(n9552), .B2(n10140), .ZN(n7576) );
  NAND2_X1 U9161 ( .A1(n7577), .A2(n7576), .ZN(n9926) );
  NAND2_X1 U9162 ( .A1(n9926), .A2(n9810), .ZN(n7578) );
  OAI211_X1 U9163 ( .C1(n9931), .C2(n9813), .A(n7579), .B(n7578), .ZN(P1_U3277) );
  XNOR2_X1 U9164 ( .A(n7677), .B(n7676), .ZN(n10025) );
  INV_X1 U9165 ( .A(n10025), .ZN(n7595) );
  OAI211_X1 U9166 ( .C1(n7584), .C2(n7583), .A(n7582), .B(n10264), .ZN(n7586)
         );
  AOI22_X1 U9167 ( .A1(n10259), .A2(n8371), .B1(n8370), .B2(n10261), .ZN(n7585) );
  NAND2_X1 U9168 ( .A1(n7586), .A2(n7585), .ZN(n10024) );
  NAND2_X1 U9169 ( .A1(n7587), .A2(n10027), .ZN(n7588) );
  INV_X1 U9170 ( .A(n7588), .ZN(n7589) );
  INV_X1 U9171 ( .A(n7607), .ZN(n10021) );
  OR2_X1 U9172 ( .A1(n7588), .A2(n7607), .ZN(n8652) );
  OAI21_X1 U9173 ( .B1(n7589), .B2(n10021), .A(n8652), .ZN(n10022) );
  INV_X1 U9174 ( .A(n7590), .ZN(n7602) );
  OAI22_X1 U9175 ( .A1(n10299), .A2(n5457), .B1(n7602), .B2(n10297), .ZN(n7591) );
  AOI21_X1 U9176 ( .B1(n7607), .B2(n10302), .A(n7591), .ZN(n7592) );
  OAI21_X1 U9177 ( .B1(n10022), .B2(n10273), .A(n7592), .ZN(n7593) );
  AOI21_X1 U9178 ( .B1(n10024), .B2(n10299), .A(n7593), .ZN(n7594) );
  OAI21_X1 U9179 ( .B1(n7595), .B2(n8639), .A(n7594), .ZN(P2_U3281) );
  INV_X1 U9180 ( .A(n7596), .ZN(n7598) );
  NAND2_X1 U9181 ( .A1(n7598), .A2(n7597), .ZN(n7599) );
  XNOR2_X1 U9182 ( .A(n7607), .B(n8165), .ZN(n8268) );
  XNOR2_X1 U9183 ( .A(n8270), .B(n8268), .ZN(n7601) );
  AOI22_X1 U9184 ( .A1(n7601), .A2(n8336), .B1(n8313), .B2(n8648), .ZN(n7610)
         );
  AND2_X1 U9185 ( .A1(n8648), .A2(n8156), .ZN(n7658) );
  NAND2_X1 U9186 ( .A1(n7601), .A2(n7658), .ZN(n8269) );
  INV_X1 U9187 ( .A(n8269), .ZN(n7609) );
  OAI22_X1 U9188 ( .A1(n8355), .A2(n7602), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5452), .ZN(n7606) );
  OAI22_X1 U9189 ( .A1(n8357), .A2(n7604), .B1(n8356), .B2(n7603), .ZN(n7605)
         );
  AOI211_X1 U9190 ( .C1(n7607), .C2(n8360), .A(n7606), .B(n7605), .ZN(n7608)
         );
  OAI21_X1 U9191 ( .B1(n7610), .B2(n7609), .A(n7608), .ZN(P2_U3243) );
  INV_X1 U9192 ( .A(n7899), .ZN(n7612) );
  OAI222_X1 U9193 ( .A1(n7611), .A2(P2_U3152), .B1(n9134), .B2(n7612), .C1(
        n8899), .C2(n9137), .ZN(P2_U3334) );
  OAI222_X1 U9194 ( .A1(n7613), .A2(P1_U3084), .B1(n9971), .B2(n7612), .C1(
        n8783), .C2(n9968), .ZN(P1_U3329) );
  XNOR2_X1 U9195 ( .A(n7614), .B(n9313), .ZN(n7616) );
  INV_X1 U9196 ( .A(n7616), .ZN(n9935) );
  NAND2_X1 U9197 ( .A1(n7616), .A2(n7615), .ZN(n7623) );
  XNOR2_X1 U9198 ( .A(n7617), .B(n9313), .ZN(n7621) );
  NAND2_X1 U9199 ( .A1(n9553), .A2(n10140), .ZN(n7618) );
  OAI21_X1 U9200 ( .B1(n7619), .B2(n9818), .A(n7618), .ZN(n7620) );
  AOI21_X1 U9201 ( .B1(n7621), .B2(n10135), .A(n7620), .ZN(n7622) );
  NAND2_X1 U9202 ( .A1(n7623), .A2(n7622), .ZN(n9937) );
  NAND2_X1 U9203 ( .A1(n9937), .A2(n9810), .ZN(n7632) );
  NAND2_X1 U9204 ( .A1(n7624), .A2(n9932), .ZN(n7625) );
  AND2_X1 U9205 ( .A1(n7626), .A2(n7625), .ZN(n9933) );
  OAI22_X1 U9206 ( .A1(n9810), .A2(n6405), .B1(n7627), .B2(n10150), .ZN(n7630)
         );
  INV_X1 U9207 ( .A(n9932), .ZN(n7628) );
  NOR2_X1 U9208 ( .A1(n7628), .A2(n9799), .ZN(n7629) );
  AOI211_X1 U9209 ( .C1(n9933), .C2(n9733), .A(n7630), .B(n7629), .ZN(n7631)
         );
  OAI211_X1 U9210 ( .C1(n9935), .C2(n7633), .A(n7632), .B(n7631), .ZN(P1_U3278) );
  AND2_X1 U9211 ( .A1(n7636), .A2(n7637), .ZN(n7634) );
  INV_X1 U9212 ( .A(n7636), .ZN(n7639) );
  INV_X1 U9213 ( .A(n7637), .ZN(n7638) );
  NAND2_X1 U9214 ( .A1(n7639), .A2(n7638), .ZN(n7640) );
  NAND2_X1 U9215 ( .A1(n9928), .A2(n8044), .ZN(n7642) );
  NAND2_X1 U9216 ( .A1(n9553), .A2(n7347), .ZN(n7641) );
  NAND2_X1 U9217 ( .A1(n7642), .A2(n7641), .ZN(n7643) );
  XNOR2_X1 U9218 ( .A(n7643), .B(n8047), .ZN(n7746) );
  AND2_X1 U9219 ( .A1(n9553), .A2(n7928), .ZN(n7644) );
  AOI21_X1 U9220 ( .B1(n9928), .B2(n7347), .A(n7644), .ZN(n7742) );
  INV_X1 U9221 ( .A(n7742), .ZN(n7747) );
  XNOR2_X1 U9222 ( .A(n7746), .B(n7747), .ZN(n7645) );
  XNOR2_X1 U9223 ( .A(n7760), .B(n7645), .ZN(n7652) );
  INV_X1 U9224 ( .A(n9552), .ZN(n7727) );
  NOR2_X1 U9225 ( .A1(n7727), .A2(n9234), .ZN(n7646) );
  AOI211_X1 U9226 ( .C1(n9236), .C2(n9554), .A(n7647), .B(n7646), .ZN(n7648)
         );
  OAI21_X1 U9227 ( .B1(n9249), .B2(n7649), .A(n7648), .ZN(n7650) );
  AOI21_X1 U9228 ( .B1(n9928), .B2(n9251), .A(n7650), .ZN(n7651) );
  OAI21_X1 U9229 ( .B1(n7652), .B2(n9253), .A(n7651), .ZN(P1_U3213) );
  XNOR2_X1 U9230 ( .A(n8110), .B(n8165), .ZN(n7653) );
  AND2_X1 U9231 ( .A1(n8647), .A2(n4486), .ZN(n7654) );
  NAND2_X1 U9232 ( .A1(n7653), .A2(n7654), .ZN(n8130) );
  INV_X1 U9233 ( .A(n7653), .ZN(n8326) );
  INV_X1 U9234 ( .A(n7654), .ZN(n7655) );
  NAND2_X1 U9235 ( .A1(n8326), .A2(n7655), .ZN(n7656) );
  AND2_X1 U9236 ( .A1(n8130), .A2(n7656), .ZN(n7665) );
  XNOR2_X1 U9237 ( .A(n10015), .B(n8165), .ZN(n8273) );
  AND2_X1 U9238 ( .A1(n8370), .A2(n8156), .ZN(n7660) );
  OAI22_X1 U9239 ( .A1(n8273), .A2(n7660), .B1(n8268), .B2(n7658), .ZN(n7657)
         );
  NAND2_X1 U9240 ( .A1(n8268), .A2(n7658), .ZN(n7659) );
  INV_X1 U9241 ( .A(n7660), .ZN(n8272) );
  NAND2_X1 U9242 ( .A1(n7659), .A2(n8272), .ZN(n7662) );
  INV_X1 U9243 ( .A(n7659), .ZN(n7661) );
  AOI22_X1 U9244 ( .A1(n8273), .A2(n7662), .B1(n7661), .B2(n7660), .ZN(n7663)
         );
  NAND2_X1 U9245 ( .A1(n7664), .A2(n7665), .ZN(n8325) );
  OAI211_X1 U9246 ( .C1(n7665), .C2(n7664), .A(n8325), .B(n8336), .ZN(n7671)
         );
  NAND2_X1 U9247 ( .A1(n8369), .A2(n10261), .ZN(n7667) );
  NAND2_X1 U9248 ( .A1(n8370), .A2(n10259), .ZN(n7666) );
  AND2_X1 U9249 ( .A1(n7667), .A2(n7666), .ZN(n7683) );
  OAI22_X1 U9250 ( .A1(n8263), .A2(n7683), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7668), .ZN(n7669) );
  AOI21_X1 U9251 ( .B1(n7686), .B2(n8342), .A(n7669), .ZN(n7670) );
  OAI211_X1 U9252 ( .C1(n10011), .C2(n8338), .A(n7671), .B(n7670), .ZN(
        P2_U3230) );
  INV_X1 U9253 ( .A(n7914), .ZN(n7675) );
  OAI222_X1 U9254 ( .A1(n9137), .A2(n7673), .B1(n9134), .B2(n7675), .C1(n7672), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9255 ( .A1(n9968), .A2(n7915), .B1(n9971), .B2(n7675), .C1(n7674), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI21_X1 U9256 ( .B1(n7679), .B2(n7678), .A(n8109), .ZN(n10014) );
  INV_X1 U9257 ( .A(n10014), .ZN(n7691) );
  NAND2_X1 U9258 ( .A1(n7680), .A2(n10264), .ZN(n7685) );
  AOI21_X1 U9259 ( .B1(n8640), .B2(n7682), .A(n7681), .ZN(n7684) );
  OAI21_X1 U9260 ( .B1(n7685), .B2(n7684), .A(n7683), .ZN(n10013) );
  OAI211_X1 U9261 ( .C1(n8654), .C2(n10011), .A(n8624), .B(n10295), .ZN(n10010) );
  AOI22_X1 U9262 ( .A1(n10308), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n7686), .B2(
        n10245), .ZN(n7688) );
  NAND2_X1 U9263 ( .A1(n8110), .A2(n10302), .ZN(n7687) );
  OAI211_X1 U9264 ( .C1(n10010), .C2(n10304), .A(n7688), .B(n7687), .ZN(n7689)
         );
  AOI21_X1 U9265 ( .B1(n10013), .B2(n10299), .A(n7689), .ZN(n7690) );
  OAI21_X1 U9266 ( .B1(n7691), .B2(n8639), .A(n7690), .ZN(P2_U3279) );
  OR2_X1 U9267 ( .A1(n9928), .A2(n9553), .ZN(n7693) );
  NAND2_X1 U9268 ( .A1(n7694), .A2(n6907), .ZN(n7696) );
  AOI22_X1 U9269 ( .A1(n7803), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10117), 
        .B2(n7802), .ZN(n7695) );
  NAND2_X1 U9270 ( .A1(n7697), .A2(n6907), .ZN(n7700) );
  AOI22_X1 U9271 ( .A1(n7803), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7698), .B2(
        n7802), .ZN(n7699) );
  NAND2_X1 U9272 ( .A1(n6431), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7708) );
  OR2_X1 U9273 ( .A1(n4476), .A2(n7068), .ZN(n7707) );
  INV_X1 U9274 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7701) );
  NAND2_X1 U9275 ( .A1(n7702), .A2(n7701), .ZN(n7703) );
  NAND2_X1 U9276 ( .A1(n7719), .A2(n7703), .ZN(n9184) );
  OR2_X1 U9277 ( .A1(n6527), .A2(n9184), .ZN(n7706) );
  OR2_X1 U9278 ( .A1(n4478), .A2(n7704), .ZN(n7705) );
  OR2_X1 U9279 ( .A1(n9916), .A2(n9817), .ZN(n9388) );
  NAND2_X1 U9280 ( .A1(n9916), .A2(n9817), .ZN(n9387) );
  OAI21_X1 U9281 ( .B1(n7710), .B2(n7709), .A(n7968), .ZN(n9918) );
  INV_X1 U9282 ( .A(n9825), .ZN(n7711) );
  INV_X1 U9283 ( .A(n9916), .ZN(n9189) );
  AOI211_X1 U9284 ( .C1(n9916), .C2(n7711), .A(n10205), .B(n9797), .ZN(n9915)
         );
  NOR2_X1 U9285 ( .A1(n9189), .A2(n9799), .ZN(n7713) );
  OAI22_X1 U9286 ( .A1(n9810), .A2(n7068), .B1(n9184), .B2(n10150), .ZN(n7712)
         );
  AOI211_X1 U9287 ( .C1(n9915), .C2(n7714), .A(n7713), .B(n7712), .ZN(n7729)
         );
  INV_X1 U9288 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7715) );
  OR2_X1 U9289 ( .A1(n6557), .A2(n7715), .ZN(n7716) );
  OAI21_X1 U9290 ( .B1(n4479), .B2(n7717), .A(n7716), .ZN(n7723) );
  NAND2_X1 U9291 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  NAND2_X1 U9292 ( .A1(n7786), .A2(n7720), .ZN(n9801) );
  NOR2_X1 U9293 ( .A1(n6527), .A2(n9801), .ZN(n7722) );
  NOR2_X1 U9294 ( .A1(n4477), .A2(n7211), .ZN(n7721) );
  OR2_X1 U9295 ( .A1(n9919), .A2(n7727), .ZN(n9382) );
  NAND2_X1 U9296 ( .A1(n9919), .A2(n7727), .ZN(n9383) );
  NAND2_X1 U9297 ( .A1(n9382), .A2(n9383), .ZN(n9814) );
  NAND2_X1 U9298 ( .A1(n7725), .A2(n9383), .ZN(n7986) );
  XOR2_X1 U9299 ( .A(n9385), .B(n7986), .Z(n7726) );
  OAI222_X1 U9300 ( .A1(n9816), .A2(n9784), .B1(n9818), .B2(n7727), .C1(n7726), 
        .C2(n9807), .ZN(n9914) );
  NAND2_X1 U9301 ( .A1(n9914), .A2(n9810), .ZN(n7728) );
  OAI211_X1 U9302 ( .C1(n9918), .C2(n9813), .A(n7729), .B(n7728), .ZN(P1_U3275) );
  NAND2_X1 U9303 ( .A1(n9136), .A2(n6907), .ZN(n7731) );
  OR2_X1 U9304 ( .A1(n8094), .A2(n9969), .ZN(n7730) );
  OR2_X1 U9305 ( .A1(n9649), .A2(n7945), .ZN(n7740) );
  NAND2_X1 U9306 ( .A1(n7921), .A2(n8938), .ZN(n7732) );
  NAND2_X1 U9307 ( .A1(n9647), .A2(n6213), .ZN(n7738) );
  INV_X1 U9308 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U9309 ( .A1(n7887), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7735) );
  INV_X1 U9310 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n7733) );
  OR2_X1 U9311 ( .A1(n4477), .A2(n7733), .ZN(n7734) );
  OAI211_X1 U9312 ( .C1(n6557), .C2(n8879), .A(n7735), .B(n7734), .ZN(n7736)
         );
  INV_X1 U9313 ( .A(n7736), .ZN(n7737) );
  NAND2_X1 U9314 ( .A1(n9546), .A2(n7928), .ZN(n7739) );
  NAND2_X1 U9315 ( .A1(n7740), .A2(n7739), .ZN(n7936) );
  OAI22_X1 U9316 ( .A1(n9649), .A2(n7946), .B1(n9671), .B2(n7945), .ZN(n7741)
         );
  XNOR2_X1 U9317 ( .A(n7741), .B(n7947), .ZN(n7935) );
  NAND2_X1 U9318 ( .A1(n7746), .A2(n7742), .ZN(n7764) );
  NAND2_X1 U9319 ( .A1(n7760), .A2(n7764), .ZN(n7750) );
  NAND2_X1 U9320 ( .A1(n9919), .A2(n8044), .ZN(n7744) );
  NAND2_X1 U9321 ( .A1(n9552), .A2(n7347), .ZN(n7743) );
  NAND2_X1 U9322 ( .A1(n7744), .A2(n7743), .ZN(n7745) );
  XNOR2_X1 U9323 ( .A(n7745), .B(n8047), .ZN(n7763) );
  INV_X1 U9324 ( .A(n7746), .ZN(n7748) );
  NAND2_X1 U9325 ( .A1(n7748), .A2(n7747), .ZN(n7761) );
  AND2_X1 U9326 ( .A1(n7763), .A2(n7761), .ZN(n7749) );
  NAND2_X1 U9327 ( .A1(n7750), .A2(n7749), .ZN(n9241) );
  NAND2_X1 U9328 ( .A1(n9919), .A2(n7347), .ZN(n7752) );
  NAND2_X1 U9329 ( .A1(n9552), .A2(n7928), .ZN(n7751) );
  NAND2_X1 U9330 ( .A1(n7752), .A2(n7751), .ZN(n9244) );
  NAND2_X1 U9331 ( .A1(n9241), .A2(n9244), .ZN(n9180) );
  NAND2_X1 U9332 ( .A1(n9916), .A2(n8044), .ZN(n7754) );
  OR2_X1 U9333 ( .A1(n9817), .A2(n7945), .ZN(n7753) );
  NAND2_X1 U9334 ( .A1(n7754), .A2(n7753), .ZN(n7755) );
  XNOR2_X1 U9335 ( .A(n7755), .B(n8047), .ZN(n7758) );
  NOR2_X1 U9336 ( .A1(n9817), .A2(n7943), .ZN(n7756) );
  AOI21_X1 U9337 ( .B1(n9916), .B2(n7347), .A(n7756), .ZN(n7757) );
  NAND2_X1 U9338 ( .A1(n7758), .A2(n7757), .ZN(n7768) );
  OR2_X1 U9339 ( .A1(n7758), .A2(n7757), .ZN(n7759) );
  AND2_X1 U9340 ( .A1(n7768), .A2(n7759), .ZN(n9179) );
  INV_X1 U9341 ( .A(n7760), .ZN(n7762) );
  NAND2_X1 U9342 ( .A1(n7762), .A2(n7761), .ZN(n7767) );
  INV_X1 U9343 ( .A(n7763), .ZN(n7765) );
  AND2_X1 U9344 ( .A1(n7765), .A2(n7764), .ZN(n7766) );
  NAND2_X1 U9345 ( .A1(n7769), .A2(n6907), .ZN(n7772) );
  AOI22_X1 U9346 ( .A1(n7770), .A2(n7802), .B1(n7803), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U9347 ( .A1(n9911), .A2(n8044), .ZN(n7774) );
  NAND2_X1 U9348 ( .A1(n9550), .A2(n7347), .ZN(n7773) );
  NAND2_X1 U9349 ( .A1(n7774), .A2(n7773), .ZN(n7775) );
  XNOR2_X1 U9350 ( .A(n7775), .B(n7947), .ZN(n7777) );
  AND2_X1 U9351 ( .A1(n9550), .A2(n7928), .ZN(n7776) );
  AOI21_X1 U9352 ( .B1(n9911), .B2(n7347), .A(n7776), .ZN(n7778) );
  XNOR2_X1 U9353 ( .A(n7777), .B(n7778), .ZN(n9192) );
  INV_X1 U9354 ( .A(n7777), .ZN(n7779) );
  NAND2_X1 U9355 ( .A1(n7779), .A2(n7778), .ZN(n7780) );
  NAND2_X1 U9356 ( .A1(n7781), .A2(n6907), .ZN(n7784) );
  AOI22_X1 U9357 ( .A1(n7782), .A2(n7802), .B1(n7803), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n7783) );
  NAND2_X1 U9358 ( .A1(n9906), .A2(n8044), .ZN(n7793) );
  NAND2_X1 U9359 ( .A1(n6431), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7791) );
  OR2_X1 U9360 ( .A1(n4479), .A2(n9583), .ZN(n7790) );
  INV_X1 U9361 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U9362 ( .A1(n7786), .A2(n7785), .ZN(n7787) );
  NAND2_X1 U9363 ( .A1(n7807), .A2(n7787), .ZN(n9788) );
  OR2_X1 U9364 ( .A1(n6527), .A2(n9788), .ZN(n7789) );
  INV_X1 U9365 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9588) );
  OR2_X1 U9366 ( .A1(n4477), .A2(n9588), .ZN(n7788) );
  OR2_X1 U9367 ( .A1(n9809), .A2(n7945), .ZN(n7792) );
  NAND2_X1 U9368 ( .A1(n7793), .A2(n7792), .ZN(n7794) );
  XNOR2_X1 U9369 ( .A(n7794), .B(n8047), .ZN(n7798) );
  NAND2_X1 U9370 ( .A1(n7797), .A2(n7798), .ZN(n9229) );
  NAND2_X1 U9371 ( .A1(n9906), .A2(n7347), .ZN(n7796) );
  OR2_X1 U9372 ( .A1(n9809), .A2(n7943), .ZN(n7795) );
  NAND2_X1 U9373 ( .A1(n7796), .A2(n7795), .ZN(n9232) );
  INV_X1 U9374 ( .A(n7798), .ZN(n7799) );
  NAND2_X1 U9375 ( .A1(n7801), .A2(n6907), .ZN(n7805) );
  AOI22_X1 U9376 ( .A1(n7803), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10148), 
        .B2(n7802), .ZN(n7804) );
  NAND2_X1 U9377 ( .A1(n9900), .A2(n8044), .ZN(n7815) );
  NAND2_X1 U9378 ( .A1(n6431), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7813) );
  INV_X1 U9379 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U9380 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND2_X1 U9381 ( .A1(n7827), .A2(n7808), .ZN(n9766) );
  OR2_X1 U9382 ( .A1(n9766), .A2(n6527), .ZN(n7812) );
  INV_X1 U9383 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7809) );
  OR2_X1 U9384 ( .A1(n4476), .A2(n7809), .ZN(n7811) );
  INV_X1 U9385 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9584) );
  OR2_X1 U9386 ( .A1(n4479), .A2(n9584), .ZN(n7810) );
  NAND4_X1 U9387 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n9549)
         );
  NAND2_X1 U9388 ( .A1(n9549), .A2(n7347), .ZN(n7814) );
  NAND2_X1 U9389 ( .A1(n7815), .A2(n7814), .ZN(n7816) );
  XNOR2_X1 U9390 ( .A(n7816), .B(n7947), .ZN(n7819) );
  NAND2_X1 U9391 ( .A1(n9900), .A2(n4480), .ZN(n7818) );
  NAND2_X1 U9392 ( .A1(n9549), .A2(n7928), .ZN(n7817) );
  NAND2_X1 U9393 ( .A1(n7818), .A2(n7817), .ZN(n7820) );
  AND2_X1 U9394 ( .A1(n7819), .A2(n7820), .ZN(n9155) );
  INV_X1 U9395 ( .A(n7819), .ZN(n7822) );
  INV_X1 U9396 ( .A(n7820), .ZN(n7821) );
  NAND2_X1 U9397 ( .A1(n7822), .A2(n7821), .ZN(n9153) );
  NAND2_X1 U9398 ( .A1(n7823), .A2(n6907), .ZN(n7826) );
  OR2_X1 U9399 ( .A1(n8094), .A2(n7824), .ZN(n7825) );
  NAND2_X1 U9400 ( .A1(n9896), .A2(n8044), .ZN(n7835) );
  INV_X1 U9401 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U9402 ( .A1(n7827), .A2(n9213), .ZN(n7828) );
  NAND2_X1 U9403 ( .A1(n7847), .A2(n7828), .ZN(n9753) );
  OR2_X1 U9404 ( .A1(n9753), .A2(n6527), .ZN(n7833) );
  INV_X1 U9405 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n7829) );
  OR2_X1 U9406 ( .A1(n6557), .A2(n7829), .ZN(n7831) );
  INV_X1 U9407 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8903) );
  OR2_X1 U9408 ( .A1(n4478), .A2(n8903), .ZN(n7830) );
  AND2_X1 U9409 ( .A1(n7831), .A2(n7830), .ZN(n7832) );
  OAI211_X1 U9410 ( .C1(n4477), .C2(n9754), .A(n7833), .B(n7832), .ZN(n9773)
         );
  NAND2_X1 U9411 ( .A1(n9773), .A2(n7347), .ZN(n7834) );
  NAND2_X1 U9412 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  XNOR2_X1 U9413 ( .A(n7836), .B(n7947), .ZN(n7838) );
  AND2_X1 U9414 ( .A1(n9773), .A2(n7928), .ZN(n7837) );
  AOI21_X1 U9415 ( .B1(n9896), .B2(n7347), .A(n7837), .ZN(n7839) );
  XNOR2_X1 U9416 ( .A(n7838), .B(n7839), .ZN(n9210) );
  INV_X1 U9417 ( .A(n7838), .ZN(n7840) );
  NAND2_X1 U9418 ( .A1(n7840), .A2(n7839), .ZN(n7841) );
  NAND2_X1 U9419 ( .A1(n7842), .A2(n6907), .ZN(n7845) );
  OR2_X1 U9420 ( .A1(n6506), .A2(n7843), .ZN(n7844) );
  NAND2_X1 U9421 ( .A1(n9889), .A2(n8044), .ZN(n7853) );
  NAND2_X1 U9422 ( .A1(n7847), .A2(n7846), .ZN(n7848) );
  AND2_X1 U9423 ( .A1(n7864), .A2(n7848), .ZN(n9742) );
  NAND2_X1 U9424 ( .A1(n9742), .A2(n6213), .ZN(n7851) );
  AOI22_X1 U9425 ( .A1(n6431), .A2(P1_REG0_REG_21__SCAN_IN), .B1(n7992), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U9426 ( .A1(n7887), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U9427 ( .A1(n9728), .A2(n7347), .ZN(n7852) );
  NAND2_X1 U9428 ( .A1(n7853), .A2(n7852), .ZN(n7854) );
  XNOR2_X1 U9429 ( .A(n7854), .B(n7947), .ZN(n7856) );
  NOR2_X1 U9430 ( .A1(n9760), .A2(n7943), .ZN(n7855) );
  AOI21_X1 U9431 ( .B1(n9889), .B2(n4480), .A(n7855), .ZN(n7857) );
  XNOR2_X1 U9432 ( .A(n7856), .B(n7857), .ZN(n9164) );
  INV_X1 U9433 ( .A(n7856), .ZN(n7858) );
  NAND2_X1 U9434 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U9435 ( .A1(n7860), .A2(n6907), .ZN(n7863) );
  OR2_X1 U9436 ( .A1(n8094), .A2(n7861), .ZN(n7862) );
  NAND2_X2 U9437 ( .A1(n7863), .A2(n7862), .ZN(n9883) );
  INV_X1 U9438 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U9439 ( .A1(n7864), .A2(n9223), .ZN(n7865) );
  NAND2_X1 U9440 ( .A1(n7885), .A2(n7865), .ZN(n9721) );
  OR2_X1 U9441 ( .A1(n9721), .A2(n6527), .ZN(n7871) );
  INV_X1 U9442 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U9443 ( .A1(n7992), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U9444 ( .A1(n6431), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7866) );
  OAI211_X1 U9445 ( .C1(n4478), .C2(n7868), .A(n7867), .B(n7866), .ZN(n7869)
         );
  INV_X1 U9446 ( .A(n7869), .ZN(n7870) );
  NAND2_X1 U9447 ( .A1(n7871), .A2(n7870), .ZN(n9738) );
  AND2_X1 U9448 ( .A1(n9738), .A2(n7928), .ZN(n7872) );
  AOI21_X1 U9449 ( .B1(n9883), .B2(n7347), .A(n7872), .ZN(n7877) );
  INV_X1 U9450 ( .A(n7877), .ZN(n7873) );
  NAND2_X1 U9451 ( .A1(n9883), .A2(n8044), .ZN(n7875) );
  NAND2_X1 U9452 ( .A1(n9738), .A2(n4480), .ZN(n7874) );
  NAND2_X1 U9453 ( .A1(n7875), .A2(n7874), .ZN(n7876) );
  XNOR2_X1 U9454 ( .A(n7876), .B(n8047), .ZN(n9221) );
  NAND2_X1 U9455 ( .A1(n9220), .A2(n9221), .ZN(n7879) );
  NAND2_X1 U9456 ( .A1(n7878), .A2(n7877), .ZN(n9219) );
  NAND2_X1 U9457 ( .A1(n7880), .A2(n6907), .ZN(n7883) );
  OR2_X1 U9458 ( .A1(n8094), .A2(n7881), .ZN(n7882) );
  NAND2_X1 U9459 ( .A1(n9878), .A2(n8044), .ZN(n7895) );
  INV_X1 U9460 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U9461 ( .A1(n7885), .A2(n7884), .ZN(n7886) );
  NAND2_X1 U9462 ( .A1(n7901), .A2(n7886), .ZN(n9703) );
  OR2_X1 U9463 ( .A1(n9703), .A2(n6527), .ZN(n7893) );
  INV_X1 U9464 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U9465 ( .A1(n7887), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U9466 ( .A1(n7992), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7888) );
  OAI211_X1 U9467 ( .C1(n6557), .C2(n7890), .A(n7889), .B(n7888), .ZN(n7891)
         );
  INV_X1 U9468 ( .A(n7891), .ZN(n7892) );
  NAND2_X1 U9469 ( .A1(n7893), .A2(n7892), .ZN(n9729) );
  NAND2_X1 U9470 ( .A1(n9729), .A2(n7347), .ZN(n7894) );
  NAND2_X1 U9471 ( .A1(n7895), .A2(n7894), .ZN(n7896) );
  XNOR2_X1 U9472 ( .A(n7896), .B(n8047), .ZN(n7897) );
  INV_X1 U9473 ( .A(n9878), .ZN(n9706) );
  OAI22_X1 U9474 ( .A1(n9706), .A2(n7945), .B1(n9688), .B2(n7943), .ZN(n9146)
         );
  NAND2_X1 U9475 ( .A1(n7898), .A2(n7897), .ZN(n9143) );
  OR2_X1 U9476 ( .A1(n6506), .A2(n8783), .ZN(n7900) );
  NAND2_X1 U9477 ( .A1(n9875), .A2(n8044), .ZN(n7909) );
  NAND2_X1 U9478 ( .A1(n7901), .A2(n9201), .ZN(n7902) );
  AND2_X1 U9479 ( .A1(n7919), .A2(n7902), .ZN(n9682) );
  INV_X1 U9480 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U9481 ( .A1(n7992), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7905) );
  INV_X1 U9482 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n7903) );
  OR2_X1 U9483 ( .A1(n6557), .A2(n7903), .ZN(n7904) );
  OAI211_X1 U9484 ( .C1(n4479), .C2(n7906), .A(n7905), .B(n7904), .ZN(n7907)
         );
  AOI21_X1 U9485 ( .B1(n9682), .B2(n6213), .A(n7907), .ZN(n9710) );
  OR2_X1 U9486 ( .A1(n9710), .A2(n7945), .ZN(n7908) );
  NAND2_X1 U9487 ( .A1(n7909), .A2(n7908), .ZN(n7910) );
  XNOR2_X1 U9488 ( .A(n7910), .B(n7947), .ZN(n7911) );
  INV_X1 U9489 ( .A(n9710), .ZN(n9548) );
  AOI22_X1 U9490 ( .A1(n9875), .A2(n7347), .B1(n7928), .B2(n9548), .ZN(n7912)
         );
  XNOR2_X1 U9491 ( .A(n7911), .B(n7912), .ZN(n9200) );
  INV_X1 U9492 ( .A(n7911), .ZN(n7913) );
  NAND2_X1 U9493 ( .A1(n7914), .A2(n6907), .ZN(n7917) );
  OR2_X1 U9494 ( .A1(n6506), .A2(n7915), .ZN(n7916) );
  INV_X1 U9495 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U9496 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  NAND2_X1 U9497 ( .A1(n7921), .A2(n7920), .ZN(n9676) );
  OR2_X1 U9498 ( .A1(n9676), .A2(n6527), .ZN(n7927) );
  INV_X1 U9499 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U9500 ( .A1(n6431), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U9501 ( .A1(n7992), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7922) );
  OAI211_X1 U9502 ( .C1(n4479), .C2(n7924), .A(n7923), .B(n7922), .ZN(n7925)
         );
  INV_X1 U9503 ( .A(n7925), .ZN(n7926) );
  AOI22_X1 U9504 ( .A1(n9667), .A2(n4480), .B1(n7928), .B2(n9547), .ZN(n7932)
         );
  NAND2_X1 U9505 ( .A1(n9667), .A2(n8044), .ZN(n7930) );
  NAND2_X1 U9506 ( .A1(n9547), .A2(n7347), .ZN(n7929) );
  NAND2_X1 U9507 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  XNOR2_X1 U9508 ( .A(n7931), .B(n7947), .ZN(n7934) );
  XOR2_X1 U9509 ( .A(n7932), .B(n7934), .Z(n9172) );
  INV_X1 U9510 ( .A(n7932), .ZN(n7933) );
  XNOR2_X1 U9511 ( .A(n7935), .B(n7936), .ZN(n8040) );
  NAND2_X1 U9512 ( .A1(n9132), .A2(n6907), .ZN(n7938) );
  OR2_X1 U9513 ( .A1(n8094), .A2(n9967), .ZN(n7937) );
  XNOR2_X1 U9514 ( .A(n7951), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9632) );
  INV_X1 U9515 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7941) );
  NAND2_X1 U9516 ( .A1(n7992), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7940) );
  NAND2_X1 U9517 ( .A1(n6431), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7939) );
  OAI211_X1 U9518 ( .C1(n4478), .C2(n7941), .A(n7940), .B(n7939), .ZN(n7942)
         );
  NOR2_X1 U9519 ( .A1(n9654), .A2(n7943), .ZN(n7944) );
  AOI21_X1 U9520 ( .B1(n9854), .B2(n7347), .A(n7944), .ZN(n8051) );
  INV_X1 U9521 ( .A(n9854), .ZN(n9634) );
  OAI22_X1 U9522 ( .A1(n9634), .A2(n7946), .B1(n9654), .B2(n7945), .ZN(n7948)
         );
  XNOR2_X1 U9523 ( .A(n7948), .B(n7947), .ZN(n8053) );
  XOR2_X1 U9524 ( .A(n8051), .B(n8053), .Z(n7949) );
  XNOR2_X1 U9525 ( .A(n8042), .B(n7949), .ZN(n7964) );
  INV_X1 U9526 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7959) );
  INV_X1 U9527 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7950) );
  OAI21_X1 U9528 ( .B1(n7951), .B2(n7959), .A(n7950), .ZN(n7952) );
  NAND2_X1 U9529 ( .A1(n7952), .A2(n7998), .ZN(n9620) );
  OR2_X1 U9530 ( .A1(n9620), .A2(n6527), .ZN(n7958) );
  INV_X1 U9531 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U9532 ( .A1(n7992), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7954) );
  NAND2_X1 U9533 ( .A1(n6431), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7953) );
  OAI211_X1 U9534 ( .C1(n4478), .C2(n7955), .A(n7954), .B(n7953), .ZN(n7956)
         );
  INV_X1 U9535 ( .A(n7956), .ZN(n7957) );
  OAI22_X1 U9536 ( .A1(n9671), .A2(n9245), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7959), .ZN(n7960) );
  AOI21_X1 U9537 ( .B1(n9632), .B2(n9203), .A(n7960), .ZN(n7961) );
  OAI21_X1 U9538 ( .B1(n9638), .B2(n9234), .A(n7961), .ZN(n7962) );
  AOI21_X1 U9539 ( .B1(n9854), .B2(n9251), .A(n7962), .ZN(n7963) );
  OAI21_X1 U9540 ( .B1(n7964), .B2(n9253), .A(n7963), .ZN(P1_U3212) );
  NAND2_X1 U9541 ( .A1(n8004), .A2(n6907), .ZN(n7966) );
  INV_X1 U9542 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8005) );
  OR2_X1 U9543 ( .A1(n8094), .A2(n8005), .ZN(n7965) );
  INV_X1 U9544 ( .A(n9849), .ZN(n9622) );
  AND2_X1 U9545 ( .A1(n9878), .A2(n9729), .ZN(n9691) );
  AND2_X1 U9546 ( .A1(n9875), .A2(n9548), .ZN(n7981) );
  OR2_X1 U9547 ( .A1(n9691), .A2(n7981), .ZN(n9661) );
  NAND2_X1 U9548 ( .A1(n9667), .A2(n9687), .ZN(n9433) );
  NAND2_X1 U9549 ( .A1(n9434), .A2(n9433), .ZN(n9665) );
  OR2_X1 U9550 ( .A1(n9661), .A2(n9668), .ZN(n7979) );
  INV_X1 U9551 ( .A(n9817), .ZN(n9551) );
  NAND2_X1 U9552 ( .A1(n9916), .A2(n9551), .ZN(n7967) );
  NAND2_X1 U9553 ( .A1(n7968), .A2(n7967), .ZN(n9796) );
  OR2_X1 U9554 ( .A1(n9911), .A2(n9550), .ZN(n7969) );
  NAND2_X1 U9555 ( .A1(n9796), .A2(n7969), .ZN(n7971) );
  NAND2_X1 U9556 ( .A1(n9911), .A2(n9550), .ZN(n7970) );
  NAND2_X1 U9557 ( .A1(n7971), .A2(n7970), .ZN(n9779) );
  OR2_X1 U9558 ( .A1(n9906), .A2(n9809), .ZN(n9401) );
  NAND2_X1 U9559 ( .A1(n9906), .A2(n9809), .ZN(n9397) );
  NAND2_X1 U9560 ( .A1(n9401), .A2(n9397), .ZN(n9781) );
  INV_X1 U9561 ( .A(n9809), .ZN(n9774) );
  NAND2_X1 U9562 ( .A1(n9906), .A2(n9774), .ZN(n7972) );
  OR2_X1 U9563 ( .A1(n9900), .A2(n9549), .ZN(n7973) );
  AND2_X1 U9564 ( .A1(n9896), .A2(n9773), .ZN(n7974) );
  OAI22_X1 U9565 ( .A1(n9750), .A2(n7974), .B1(n9773), .B2(n9896), .ZN(n9745)
         );
  INV_X1 U9566 ( .A(n9745), .ZN(n7976) );
  OR2_X1 U9567 ( .A1(n9889), .A2(n9760), .ZN(n9416) );
  NAND2_X1 U9568 ( .A1(n9889), .A2(n9760), .ZN(n9725) );
  NAND2_X1 U9569 ( .A1(n9889), .A2(n9728), .ZN(n7977) );
  OR2_X1 U9570 ( .A1(n9883), .A2(n9738), .ZN(n7978) );
  NOR2_X1 U9571 ( .A1(n7979), .A2(n9700), .ZN(n7983) );
  NAND2_X1 U9572 ( .A1(n9875), .A2(n9710), .ZN(n9426) );
  INV_X1 U9573 ( .A(n9695), .ZN(n7980) );
  OR2_X1 U9574 ( .A1(n9878), .A2(n9729), .ZN(n9693) );
  NAND2_X1 U9575 ( .A1(n9854), .A2(n9654), .ZN(n9442) );
  NAND2_X1 U9576 ( .A1(n9849), .A2(n9638), .ZN(n9451) );
  NAND2_X1 U9577 ( .A1(n9125), .A2(n6907), .ZN(n7985) );
  OR2_X1 U9578 ( .A1(n8094), .A2(n9965), .ZN(n7984) );
  NAND2_X1 U9579 ( .A1(n9844), .A2(n9616), .ZN(n9521) );
  NAND2_X1 U9580 ( .A1(n7986), .A2(n9388), .ZN(n7987) );
  OR2_X1 U9581 ( .A1(n9911), .A2(n9784), .ZN(n9260) );
  NAND2_X1 U9582 ( .A1(n9911), .A2(n9784), .ZN(n9262) );
  NAND2_X1 U9583 ( .A1(n9260), .A2(n9262), .ZN(n9805) );
  OR2_X1 U9584 ( .A1(n9900), .A2(n9783), .ZN(n9400) );
  NAND2_X1 U9585 ( .A1(n9900), .A2(n9783), .ZN(n9404) );
  NAND2_X1 U9586 ( .A1(n9771), .A2(n9772), .ZN(n9770) );
  INV_X1 U9587 ( .A(n9773), .ZN(n9159) );
  NAND2_X1 U9588 ( .A1(n9896), .A2(n9159), .ZN(n9403) );
  NAND2_X1 U9589 ( .A1(n9415), .A2(n9403), .ZN(n9757) );
  INV_X1 U9590 ( .A(n9738), .ZN(n9709) );
  NAND2_X1 U9591 ( .A1(n9883), .A2(n9709), .ZN(n9296) );
  AND2_X1 U9592 ( .A1(n9296), .A2(n9725), .ZN(n9421) );
  NAND2_X1 U9593 ( .A1(n7988), .A2(n9418), .ZN(n9707) );
  NAND2_X1 U9594 ( .A1(n9878), .A2(n9688), .ZN(n9507) );
  AND2_X1 U9595 ( .A1(n9424), .A2(n9684), .ZN(n9511) );
  INV_X1 U9596 ( .A(n9433), .ZN(n7989) );
  NAND2_X1 U9597 ( .A1(n7990), .A2(n9434), .ZN(n9650) );
  NAND2_X1 U9598 ( .A1(n9859), .A2(n9671), .ZN(n9441) );
  NAND2_X1 U9599 ( .A1(n9656), .A2(n9440), .ZN(n9635) );
  XNOR2_X1 U9600 ( .A(n7991), .B(n9456), .ZN(n7997) );
  INV_X1 U9601 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U9602 ( .A1(n6431), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U9603 ( .A1(n7992), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7993) );
  OAI211_X1 U9604 ( .C1(n4479), .C2(n8901), .A(n7994), .B(n7993), .ZN(n9544)
         );
  NAND2_X1 U9605 ( .A1(n7995), .A2(P1_B_REG_SCAN_IN), .ZN(n7996) );
  AND2_X1 U9606 ( .A1(n10140), .A2(n7996), .ZN(n8103) );
  OAI21_X1 U9607 ( .B1(n7998), .B2(n10150), .A(n9847), .ZN(n8002) );
  INV_X1 U9608 ( .A(n9667), .ZN(n9866) );
  INV_X1 U9609 ( .A(n9883), .ZN(n9724) );
  INV_X1 U9610 ( .A(n9889), .ZN(n9736) );
  INV_X1 U9611 ( .A(n9906), .ZN(n9793) );
  INV_X1 U9612 ( .A(n9911), .ZN(n9800) );
  NAND2_X1 U9613 ( .A1(n9793), .A2(n9798), .ZN(n9785) );
  NAND2_X1 U9614 ( .A1(n9866), .A2(n9681), .ZN(n9675) );
  NAND2_X1 U9615 ( .A1(n9622), .A2(n9631), .ZN(n9623) );
  NOR2_X2 U9616 ( .A1(n9623), .A2(n9844), .ZN(n9606) );
  AOI21_X1 U9617 ( .B1(n9844), .B2(n9623), .A(n9606), .ZN(n9845) );
  INV_X1 U9618 ( .A(n9845), .ZN(n8000) );
  AOI22_X1 U9619 ( .A1(n9844), .A2(n9830), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10157), .ZN(n7999) );
  OAI21_X1 U9620 ( .B1(n8000), .B2(n9832), .A(n7999), .ZN(n8001) );
  AOI21_X1 U9621 ( .B1(n8002), .B2(n9810), .A(n8001), .ZN(n8003) );
  OAI21_X1 U9622 ( .B1(n9848), .B2(n9813), .A(n8003), .ZN(P1_U3355) );
  INV_X1 U9623 ( .A(n8004), .ZN(n9131) );
  OAI222_X1 U9624 ( .A1(n9968), .A2(n8005), .B1(P1_U3084), .B2(n5956), .C1(
        n9971), .C2(n9131), .ZN(P1_U3325) );
  INV_X1 U9625 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10469) );
  NOR2_X1 U9626 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8006) );
  AOI21_X1 U9627 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n8006), .ZN(n10439) );
  NOR2_X1 U9628 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8007) );
  AOI21_X1 U9629 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n8007), .ZN(n10442) );
  NOR2_X1 U9630 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8008) );
  AOI21_X1 U9631 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n8008), .ZN(n10445) );
  NOR2_X1 U9632 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8009) );
  AOI21_X1 U9633 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n8009), .ZN(n10448) );
  NOR2_X1 U9634 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8010) );
  AOI21_X1 U9635 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n8010), .ZN(n10451) );
  NOR2_X1 U9636 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8017) );
  XNOR2_X1 U9637 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10479) );
  NAND2_X1 U9638 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n8015) );
  XOR2_X1 U9639 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10477) );
  NAND2_X1 U9640 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n8013) );
  XOR2_X1 U9641 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10463) );
  AOI21_X1 U9642 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10431) );
  INV_X1 U9643 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8011) );
  NAND3_X1 U9644 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10433) );
  OAI21_X1 U9645 ( .B1(n10431), .B2(n8011), .A(n10433), .ZN(n10462) );
  NAND2_X1 U9646 ( .A1(n10463), .A2(n10462), .ZN(n8012) );
  NAND2_X1 U9647 ( .A1(n8013), .A2(n8012), .ZN(n10476) );
  NAND2_X1 U9648 ( .A1(n10477), .A2(n10476), .ZN(n8014) );
  NAND2_X1 U9649 ( .A1(n8015), .A2(n8014), .ZN(n10478) );
  NOR2_X1 U9650 ( .A1(n10479), .A2(n10478), .ZN(n8016) );
  NOR2_X1 U9651 ( .A1(n8017), .A2(n8016), .ZN(n8018) );
  NOR2_X1 U9652 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n8018), .ZN(n10465) );
  AND2_X1 U9653 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n8018), .ZN(n10464) );
  NOR2_X1 U9654 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10464), .ZN(n8019) );
  NOR2_X1 U9655 ( .A1(n10465), .A2(n8019), .ZN(n8020) );
  NAND2_X1 U9656 ( .A1(n8020), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n8022) );
  XOR2_X1 U9657 ( .A(n8020), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10461) );
  NAND2_X1 U9658 ( .A1(n10461), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U9659 ( .A1(n8022), .A2(n8021), .ZN(n8023) );
  NAND2_X1 U9660 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8023), .ZN(n8025) );
  XOR2_X1 U9661 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8023), .Z(n10474) );
  NAND2_X1 U9662 ( .A1(n10474), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U9663 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  NAND2_X1 U9664 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8026), .ZN(n8028) );
  XOR2_X1 U9665 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n8026), .Z(n10475) );
  NAND2_X1 U9666 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10475), .ZN(n8027) );
  NAND2_X1 U9667 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  AND2_X1 U9668 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n8029), .ZN(n8030) );
  INV_X1 U9669 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10473) );
  XNOR2_X1 U9670 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n8029), .ZN(n10472) );
  NOR2_X1 U9671 ( .A1(n10473), .A2(n10472), .ZN(n10471) );
  NAND2_X1 U9672 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n8031) );
  OAI21_X1 U9673 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n8031), .ZN(n10459) );
  NAND2_X1 U9674 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n8032) );
  OAI21_X1 U9675 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8032), .ZN(n10456) );
  NOR2_X1 U9676 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8033) );
  AOI21_X1 U9677 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n8033), .ZN(n10453) );
  NAND2_X1 U9678 ( .A1(n10454), .A2(n10453), .ZN(n10452) );
  NAND2_X1 U9679 ( .A1(n10451), .A2(n10450), .ZN(n10449) );
  NAND2_X1 U9680 ( .A1(n10448), .A2(n10447), .ZN(n10446) );
  OAI21_X1 U9681 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10446), .ZN(n10444) );
  NAND2_X1 U9682 ( .A1(n10445), .A2(n10444), .ZN(n10443) );
  OAI21_X1 U9683 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10443), .ZN(n10441) );
  NAND2_X1 U9684 ( .A1(n10442), .A2(n10441), .ZN(n10440) );
  OAI21_X1 U9685 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10440), .ZN(n10438) );
  NAND2_X1 U9686 ( .A1(n10439), .A2(n10438), .ZN(n10437) );
  OAI21_X1 U9687 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10437), .ZN(n10468) );
  NOR2_X1 U9688 ( .A1(n10469), .A2(n10468), .ZN(n8034) );
  NAND2_X1 U9689 ( .A1(n10469), .A2(n10468), .ZN(n10467) );
  OAI21_X1 U9690 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n8034), .A(n10467), .ZN(
        n8036) );
  XNOR2_X1 U9691 ( .A(n4737), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n8035) );
  XNOR2_X1 U9692 ( .A(n8036), .B(n8035), .ZN(ADD_1071_U4) );
  AOI22_X1 U9693 ( .A1(n9647), .A2(n9203), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8038) );
  NAND2_X1 U9694 ( .A1(n9547), .A2(n9236), .ZN(n8037) );
  OAI211_X1 U9695 ( .C1(n9654), .C2(n9234), .A(n8038), .B(n8037), .ZN(n8041)
         );
  INV_X1 U9696 ( .A(n8053), .ZN(n8043) );
  NAND2_X1 U9697 ( .A1(n9849), .A2(n8044), .ZN(n8046) );
  NAND2_X1 U9698 ( .A1(n9545), .A2(n4480), .ZN(n8045) );
  NAND2_X1 U9699 ( .A1(n8046), .A2(n8045), .ZN(n8048) );
  XNOR2_X1 U9700 ( .A(n8048), .B(n8047), .ZN(n8050) );
  AOI22_X1 U9701 ( .A1(n9849), .A2(n7347), .B1(n7928), .B2(n9545), .ZN(n8049)
         );
  XNOR2_X1 U9702 ( .A(n8050), .B(n8049), .ZN(n8054) );
  INV_X1 U9703 ( .A(n8054), .ZN(n8059) );
  INV_X1 U9704 ( .A(n8051), .ZN(n8052) );
  NAND2_X1 U9705 ( .A1(n8053), .A2(n8052), .ZN(n8058) );
  NAND3_X1 U9706 ( .A1(n8059), .A2(n9211), .A3(n8058), .ZN(n8064) );
  NAND3_X1 U9707 ( .A1(n8065), .A2(n9211), .A3(n8054), .ZN(n8063) );
  NAND2_X1 U9708 ( .A1(n4778), .A2(n9236), .ZN(n8057) );
  INV_X1 U9709 ( .A(n9620), .ZN(n8055) );
  AOI22_X1 U9710 ( .A1(n8055), .A2(n9203), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8056) );
  OAI211_X1 U9711 ( .C1(n9616), .C2(n9234), .A(n8057), .B(n8056), .ZN(n8061)
         );
  NOR3_X1 U9712 ( .A1(n8059), .A2(n9253), .A3(n8058), .ZN(n8060) );
  AOI211_X1 U9713 ( .C1(n9849), .C2(n9251), .A(n8061), .B(n8060), .ZN(n8062)
         );
  OAI211_X1 U9714 ( .C1(n8065), .C2(n8064), .A(n8063), .B(n8062), .ZN(P1_U3218) );
  XNOR2_X1 U9715 ( .A(n8421), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n8429) );
  NOR2_X1 U9716 ( .A1(n8429), .A2(n8430), .ZN(n8428) );
  NAND2_X1 U9717 ( .A1(n8067), .A2(n8444), .ZN(n8068) );
  NAND2_X1 U9718 ( .A1(n8068), .A2(n8435), .ZN(n8069) );
  XNOR2_X1 U9719 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8069), .ZN(n8085) );
  INV_X1 U9720 ( .A(n8085), .ZN(n8083) );
  INV_X1 U9721 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8081) );
  INV_X1 U9722 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8079) );
  INV_X1 U9723 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8070) );
  MUX2_X1 U9724 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8070), .S(n8421), .Z(n8076)
         );
  OR2_X1 U9725 ( .A1(n8071), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8074) );
  INV_X1 U9726 ( .A(n8072), .ZN(n8073) );
  NAND2_X1 U9727 ( .A1(n8074), .A2(n8073), .ZN(n8425) );
  INV_X1 U9728 ( .A(n8425), .ZN(n8075) );
  NAND2_X1 U9729 ( .A1(n8076), .A2(n8075), .ZN(n8422) );
  NAND2_X1 U9730 ( .A1(n8421), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U9731 ( .A1(n8422), .A2(n8077), .ZN(n8439) );
  AOI22_X1 U9732 ( .A1(n8078), .A2(n8079), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8444), .ZN(n8438) );
  NOR2_X1 U9733 ( .A1(n8439), .A2(n8438), .ZN(n8441) );
  AOI21_X1 U9734 ( .B1(n8444), .B2(n8079), .A(n8441), .ZN(n8080) );
  XNOR2_X1 U9735 ( .A(n8081), .B(n8080), .ZN(n8084) );
  OAI21_X1 U9736 ( .B1(n8084), .B2(n10229), .A(n10227), .ZN(n8082) );
  AOI21_X1 U9737 ( .B1(n8083), .B2(n10226), .A(n8082), .ZN(n8088) );
  AOI22_X1 U9738 ( .A1(n8085), .A2(n10226), .B1(n10224), .B2(n8084), .ZN(n8087) );
  NAND2_X1 U9739 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8089) );
  OAI211_X1 U9740 ( .C1(n4737), .C2(n8091), .A(n8090), .B(n8089), .ZN(P2_U3264) );
  NAND2_X1 U9741 ( .A1(n8092), .A2(n6907), .ZN(n8093) );
  NAND2_X1 U9742 ( .A1(n8106), .A2(n6907), .ZN(n8096) );
  INV_X1 U9743 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8108) );
  OR2_X1 U9744 ( .A1(n8094), .A2(n8108), .ZN(n8095) );
  NAND2_X1 U9745 ( .A1(n9607), .A2(n9606), .ZN(n9605) );
  XNOR2_X1 U9746 ( .A(n9839), .B(n9605), .ZN(n9837) );
  NAND2_X1 U9747 ( .A1(n9837), .A2(n9733), .ZN(n8105) );
  INV_X1 U9748 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8097) );
  NOR2_X1 U9749 ( .A1(n4478), .A2(n8097), .ZN(n8102) );
  INV_X1 U9750 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8098) );
  NOR2_X1 U9751 ( .A1(n4476), .A2(n8098), .ZN(n8101) );
  INV_X1 U9752 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8099) );
  NOR2_X1 U9753 ( .A1(n6557), .A2(n8099), .ZN(n8100) );
  OR3_X1 U9754 ( .A1(n8102), .A2(n8101), .A3(n8100), .ZN(n9543) );
  NAND2_X1 U9755 ( .A1(n9543), .A2(n8103), .ZN(n9842) );
  NOR2_X1 U9756 ( .A1(n10157), .A2(n9842), .ZN(n9609) );
  AOI21_X1 U9757 ( .B1(n10157), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9609), .ZN(
        n8104) );
  OAI211_X1 U9758 ( .C1(n9839), .C2(n9799), .A(n8105), .B(n8104), .ZN(P1_U3261) );
  INV_X1 U9759 ( .A(n8106), .ZN(n9124) );
  OAI222_X1 U9760 ( .A1(n9968), .A2(n8108), .B1(n9971), .B2(n9124), .C1(n8107), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  INV_X1 U9761 ( .A(n8539), .ZN(n8499) );
  INV_X1 U9762 ( .A(n9094), .ZN(n8614) );
  NOR2_X1 U9763 ( .A1(n9098), .A2(n8369), .ZN(n8112) );
  INV_X1 U9764 ( .A(n9098), .ZN(n8628) );
  INV_X1 U9765 ( .A(n9081), .ZN(n8583) );
  NAND2_X1 U9766 ( .A1(n8583), .A2(n8593), .ZN(n8113) );
  INV_X1 U9767 ( .A(n8569), .ZN(n8114) );
  INV_X1 U9768 ( .A(n9076), .ZN(n8567) );
  OAI21_X1 U9769 ( .B1(n9063), .B2(n8499), .A(n8511), .ZN(n8493) );
  NAND2_X1 U9770 ( .A1(n8493), .A2(n8492), .ZN(n8491) );
  INV_X1 U9771 ( .A(n8477), .ZN(n8368) );
  NAND2_X1 U9772 ( .A1(n8491), .A2(n8115), .ZN(n8483) );
  NAND2_X1 U9773 ( .A1(n8483), .A2(n8482), .ZN(n8481) );
  INV_X1 U9774 ( .A(n8498), .ZN(n8367) );
  NAND2_X1 U9775 ( .A1(n8481), .A2(n8117), .ZN(n8465) );
  NAND2_X1 U9776 ( .A1(n8465), .A2(n8464), .ZN(n8463) );
  INV_X1 U9777 ( .A(n9063), .ZN(n8518) );
  INV_X1 U9778 ( .A(n8602), .ZN(n8611) );
  NAND2_X1 U9779 ( .A1(n8518), .A2(n8531), .ZN(n8515) );
  AOI21_X1 U9780 ( .B1(n9037), .B2(n8466), .A(n8452), .ZN(n9038) );
  INV_X1 U9781 ( .A(n9037), .ZN(n8121) );
  INV_X1 U9782 ( .A(n8118), .ZN(n8119) );
  AOI22_X1 U9783 ( .A1(n10308), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8119), .B2(
        n10245), .ZN(n8120) );
  OAI21_X1 U9784 ( .B1(n8121), .B2(n8627), .A(n8120), .ZN(n8122) );
  AOI21_X1 U9785 ( .B1(n9038), .B2(n8637), .A(n8122), .ZN(n8129) );
  XNOR2_X1 U9786 ( .A(n8124), .B(n8123), .ZN(n8127) );
  INV_X1 U9787 ( .A(P2_B_REG_SCAN_IN), .ZN(n8125) );
  NOR2_X1 U9788 ( .A1(n9133), .A2(n8125), .ZN(n8126) );
  NOR2_X1 U9789 ( .A1(n10284), .A2(n8126), .ZN(n8448) );
  OR2_X1 U9790 ( .A1(n9040), .A2(n10308), .ZN(n8128) );
  OAI211_X1 U9791 ( .C1(n9041), .C2(n8639), .A(n8129), .B(n8128), .ZN(P2_U3267) );
  XNOR2_X1 U9792 ( .A(n9066), .B(n8212), .ZN(n8158) );
  NAND2_X1 U9793 ( .A1(n8558), .A2(n4486), .ZN(n8299) );
  NAND2_X1 U9794 ( .A1(n8325), .A2(n8130), .ZN(n8135) );
  XNOR2_X1 U9795 ( .A(n9098), .B(n8165), .ZN(n8194) );
  AND2_X1 U9796 ( .A1(n8369), .A2(n8156), .ZN(n8131) );
  NAND2_X1 U9797 ( .A1(n8194), .A2(n8131), .ZN(n8136) );
  INV_X1 U9798 ( .A(n8194), .ZN(n8133) );
  INV_X1 U9799 ( .A(n8131), .ZN(n8132) );
  NAND2_X1 U9800 ( .A1(n8133), .A2(n8132), .ZN(n8134) );
  AND2_X1 U9801 ( .A1(n8136), .A2(n8134), .ZN(n8323) );
  XNOR2_X1 U9802 ( .A(n9094), .B(n8165), .ZN(n8137) );
  NAND2_X1 U9803 ( .A1(n8632), .A2(n4486), .ZN(n8138) );
  XNOR2_X1 U9804 ( .A(n8137), .B(n8138), .ZN(n8196) );
  INV_X1 U9805 ( .A(n8137), .ZN(n8139) );
  NAND2_X1 U9806 ( .A1(n8139), .A2(n8138), .ZN(n8140) );
  XNOR2_X1 U9807 ( .A(n9088), .B(n8165), .ZN(n8141) );
  AND2_X1 U9808 ( .A1(n8586), .A2(n8156), .ZN(n8142) );
  NAND2_X1 U9809 ( .A1(n8141), .A2(n8142), .ZN(n8147) );
  INV_X1 U9810 ( .A(n8141), .ZN(n8244) );
  INV_X1 U9811 ( .A(n8142), .ZN(n8143) );
  NAND2_X1 U9812 ( .A1(n8244), .A2(n8143), .ZN(n8144) );
  NAND2_X1 U9813 ( .A1(n8147), .A2(n8144), .ZN(n8308) );
  XNOR2_X1 U9814 ( .A(n9081), .B(n8165), .ZN(n8150) );
  NAND2_X1 U9815 ( .A1(n8571), .A2(n4486), .ZN(n8148) );
  XNOR2_X1 U9816 ( .A(n8150), .B(n8148), .ZN(n8241) );
  INV_X1 U9817 ( .A(n8148), .ZN(n8149) );
  XNOR2_X1 U9818 ( .A(n9076), .B(n8212), .ZN(n8151) );
  NAND2_X1 U9819 ( .A1(n8587), .A2(n8156), .ZN(n8314) );
  INV_X1 U9820 ( .A(n8151), .ZN(n8152) );
  NAND2_X1 U9821 ( .A1(n8572), .A2(n8156), .ZN(n8175) );
  AOI21_X1 U9822 ( .B1(n8158), .B2(n8297), .A(n8175), .ZN(n8157) );
  INV_X1 U9823 ( .A(n8158), .ZN(n8295) );
  INV_X1 U9824 ( .A(n8299), .ZN(n8159) );
  NAND2_X1 U9825 ( .A1(n8295), .A2(n8159), .ZN(n8160) );
  XNOR2_X1 U9826 ( .A(n9063), .B(n8165), .ZN(n8161) );
  NOR2_X1 U9827 ( .A1(n8539), .A2(n8211), .ZN(n8162) );
  AND2_X1 U9828 ( .A1(n8161), .A2(n8162), .ZN(n8253) );
  INV_X1 U9829 ( .A(n8161), .ZN(n8254) );
  INV_X1 U9830 ( .A(n8162), .ZN(n8163) );
  NAND2_X1 U9831 ( .A1(n8254), .A2(n8163), .ZN(n8252) );
  NAND2_X1 U9832 ( .A1(n8164), .A2(n8252), .ZN(n8352) );
  XNOR2_X1 U9833 ( .A(n9056), .B(n8165), .ZN(n8167) );
  NOR2_X1 U9834 ( .A1(n8477), .A2(n8211), .ZN(n8166) );
  XNOR2_X1 U9835 ( .A(n8167), .B(n8166), .ZN(n8351) );
  NAND2_X1 U9836 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  XNOR2_X1 U9837 ( .A(n9049), .B(n8212), .ZN(n8206) );
  NOR2_X1 U9838 ( .A1(n8498), .A2(n8211), .ZN(n8207) );
  XNOR2_X1 U9839 ( .A(n8206), .B(n8207), .ZN(n8209) );
  XNOR2_X1 U9840 ( .A(n8210), .B(n8209), .ZN(n8174) );
  INV_X1 U9841 ( .A(n8486), .ZN(n8170) );
  OAI22_X1 U9842 ( .A1(n8355), .A2(n8170), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8169), .ZN(n8172) );
  OAI22_X1 U9843 ( .A1(n8357), .A2(n8478), .B1(n8356), .B2(n8477), .ZN(n8171)
         );
  AOI211_X1 U9844 ( .C1(n9049), .C2(n8360), .A(n8172), .B(n8171), .ZN(n8173)
         );
  OAI21_X1 U9845 ( .B1(n8174), .B2(n8362), .A(n8173), .ZN(P2_U3216) );
  AOI22_X1 U9846 ( .A1(n8177), .A2(n8336), .B1(n8313), .B2(n8572), .ZN(n8184)
         );
  INV_X1 U9847 ( .A(n8175), .ZN(n8176) );
  NAND2_X1 U9848 ( .A1(n8177), .A2(n8176), .ZN(n8294) );
  INV_X1 U9849 ( .A(n8294), .ZN(n8183) );
  OAI22_X1 U9850 ( .A1(n8355), .A2(n8551), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8178), .ZN(n8181) );
  OAI22_X1 U9851 ( .A1(n8357), .A2(n8297), .B1(n8356), .B2(n8179), .ZN(n8180)
         );
  AOI211_X1 U9852 ( .C1(n9071), .C2(n8360), .A(n8181), .B(n8180), .ZN(n8182)
         );
  OAI21_X1 U9853 ( .B1(n8184), .B2(n8183), .A(n8182), .ZN(P2_U3218) );
  OAI211_X1 U9854 ( .C1(n8187), .C2(n8186), .A(n8185), .B(n8336), .ZN(n8193)
         );
  AOI22_X1 U9855 ( .A1(n8342), .A2(n8188), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n8192) );
  AOI22_X1 U9856 ( .A1(n8318), .A2(n8374), .B1(n8346), .B2(n8376), .ZN(n8191)
         );
  NAND2_X1 U9857 ( .A1(n8189), .A2(n8360), .ZN(n8190) );
  NAND4_X1 U9858 ( .A1(n8193), .A2(n8192), .A3(n8191), .A4(n8190), .ZN(
        P2_U3219) );
  NAND3_X1 U9859 ( .A1(n8194), .A2(n8313), .A3(n8369), .ZN(n8195) );
  OAI21_X1 U9860 ( .B1(n8327), .B2(n8362), .A(n8195), .ZN(n8203) );
  INV_X1 U9861 ( .A(n8196), .ZN(n8202) );
  NAND2_X1 U9862 ( .A1(n8586), .A2(n10261), .ZN(n8198) );
  NAND2_X1 U9863 ( .A1(n8369), .A2(n10259), .ZN(n8197) );
  NAND2_X1 U9864 ( .A1(n8198), .A2(n8197), .ZN(n8617) );
  AOI22_X1 U9865 ( .A1(n8287), .A2(n8617), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8200) );
  NAND2_X1 U9866 ( .A1(n8342), .A2(n8612), .ZN(n8199) );
  OAI211_X1 U9867 ( .C1(n8614), .C2(n8338), .A(n8200), .B(n8199), .ZN(n8201)
         );
  AOI21_X1 U9868 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8204) );
  OAI21_X1 U9869 ( .B1(n8205), .B2(n8362), .A(n8204), .ZN(P2_U3221) );
  INV_X1 U9870 ( .A(n8206), .ZN(n8208) );
  NOR2_X1 U9871 ( .A1(n8478), .A2(n8211), .ZN(n8213) );
  XNOR2_X1 U9872 ( .A(n8213), .B(n8212), .ZN(n8215) );
  INV_X1 U9873 ( .A(n8215), .ZN(n8216) );
  NOR3_X1 U9874 ( .A1(n8471), .A2(n8216), .A3(n8360), .ZN(n8214) );
  AOI21_X1 U9875 ( .B1(n8471), .B2(n8216), .A(n8214), .ZN(n8221) );
  NOR3_X1 U9876 ( .A1(n8471), .A2(n8215), .A3(n8360), .ZN(n8218) );
  NOR2_X1 U9877 ( .A1(n9043), .A2(n8216), .ZN(n8217) );
  OAI21_X1 U9878 ( .B1(n8471), .B2(n8338), .A(n8362), .ZN(n8220) );
  INV_X1 U9879 ( .A(n8222), .ZN(n8469) );
  AOI22_X1 U9880 ( .A1(n8342), .A2(n8469), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8224) );
  INV_X1 U9881 ( .A(n8460), .ZN(n8365) );
  AOI22_X1 U9882 ( .A1(n8318), .A2(n8365), .B1(n8367), .B2(n8346), .ZN(n8223)
         );
  NAND3_X1 U9883 ( .A1(n8225), .A2(n8224), .A3(n8223), .ZN(P2_U3222) );
  INV_X1 U9884 ( .A(n8226), .ZN(n8227) );
  AOI21_X1 U9885 ( .B1(n8228), .B2(n8227), .A(n8362), .ZN(n8232) );
  NOR3_X1 U9886 ( .A1(n8345), .A2(n8339), .A3(n8229), .ZN(n8231) );
  OAI21_X1 U9887 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(n8240) );
  NAND2_X1 U9888 ( .A1(n8376), .A2(n10261), .ZN(n8234) );
  NAND2_X1 U9889 ( .A1(n10262), .A2(n10259), .ZN(n8233) );
  AND2_X1 U9890 ( .A1(n8234), .A2(n8233), .ZN(n10240) );
  OAI22_X1 U9891 ( .A1(n8263), .A2(n10240), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8235), .ZN(n8236) );
  INV_X1 U9892 ( .A(n8236), .ZN(n8239) );
  NAND2_X1 U9893 ( .A1(n8360), .A2(n10375), .ZN(n8238) );
  NAND2_X1 U9894 ( .A1(n8342), .A2(n10244), .ZN(n8237) );
  NAND4_X1 U9895 ( .A1(n8240), .A2(n8239), .A3(n8238), .A4(n8237), .ZN(
        P2_U3223) );
  INV_X1 U9896 ( .A(n8241), .ZN(n8242) );
  AOI21_X1 U9897 ( .B1(n8305), .B2(n8242), .A(n8362), .ZN(n8247) );
  NOR3_X1 U9898 ( .A1(n8244), .A2(n8243), .A3(n8345), .ZN(n8246) );
  OAI21_X1 U9899 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8251) );
  AOI22_X1 U9900 ( .A1(n8342), .A2(n8581), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8250) );
  AOI22_X1 U9901 ( .A1(n8318), .A2(n8587), .B1(n8346), .B2(n8586), .ZN(n8249)
         );
  NAND2_X1 U9902 ( .A1(n9081), .A2(n8360), .ZN(n8248) );
  NAND4_X1 U9903 ( .A1(n8251), .A2(n8250), .A3(n8249), .A4(n8248), .ZN(
        P2_U3225) );
  INV_X1 U9904 ( .A(n8252), .ZN(n8256) );
  OR3_X1 U9905 ( .A1(n8253), .A2(n8256), .A3(n8362), .ZN(n8259) );
  NOR3_X1 U9906 ( .A1(n8254), .A2(n8539), .A3(n8345), .ZN(n8255) );
  AOI21_X1 U9907 ( .B1(n8336), .B2(n8256), .A(n8255), .ZN(n8258) );
  MUX2_X1 U9908 ( .A(n8259), .B(n8258), .S(n8257), .Z(n8267) );
  INV_X1 U9909 ( .A(n8519), .ZN(n8265) );
  OR2_X1 U9910 ( .A1(n8477), .A2(n10284), .ZN(n8261) );
  NAND2_X1 U9911 ( .A1(n8558), .A2(n10259), .ZN(n8260) );
  AND2_X1 U9912 ( .A1(n8261), .A2(n8260), .ZN(n8526) );
  OAI22_X1 U9913 ( .A1(n8526), .A2(n8263), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8262), .ZN(n8264) );
  AOI21_X1 U9914 ( .B1(n8265), .B2(n8342), .A(n8264), .ZN(n8266) );
  OAI211_X1 U9915 ( .C1(n8518), .C2(n8338), .A(n8267), .B(n8266), .ZN(P2_U3227) );
  INV_X1 U9916 ( .A(n8268), .ZN(n8271) );
  OAI21_X1 U9917 ( .B1(n8271), .B2(n8270), .A(n8269), .ZN(n8275) );
  XNOR2_X1 U9918 ( .A(n8273), .B(n8272), .ZN(n8274) );
  XNOR2_X1 U9919 ( .A(n8275), .B(n8274), .ZN(n8282) );
  INV_X1 U9920 ( .A(n8655), .ZN(n8277) );
  OAI22_X1 U9921 ( .A1(n8355), .A2(n8277), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8276), .ZN(n8280) );
  OAI22_X1 U9922 ( .A1(n8357), .A2(n8330), .B1(n8356), .B2(n8278), .ZN(n8279)
         );
  AOI211_X1 U9923 ( .C1(n10015), .C2(n8360), .A(n8280), .B(n8279), .ZN(n8281)
         );
  OAI21_X1 U9924 ( .B1(n8282), .B2(n8362), .A(n8281), .ZN(P2_U3228) );
  AOI21_X1 U9925 ( .B1(n8284), .B2(n8283), .A(n8362), .ZN(n8285) );
  NAND2_X1 U9926 ( .A1(n8285), .A2(n8335), .ZN(n8292) );
  AOI22_X1 U9927 ( .A1(n8287), .A2(n8286), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n8291) );
  AOI22_X1 U9928 ( .A1(n8360), .A2(n8289), .B1(n8342), .B2(n8288), .ZN(n8290)
         );
  NAND3_X1 U9929 ( .A1(n8292), .A2(n8291), .A3(n8290), .ZN(P2_U3229) );
  INV_X1 U9930 ( .A(n9066), .ZN(n8535) );
  NAND2_X1 U9931 ( .A1(n8294), .A2(n8293), .ZN(n8296) );
  XNOR2_X1 U9932 ( .A(n8296), .B(n8295), .ZN(n8300) );
  OAI22_X1 U9933 ( .A1(n8300), .A2(n8362), .B1(n8297), .B2(n8345), .ZN(n8298)
         );
  OAI21_X1 U9934 ( .B1(n8300), .B2(n8299), .A(n8298), .ZN(n8304) );
  NOR2_X1 U9935 ( .A1(n8355), .A2(n8532), .ZN(n8302) );
  OAI22_X1 U9936 ( .A1(n8357), .A2(n8539), .B1(n8356), .B2(n8538), .ZN(n8301)
         );
  AOI211_X1 U9937 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3152), .A(n8302), 
        .B(n8301), .ZN(n8303) );
  OAI211_X1 U9938 ( .C1(n8535), .C2(n8338), .A(n8304), .B(n8303), .ZN(P2_U3231) );
  INV_X1 U9939 ( .A(n8305), .ZN(n8306) );
  AOI211_X1 U9940 ( .C1(n8308), .C2(n8307), .A(n8362), .B(n8306), .ZN(n8312)
         );
  AOI22_X1 U9941 ( .A1(n8342), .A2(n8603), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8310) );
  AOI22_X1 U9942 ( .A1(n8318), .A2(n8571), .B1(n8346), .B2(n8632), .ZN(n8309)
         );
  OAI211_X1 U9943 ( .C1(n8605), .C2(n8338), .A(n8310), .B(n8309), .ZN(n8311)
         );
  OR2_X1 U9944 ( .A1(n8312), .A2(n8311), .ZN(P2_U3235) );
  NAND2_X1 U9945 ( .A1(n8313), .A2(n8587), .ZN(n8317) );
  NAND2_X1 U9946 ( .A1(n8336), .A2(n8314), .ZN(n8316) );
  MUX2_X1 U9947 ( .A(n8317), .B(n8316), .S(n8315), .Z(n8322) );
  AOI22_X1 U9948 ( .A1(n8342), .A2(n8565), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8321) );
  AOI22_X1 U9949 ( .A1(n8318), .A2(n8572), .B1(n8346), .B2(n8571), .ZN(n8320)
         );
  NAND2_X1 U9950 ( .A1(n9076), .A2(n8360), .ZN(n8319) );
  NAND4_X1 U9951 ( .A1(n8322), .A2(n8321), .A3(n8320), .A4(n8319), .ZN(
        P2_U3237) );
  INV_X1 U9952 ( .A(n8323), .ZN(n8324) );
  AOI21_X1 U9953 ( .B1(n8325), .B2(n8324), .A(n8362), .ZN(n8329) );
  NOR3_X1 U9954 ( .A1(n8326), .A2(n8330), .A3(n8345), .ZN(n8328) );
  OAI21_X1 U9955 ( .B1(n8329), .B2(n8328), .A(n8327), .ZN(n8333) );
  AND2_X1 U9956 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8437) );
  OAI22_X1 U9957 ( .A1(n8357), .A2(n8594), .B1(n8356), .B2(n8330), .ZN(n8331)
         );
  AOI211_X1 U9958 ( .C1(n8342), .C2(n8625), .A(n8437), .B(n8331), .ZN(n8332)
         );
  OAI211_X1 U9959 ( .C1(n8628), .C2(n8338), .A(n8333), .B(n8332), .ZN(P2_U3240) );
  OAI21_X1 U9960 ( .B1(n8344), .B2(n8335), .A(n8334), .ZN(n8337) );
  NAND2_X1 U9961 ( .A1(n8337), .A2(n8336), .ZN(n8350) );
  OAI22_X1 U9962 ( .A1(n8357), .A2(n8339), .B1(n10361), .B2(n8338), .ZN(n8340)
         );
  AOI211_X1 U9963 ( .C1(n10268), .C2(n8342), .A(n8341), .B(n8340), .ZN(n8349)
         );
  NOR3_X1 U9964 ( .A1(n8345), .A2(n8344), .A3(n8343), .ZN(n8347) );
  OAI21_X1 U9965 ( .B1(n8347), .B2(n8346), .A(n10260), .ZN(n8348) );
  NAND3_X1 U9966 ( .A1(n8350), .A2(n8349), .A3(n8348), .ZN(P2_U3241) );
  XNOR2_X1 U9967 ( .A(n8352), .B(n8351), .ZN(n8363) );
  INV_X1 U9968 ( .A(n8502), .ZN(n8354) );
  OAI22_X1 U9969 ( .A1(n8355), .A2(n8354), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8353), .ZN(n8359) );
  OAI22_X1 U9970 ( .A1(n8357), .A2(n8498), .B1(n8356), .B2(n8539), .ZN(n8358)
         );
  AOI211_X1 U9971 ( .C1(n9056), .C2(n8360), .A(n8359), .B(n8358), .ZN(n8361)
         );
  OAI21_X1 U9972 ( .B1(n8363), .B2(n8362), .A(n8361), .ZN(P2_U3242) );
  MUX2_X1 U9973 ( .A(n8364), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8383), .Z(
        P2_U3582) );
  MUX2_X1 U9974 ( .A(n8365), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8383), .Z(
        P2_U3581) );
  MUX2_X1 U9975 ( .A(n8366), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8383), .Z(
        P2_U3580) );
  MUX2_X1 U9976 ( .A(n8367), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8383), .Z(
        P2_U3579) );
  MUX2_X1 U9977 ( .A(n8368), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8383), .Z(
        P2_U3578) );
  MUX2_X1 U9978 ( .A(n8499), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8383), .Z(
        P2_U3577) );
  MUX2_X1 U9979 ( .A(n8558), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8383), .Z(
        P2_U3576) );
  MUX2_X1 U9980 ( .A(n8572), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8383), .Z(
        P2_U3575) );
  MUX2_X1 U9981 ( .A(n8587), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8383), .Z(
        P2_U3574) );
  MUX2_X1 U9982 ( .A(n8571), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8383), .Z(
        P2_U3573) );
  MUX2_X1 U9983 ( .A(n8586), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8383), .Z(
        P2_U3572) );
  MUX2_X1 U9984 ( .A(n8632), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8383), .Z(
        P2_U3571) );
  MUX2_X1 U9985 ( .A(n8369), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8383), .Z(
        P2_U3570) );
  MUX2_X1 U9986 ( .A(n8647), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8383), .Z(
        P2_U3569) );
  MUX2_X1 U9987 ( .A(n8370), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8383), .Z(
        P2_U3568) );
  MUX2_X1 U9988 ( .A(n8648), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8383), .Z(
        P2_U3567) );
  MUX2_X1 U9989 ( .A(n8371), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8379), .Z(
        P2_U3566) );
  MUX2_X1 U9990 ( .A(n8372), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8379), .Z(
        P2_U3565) );
  MUX2_X1 U9991 ( .A(n8373), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8379), .Z(
        P2_U3564) );
  MUX2_X1 U9992 ( .A(n8374), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8379), .Z(
        P2_U3563) );
  MUX2_X1 U9993 ( .A(n8375), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8379), .Z(
        P2_U3562) );
  MUX2_X1 U9994 ( .A(n8376), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8379), .Z(
        P2_U3561) );
  MUX2_X1 U9995 ( .A(n8377), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8379), .Z(
        P2_U3560) );
  MUX2_X1 U9996 ( .A(n10262), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8379), .Z(
        P2_U3559) );
  MUX2_X1 U9997 ( .A(n8378), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8379), .Z(
        P2_U3558) );
  MUX2_X1 U9998 ( .A(n10260), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8379), .Z(
        P2_U3557) );
  MUX2_X1 U9999 ( .A(n8380), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8383), .Z(
        P2_U3556) );
  MUX2_X1 U10000 ( .A(n8381), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8383), .Z(
        P2_U3555) );
  MUX2_X1 U10001 ( .A(n8382), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8383), .Z(
        P2_U3554) );
  MUX2_X1 U10002 ( .A(n6578), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8383), .Z(
        P2_U3553) );
  NAND2_X1 U10003 ( .A1(n9992), .A2(n8384), .ZN(n8395) );
  OAI211_X1 U10004 ( .C1(n8387), .C2(n8386), .A(n10226), .B(n8385), .ZN(n8394)
         );
  AND2_X1 U10005 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8388) );
  AOI21_X1 U10006 ( .B1(n10231), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8388), .ZN(
        n8393) );
  OAI211_X1 U10007 ( .C1(n8391), .C2(n8390), .A(n10224), .B(n8389), .ZN(n8392)
         );
  NAND4_X1 U10008 ( .A1(n8395), .A2(n8394), .A3(n8393), .A4(n8392), .ZN(
        P2_U3254) );
  NAND2_X1 U10009 ( .A1(n9992), .A2(n8396), .ZN(n8407) );
  OAI211_X1 U10010 ( .C1(n8399), .C2(n8398), .A(n10226), .B(n8397), .ZN(n8406)
         );
  NOR2_X1 U10011 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8830), .ZN(n8400) );
  AOI21_X1 U10012 ( .B1(n10231), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8400), .ZN(
        n8405) );
  OAI211_X1 U10013 ( .C1(n8403), .C2(n8402), .A(n10224), .B(n8401), .ZN(n8404)
         );
  NAND4_X1 U10014 ( .A1(n8407), .A2(n8406), .A3(n8405), .A4(n8404), .ZN(
        P2_U3255) );
  NOR2_X1 U10015 ( .A1(n8409), .A2(n8408), .ZN(n8411) );
  OAI21_X1 U10016 ( .B1(n8411), .B2(n8410), .A(n10224), .ZN(n8420) );
  AOI21_X1 U10017 ( .B1(n10231), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8412), .ZN(
        n8419) );
  OAI211_X1 U10018 ( .C1(n8415), .C2(n8414), .A(n10226), .B(n8413), .ZN(n8418)
         );
  OR2_X1 U10019 ( .A1(n10227), .A2(n8416), .ZN(n8417) );
  NAND4_X1 U10020 ( .A1(n8420), .A2(n8419), .A3(n8418), .A4(n8417), .ZN(
        P2_U3257) );
  INV_X1 U10021 ( .A(n8421), .ZN(n8434) );
  AND2_X1 U10022 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8427) );
  MUX2_X1 U10023 ( .A(n8070), .B(P2_REG1_REG_17__SCAN_IN), .S(n8421), .Z(n8424) );
  INV_X1 U10024 ( .A(n8422), .ZN(n8423) );
  AOI211_X1 U10025 ( .C1(n8425), .C2(n8424), .A(n8423), .B(n10229), .ZN(n8426)
         );
  AOI211_X1 U10026 ( .C1(n10231), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8427), .B(
        n8426), .ZN(n8433) );
  AOI211_X1 U10027 ( .C1(n8430), .C2(n8429), .A(n8428), .B(n9986), .ZN(n8431)
         );
  INV_X1 U10028 ( .A(n8431), .ZN(n8432) );
  OAI211_X1 U10029 ( .C1(n10227), .C2(n8434), .A(n8433), .B(n8432), .ZN(
        P2_U3262) );
  OAI21_X1 U10030 ( .B1(n8436), .B2(n5505), .A(n8435), .ZN(n8446) );
  AOI21_X1 U10031 ( .B1(n10231), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8437), .ZN(
        n8443) );
  AND2_X1 U10032 ( .A1(n8439), .A2(n8438), .ZN(n8440) );
  OAI21_X1 U10033 ( .B1(n8441), .B2(n8440), .A(n10224), .ZN(n8442) );
  OAI211_X1 U10034 ( .C1(n10227), .C2(n8444), .A(n8443), .B(n8442), .ZN(n8445)
         );
  AOI21_X1 U10035 ( .B1(n8446), .B2(n10226), .A(n8445), .ZN(n8447) );
  INV_X1 U10036 ( .A(n8447), .ZN(P2_U3263) );
  NAND2_X1 U10037 ( .A1(n9034), .A2(n8452), .ZN(n9030) );
  XNOR2_X1 U10038 ( .A(n9030), .B(n9022), .ZN(n9024) );
  NAND2_X1 U10039 ( .A1(n8449), .A2(n8448), .ZN(n9032) );
  NOR2_X1 U10040 ( .A1(n10308), .A2(n9032), .ZN(n8455) );
  AOI21_X1 U10041 ( .B1(n10308), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8455), .ZN(
        n8451) );
  NAND2_X1 U10042 ( .A1(n9022), .A2(n10302), .ZN(n8450) );
  OAI211_X1 U10043 ( .C1(n9024), .C2(n10273), .A(n8451), .B(n8450), .ZN(
        P2_U3265) );
  INV_X1 U10044 ( .A(n8452), .ZN(n8453) );
  NAND2_X1 U10045 ( .A1(n8454), .A2(n8453), .ZN(n9031) );
  NAND3_X1 U10046 ( .A1(n9031), .A2(n8637), .A3(n9030), .ZN(n8457) );
  AOI21_X1 U10047 ( .B1(n10308), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8455), .ZN(
        n8456) );
  OAI211_X1 U10048 ( .C1(n9034), .C2(n8627), .A(n8457), .B(n8456), .ZN(
        P2_U3266) );
  AOI211_X1 U10049 ( .C1(n8459), .C2(n8464), .A(n10281), .B(n8458), .ZN(n8462)
         );
  OAI22_X1 U10050 ( .A1(n8498), .A2(n10286), .B1(n8460), .B2(n10284), .ZN(
        n8461) );
  NOR2_X1 U10051 ( .A1(n8462), .A2(n8461), .ZN(n9046) );
  OAI21_X1 U10052 ( .B1(n8465), .B2(n8464), .A(n8463), .ZN(n9042) );
  NAND2_X1 U10053 ( .A1(n9042), .A2(n10306), .ZN(n8474) );
  INV_X1 U10054 ( .A(n8485), .ZN(n8468) );
  INV_X1 U10055 ( .A(n8466), .ZN(n8467) );
  AOI21_X1 U10056 ( .B1(n9043), .B2(n8468), .A(n8467), .ZN(n9044) );
  AOI22_X1 U10057 ( .A1(n10308), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8469), 
        .B2(n10245), .ZN(n8470) );
  OAI21_X1 U10058 ( .B1(n8471), .B2(n8627), .A(n8470), .ZN(n8472) );
  AOI21_X1 U10059 ( .B1(n9044), .B2(n8637), .A(n8472), .ZN(n8473) );
  OAI211_X1 U10060 ( .C1(n10308), .C2(n9046), .A(n8474), .B(n8473), .ZN(
        P2_U3268) );
  AOI211_X1 U10061 ( .C1(n8482), .C2(n8476), .A(n10281), .B(n8475), .ZN(n8480)
         );
  OAI22_X1 U10062 ( .A1(n8478), .A2(n10284), .B1(n8477), .B2(n10286), .ZN(
        n8479) );
  NOR2_X1 U10063 ( .A1(n8480), .A2(n8479), .ZN(n9052) );
  OAI21_X1 U10064 ( .B1(n8483), .B2(n8482), .A(n8481), .ZN(n9048) );
  AND2_X1 U10065 ( .A1(n9049), .A2(n4506), .ZN(n8484) );
  NOR2_X1 U10066 ( .A1(n8485), .A2(n8484), .ZN(n9050) );
  NAND2_X1 U10067 ( .A1(n9050), .A2(n8637), .ZN(n8488) );
  AOI22_X1 U10068 ( .A1(n10308), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8486), 
        .B2(n10245), .ZN(n8487) );
  OAI211_X1 U10069 ( .C1(n8116), .C2(n8627), .A(n8488), .B(n8487), .ZN(n8489)
         );
  AOI21_X1 U10070 ( .B1(n9048), .B2(n10306), .A(n8489), .ZN(n8490) );
  OAI21_X1 U10071 ( .B1(n10308), .B2(n9052), .A(n8490), .ZN(P2_U3269) );
  OAI21_X1 U10072 ( .B1(n8493), .B2(n8492), .A(n8491), .ZN(n9054) );
  INV_X1 U10073 ( .A(n9054), .ZN(n8510) );
  AOI22_X1 U10074 ( .A1(n9056), .A2(n10302), .B1(n10308), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8509) );
  OAI21_X1 U10075 ( .B1(n8495), .B2(n4540), .A(n8494), .ZN(n8496) );
  NAND2_X1 U10076 ( .A1(n8496), .A2(n10264), .ZN(n9058) );
  INV_X1 U10077 ( .A(n9058), .ZN(n8507) );
  AOI21_X1 U10078 ( .B1(n9056), .B2(n8515), .A(n10402), .ZN(n8497) );
  NAND2_X1 U10079 ( .A1(n8497), .A2(n4506), .ZN(n9057) );
  OR2_X1 U10080 ( .A1(n8498), .A2(n10284), .ZN(n8501) );
  NAND2_X1 U10081 ( .A1(n8499), .A2(n10259), .ZN(n8500) );
  NAND2_X1 U10082 ( .A1(n8501), .A2(n8500), .ZN(n9055) );
  INV_X1 U10083 ( .A(n9055), .ZN(n8504) );
  NAND2_X1 U10084 ( .A1(n10245), .A2(n8502), .ZN(n8503) );
  OAI211_X1 U10085 ( .C1(n9057), .C2(n4573), .A(n8504), .B(n8503), .ZN(n8506)
         );
  OAI21_X1 U10086 ( .B1(n8507), .B2(n8506), .A(n10299), .ZN(n8508) );
  OAI211_X1 U10087 ( .C1(n8510), .C2(n8639), .A(n8509), .B(n8508), .ZN(
        P2_U3270) );
  OAI21_X1 U10088 ( .B1(n8513), .B2(n8512), .A(n8511), .ZN(n8514) );
  INV_X1 U10089 ( .A(n8514), .ZN(n9065) );
  INV_X1 U10090 ( .A(n8531), .ZN(n8517) );
  INV_X1 U10091 ( .A(n8515), .ZN(n8516) );
  AOI211_X1 U10092 ( .C1(n9063), .C2(n8517), .A(n10402), .B(n8516), .ZN(n9062)
         );
  INV_X1 U10093 ( .A(n10304), .ZN(n10250) );
  NOR2_X1 U10094 ( .A1(n8518), .A2(n8627), .ZN(n8522) );
  INV_X1 U10095 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8520) );
  OAI22_X1 U10096 ( .A1(n10299), .A2(n8520), .B1(n8519), .B2(n10297), .ZN(
        n8521) );
  AOI211_X1 U10097 ( .C1(n9062), .C2(n10250), .A(n8522), .B(n8521), .ZN(n8529)
         );
  OAI211_X1 U10098 ( .C1(n8525), .C2(n8524), .A(n8523), .B(n10264), .ZN(n8527)
         );
  NAND2_X1 U10099 ( .A1(n8527), .A2(n8526), .ZN(n9061) );
  NAND2_X1 U10100 ( .A1(n9061), .A2(n10299), .ZN(n8528) );
  OAI211_X1 U10101 ( .C1(n9065), .C2(n8639), .A(n8529), .B(n8528), .ZN(
        P2_U3271) );
  XNOR2_X1 U10102 ( .A(n8530), .B(n8537), .ZN(n9070) );
  AOI21_X1 U10103 ( .B1(n9066), .B2(n8549), .A(n8531), .ZN(n9067) );
  INV_X1 U10104 ( .A(n8532), .ZN(n8533) );
  AOI22_X1 U10105 ( .A1(n10308), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8533), 
        .B2(n10245), .ZN(n8534) );
  OAI21_X1 U10106 ( .B1(n8535), .B2(n8627), .A(n8534), .ZN(n8544) );
  AOI21_X1 U10107 ( .B1(n8536), .B2(n8537), .A(n10281), .ZN(n8542) );
  OAI22_X1 U10108 ( .A1(n8539), .A2(n10284), .B1(n8538), .B2(n10286), .ZN(
        n8540) );
  AOI21_X1 U10109 ( .B1(n8542), .B2(n8541), .A(n8540), .ZN(n9069) );
  NOR2_X1 U10110 ( .A1(n9069), .A2(n10308), .ZN(n8543) );
  AOI211_X1 U10111 ( .C1(n9067), .C2(n8637), .A(n8544), .B(n8543), .ZN(n8545)
         );
  OAI21_X1 U10112 ( .B1(n9070), .B2(n8639), .A(n8545), .ZN(P2_U3272) );
  OAI21_X1 U10113 ( .B1(n8548), .B2(n8547), .A(n8546), .ZN(n9075) );
  INV_X1 U10114 ( .A(n8549), .ZN(n8550) );
  AOI21_X1 U10115 ( .B1(n9071), .B2(n8563), .A(n8550), .ZN(n9072) );
  NOR2_X1 U10116 ( .A1(n4728), .A2(n8627), .ZN(n8554) );
  INV_X1 U10117 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8552) );
  OAI22_X1 U10118 ( .A1(n10299), .A2(n8552), .B1(n8551), .B2(n10297), .ZN(
        n8553) );
  AOI211_X1 U10119 ( .C1(n9072), .C2(n8637), .A(n8554), .B(n8553), .ZN(n8561)
         );
  OAI21_X1 U10120 ( .B1(n8557), .B2(n8556), .A(n8555), .ZN(n8559) );
  AOI222_X1 U10121 ( .A1(n10264), .A2(n8559), .B1(n8558), .B2(n10261), .C1(
        n8587), .C2(n10259), .ZN(n9074) );
  OR2_X1 U10122 ( .A1(n9074), .A2(n10308), .ZN(n8560) );
  OAI211_X1 U10123 ( .C1(n9075), .C2(n8639), .A(n8561), .B(n8560), .ZN(
        P2_U3273) );
  XNOR2_X1 U10124 ( .A(n8562), .B(n8569), .ZN(n9080) );
  INV_X1 U10125 ( .A(n8563), .ZN(n8564) );
  AOI21_X1 U10126 ( .B1(n9076), .B2(n4732), .A(n8564), .ZN(n9077) );
  AOI22_X1 U10127 ( .A1(n10308), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8565), 
        .B2(n10245), .ZN(n8566) );
  OAI21_X1 U10128 ( .B1(n8567), .B2(n8627), .A(n8566), .ZN(n8576) );
  OAI211_X1 U10129 ( .C1(n8570), .C2(n8569), .A(n8568), .B(n10264), .ZN(n8574)
         );
  AOI22_X1 U10130 ( .A1(n8572), .A2(n10261), .B1(n8571), .B2(n10259), .ZN(
        n8573) );
  AND2_X1 U10131 ( .A1(n8574), .A2(n8573), .ZN(n9079) );
  NOR2_X1 U10132 ( .A1(n9079), .A2(n10308), .ZN(n8575) );
  AOI211_X1 U10133 ( .C1(n9077), .C2(n8637), .A(n8576), .B(n8575), .ZN(n8577)
         );
  OAI21_X1 U10134 ( .B1(n9080), .B2(n8639), .A(n8577), .ZN(P2_U3274) );
  XNOR2_X1 U10135 ( .A(n8579), .B(n8578), .ZN(n9085) );
  AOI21_X1 U10136 ( .B1(n9081), .B2(n8600), .A(n8580), .ZN(n9082) );
  AOI22_X1 U10137 ( .A1(n10308), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8581), 
        .B2(n10245), .ZN(n8582) );
  OAI21_X1 U10138 ( .B1(n8583), .B2(n8627), .A(n8582), .ZN(n8590) );
  OAI21_X1 U10139 ( .B1(n8585), .B2(n5549), .A(n8584), .ZN(n8588) );
  AOI222_X1 U10140 ( .A1(n10264), .A2(n8588), .B1(n8587), .B2(n10261), .C1(
        n8586), .C2(n10259), .ZN(n9084) );
  NOR2_X1 U10141 ( .A1(n9084), .A2(n10308), .ZN(n8589) );
  AOI211_X1 U10142 ( .C1(n9082), .C2(n8637), .A(n8590), .B(n8589), .ZN(n8591)
         );
  OAI21_X1 U10143 ( .B1(n9085), .B2(n8639), .A(n8591), .ZN(P2_U3275) );
  AOI21_X1 U10144 ( .B1(n8592), .B2(n8598), .A(n10281), .ZN(n8597) );
  OAI22_X1 U10145 ( .A1(n8594), .A2(n10286), .B1(n8593), .B2(n10284), .ZN(
        n8595) );
  AOI21_X1 U10146 ( .B1(n8597), .B2(n8596), .A(n8595), .ZN(n9091) );
  OR2_X1 U10147 ( .A1(n8599), .A2(n8598), .ZN(n9087) );
  NAND3_X1 U10148 ( .A1(n9087), .A2(n9086), .A3(n10306), .ZN(n8608) );
  INV_X1 U10149 ( .A(n8600), .ZN(n8601) );
  AOI21_X1 U10150 ( .B1(n9088), .B2(n8602), .A(n8601), .ZN(n9089) );
  AOI22_X1 U10151 ( .A1(n10308), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8603), 
        .B2(n10245), .ZN(n8604) );
  OAI21_X1 U10152 ( .B1(n8605), .B2(n8627), .A(n8604), .ZN(n8606) );
  AOI21_X1 U10153 ( .B1(n9089), .B2(n8637), .A(n8606), .ZN(n8607) );
  OAI211_X1 U10154 ( .C1(n10308), .C2(n9091), .A(n8608), .B(n8607), .ZN(
        P2_U3276) );
  XNOR2_X1 U10155 ( .A(n8610), .B(n8609), .ZN(n9097) );
  AOI211_X1 U10156 ( .C1(n9094), .C2(n8623), .A(n10402), .B(n8611), .ZN(n9093)
         );
  AOI22_X1 U10157 ( .A1(n10308), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8612), 
        .B2(n10245), .ZN(n8613) );
  OAI21_X1 U10158 ( .B1(n8614), .B2(n8627), .A(n8613), .ZN(n8620) );
  OAI21_X1 U10159 ( .B1(n8616), .B2(n5523), .A(n8615), .ZN(n8618) );
  AOI21_X1 U10160 ( .B1(n8618), .B2(n10264), .A(n8617), .ZN(n9096) );
  NOR2_X1 U10161 ( .A1(n9096), .A2(n10308), .ZN(n8619) );
  AOI211_X1 U10162 ( .C1(n9093), .C2(n10250), .A(n8620), .B(n8619), .ZN(n8621)
         );
  OAI21_X1 U10163 ( .B1(n9097), .B2(n8639), .A(n8621), .ZN(P2_U3277) );
  XNOR2_X1 U10164 ( .A(n8622), .B(n8630), .ZN(n9102) );
  AOI21_X1 U10165 ( .B1(n9098), .B2(n8624), .A(n4733), .ZN(n9099) );
  AOI22_X1 U10166 ( .A1(n10308), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8625), 
        .B2(n10245), .ZN(n8626) );
  OAI21_X1 U10167 ( .B1(n8628), .B2(n8627), .A(n8626), .ZN(n8636) );
  OAI211_X1 U10168 ( .C1(n8631), .C2(n8630), .A(n8629), .B(n10264), .ZN(n8634)
         );
  AOI22_X1 U10169 ( .A1(n10259), .A2(n8647), .B1(n8632), .B2(n10261), .ZN(
        n8633) );
  AND2_X1 U10170 ( .A1(n8634), .A2(n8633), .ZN(n9101) );
  NOR2_X1 U10171 ( .A1(n9101), .A2(n10308), .ZN(n8635) );
  AOI211_X1 U10172 ( .C1(n9099), .C2(n8637), .A(n8636), .B(n8635), .ZN(n8638)
         );
  OAI21_X1 U10173 ( .B1(n9102), .B2(n8639), .A(n8638), .ZN(P2_U3278) );
  INV_X1 U10174 ( .A(n8640), .ZN(n8641) );
  AOI21_X1 U10175 ( .B1(n8643), .B2(n8642), .A(n8641), .ZN(n8651) );
  XNOR2_X1 U10176 ( .A(n8645), .B(n8644), .ZN(n10020) );
  NAND2_X1 U10177 ( .A1(n10020), .A2(n8646), .ZN(n8650) );
  AOI22_X1 U10178 ( .A1(n10259), .A2(n8648), .B1(n8647), .B2(n10261), .ZN(
        n8649) );
  OAI211_X1 U10179 ( .C1(n10281), .C2(n8651), .A(n8650), .B(n8649), .ZN(n10018) );
  INV_X1 U10180 ( .A(n10018), .ZN(n8660) );
  AND2_X1 U10181 ( .A1(n8652), .A2(n10015), .ZN(n8653) );
  OR2_X1 U10182 ( .A1(n8654), .A2(n8653), .ZN(n10017) );
  AOI22_X1 U10183 ( .A1(n10308), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8655), 
        .B2(n10245), .ZN(n8657) );
  NAND2_X1 U10184 ( .A1(n10015), .A2(n10302), .ZN(n8656) );
  OAI211_X1 U10185 ( .C1(n10017), .C2(n10273), .A(n8657), .B(n8656), .ZN(n8658) );
  AOI21_X1 U10186 ( .B1(n10020), .B2(n10251), .A(n8658), .ZN(n8659) );
  OAI21_X1 U10187 ( .B1(n8660), .B2(n10308), .A(n8659), .ZN(P2_U3280) );
  OAI22_X1 U10188 ( .A1(SI_18_), .A2(keyinput28), .B1(P1_REG0_REG_7__SCAN_IN), 
        .B2(keyinput67), .ZN(n8661) );
  AOI221_X1 U10189 ( .B1(SI_18_), .B2(keyinput28), .C1(keyinput67), .C2(
        P1_REG0_REG_7__SCAN_IN), .A(n8661), .ZN(n8668) );
  OAI22_X1 U10190 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(keyinput105), .B1(
        P1_REG1_REG_18__SCAN_IN), .B2(keyinput8), .ZN(n8662) );
  AOI221_X1 U10191 ( .B1(P1_REG3_REG_14__SCAN_IN), .B2(keyinput105), .C1(
        keyinput8), .C2(P1_REG1_REG_18__SCAN_IN), .A(n8662), .ZN(n8667) );
  OAI22_X1 U10192 ( .A1(P1_D_REG_30__SCAN_IN), .A2(keyinput56), .B1(
        P2_D_REG_4__SCAN_IN), .B2(keyinput5), .ZN(n8663) );
  AOI221_X1 U10193 ( .B1(P1_D_REG_30__SCAN_IN), .B2(keyinput56), .C1(keyinput5), .C2(P2_D_REG_4__SCAN_IN), .A(n8663), .ZN(n8666) );
  OAI22_X1 U10194 ( .A1(SI_27_), .A2(keyinput85), .B1(keyinput24), .B2(
        P1_ADDR_REG_2__SCAN_IN), .ZN(n8664) );
  AOI221_X1 U10195 ( .B1(SI_27_), .B2(keyinput85), .C1(P1_ADDR_REG_2__SCAN_IN), 
        .C2(keyinput24), .A(n8664), .ZN(n8665) );
  NAND4_X1 U10196 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8665), .ZN(n8696)
         );
  OAI22_X1 U10197 ( .A1(P1_D_REG_26__SCAN_IN), .A2(keyinput20), .B1(keyinput14), .B2(P2_REG0_REG_12__SCAN_IN), .ZN(n8669) );
  AOI221_X1 U10198 ( .B1(P1_D_REG_26__SCAN_IN), .B2(keyinput20), .C1(
        P2_REG0_REG_12__SCAN_IN), .C2(keyinput14), .A(n8669), .ZN(n8676) );
  OAI22_X1 U10199 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(keyinput61), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput36), .ZN(n8670) );
  AOI221_X1 U10200 ( .B1(P1_DATAO_REG_10__SCAN_IN), .B2(keyinput61), .C1(
        keyinput36), .C2(P2_REG3_REG_4__SCAN_IN), .A(n8670), .ZN(n8675) );
  OAI22_X1 U10201 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput99), .B1(
        P2_D_REG_3__SCAN_IN), .B2(keyinput74), .ZN(n8671) );
  AOI221_X1 U10202 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput99), .C1(
        keyinput74), .C2(P2_D_REG_3__SCAN_IN), .A(n8671), .ZN(n8674) );
  OAI22_X1 U10203 ( .A1(P1_REG0_REG_14__SCAN_IN), .A2(keyinput17), .B1(
        keyinput94), .B2(P2_D_REG_19__SCAN_IN), .ZN(n8672) );
  AOI221_X1 U10204 ( .B1(P1_REG0_REG_14__SCAN_IN), .B2(keyinput17), .C1(
        P2_D_REG_19__SCAN_IN), .C2(keyinput94), .A(n8672), .ZN(n8673) );
  NAND4_X1 U10205 ( .A1(n8676), .A2(n8675), .A3(n8674), .A4(n8673), .ZN(n8695)
         );
  OAI22_X1 U10206 ( .A1(P1_D_REG_21__SCAN_IN), .A2(keyinput59), .B1(keyinput30), .B2(P2_REG2_REG_20__SCAN_IN), .ZN(n8677) );
  AOI221_X1 U10207 ( .B1(P1_D_REG_21__SCAN_IN), .B2(keyinput59), .C1(
        P2_REG2_REG_20__SCAN_IN), .C2(keyinput30), .A(n8677), .ZN(n8684) );
  OAI22_X1 U10208 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput101), .B1(keyinput75), .B2(P1_REG3_REG_25__SCAN_IN), .ZN(n8678) );
  AOI221_X1 U10209 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput101), .C1(
        P1_REG3_REG_25__SCAN_IN), .C2(keyinput75), .A(n8678), .ZN(n8683) );
  OAI22_X1 U10210 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput41), .B1(
        P2_REG1_REG_14__SCAN_IN), .B2(keyinput19), .ZN(n8679) );
  AOI221_X1 U10211 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput41), .C1(
        keyinput19), .C2(P2_REG1_REG_14__SCAN_IN), .A(n8679), .ZN(n8682) );
  OAI22_X1 U10212 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput106), .B1(
        P1_REG0_REG_24__SCAN_IN), .B2(keyinput97), .ZN(n8680) );
  AOI221_X1 U10213 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput106), .C1(
        keyinput97), .C2(P1_REG0_REG_24__SCAN_IN), .A(n8680), .ZN(n8681) );
  NAND4_X1 U10214 ( .A1(n8684), .A2(n8683), .A3(n8682), .A4(n8681), .ZN(n8694)
         );
  OAI22_X1 U10215 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput98), .B1(
        keyinput57), .B2(P1_IR_REG_30__SCAN_IN), .ZN(n8685) );
  AOI221_X1 U10216 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput98), .C1(
        P1_IR_REG_30__SCAN_IN), .C2(keyinput57), .A(n8685), .ZN(n8692) );
  OAI22_X1 U10217 ( .A1(P2_REG1_REG_21__SCAN_IN), .A2(keyinput1), .B1(
        keyinput6), .B2(P2_REG1_REG_15__SCAN_IN), .ZN(n8686) );
  AOI221_X1 U10218 ( .B1(P2_REG1_REG_21__SCAN_IN), .B2(keyinput1), .C1(
        P2_REG1_REG_15__SCAN_IN), .C2(keyinput6), .A(n8686), .ZN(n8691) );
  OAI22_X1 U10219 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput116), .B1(
        keyinput86), .B2(P1_REG1_REG_27__SCAN_IN), .ZN(n8687) );
  AOI221_X1 U10220 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput116), .C1(
        P1_REG1_REG_27__SCAN_IN), .C2(keyinput86), .A(n8687), .ZN(n8690) );
  OAI22_X1 U10221 ( .A1(P1_REG0_REG_0__SCAN_IN), .A2(keyinput39), .B1(
        keyinput60), .B2(P2_IR_REG_0__SCAN_IN), .ZN(n8688) );
  AOI221_X1 U10222 ( .B1(P1_REG0_REG_0__SCAN_IN), .B2(keyinput39), .C1(
        P2_IR_REG_0__SCAN_IN), .C2(keyinput60), .A(n8688), .ZN(n8689) );
  NAND4_X1 U10223 ( .A1(n8692), .A2(n8691), .A3(n8690), .A4(n8689), .ZN(n8693)
         );
  NOR4_X1 U10224 ( .A1(n8696), .A2(n8695), .A3(n8694), .A4(n8693), .ZN(n9003)
         );
  AOI22_X1 U10225 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput238), .B1(
        P1_REG0_REG_7__SCAN_IN), .B2(keyinput195), .ZN(n8697) );
  OAI221_X1 U10226 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput238), .C1(
        P1_REG0_REG_7__SCAN_IN), .C2(keyinput195), .A(n8697), .ZN(n8704) );
  AOI22_X1 U10227 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(keyinput134), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(keyinput217), .ZN(n8698) );
  OAI221_X1 U10228 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(keyinput134), .C1(
        P1_DATAO_REG_2__SCAN_IN), .C2(keyinput217), .A(n8698), .ZN(n8703) );
  AOI22_X1 U10229 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(keyinput198), .B1(
        P2_REG0_REG_5__SCAN_IN), .B2(keyinput154), .ZN(n8699) );
  OAI221_X1 U10230 ( .B1(P1_DATAO_REG_29__SCAN_IN), .B2(keyinput198), .C1(
        P2_REG0_REG_5__SCAN_IN), .C2(keyinput154), .A(n8699), .ZN(n8702) );
  AOI22_X1 U10231 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(keyinput201), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput164), .ZN(n8700) );
  OAI221_X1 U10232 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(keyinput201), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput164), .A(n8700), .ZN(n8701) );
  NOR4_X1 U10233 ( .A1(n8704), .A2(n8703), .A3(n8702), .A4(n8701), .ZN(n8732)
         );
  AOI22_X1 U10234 ( .A1(P2_REG0_REG_19__SCAN_IN), .A2(keyinput245), .B1(
        P2_D_REG_21__SCAN_IN), .B2(keyinput146), .ZN(n8705) );
  OAI221_X1 U10235 ( .B1(P2_REG0_REG_19__SCAN_IN), .B2(keyinput245), .C1(
        P2_D_REG_21__SCAN_IN), .C2(keyinput146), .A(n8705), .ZN(n8712) );
  AOI22_X1 U10236 ( .A1(P1_D_REG_16__SCAN_IN), .A2(keyinput191), .B1(
        P1_D_REG_26__SCAN_IN), .B2(keyinput148), .ZN(n8706) );
  OAI221_X1 U10237 ( .B1(P1_D_REG_16__SCAN_IN), .B2(keyinput191), .C1(
        P1_D_REG_26__SCAN_IN), .C2(keyinput148), .A(n8706), .ZN(n8711) );
  AOI22_X1 U10238 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(keyinput232), .B1(
        P2_REG2_REG_20__SCAN_IN), .B2(keyinput158), .ZN(n8707) );
  OAI221_X1 U10239 ( .B1(P2_REG0_REG_22__SCAN_IN), .B2(keyinput232), .C1(
        P2_REG2_REG_20__SCAN_IN), .C2(keyinput158), .A(n8707), .ZN(n8710) );
  AOI22_X1 U10240 ( .A1(P1_REG0_REG_5__SCAN_IN), .A2(keyinput160), .B1(
        P1_REG0_REG_14__SCAN_IN), .B2(keyinput145), .ZN(n8708) );
  OAI221_X1 U10241 ( .B1(P1_REG0_REG_5__SCAN_IN), .B2(keyinput160), .C1(
        P1_REG0_REG_14__SCAN_IN), .C2(keyinput145), .A(n8708), .ZN(n8709) );
  NOR4_X1 U10242 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), .ZN(n8731)
         );
  AOI22_X1 U10243 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(keyinput209), .B1(
        P1_REG2_REG_3__SCAN_IN), .B2(keyinput207), .ZN(n8713) );
  OAI221_X1 U10244 ( .B1(P1_REG1_REG_30__SCAN_IN), .B2(keyinput209), .C1(
        P1_REG2_REG_3__SCAN_IN), .C2(keyinput207), .A(n8713), .ZN(n8720) );
  AOI22_X1 U10245 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(keyinput194), .B1(
        P1_REG0_REG_9__SCAN_IN), .B2(keyinput177), .ZN(n8714) );
  OAI221_X1 U10246 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(keyinput194), .C1(
        P1_REG0_REG_9__SCAN_IN), .C2(keyinput177), .A(n8714), .ZN(n8719) );
  AOI22_X1 U10247 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(keyinput200), .B1(
        P1_REG0_REG_26__SCAN_IN), .B2(keyinput180), .ZN(n8715) );
  OAI221_X1 U10248 ( .B1(P1_REG1_REG_24__SCAN_IN), .B2(keyinput200), .C1(
        P1_REG0_REG_26__SCAN_IN), .C2(keyinput180), .A(n8715), .ZN(n8718) );
  AOI22_X1 U10249 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput203), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(keyinput228), .ZN(n8716) );
  OAI221_X1 U10250 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput203), .C1(
        P1_DATAO_REG_18__SCAN_IN), .C2(keyinput228), .A(n8716), .ZN(n8717) );
  NOR4_X1 U10251 ( .A1(n8720), .A2(n8719), .A3(n8718), .A4(n8717), .ZN(n8730)
         );
  AOI22_X1 U10252 ( .A1(P2_REG0_REG_23__SCAN_IN), .A2(keyinput212), .B1(SI_27_), .B2(keyinput213), .ZN(n8721) );
  OAI221_X1 U10253 ( .B1(P2_REG0_REG_23__SCAN_IN), .B2(keyinput212), .C1(
        SI_27_), .C2(keyinput213), .A(n8721), .ZN(n8728) );
  AOI22_X1 U10254 ( .A1(P2_D_REG_19__SCAN_IN), .A2(keyinput222), .B1(
        P1_REG2_REG_26__SCAN_IN), .B2(keyinput205), .ZN(n8722) );
  OAI221_X1 U10255 ( .B1(P2_D_REG_19__SCAN_IN), .B2(keyinput222), .C1(
        P1_REG2_REG_26__SCAN_IN), .C2(keyinput205), .A(n8722), .ZN(n8727) );
  AOI22_X1 U10256 ( .A1(P2_REG0_REG_12__SCAN_IN), .A2(keyinput142), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput252), .ZN(n8723) );
  OAI221_X1 U10257 ( .B1(P2_REG0_REG_12__SCAN_IN), .B2(keyinput142), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput252), .A(n8723), .ZN(n8726) );
  AOI22_X1 U10258 ( .A1(P1_REG0_REG_23__SCAN_IN), .A2(keyinput130), .B1(SI_18_), .B2(keyinput156), .ZN(n8724) );
  OAI221_X1 U10259 ( .B1(P1_REG0_REG_23__SCAN_IN), .B2(keyinput130), .C1(
        SI_18_), .C2(keyinput156), .A(n8724), .ZN(n8725) );
  NOR4_X1 U10260 ( .A1(n8728), .A2(n8727), .A3(n8726), .A4(n8725), .ZN(n8729)
         );
  NAND4_X1 U10261 ( .A1(n8732), .A2(n8731), .A3(n8730), .A4(n8729), .ZN(n8861)
         );
  AOI22_X1 U10262 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(keyinput233), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(keyinput151), .ZN(n8733) );
  OAI221_X1 U10263 ( .B1(P1_REG3_REG_14__SCAN_IN), .B2(keyinput233), .C1(
        P1_DATAO_REG_24__SCAN_IN), .C2(keyinput151), .A(n8733), .ZN(n8740) );
  AOI22_X1 U10264 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(keyinput144), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(keyinput255), .ZN(n8734) );
  OAI221_X1 U10265 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(keyinput144), .C1(
        P1_DATAO_REG_0__SCAN_IN), .C2(keyinput255), .A(n8734), .ZN(n8739) );
  AOI22_X1 U10266 ( .A1(P2_D_REG_16__SCAN_IN), .A2(keyinput192), .B1(
        P1_REG1_REG_12__SCAN_IN), .B2(keyinput236), .ZN(n8735) );
  OAI221_X1 U10267 ( .B1(P2_D_REG_16__SCAN_IN), .B2(keyinput192), .C1(
        P1_REG1_REG_12__SCAN_IN), .C2(keyinput236), .A(n8735), .ZN(n8738) );
  AOI22_X1 U10268 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(keyinput137), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(keyinput239), .ZN(n8736) );
  OAI221_X1 U10269 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(keyinput137), .C1(
        P1_ADDR_REG_17__SCAN_IN), .C2(keyinput239), .A(n8736), .ZN(n8737) );
  NOR4_X1 U10270 ( .A1(n8740), .A2(n8739), .A3(n8738), .A4(n8737), .ZN(n8768)
         );
  AOI22_X1 U10271 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput162), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput131), .ZN(n8741) );
  OAI221_X1 U10272 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput162), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput131), .A(n8741), .ZN(n8748) );
  AOI22_X1 U10273 ( .A1(P2_D_REG_3__SCAN_IN), .A2(keyinput202), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(keyinput234), .ZN(n8742) );
  OAI221_X1 U10274 ( .B1(P2_D_REG_3__SCAN_IN), .B2(keyinput202), .C1(
        P1_REG3_REG_3__SCAN_IN), .C2(keyinput234), .A(n8742), .ZN(n8747) );
  AOI22_X1 U10275 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput139), .B1(
        P1_REG1_REG_20__SCAN_IN), .B2(keyinput150), .ZN(n8743) );
  OAI221_X1 U10276 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput139), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput150), .A(n8743), .ZN(n8746) );
  AOI22_X1 U10277 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(keyinput208), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput149), .ZN(n8744) );
  OAI221_X1 U10278 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(keyinput208), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput149), .A(n8744), .ZN(n8745) );
  NOR4_X1 U10279 ( .A1(n8748), .A2(n8747), .A3(n8746), .A4(n8745), .ZN(n8767)
         );
  AOI22_X1 U10280 ( .A1(P2_REG0_REG_20__SCAN_IN), .A2(keyinput253), .B1(
        P1_REG0_REG_6__SCAN_IN), .B2(keyinput230), .ZN(n8749) );
  OAI221_X1 U10281 ( .B1(P2_REG0_REG_20__SCAN_IN), .B2(keyinput253), .C1(
        P1_REG0_REG_6__SCAN_IN), .C2(keyinput230), .A(n8749), .ZN(n8756) );
  AOI22_X1 U10282 ( .A1(P2_REG1_REG_26__SCAN_IN), .A2(keyinput175), .B1(
        P2_D_REG_27__SCAN_IN), .B2(keyinput242), .ZN(n8750) );
  OAI221_X1 U10283 ( .B1(P2_REG1_REG_26__SCAN_IN), .B2(keyinput175), .C1(
        P2_D_REG_27__SCAN_IN), .C2(keyinput242), .A(n8750), .ZN(n8755) );
  AOI22_X1 U10284 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(keyinput214), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(keyinput251), .ZN(n8751) );
  OAI221_X1 U10285 ( .B1(P1_REG1_REG_27__SCAN_IN), .B2(keyinput214), .C1(
        P1_DATAO_REG_3__SCAN_IN), .C2(keyinput251), .A(n8751), .ZN(n8754) );
  AOI22_X1 U10286 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(keyinput249), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(keyinput189), .ZN(n8752) );
  OAI221_X1 U10287 ( .B1(P2_REG2_REG_27__SCAN_IN), .B2(keyinput249), .C1(
        P1_DATAO_REG_10__SCAN_IN), .C2(keyinput189), .A(n8752), .ZN(n8753) );
  NOR4_X1 U10288 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), .ZN(n8766)
         );
  AOI22_X1 U10289 ( .A1(P2_REG0_REG_15__SCAN_IN), .A2(keyinput247), .B1(
        P2_IR_REG_4__SCAN_IN), .B2(keyinput178), .ZN(n8757) );
  OAI221_X1 U10290 ( .B1(P2_REG0_REG_15__SCAN_IN), .B2(keyinput247), .C1(
        P2_IR_REG_4__SCAN_IN), .C2(keyinput178), .A(n8757), .ZN(n8764) );
  AOI22_X1 U10291 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(keyinput216), .B1(
        P2_REG1_REG_30__SCAN_IN), .B2(keyinput193), .ZN(n8758) );
  OAI221_X1 U10292 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(keyinput216), .C1(
        P2_REG1_REG_30__SCAN_IN), .C2(keyinput193), .A(n8758), .ZN(n8763) );
  AOI22_X1 U10293 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(keyinput188), .B1(
        P2_IR_REG_16__SCAN_IN), .B2(keyinput211), .ZN(n8759) );
  OAI221_X1 U10294 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(keyinput188), .C1(
        P2_IR_REG_16__SCAN_IN), .C2(keyinput211), .A(n8759), .ZN(n8762) );
  AOI22_X1 U10295 ( .A1(P1_REG2_REG_31__SCAN_IN), .A2(keyinput240), .B1(SI_21_), .B2(keyinput171), .ZN(n8760) );
  OAI221_X1 U10296 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(keyinput240), .C1(
        SI_21_), .C2(keyinput171), .A(n8760), .ZN(n8761) );
  NOR4_X1 U10297 ( .A1(n8764), .A2(n8763), .A3(n8762), .A4(n8761), .ZN(n8765)
         );
  NAND4_X1 U10298 ( .A1(n8768), .A2(n8767), .A3(n8766), .A4(n8765), .ZN(n8860)
         );
  AOI22_X1 U10299 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(keyinput155), .B1(
        P2_D_REG_23__SCAN_IN), .B2(keyinput210), .ZN(n8769) );
  OAI221_X1 U10300 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(keyinput155), .C1(
        P2_D_REG_23__SCAN_IN), .C2(keyinput210), .A(n8769), .ZN(n8778) );
  AOI22_X1 U10301 ( .A1(n7950), .A2(keyinput161), .B1(keyinput140), .B2(n8771), 
        .ZN(n8770) );
  OAI221_X1 U10302 ( .B1(n7950), .B2(keyinput161), .C1(n8771), .C2(keyinput140), .A(n8770), .ZN(n8777) );
  INV_X1 U10303 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U10304 ( .A1(n7443), .A2(keyinput243), .B1(n10163), .B2(keyinput187), .ZN(n8772) );
  OAI221_X1 U10305 ( .B1(n7443), .B2(keyinput243), .C1(n10163), .C2(
        keyinput187), .A(n8772), .ZN(n8776) );
  INV_X1 U10306 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8774) );
  AOI22_X1 U10307 ( .A1(n5269), .A2(keyinput172), .B1(n8774), .B2(keyinput185), 
        .ZN(n8773) );
  OAI221_X1 U10308 ( .B1(n5269), .B2(keyinput172), .C1(n8774), .C2(keyinput185), .A(n8773), .ZN(n8775) );
  NOR4_X1 U10309 ( .A1(n8778), .A2(n8777), .A3(n8776), .A4(n8775), .ZN(n8814)
         );
  INV_X1 U10310 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U10311 ( .A1(n10162), .A2(keyinput159), .B1(keyinput167), .B2(n6192), .ZN(n8779) );
  OAI221_X1 U10312 ( .B1(n10162), .B2(keyinput159), .C1(n6192), .C2(
        keyinput167), .A(n8779), .ZN(n8789) );
  INV_X1 U10313 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8781) );
  AOI22_X1 U10314 ( .A1(n7559), .A2(keyinput179), .B1(keyinput129), .B2(n8781), 
        .ZN(n8780) );
  OAI221_X1 U10315 ( .B1(n7559), .B2(keyinput179), .C1(n8781), .C2(keyinput129), .A(n8780), .ZN(n8788) );
  INV_X1 U10316 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U10317 ( .A1(n10160), .A2(keyinput184), .B1(keyinput170), .B2(n8783), .ZN(n8782) );
  OAI221_X1 U10318 ( .B1(n10160), .B2(keyinput184), .C1(n8783), .C2(
        keyinput170), .A(n8782), .ZN(n8787) );
  XNOR2_X1 U10319 ( .A(P1_REG0_REG_24__SCAN_IN), .B(keyinput225), .ZN(n8785)
         );
  XNOR2_X1 U10320 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput248), .ZN(n8784) );
  NAND2_X1 U10321 ( .A1(n8785), .A2(n8784), .ZN(n8786) );
  NOR4_X1 U10322 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n8813)
         );
  AOI22_X1 U10323 ( .A1(n10428), .A2(keyinput174), .B1(n8880), .B2(keyinput186), .ZN(n8790) );
  OAI221_X1 U10324 ( .B1(n10428), .B2(keyinput174), .C1(n8880), .C2(
        keyinput186), .A(n8790), .ZN(n8800) );
  INV_X1 U10325 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8793) );
  INV_X1 U10326 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8792) );
  AOI22_X1 U10327 ( .A1(n8793), .A2(keyinput152), .B1(n8792), .B2(keyinput153), 
        .ZN(n8791) );
  OAI221_X1 U10328 ( .B1(n8793), .B2(keyinput152), .C1(n8792), .C2(keyinput153), .A(n8791), .ZN(n8799) );
  AOI22_X1 U10329 ( .A1(n8938), .A2(keyinput181), .B1(n8947), .B2(keyinput221), 
        .ZN(n8794) );
  OAI221_X1 U10330 ( .B1(n8938), .B2(keyinput181), .C1(n8947), .C2(keyinput221), .A(n8794), .ZN(n8798) );
  XNOR2_X1 U10331 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput244), .ZN(n8796) );
  XNOR2_X1 U10332 ( .A(SI_1_), .B(keyinput199), .ZN(n8795) );
  NAND2_X1 U10333 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  NOR4_X1 U10334 ( .A1(n8800), .A2(n8799), .A3(n8798), .A4(n8797), .ZN(n8812)
         );
  INV_X1 U10335 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U10336 ( .A1(n10166), .A2(keyinput229), .B1(keyinput254), .B2(n5452), .ZN(n8801) );
  OAI221_X1 U10337 ( .B1(n10166), .B2(keyinput229), .C1(n5452), .C2(
        keyinput254), .A(n8801), .ZN(n8810) );
  INV_X1 U10338 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10313) );
  INV_X1 U10339 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10008) );
  AOI22_X1 U10340 ( .A1(n10313), .A2(keyinput235), .B1(n10008), .B2(
        keyinput135), .ZN(n8802) );
  OAI221_X1 U10341 ( .B1(n10313), .B2(keyinput235), .C1(n10008), .C2(
        keyinput135), .A(n8802), .ZN(n8809) );
  INV_X1 U10342 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10167) );
  INV_X1 U10343 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8804) );
  AOI22_X1 U10344 ( .A1(n10167), .A2(keyinput246), .B1(keyinput197), .B2(n8804), .ZN(n8803) );
  OAI221_X1 U10345 ( .B1(n10167), .B2(keyinput246), .C1(n8804), .C2(
        keyinput197), .A(n8803), .ZN(n8808) );
  XNOR2_X1 U10346 ( .A(P2_REG0_REG_24__SCAN_IN), .B(keyinput237), .ZN(n8806)
         );
  XNOR2_X1 U10347 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput157), .ZN(n8805) );
  NAND2_X1 U10348 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  NOR4_X1 U10349 ( .A1(n8810), .A2(n8809), .A3(n8808), .A4(n8807), .ZN(n8811)
         );
  NAND4_X1 U10350 ( .A1(n8814), .A2(n8813), .A3(n8812), .A4(n8811), .ZN(n8859)
         );
  INV_X1 U10351 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U10352 ( .A1(n10316), .A2(keyinput132), .B1(n10071), .B2(
        keyinput165), .ZN(n8815) );
  OAI221_X1 U10353 ( .B1(n10316), .B2(keyinput132), .C1(n10071), .C2(
        keyinput165), .A(n8815), .ZN(n8823) );
  AOI22_X1 U10354 ( .A1(n8917), .A2(keyinput182), .B1(n8817), .B2(keyinput226), 
        .ZN(n8816) );
  OAI221_X1 U10355 ( .B1(n8917), .B2(keyinput182), .C1(n8817), .C2(keyinput226), .A(n8816), .ZN(n8822) );
  INV_X1 U10356 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8874) );
  AOI22_X1 U10357 ( .A1(n8874), .A2(keyinput138), .B1(n5457), .B2(keyinput219), 
        .ZN(n8818) );
  OAI221_X1 U10358 ( .B1(n8874), .B2(keyinput138), .C1(n5457), .C2(keyinput219), .A(n8818), .ZN(n8821) );
  INV_X1 U10359 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8949) );
  AOI22_X1 U10360 ( .A1(n5341), .A2(keyinput163), .B1(keyinput141), .B2(n8949), 
        .ZN(n8819) );
  OAI221_X1 U10361 ( .B1(n5341), .B2(keyinput163), .C1(n8949), .C2(keyinput141), .A(n8819), .ZN(n8820) );
  NOR4_X1 U10362 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n8857)
         );
  INV_X1 U10363 ( .A(SI_7_), .ZN(n8826) );
  AOI22_X1 U10364 ( .A1(n8826), .A2(keyinput218), .B1(keyinput220), .B2(n8825), 
        .ZN(n8824) );
  OAI221_X1 U10365 ( .B1(n8826), .B2(keyinput218), .C1(n8825), .C2(keyinput220), .A(n8824), .ZN(n8835) );
  AOI22_X1 U10366 ( .A1(n8828), .A2(keyinput215), .B1(n8865), .B2(keyinput166), 
        .ZN(n8827) );
  OAI221_X1 U10367 ( .B1(n8828), .B2(keyinput215), .C1(n8865), .C2(keyinput166), .A(n8827), .ZN(n8834) );
  AOI22_X1 U10368 ( .A1(n8830), .A2(keyinput169), .B1(n5515), .B2(keyinput224), 
        .ZN(n8829) );
  OAI221_X1 U10369 ( .B1(n8830), .B2(keyinput169), .C1(n5515), .C2(keyinput224), .A(n8829), .ZN(n8833) );
  AOI22_X1 U10370 ( .A1(n4911), .A2(keyinput227), .B1(keyinput241), .B2(n8951), 
        .ZN(n8831) );
  OAI221_X1 U10371 ( .B1(n4911), .B2(keyinput227), .C1(n8951), .C2(keyinput241), .A(n8831), .ZN(n8832) );
  NOR4_X1 U10372 ( .A1(n8835), .A2(n8834), .A3(n8833), .A4(n8832), .ZN(n8856)
         );
  INV_X1 U10373 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U10374 ( .A1(n8929), .A2(keyinput183), .B1(n10317), .B2(keyinput133), .ZN(n8836) );
  OAI221_X1 U10375 ( .B1(n8929), .B2(keyinput183), .C1(n10317), .C2(
        keyinput133), .A(n8836), .ZN(n8844) );
  AOI22_X1 U10376 ( .A1(n8891), .A2(keyinput128), .B1(keyinput136), .B2(n9583), 
        .ZN(n8837) );
  OAI221_X1 U10377 ( .B1(n8891), .B2(keyinput128), .C1(n9583), .C2(keyinput136), .A(n8837), .ZN(n8843) );
  AOI22_X1 U10378 ( .A1(n8941), .A2(keyinput168), .B1(n8915), .B2(keyinput143), 
        .ZN(n8838) );
  OAI221_X1 U10379 ( .B1(n8941), .B2(keyinput168), .C1(n8915), .C2(keyinput143), .A(n8838), .ZN(n8842) );
  XOR2_X1 U10380 ( .A(n10032), .B(keyinput147), .Z(n8840) );
  XNOR2_X1 U10381 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput223), .ZN(n8839) );
  NAND2_X1 U10382 ( .A1(n8840), .A2(n8839), .ZN(n8841) );
  NOR4_X1 U10383 ( .A1(n8844), .A2(n8843), .A3(n8842), .A4(n8841), .ZN(n8855)
         );
  INV_X1 U10384 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U10385 ( .A1(n8864), .A2(keyinput173), .B1(keyinput231), .B2(n10314), .ZN(n8845) );
  OAI221_X1 U10386 ( .B1(n8864), .B2(keyinput173), .C1(n10314), .C2(
        keyinput231), .A(n8845), .ZN(n8853) );
  INV_X1 U10387 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U10388 ( .A1(n10161), .A2(keyinput196), .B1(keyinput204), .B2(n8867), .ZN(n8846) );
  OAI221_X1 U10389 ( .B1(n10161), .B2(keyinput196), .C1(n8867), .C2(
        keyinput204), .A(n8846), .ZN(n8849) );
  INV_X1 U10390 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10318) );
  XNOR2_X1 U10391 ( .A(n10318), .B(keyinput176), .ZN(n8848) );
  XOR2_X1 U10392 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput250), .Z(n8847) );
  OR3_X1 U10393 ( .A1(n8849), .A2(n8848), .A3(n8847), .ZN(n8852) );
  INV_X1 U10394 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8888) );
  INV_X1 U10395 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U10396 ( .A1(n8888), .A2(keyinput206), .B1(n10315), .B2(keyinput190), .ZN(n8850) );
  OAI221_X1 U10397 ( .B1(n8888), .B2(keyinput206), .C1(n10315), .C2(
        keyinput190), .A(n8850), .ZN(n8851) );
  NOR3_X1 U10398 ( .A1(n8853), .A2(n8852), .A3(n8851), .ZN(n8854) );
  NAND4_X1 U10399 ( .A1(n8857), .A2(n8856), .A3(n8855), .A4(n8854), .ZN(n8858)
         );
  NOR4_X1 U10400 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(n8964)
         );
  AOI22_X1 U10401 ( .A1(n6558), .A2(keyinput32), .B1(n10050), .B2(keyinput108), 
        .ZN(n8862) );
  OAI221_X1 U10402 ( .B1(n6558), .B2(keyinput32), .C1(n10050), .C2(keyinput108), .A(n8862), .ZN(n8872) );
  AOI22_X1 U10403 ( .A1(n8865), .A2(keyinput38), .B1(keyinput45), .B2(n8864), 
        .ZN(n8863) );
  OAI221_X1 U10404 ( .B1(n8865), .B2(keyinput38), .C1(n8864), .C2(keyinput45), 
        .A(n8863), .ZN(n8871) );
  AOI22_X1 U10405 ( .A1(n5457), .A2(keyinput91), .B1(n8867), .B2(keyinput76), 
        .ZN(n8866) );
  OAI221_X1 U10406 ( .B1(n5457), .B2(keyinput91), .C1(n8867), .C2(keyinput76), 
        .A(n8866), .ZN(n8870) );
  AOI22_X1 U10407 ( .A1(n10162), .A2(keyinput31), .B1(keyinput112), .B2(n8098), 
        .ZN(n8868) );
  OAI221_X1 U10408 ( .B1(n10162), .B2(keyinput31), .C1(n8098), .C2(keyinput112), .A(n8868), .ZN(n8869) );
  NOR4_X1 U10409 ( .A1(n8872), .A2(n8871), .A3(n8870), .A4(n8869), .ZN(n8913)
         );
  AOI22_X1 U10410 ( .A1(n5515), .A2(keyinput96), .B1(keyinput10), .B2(n8874), 
        .ZN(n8873) );
  OAI221_X1 U10411 ( .B1(n5515), .B2(keyinput96), .C1(n8874), .C2(keyinput10), 
        .A(n8873), .ZN(n8886) );
  INV_X1 U10412 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U10413 ( .A1(n8876), .A2(keyinput123), .B1(keyinput114), .B2(n10311), .ZN(n8875) );
  OAI221_X1 U10414 ( .B1(n8876), .B2(keyinput123), .C1(n10311), .C2(
        keyinput114), .A(n8875), .ZN(n8885) );
  AOI22_X1 U10415 ( .A1(n8879), .A2(keyinput52), .B1(keyinput117), .B2(n8878), 
        .ZN(n8877) );
  OAI221_X1 U10416 ( .B1(n8879), .B2(keyinput52), .C1(n8878), .C2(keyinput117), 
        .A(n8877), .ZN(n8884) );
  XOR2_X1 U10417 ( .A(n8880), .B(keyinput58), .Z(n8882) );
  XNOR2_X1 U10418 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput21), .ZN(n8881) );
  NAND2_X1 U10419 ( .A1(n8882), .A2(n8881), .ZN(n8883) );
  NOR4_X1 U10420 ( .A1(n8886), .A2(n8885), .A3(n8884), .A4(n8883), .ZN(n8912)
         );
  INV_X1 U10421 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U10422 ( .A1(n8888), .A2(keyinput78), .B1(keyinput9), .B2(n10435), 
        .ZN(n8887) );
  OAI221_X1 U10423 ( .B1(n8888), .B2(keyinput78), .C1(n10435), .C2(keyinput9), 
        .A(n8887), .ZN(n8897) );
  AOI22_X1 U10424 ( .A1(n6781), .A2(keyinput102), .B1(keyinput79), .B2(n6465), 
        .ZN(n8889) );
  OAI221_X1 U10425 ( .B1(n6781), .B2(keyinput102), .C1(n6465), .C2(keyinput79), 
        .A(n8889), .ZN(n8896) );
  AOI22_X1 U10426 ( .A1(n8891), .A2(keyinput0), .B1(keyinput121), .B2(n5612), 
        .ZN(n8890) );
  OAI221_X1 U10427 ( .B1(n8891), .B2(keyinput0), .C1(n5612), .C2(keyinput121), 
        .A(n8890), .ZN(n8895) );
  XNOR2_X1 U10428 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput120), .ZN(n8893) );
  XNOR2_X1 U10429 ( .A(SI_21_), .B(keyinput43), .ZN(n8892) );
  NAND2_X1 U10430 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  NOR4_X1 U10431 ( .A1(n8897), .A2(n8896), .A3(n8895), .A4(n8894), .ZN(n8911)
         );
  INV_X1 U10432 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U10433 ( .A1(n8899), .A2(keyinput23), .B1(n10164), .B2(keyinput63), 
        .ZN(n8898) );
  OAI221_X1 U10434 ( .B1(n8899), .B2(keyinput23), .C1(n10164), .C2(keyinput63), 
        .A(n8898), .ZN(n8909) );
  AOI22_X1 U10435 ( .A1(n10315), .A2(keyinput62), .B1(keyinput81), .B2(n8901), 
        .ZN(n8900) );
  OAI221_X1 U10436 ( .B1(n10315), .B2(keyinput62), .C1(n8901), .C2(keyinput81), 
        .A(n8900), .ZN(n8908) );
  AOI22_X1 U10437 ( .A1(n5452), .A2(keyinput126), .B1(n8903), .B2(keyinput22), 
        .ZN(n8902) );
  OAI221_X1 U10438 ( .B1(n5452), .B2(keyinput126), .C1(n8903), .C2(keyinput22), 
        .A(n8902), .ZN(n8907) );
  AOI22_X1 U10439 ( .A1(n8905), .A2(keyinput125), .B1(n6080), .B2(keyinput124), 
        .ZN(n8904) );
  OAI221_X1 U10440 ( .B1(n8905), .B2(keyinput125), .C1(n6080), .C2(keyinput124), .A(n8904), .ZN(n8906) );
  NOR4_X1 U10441 ( .A1(n8909), .A2(n8908), .A3(n8907), .A4(n8906), .ZN(n8910)
         );
  NAND4_X1 U10442 ( .A1(n8913), .A2(n8912), .A3(n8911), .A4(n8910), .ZN(n8963)
         );
  AOI22_X1 U10443 ( .A1(n5269), .A2(keyinput44), .B1(n8915), .B2(keyinput15), 
        .ZN(n8914) );
  OAI221_X1 U10444 ( .B1(n5269), .B2(keyinput44), .C1(n8915), .C2(keyinput15), 
        .A(n8914), .ZN(n8925) );
  AOI22_X1 U10445 ( .A1(n8917), .A2(keyinput54), .B1(n5213), .B2(keyinput110), 
        .ZN(n8916) );
  OAI221_X1 U10446 ( .B1(n8917), .B2(keyinput54), .C1(n5213), .C2(keyinput110), 
        .A(n8916), .ZN(n8924) );
  AOI22_X1 U10447 ( .A1(n7950), .A2(keyinput33), .B1(keyinput104), .B2(n8919), 
        .ZN(n8918) );
  OAI221_X1 U10448 ( .B1(n7950), .B2(keyinput33), .C1(n8919), .C2(keyinput104), 
        .A(n8918), .ZN(n8923) );
  XNOR2_X1 U10449 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput83), .ZN(n8921) );
  XNOR2_X1 U10450 ( .A(P1_REG0_REG_23__SCAN_IN), .B(keyinput2), .ZN(n8920) );
  NAND2_X1 U10451 ( .A1(n8921), .A2(n8920), .ZN(n8922) );
  NOR4_X1 U10452 ( .A1(n8925), .A2(n8924), .A3(n8923), .A4(n8922), .ZN(n8961)
         );
  AOI22_X1 U10453 ( .A1(n9127), .A2(keyinput70), .B1(n7559), .B2(keyinput51), 
        .ZN(n8926) );
  OAI221_X1 U10454 ( .B1(n9127), .B2(keyinput70), .C1(n7559), .C2(keyinput51), 
        .A(n8926), .ZN(n8935) );
  INV_X1 U10455 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U10456 ( .A1(n8520), .A2(keyinput27), .B1(n10312), .B2(keyinput82), 
        .ZN(n8927) );
  OAI221_X1 U10457 ( .B1(n8520), .B2(keyinput27), .C1(n10312), .C2(keyinput82), 
        .A(n8927), .ZN(n8934) );
  AOI22_X1 U10458 ( .A1(n10008), .A2(keyinput7), .B1(keyinput55), .B2(n8929), 
        .ZN(n8928) );
  OAI221_X1 U10459 ( .B1(n10008), .B2(keyinput7), .C1(n8929), .C2(keyinput55), 
        .A(n8928), .ZN(n8933) );
  XNOR2_X1 U10460 ( .A(P2_REG1_REG_18__SCAN_IN), .B(keyinput66), .ZN(n8931) );
  XNOR2_X1 U10461 ( .A(SI_1_), .B(keyinput71), .ZN(n8930) );
  NAND2_X1 U10462 ( .A1(n8931), .A2(n8930), .ZN(n8932) );
  NOR4_X1 U10463 ( .A1(n8935), .A2(n8934), .A3(n8933), .A4(n8932), .ZN(n8960)
         );
  AOI22_X1 U10464 ( .A1(n10313), .A2(keyinput107), .B1(keyinput46), .B2(n10428), .ZN(n8936) );
  OAI221_X1 U10465 ( .B1(n10313), .B2(keyinput107), .C1(n10428), .C2(
        keyinput46), .A(n8936), .ZN(n8945) );
  AOI22_X1 U10466 ( .A1(n8938), .A2(keyinput53), .B1(keyinput80), .B2(n7496), 
        .ZN(n8937) );
  OAI221_X1 U10467 ( .B1(n8938), .B2(keyinput53), .C1(n7496), .C2(keyinput80), 
        .A(n8937), .ZN(n8944) );
  AOI22_X1 U10468 ( .A1(n7733), .A2(keyinput77), .B1(keyinput35), .B2(n5341), 
        .ZN(n8939) );
  OAI221_X1 U10469 ( .B1(n7733), .B2(keyinput77), .C1(n5341), .C2(keyinput35), 
        .A(n8939), .ZN(n8943) );
  AOI22_X1 U10470 ( .A1(n7443), .A2(keyinput115), .B1(n8941), .B2(keyinput40), 
        .ZN(n8940) );
  OAI221_X1 U10471 ( .B1(n7443), .B2(keyinput115), .C1(n8941), .C2(keyinput40), 
        .A(n8940), .ZN(n8942) );
  NOR4_X1 U10472 ( .A1(n8945), .A2(n8944), .A3(n8943), .A4(n8942), .ZN(n8959)
         );
  AOI22_X1 U10473 ( .A1(n5456), .A2(keyinput119), .B1(n8947), .B2(keyinput93), 
        .ZN(n8946) );
  OAI221_X1 U10474 ( .B1(n5456), .B2(keyinput119), .C1(n8947), .C2(keyinput93), 
        .A(n8946), .ZN(n8957) );
  AOI22_X1 U10475 ( .A1(n8949), .A2(keyinput13), .B1(n5601), .B2(keyinput34), 
        .ZN(n8948) );
  OAI221_X1 U10476 ( .B1(n8949), .B2(keyinput13), .C1(n5601), .C2(keyinput34), 
        .A(n8948), .ZN(n8956) );
  AOI22_X1 U10477 ( .A1(n7206), .A2(keyinput111), .B1(n8951), .B2(keyinput113), 
        .ZN(n8950) );
  OAI221_X1 U10478 ( .B1(n7206), .B2(keyinput111), .C1(n8951), .C2(keyinput113), .A(n8950), .ZN(n8955) );
  AOI22_X1 U10479 ( .A1(n10316), .A2(keyinput4), .B1(keyinput84), .B2(n8953), 
        .ZN(n8952) );
  OAI221_X1 U10480 ( .B1(n10316), .B2(keyinput4), .C1(n8953), .C2(keyinput84), 
        .A(n8952), .ZN(n8954) );
  NOR4_X1 U10481 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n8958)
         );
  NAND4_X1 U10482 ( .A1(n8961), .A2(n8960), .A3(n8959), .A4(n8958), .ZN(n8962)
         );
  NOR3_X1 U10483 ( .A1(n8964), .A2(n8963), .A3(n8962), .ZN(n9002) );
  OAI22_X1 U10484 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput95), .B1(
        P1_D_REG_28__SCAN_IN), .B2(keyinput68), .ZN(n8965) );
  AOI221_X1 U10485 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput95), .C1(
        keyinput68), .C2(P1_D_REG_28__SCAN_IN), .A(n8965), .ZN(n8972) );
  OAI22_X1 U10486 ( .A1(SI_20_), .A2(keyinput87), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(keyinput11), .ZN(n8966) );
  AOI221_X1 U10487 ( .B1(SI_20_), .B2(keyinput87), .C1(keyinput11), .C2(
        P2_REG3_REG_0__SCAN_IN), .A(n8966), .ZN(n8971) );
  OAI22_X1 U10488 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput118), .B1(
        keyinput100), .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8967) );
  AOI221_X1 U10489 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput118), .C1(
        P1_DATAO_REG_18__SCAN_IN), .C2(keyinput100), .A(n8967), .ZN(n8970) );
  OAI22_X1 U10490 ( .A1(P1_REG0_REG_21__SCAN_IN), .A2(keyinput69), .B1(
        keyinput25), .B2(P2_REG1_REG_24__SCAN_IN), .ZN(n8968) );
  AOI221_X1 U10491 ( .B1(P1_REG0_REG_21__SCAN_IN), .B2(keyinput69), .C1(
        P2_REG1_REG_24__SCAN_IN), .C2(keyinput25), .A(n8968), .ZN(n8969) );
  NAND4_X1 U10492 ( .A1(n8972), .A2(n8971), .A3(n8970), .A4(n8969), .ZN(n9000)
         );
  OAI22_X1 U10493 ( .A1(P2_D_REG_12__SCAN_IN), .A2(keyinput103), .B1(
        P2_REG1_REG_30__SCAN_IN), .B2(keyinput65), .ZN(n8973) );
  AOI221_X1 U10494 ( .B1(P2_D_REG_12__SCAN_IN), .B2(keyinput103), .C1(
        keyinput65), .C2(P2_REG1_REG_30__SCAN_IN), .A(n8973), .ZN(n8980) );
  OAI22_X1 U10495 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(keyinput16), .B1(
        keyinput109), .B2(P2_REG0_REG_24__SCAN_IN), .ZN(n8974) );
  AOI221_X1 U10496 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(keyinput16), .C1(
        P2_REG0_REG_24__SCAN_IN), .C2(keyinput109), .A(n8974), .ZN(n8979) );
  OAI22_X1 U10497 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput122), .B1(
        keyinput26), .B2(P2_REG0_REG_5__SCAN_IN), .ZN(n8975) );
  AOI221_X1 U10498 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput122), .C1(
        P2_REG0_REG_5__SCAN_IN), .C2(keyinput26), .A(n8975), .ZN(n8978) );
  OAI22_X1 U10499 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput42), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput92), .ZN(n8976) );
  AOI221_X1 U10500 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput42), .C1(
        keyinput92), .C2(P2_REG3_REG_18__SCAN_IN), .A(n8976), .ZN(n8977) );
  NAND4_X1 U10501 ( .A1(n8980), .A2(n8979), .A3(n8978), .A4(n8977), .ZN(n8999)
         );
  OAI22_X1 U10502 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(keyinput89), .B1(
        P2_ADDR_REG_14__SCAN_IN), .B2(keyinput73), .ZN(n8981) );
  AOI221_X1 U10503 ( .B1(P1_DATAO_REG_2__SCAN_IN), .B2(keyinput89), .C1(
        keyinput73), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8981), .ZN(n8988) );
  OAI22_X1 U10504 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput3), .B1(
        P2_D_REG_21__SCAN_IN), .B2(keyinput18), .ZN(n8982) );
  AOI221_X1 U10505 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput3), .C1(
        keyinput18), .C2(P2_D_REG_21__SCAN_IN), .A(n8982), .ZN(n8987) );
  OAI22_X1 U10506 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(keyinput72), .B1(
        keyinput49), .B2(P1_REG0_REG_9__SCAN_IN), .ZN(n8983) );
  AOI221_X1 U10507 ( .B1(P1_REG1_REG_24__SCAN_IN), .B2(keyinput72), .C1(
        P1_REG0_REG_9__SCAN_IN), .C2(keyinput49), .A(n8983), .ZN(n8986) );
  OAI22_X1 U10508 ( .A1(SI_7_), .A2(keyinput90), .B1(keyinput50), .B2(
        P2_IR_REG_4__SCAN_IN), .ZN(n8984) );
  AOI221_X1 U10509 ( .B1(SI_7_), .B2(keyinput90), .C1(P2_IR_REG_4__SCAN_IN), 
        .C2(keyinput50), .A(n8984), .ZN(n8985) );
  NAND4_X1 U10510 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n8998)
         );
  OAI22_X1 U10511 ( .A1(P2_D_REG_2__SCAN_IN), .A2(keyinput48), .B1(
        P2_REG1_REG_26__SCAN_IN), .B2(keyinput47), .ZN(n8989) );
  AOI221_X1 U10512 ( .B1(P2_D_REG_2__SCAN_IN), .B2(keyinput48), .C1(keyinput47), .C2(P2_REG1_REG_26__SCAN_IN), .A(n8989), .ZN(n8996) );
  OAI22_X1 U10513 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput29), .B1(
        P1_REG0_REG_13__SCAN_IN), .B2(keyinput12), .ZN(n8990) );
  AOI221_X1 U10514 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput29), .C1(
        keyinput12), .C2(P1_REG0_REG_13__SCAN_IN), .A(n8990), .ZN(n8995) );
  OAI22_X1 U10515 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput127), .B1(
        P2_D_REG_16__SCAN_IN), .B2(keyinput64), .ZN(n8991) );
  AOI221_X1 U10516 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput127), .C1(
        keyinput64), .C2(P2_D_REG_16__SCAN_IN), .A(n8991), .ZN(n8994) );
  OAI22_X1 U10517 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(keyinput37), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(keyinput88), .ZN(n8992) );
  AOI221_X1 U10518 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(keyinput37), .C1(
        keyinput88), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n8992), .ZN(n8993) );
  NAND4_X1 U10519 ( .A1(n8996), .A2(n8995), .A3(n8994), .A4(n8993), .ZN(n8997)
         );
  NOR4_X1 U10520 ( .A1(n9000), .A2(n8999), .A3(n8998), .A4(n8997), .ZN(n9001)
         );
  NAND3_X1 U10521 ( .A1(n9003), .A2(n9002), .A3(n9001), .ZN(n9021) );
  XNOR2_X1 U10522 ( .A(n9004), .B(n9005), .ZN(n10370) );
  AOI21_X1 U10523 ( .B1(n9006), .B2(n9012), .A(n10402), .ZN(n9007) );
  NAND2_X1 U10524 ( .A1(n9007), .A2(n10246), .ZN(n10369) );
  INV_X1 U10525 ( .A(n9008), .ZN(n9009) );
  OAI22_X1 U10526 ( .A1(n10299), .A2(n9010), .B1(n9009), .B2(n10297), .ZN(
        n9011) );
  AOI21_X1 U10527 ( .B1(n10302), .B2(n9012), .A(n9011), .ZN(n9013) );
  OAI21_X1 U10528 ( .B1(n10304), .B2(n10369), .A(n9013), .ZN(n9019) );
  XNOR2_X1 U10529 ( .A(n9015), .B(n9014), .ZN(n9017) );
  AOI21_X1 U10530 ( .B1(n9017), .B2(n10264), .A(n9016), .ZN(n10373) );
  NOR2_X1 U10531 ( .A1(n10373), .A2(n10308), .ZN(n9018) );
  AOI211_X1 U10532 ( .C1(n10306), .C2(n10370), .A(n9019), .B(n9018), .ZN(n9020) );
  XOR2_X1 U10533 ( .A(n9021), .B(n9020), .Z(P2_U3289) );
  NAND2_X1 U10534 ( .A1(n9022), .A2(n10376), .ZN(n9023) );
  OAI211_X1 U10535 ( .C1(n9024), .C2(n10402), .A(n9023), .B(n9032), .ZN(n9106)
         );
  NAND3_X1 U10536 ( .A1(n9027), .A2(n9026), .A3(n9025), .ZN(n9029) );
  MUX2_X1 U10537 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9106), .S(n10430), .Z(
        P2_U3551) );
  NAND3_X1 U10538 ( .A1(n9031), .A2(n10295), .A3(n9030), .ZN(n9033) );
  OAI211_X1 U10539 ( .C1(n9034), .C2(n10400), .A(n9033), .B(n9032), .ZN(n9107)
         );
  MUX2_X1 U10540 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9107), .S(n10430), .Z(
        P2_U3550) );
  NAND2_X1 U10541 ( .A1(n9036), .A2(n9035), .ZN(n10380) );
  AOI22_X1 U10542 ( .A1(n9038), .A2(n10295), .B1(n10376), .B2(n9037), .ZN(
        n9039) );
  INV_X1 U10543 ( .A(n9042), .ZN(n9047) );
  AOI22_X1 U10544 ( .A1(n9044), .A2(n10295), .B1(n10376), .B2(n9043), .ZN(
        n9045) );
  OAI211_X1 U10545 ( .C1(n9047), .C2(n10327), .A(n9046), .B(n9045), .ZN(n9108)
         );
  MUX2_X1 U10546 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9108), .S(n10430), .Z(
        P2_U3548) );
  INV_X1 U10547 ( .A(n9048), .ZN(n9053) );
  AOI22_X1 U10548 ( .A1(n9050), .A2(n10295), .B1(n10376), .B2(n9049), .ZN(
        n9051) );
  OAI211_X1 U10549 ( .C1(n9053), .C2(n10327), .A(n9052), .B(n9051), .ZN(n9109)
         );
  MUX2_X1 U10550 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9109), .S(n10430), .Z(
        P2_U3547) );
  NAND2_X1 U10551 ( .A1(n9054), .A2(n10407), .ZN(n9060) );
  AOI21_X1 U10552 ( .B1(n9056), .B2(n10376), .A(n9055), .ZN(n9059) );
  NAND4_X1 U10553 ( .A1(n9060), .A2(n9059), .A3(n9058), .A4(n9057), .ZN(n9110)
         );
  MUX2_X1 U10554 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9110), .S(n10430), .Z(
        P2_U3546) );
  AOI211_X1 U10555 ( .C1(n10376), .C2(n9063), .A(n9062), .B(n9061), .ZN(n9064)
         );
  OAI21_X1 U10556 ( .B1(n9065), .B2(n10327), .A(n9064), .ZN(n9111) );
  MUX2_X1 U10557 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9111), .S(n10430), .Z(
        P2_U3545) );
  AOI22_X1 U10558 ( .A1(n9067), .A2(n10295), .B1(n10376), .B2(n9066), .ZN(
        n9068) );
  OAI211_X1 U10559 ( .C1(n9070), .C2(n10327), .A(n9069), .B(n9068), .ZN(n9112)
         );
  MUX2_X1 U10560 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9112), .S(n10430), .Z(
        P2_U3544) );
  AOI22_X1 U10561 ( .A1(n9072), .A2(n10295), .B1(n10376), .B2(n9071), .ZN(
        n9073) );
  OAI211_X1 U10562 ( .C1(n9075), .C2(n10327), .A(n9074), .B(n9073), .ZN(n9113)
         );
  MUX2_X1 U10563 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9113), .S(n10430), .Z(
        P2_U3543) );
  AOI22_X1 U10564 ( .A1(n9077), .A2(n10295), .B1(n10376), .B2(n9076), .ZN(
        n9078) );
  OAI211_X1 U10565 ( .C1(n9080), .C2(n10327), .A(n9079), .B(n9078), .ZN(n9114)
         );
  MUX2_X1 U10566 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9114), .S(n10430), .Z(
        P2_U3542) );
  AOI22_X1 U10567 ( .A1(n9082), .A2(n10295), .B1(n10376), .B2(n9081), .ZN(
        n9083) );
  OAI211_X1 U10568 ( .C1(n9085), .C2(n10327), .A(n9084), .B(n9083), .ZN(n9115)
         );
  MUX2_X1 U10569 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9115), .S(n10430), .Z(
        P2_U3541) );
  NAND3_X1 U10570 ( .A1(n9087), .A2(n9086), .A3(n10407), .ZN(n9092) );
  AOI22_X1 U10571 ( .A1(n9089), .A2(n10295), .B1(n10376), .B2(n9088), .ZN(
        n9090) );
  NAND3_X1 U10572 ( .A1(n9092), .A2(n9091), .A3(n9090), .ZN(n9116) );
  MUX2_X1 U10573 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9116), .S(n10430), .Z(
        P2_U3540) );
  AOI21_X1 U10574 ( .B1(n10376), .B2(n9094), .A(n9093), .ZN(n9095) );
  OAI211_X1 U10575 ( .C1(n9097), .C2(n10327), .A(n9096), .B(n9095), .ZN(n9117)
         );
  MUX2_X1 U10576 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9117), .S(n10430), .Z(
        P2_U3539) );
  AOI22_X1 U10577 ( .A1(n9099), .A2(n10295), .B1(n10376), .B2(n9098), .ZN(
        n9100) );
  OAI211_X1 U10578 ( .C1(n9102), .C2(n10327), .A(n9101), .B(n9100), .ZN(n9118)
         );
  MUX2_X1 U10579 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9118), .S(n10430), .Z(
        P2_U3538) );
  INV_X1 U10580 ( .A(n9103), .ZN(n9104) );
  MUX2_X1 U10581 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9106), .S(n10409), .Z(
        P2_U3519) );
  MUX2_X1 U10582 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9107), .S(n10409), .Z(
        P2_U3518) );
  MUX2_X1 U10583 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9108), .S(n10409), .Z(
        P2_U3516) );
  MUX2_X1 U10584 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9109), .S(n10409), .Z(
        P2_U3515) );
  MUX2_X1 U10585 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9110), .S(n10409), .Z(
        P2_U3514) );
  MUX2_X1 U10586 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9111), .S(n10409), .Z(
        P2_U3513) );
  MUX2_X1 U10587 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9112), .S(n10409), .Z(
        P2_U3512) );
  MUX2_X1 U10588 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9113), .S(n10409), .Z(
        P2_U3511) );
  MUX2_X1 U10589 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9114), .S(n10409), .Z(
        P2_U3510) );
  MUX2_X1 U10590 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9115), .S(n10409), .Z(
        P2_U3509) );
  MUX2_X1 U10591 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9116), .S(n10409), .Z(
        P2_U3508) );
  MUX2_X1 U10592 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9117), .S(n10409), .Z(
        P2_U3507) );
  MUX2_X1 U10593 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9118), .S(n10409), .Z(
        P2_U3505) );
  INV_X1 U10594 ( .A(n8092), .ZN(n9121) );
  NOR4_X1 U10595 ( .A1(n5220), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5479), .A4(
        P2_U3152), .ZN(n9119) );
  AOI21_X1 U10596 ( .B1(n9129), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9119), .ZN(
        n9120) );
  OAI21_X1 U10597 ( .B1(n9121), .B2(n9134), .A(n9120), .ZN(P2_U3327) );
  AOI22_X1 U10598 ( .A1(n9122), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9129), .ZN(n9123) );
  OAI21_X1 U10599 ( .B1(n9124), .B2(n9134), .A(n9123), .ZN(P2_U3328) );
  INV_X1 U10600 ( .A(n9125), .ZN(n9963) );
  OAI222_X1 U10601 ( .A1(n9137), .A2(n9127), .B1(n9134), .B2(n9963), .C1(n9126), .C2(P2_U3152), .ZN(P2_U3329) );
  AOI21_X1 U10602 ( .B1(n9129), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9128), .ZN(
        n9130) );
  OAI21_X1 U10603 ( .B1(n9131), .B2(n9134), .A(n9130), .ZN(P2_U3330) );
  INV_X1 U10604 ( .A(n9132), .ZN(n9966) );
  OAI222_X1 U10605 ( .A1(n9137), .A2(n9135), .B1(n9134), .B2(n9966), .C1(n9133), .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U10606 ( .A(n9136), .ZN(n9970) );
  OAI222_X1 U10607 ( .A1(n9141), .A2(P2_U3152), .B1(n9139), .B2(n9970), .C1(
        n9138), .C2(n9137), .ZN(P2_U3332) );
  MUX2_X1 U10608 ( .A(n9142), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10609 ( .A(n9143), .ZN(n9144) );
  NOR2_X1 U10610 ( .A1(n9145), .A2(n9144), .ZN(n9147) );
  XNOR2_X1 U10611 ( .A(n9147), .B(n9146), .ZN(n9152) );
  NOR2_X1 U10612 ( .A1(n9249), .A2(n9703), .ZN(n9150) );
  AOI22_X1 U10613 ( .A1(n9738), .A2(n9236), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9148) );
  OAI21_X1 U10614 ( .B1(n9710), .B2(n9234), .A(n9148), .ZN(n9149) );
  AOI211_X1 U10615 ( .C1(n9878), .C2(n9251), .A(n9150), .B(n9149), .ZN(n9151)
         );
  OAI21_X1 U10616 ( .B1(n9152), .B2(n9253), .A(n9151), .ZN(P1_U3214) );
  INV_X1 U10617 ( .A(n9900), .ZN(n9769) );
  OAI21_X1 U10618 ( .B1(n9155), .B2(n4706), .A(n9154), .ZN(n9156) );
  OAI21_X1 U10619 ( .B1(n9157), .B2(n4706), .A(n9156), .ZN(n9158) );
  NAND2_X1 U10620 ( .A1(n9158), .A2(n9211), .ZN(n9163) );
  NAND2_X1 U10621 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9601) );
  OAI21_X1 U10622 ( .B1(n9159), .B2(n9234), .A(n9601), .ZN(n9161) );
  NOR2_X1 U10623 ( .A1(n9249), .A2(n9766), .ZN(n9160) );
  AOI211_X1 U10624 ( .C1(n9236), .C2(n9774), .A(n9161), .B(n9160), .ZN(n9162)
         );
  OAI211_X1 U10625 ( .C1(n9769), .C2(n9218), .A(n9163), .B(n9162), .ZN(
        P1_U3217) );
  XOR2_X1 U10626 ( .A(n9165), .B(n9164), .Z(n9170) );
  AOI22_X1 U10627 ( .A1(n9236), .A2(n9773), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9167) );
  NAND2_X1 U10628 ( .A1(n9203), .A2(n9742), .ZN(n9166) );
  OAI211_X1 U10629 ( .C1(n9709), .C2(n9234), .A(n9167), .B(n9166), .ZN(n9168)
         );
  AOI21_X1 U10630 ( .B1(n9889), .B2(n9251), .A(n9168), .ZN(n9169) );
  OAI21_X1 U10631 ( .B1(n9170), .B2(n9253), .A(n9169), .ZN(P1_U3221) );
  XOR2_X1 U10632 ( .A(n9172), .B(n9171), .Z(n9177) );
  NOR2_X1 U10633 ( .A1(n9671), .A2(n9234), .ZN(n9175) );
  AOI22_X1 U10634 ( .A1(n9548), .A2(n9236), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9173) );
  OAI21_X1 U10635 ( .B1(n9249), .B2(n9676), .A(n9173), .ZN(n9174) );
  AOI211_X1 U10636 ( .C1(n9667), .C2(n9251), .A(n9175), .B(n9174), .ZN(n9176)
         );
  OAI21_X1 U10637 ( .B1(n9177), .B2(n9253), .A(n9176), .ZN(P1_U3223) );
  INV_X1 U10638 ( .A(n9178), .ZN(n9182) );
  AOI21_X1 U10639 ( .B1(n9180), .B2(n9242), .A(n9179), .ZN(n9181) );
  OAI21_X1 U10640 ( .B1(n9182), .B2(n9181), .A(n9211), .ZN(n9188) );
  OAI21_X1 U10641 ( .B1(n9784), .B2(n9234), .A(n9183), .ZN(n9186) );
  NOR2_X1 U10642 ( .A1(n9249), .A2(n9184), .ZN(n9185) );
  AOI211_X1 U10643 ( .C1(n9236), .C2(n9552), .A(n9186), .B(n9185), .ZN(n9187)
         );
  OAI211_X1 U10644 ( .C1(n9189), .C2(n9218), .A(n9188), .B(n9187), .ZN(
        P1_U3224) );
  OAI21_X1 U10645 ( .B1(n9192), .B2(n9191), .A(n9190), .ZN(n9193) );
  NAND2_X1 U10646 ( .A1(n9193), .A2(n9211), .ZN(n9198) );
  OAI21_X1 U10647 ( .B1(n9809), .B2(n9234), .A(n9194), .ZN(n9196) );
  NOR2_X1 U10648 ( .A1(n9249), .A2(n9801), .ZN(n9195) );
  AOI211_X1 U10649 ( .C1(n9236), .C2(n9551), .A(n9196), .B(n9195), .ZN(n9197)
         );
  OAI211_X1 U10650 ( .C1(n9800), .C2(n9218), .A(n9198), .B(n9197), .ZN(
        P1_U3226) );
  XOR2_X1 U10651 ( .A(n9200), .B(n9199), .Z(n9207) );
  OAI22_X1 U10652 ( .A1(n9688), .A2(n9245), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9201), .ZN(n9202) );
  AOI21_X1 U10653 ( .B1(n9682), .B2(n9203), .A(n9202), .ZN(n9204) );
  OAI21_X1 U10654 ( .B1(n9687), .B2(n9234), .A(n9204), .ZN(n9205) );
  AOI21_X1 U10655 ( .B1(n9875), .B2(n9251), .A(n9205), .ZN(n9206) );
  OAI21_X1 U10656 ( .B1(n9207), .B2(n9253), .A(n9206), .ZN(P1_U3227) );
  INV_X1 U10657 ( .A(n9896), .ZN(n9752) );
  OAI21_X1 U10658 ( .B1(n9210), .B2(n9209), .A(n9208), .ZN(n9212) );
  NAND2_X1 U10659 ( .A1(n9212), .A2(n9211), .ZN(n9217) );
  OAI22_X1 U10660 ( .A1(n9783), .A2(n9245), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9213), .ZN(n9215) );
  NOR2_X1 U10661 ( .A1(n9249), .A2(n9753), .ZN(n9214) );
  AOI211_X1 U10662 ( .C1(n9247), .C2(n9728), .A(n9215), .B(n9214), .ZN(n9216)
         );
  OAI211_X1 U10663 ( .C1(n9752), .C2(n9218), .A(n9217), .B(n9216), .ZN(
        P1_U3231) );
  NAND2_X1 U10664 ( .A1(n9220), .A2(n9219), .ZN(n9222) );
  XNOR2_X1 U10665 ( .A(n9222), .B(n9221), .ZN(n9228) );
  OAI22_X1 U10666 ( .A1(n9760), .A2(n9245), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9223), .ZN(n9224) );
  AOI21_X1 U10667 ( .B1(n9247), .B2(n9729), .A(n9224), .ZN(n9225) );
  OAI21_X1 U10668 ( .B1(n9249), .B2(n9721), .A(n9225), .ZN(n9226) );
  AOI21_X1 U10669 ( .B1(n9883), .B2(n9251), .A(n9226), .ZN(n9227) );
  OAI21_X1 U10670 ( .B1(n9228), .B2(n9253), .A(n9227), .ZN(P1_U3233) );
  NAND2_X1 U10671 ( .A1(n9230), .A2(n9229), .ZN(n9231) );
  XOR2_X1 U10672 ( .A(n9232), .B(n9231), .Z(n9240) );
  OAI21_X1 U10673 ( .B1(n9783), .B2(n9234), .A(n9233), .ZN(n9235) );
  AOI21_X1 U10674 ( .B1(n9236), .B2(n9550), .A(n9235), .ZN(n9237) );
  OAI21_X1 U10675 ( .B1(n9249), .B2(n9788), .A(n9237), .ZN(n9238) );
  AOI21_X1 U10676 ( .B1(n9906), .B2(n9251), .A(n9238), .ZN(n9239) );
  OAI21_X1 U10677 ( .B1(n9240), .B2(n9253), .A(n9239), .ZN(P1_U3236) );
  NAND2_X1 U10678 ( .A1(n9242), .A2(n9241), .ZN(n9243) );
  XOR2_X1 U10679 ( .A(n9244), .B(n9243), .Z(n9254) );
  NAND2_X1 U10680 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10115)
         );
  OAI21_X1 U10681 ( .B1(n9819), .B2(n9245), .A(n10115), .ZN(n9246) );
  AOI21_X1 U10682 ( .B1(n9247), .B2(n9551), .A(n9246), .ZN(n9248) );
  OAI21_X1 U10683 ( .B1(n9249), .B2(n9827), .A(n9248), .ZN(n9250) );
  AOI21_X1 U10684 ( .B1(n9919), .B2(n9251), .A(n9250), .ZN(n9252) );
  OAI21_X1 U10685 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(P1_U3239) );
  INV_X1 U10686 ( .A(n9544), .ZN(n9295) );
  OR2_X1 U10687 ( .A1(n9840), .A2(n9295), .ZN(n9294) );
  NAND2_X1 U10688 ( .A1(n9294), .A2(n9543), .ZN(n9255) );
  NAND2_X1 U10689 ( .A1(n9255), .A2(n9293), .ZN(n9458) );
  AND2_X1 U10690 ( .A1(n9415), .A2(n9400), .ZN(n9399) );
  INV_X1 U10691 ( .A(n9403), .ZN(n9256) );
  NAND2_X1 U10692 ( .A1(n9416), .A2(n9256), .ZN(n9257) );
  NAND2_X1 U10693 ( .A1(n9421), .A2(n9257), .ZN(n9408) );
  OR2_X1 U10694 ( .A1(n9408), .A2(n9416), .ZN(n9258) );
  AND2_X1 U10695 ( .A1(n9258), .A2(n9418), .ZN(n9331) );
  INV_X1 U10696 ( .A(n9404), .ZN(n9259) );
  OR2_X1 U10697 ( .A1(n9408), .A2(n9259), .ZN(n9506) );
  AND2_X1 U10698 ( .A1(n9401), .A2(n9260), .ZN(n9391) );
  OR3_X1 U10699 ( .A1(n9506), .A2(n4933), .A3(n9391), .ZN(n9261) );
  OAI211_X1 U10700 ( .C1(n9399), .C2(n9408), .A(n9331), .B(n9261), .ZN(n9509)
         );
  NAND2_X1 U10701 ( .A1(n9397), .A2(n9262), .ZN(n9393) );
  INV_X1 U10702 ( .A(n9387), .ZN(n9279) );
  INV_X1 U10703 ( .A(n9263), .ZN(n9264) );
  AND2_X1 U10704 ( .A1(n9363), .A2(n9264), .ZN(n9368) );
  NAND2_X1 U10705 ( .A1(n9357), .A2(n9265), .ZN(n9346) );
  NAND2_X1 U10706 ( .A1(n9346), .A2(n9348), .ZN(n9266) );
  AND3_X1 U10707 ( .A1(n9367), .A2(n9368), .A3(n9266), .ZN(n9268) );
  NAND3_X1 U10708 ( .A1(n9383), .A2(n9268), .A3(n9377), .ZN(n9267) );
  OR3_X1 U10709 ( .A1(n9393), .A2(n9279), .A3(n9267), .ZN(n9503) );
  INV_X1 U10710 ( .A(n9268), .ZN(n9274) );
  AND2_X1 U10711 ( .A1(n9356), .A2(n9351), .ZN(n9273) );
  INV_X1 U10712 ( .A(n9363), .ZN(n9269) );
  OR2_X1 U10713 ( .A1(n9270), .A2(n9269), .ZN(n9365) );
  INV_X1 U10714 ( .A(n9367), .ZN(n9271) );
  OR2_X1 U10715 ( .A1(n9365), .A2(n9271), .ZN(n9272) );
  OAI21_X1 U10716 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(n9276) );
  NAND2_X1 U10717 ( .A1(n9375), .A2(n9275), .ZN(n9378) );
  OAI211_X1 U10718 ( .C1(n9276), .C2(n9378), .A(n9383), .B(n9377), .ZN(n9277)
         );
  AND3_X1 U10719 ( .A1(n9388), .A2(n9382), .A3(n9277), .ZN(n9278) );
  OR3_X1 U10720 ( .A1(n9393), .A2(n9279), .A3(n9278), .ZN(n9501) );
  OAI21_X1 U10721 ( .B1(n9503), .B2(n9280), .A(n9501), .ZN(n9281) );
  INV_X1 U10722 ( .A(n9281), .ZN(n9282) );
  NOR2_X1 U10723 ( .A1(n9506), .A2(n9282), .ZN(n9283) );
  OAI21_X1 U10724 ( .B1(n9509), .B2(n9283), .A(n9507), .ZN(n9284) );
  NAND2_X1 U10725 ( .A1(n9433), .A2(n9426), .ZN(n9510) );
  AOI21_X1 U10726 ( .B1(n9284), .B2(n9511), .A(n9510), .ZN(n9285) );
  NAND2_X1 U10727 ( .A1(n9440), .A2(n9434), .ZN(n9513) );
  NOR2_X1 U10728 ( .A1(n9285), .A2(n9513), .ZN(n9288) );
  NAND2_X1 U10729 ( .A1(n9451), .A2(n9442), .ZN(n9443) );
  INV_X1 U10730 ( .A(n9441), .ZN(n9286) );
  AND2_X1 U10731 ( .A1(n9444), .A2(n9286), .ZN(n9287) );
  OR2_X1 U10732 ( .A1(n9443), .A2(n9287), .ZN(n9518) );
  AOI21_X1 U10733 ( .B1(n9288), .B2(n9444), .A(n9518), .ZN(n9290) );
  NAND2_X1 U10734 ( .A1(n9454), .A2(n9450), .ZN(n9516) );
  NAND2_X1 U10735 ( .A1(n9544), .A2(n9543), .ZN(n9289) );
  NAND2_X1 U10736 ( .A1(n9840), .A2(n9289), .ZN(n9461) );
  OAI211_X1 U10737 ( .C1(n9290), .C2(n9516), .A(n9461), .B(n9521), .ZN(n9291)
         );
  AND2_X1 U10738 ( .A1(n9839), .A2(n9543), .ZN(n9474) );
  AOI211_X1 U10739 ( .C1(n9458), .C2(n9291), .A(n9472), .B(n9474), .ZN(n9330)
         );
  INV_X1 U10740 ( .A(n9543), .ZN(n9292) );
  NAND2_X1 U10741 ( .A1(n9463), .A2(n9294), .ZN(n9524) );
  NAND2_X1 U10742 ( .A1(n9840), .A2(n9295), .ZN(n9522) );
  INV_X1 U10743 ( .A(n9456), .ZN(n9326) );
  INV_X1 U10744 ( .A(n9613), .ZN(n9325) );
  INV_X1 U10745 ( .A(n9781), .ZN(n9319) );
  INV_X1 U10746 ( .A(n9814), .ZN(n9820) );
  INV_X1 U10747 ( .A(n9297), .ZN(n9312) );
  NOR3_X1 U10748 ( .A1(n9300), .A2(n9299), .A3(n9298), .ZN(n9305) );
  NOR2_X1 U10749 ( .A1(n9301), .A2(n10132), .ZN(n9302) );
  NAND4_X1 U10750 ( .A1(n9305), .A2(n9304), .A3(n9303), .A4(n9302), .ZN(n9308)
         );
  OR4_X1 U10751 ( .A1(n9308), .A2(n9307), .A3(n7095), .A4(n9306), .ZN(n9309)
         );
  NOR2_X1 U10752 ( .A1(n9310), .A2(n9309), .ZN(n9311) );
  NAND4_X1 U10753 ( .A1(n9313), .A2(n9312), .A3(n9311), .A4(n9361), .ZN(n9314)
         );
  NOR2_X1 U10754 ( .A1(n9315), .A2(n9314), .ZN(n9316) );
  NAND3_X1 U10755 ( .A1(n9385), .A2(n9820), .A3(n9316), .ZN(n9317) );
  NOR2_X1 U10756 ( .A1(n9805), .A2(n9317), .ZN(n9318) );
  NAND3_X1 U10757 ( .A1(n9772), .A2(n9319), .A3(n9318), .ZN(n9320) );
  NOR2_X1 U10758 ( .A1(n9757), .A2(n9320), .ZN(n9321) );
  AND4_X1 U10759 ( .A1(n9708), .A2(n9726), .A3(n9744), .A4(n9321), .ZN(n9322)
         );
  NAND4_X1 U10760 ( .A1(n9651), .A2(n9695), .A3(n9668), .A4(n9322), .ZN(n9323)
         );
  NOR2_X1 U10761 ( .A1(n9636), .A2(n9323), .ZN(n9324) );
  NAND4_X1 U10762 ( .A1(n9522), .A2(n9326), .A3(n9325), .A4(n9324), .ZN(n9327)
         );
  NOR2_X1 U10763 ( .A1(n9330), .A2(n9329), .ZN(n9471) );
  INV_X1 U10764 ( .A(n9460), .ZN(n9462) );
  INV_X1 U10765 ( .A(n9331), .ZN(n9410) );
  NAND2_X1 U10766 ( .A1(n9333), .A2(n9332), .ZN(n9335) );
  NAND2_X1 U10767 ( .A1(n9335), .A2(n9334), .ZN(n9337) );
  NAND2_X1 U10768 ( .A1(n9337), .A2(n9336), .ZN(n9340) );
  AND2_X1 U10769 ( .A1(n9338), .A2(n9460), .ZN(n9339) );
  NAND2_X1 U10770 ( .A1(n9340), .A2(n9339), .ZN(n9344) );
  NAND2_X1 U10771 ( .A1(n9341), .A2(n9497), .ZN(n9342) );
  NAND3_X1 U10772 ( .A1(n9342), .A2(n9462), .A3(n9499), .ZN(n9343) );
  NAND2_X1 U10773 ( .A1(n9344), .A2(n9343), .ZN(n9352) );
  NAND2_X1 U10774 ( .A1(n9345), .A2(n9351), .ZN(n9347) );
  INV_X1 U10775 ( .A(n9346), .ZN(n9354) );
  OAI21_X1 U10776 ( .B1(n9352), .B2(n9347), .A(n9354), .ZN(n9349) );
  NAND3_X1 U10777 ( .A1(n9349), .A2(n9348), .A3(n9369), .ZN(n9350) );
  NAND2_X1 U10778 ( .A1(n9350), .A2(n9462), .ZN(n9364) );
  NAND2_X1 U10779 ( .A1(n9352), .A2(n9351), .ZN(n9355) );
  NAND3_X1 U10780 ( .A1(n9355), .A2(n9354), .A3(n9353), .ZN(n9360) );
  INV_X1 U10781 ( .A(n9356), .ZN(n9358) );
  AOI21_X1 U10782 ( .B1(n9358), .B2(n9357), .A(n9462), .ZN(n9359) );
  NAND2_X1 U10783 ( .A1(n9360), .A2(n9359), .ZN(n9362) );
  NAND4_X1 U10784 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n9374)
         );
  INV_X1 U10785 ( .A(n9365), .ZN(n9366) );
  OAI21_X1 U10786 ( .B1(n9378), .B2(n9366), .A(n9460), .ZN(n9373) );
  NAND2_X1 U10787 ( .A1(n9377), .A2(n9367), .ZN(n9376) );
  INV_X1 U10788 ( .A(n9368), .ZN(n9370) );
  AND2_X1 U10789 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  OAI21_X1 U10790 ( .B1(n9376), .B2(n9371), .A(n9462), .ZN(n9372) );
  NAND3_X1 U10791 ( .A1(n9374), .A2(n9373), .A3(n9372), .ZN(n9381) );
  NAND3_X1 U10792 ( .A1(n9376), .A2(n9375), .A3(n9460), .ZN(n9380) );
  NAND3_X1 U10793 ( .A1(n9378), .A2(n9462), .A3(n9377), .ZN(n9379) );
  NAND4_X1 U10794 ( .A1(n9381), .A2(n9820), .A3(n9380), .A4(n9379), .ZN(n9386)
         );
  MUX2_X1 U10795 ( .A(n9383), .B(n9382), .S(n9460), .Z(n9384) );
  NAND3_X1 U10796 ( .A1(n9386), .A2(n9385), .A3(n9384), .ZN(n9390) );
  MUX2_X1 U10797 ( .A(n9388), .B(n9387), .S(n9460), .Z(n9389) );
  NAND2_X1 U10798 ( .A1(n9390), .A2(n9389), .ZN(n9396) );
  INV_X1 U10799 ( .A(n9391), .ZN(n9392) );
  NAND2_X1 U10800 ( .A1(n9392), .A2(n9460), .ZN(n9395) );
  NAND2_X1 U10801 ( .A1(n9393), .A2(n9462), .ZN(n9394) );
  OAI211_X1 U10802 ( .C1(n9805), .C2(n9396), .A(n9395), .B(n9394), .ZN(n9402)
         );
  NAND3_X1 U10803 ( .A1(n9402), .A2(n9397), .A3(n9404), .ZN(n9398) );
  NAND3_X1 U10804 ( .A1(n9399), .A2(n9460), .A3(n9398), .ZN(n9407) );
  NAND3_X1 U10805 ( .A1(n9402), .A2(n9401), .A3(n9400), .ZN(n9405) );
  NAND4_X1 U10806 ( .A1(n9405), .A2(n9462), .A3(n9404), .A4(n9403), .ZN(n9406)
         );
  NAND2_X1 U10807 ( .A1(n9407), .A2(n9406), .ZN(n9414) );
  NOR2_X1 U10808 ( .A1(n9408), .A2(n9414), .ZN(n9409) );
  OAI21_X1 U10809 ( .B1(n9410), .B2(n9409), .A(n9507), .ZN(n9411) );
  NAND2_X1 U10810 ( .A1(n9411), .A2(n9460), .ZN(n9413) );
  INV_X1 U10811 ( .A(n9424), .ZN(n9412) );
  AOI21_X1 U10812 ( .B1(n9413), .B2(n9684), .A(n9412), .ZN(n9432) );
  INV_X1 U10813 ( .A(n9414), .ZN(n9417) );
  NAND3_X1 U10814 ( .A1(n9417), .A2(n9416), .A3(n9415), .ZN(n9420) );
  INV_X1 U10815 ( .A(n9418), .ZN(n9419) );
  AOI21_X1 U10816 ( .B1(n9421), .B2(n9420), .A(n9419), .ZN(n9422) );
  AOI22_X1 U10817 ( .A1(n9695), .A2(n9422), .B1(n9426), .B2(n9460), .ZN(n9431)
         );
  INV_X1 U10818 ( .A(n9507), .ZN(n9423) );
  AND2_X1 U10819 ( .A1(n9424), .A2(n9423), .ZN(n9425) );
  OAI21_X1 U10820 ( .B1(n9510), .B2(n9425), .A(n9462), .ZN(n9430) );
  INV_X1 U10821 ( .A(n9426), .ZN(n9427) );
  OAI21_X1 U10822 ( .B1(n9427), .B2(n9684), .A(n9434), .ZN(n9428) );
  NAND2_X1 U10823 ( .A1(n9428), .A2(n9460), .ZN(n9429) );
  OAI211_X1 U10824 ( .C1(n9432), .C2(n9431), .A(n9430), .B(n9429), .ZN(n9438)
         );
  OR2_X1 U10825 ( .A1(n9433), .A2(n9462), .ZN(n9437) );
  INV_X1 U10826 ( .A(n9434), .ZN(n9435) );
  NAND2_X1 U10827 ( .A1(n9435), .A2(n9462), .ZN(n9436) );
  NAND4_X1 U10828 ( .A1(n9438), .A2(n9651), .A3(n9437), .A4(n9436), .ZN(n9439)
         );
  OAI211_X1 U10829 ( .C1(n9462), .C2(n9440), .A(n9439), .B(n9444), .ZN(n9449)
         );
  AOI21_X1 U10830 ( .B1(n9442), .B2(n9441), .A(n9460), .ZN(n9448) );
  NAND2_X1 U10831 ( .A1(n9443), .A2(n9460), .ZN(n9447) );
  NAND2_X1 U10832 ( .A1(n9450), .A2(n9444), .ZN(n9445) );
  NAND2_X1 U10833 ( .A1(n9445), .A2(n9462), .ZN(n9446) );
  OAI211_X1 U10834 ( .C1(n9449), .C2(n9448), .A(n9447), .B(n9446), .ZN(n9453)
         );
  MUX2_X1 U10835 ( .A(n9451), .B(n9450), .S(n9460), .Z(n9452) );
  AND2_X1 U10836 ( .A1(n9453), .A2(n9452), .ZN(n9457) );
  MUX2_X1 U10837 ( .A(n9521), .B(n9454), .S(n9460), .Z(n9455) );
  OAI211_X1 U10838 ( .C1(n9457), .C2(n9456), .A(n9461), .B(n9455), .ZN(n9459)
         );
  MUX2_X1 U10839 ( .A(n9460), .B(n9459), .S(n9458), .Z(n9466) );
  INV_X1 U10840 ( .A(n9474), .ZN(n9525) );
  OAI21_X1 U10841 ( .B1(n9462), .B2(n9461), .A(n9525), .ZN(n9464) );
  NAND2_X1 U10842 ( .A1(n9464), .A2(n9463), .ZN(n9465) );
  NAND2_X1 U10843 ( .A1(n9466), .A2(n9465), .ZN(n9476) );
  INV_X1 U10844 ( .A(n9467), .ZN(n9469) );
  OAI21_X1 U10845 ( .B1(n9476), .B2(n9469), .A(n9468), .ZN(n9470) );
  NOR3_X1 U10846 ( .A1(n9474), .A2(n9473), .A3(n9472), .ZN(n9475) );
  NAND2_X1 U10847 ( .A1(n9476), .A2(n9475), .ZN(n9477) );
  INV_X1 U10848 ( .A(n9478), .ZN(n9481) );
  NAND2_X1 U10849 ( .A1(n9564), .A2(n10171), .ZN(n9479) );
  NAND3_X1 U10850 ( .A1(n9481), .A2(n9480), .A3(n9479), .ZN(n9483) );
  NAND2_X1 U10851 ( .A1(n9483), .A2(n9482), .ZN(n9486) );
  OAI22_X1 U10852 ( .A1(n9487), .A2(n9486), .B1(n9485), .B2(n9484), .ZN(n9489)
         );
  NAND2_X1 U10853 ( .A1(n9489), .A2(n9488), .ZN(n9492) );
  NAND3_X1 U10854 ( .A1(n9492), .A2(n9491), .A3(n9490), .ZN(n9494) );
  NAND2_X1 U10855 ( .A1(n9494), .A2(n9493), .ZN(n9498) );
  INV_X1 U10856 ( .A(n9495), .ZN(n9496) );
  NAND3_X1 U10857 ( .A1(n9498), .A2(n9497), .A3(n9496), .ZN(n9500) );
  NAND2_X1 U10858 ( .A1(n9500), .A2(n9499), .ZN(n9502) );
  OAI21_X1 U10859 ( .B1(n9503), .B2(n9502), .A(n9501), .ZN(n9504) );
  INV_X1 U10860 ( .A(n9504), .ZN(n9505) );
  NOR2_X1 U10861 ( .A1(n9506), .A2(n9505), .ZN(n9508) );
  OAI21_X1 U10862 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(n9512) );
  AOI21_X1 U10863 ( .B1(n9512), .B2(n9511), .A(n9510), .ZN(n9514) );
  OR2_X1 U10864 ( .A1(n9514), .A2(n9513), .ZN(n9515) );
  NOR2_X1 U10865 ( .A1(n9636), .A2(n9515), .ZN(n9519) );
  INV_X1 U10866 ( .A(n9516), .ZN(n9517) );
  OAI21_X1 U10867 ( .B1(n9519), .B2(n9518), .A(n9517), .ZN(n9520) );
  AND3_X1 U10868 ( .A1(n9522), .A2(n9521), .A3(n9520), .ZN(n9523) );
  OR2_X1 U10869 ( .A1(n9524), .A2(n9523), .ZN(n9526) );
  NOR2_X1 U10870 ( .A1(n9533), .A2(n9690), .ZN(n9529) );
  INV_X1 U10871 ( .A(n9533), .ZN(n9535) );
  OAI21_X1 U10872 ( .B1(n9535), .B2(n9534), .A(n9537), .ZN(n9541) );
  NAND2_X1 U10873 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  OAI211_X1 U10874 ( .C1(n9539), .C2(n10065), .A(P1_B_REG_SCAN_IN), .B(n9538), 
        .ZN(n9540) );
  OAI21_X1 U10875 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(P1_U3240) );
  MUX2_X1 U10876 ( .A(n9543), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9563), .Z(
        P1_U3586) );
  MUX2_X1 U10877 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9544), .S(n9562), .Z(
        P1_U3585) );
  MUX2_X1 U10878 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9545), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10879 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n4778), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10880 ( .A(n9546), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9563), .Z(
        P1_U3581) );
  MUX2_X1 U10881 ( .A(n9547), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9563), .Z(
        P1_U3580) );
  MUX2_X1 U10882 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9548), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10883 ( .A(n9729), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9563), .Z(
        P1_U3578) );
  MUX2_X1 U10884 ( .A(n9738), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9563), .Z(
        P1_U3577) );
  MUX2_X1 U10885 ( .A(n9728), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9563), .Z(
        P1_U3576) );
  MUX2_X1 U10886 ( .A(n9773), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9563), .Z(
        P1_U3575) );
  MUX2_X1 U10887 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9549), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10888 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9774), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10889 ( .A(n9550), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9563), .Z(
        P1_U3572) );
  MUX2_X1 U10890 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9551), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10891 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9552), .S(n9562), .Z(
        P1_U3570) );
  MUX2_X1 U10892 ( .A(n9553), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9563), .Z(
        P1_U3569) );
  MUX2_X1 U10893 ( .A(n9554), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9563), .Z(
        P1_U3568) );
  MUX2_X1 U10894 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9555), .S(n9562), .Z(
        P1_U3566) );
  MUX2_X1 U10895 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9556), .S(n9562), .Z(
        P1_U3564) );
  MUX2_X1 U10896 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9557), .S(n9562), .Z(
        P1_U3562) );
  MUX2_X1 U10897 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9558), .S(n9562), .Z(
        P1_U3561) );
  MUX2_X1 U10898 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9559), .S(n9562), .Z(
        P1_U3560) );
  MUX2_X1 U10899 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9560), .S(n9562), .Z(
        P1_U3559) );
  MUX2_X1 U10900 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9561), .S(n9562), .Z(
        P1_U3558) );
  MUX2_X1 U10901 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10139), .S(n9562), .Z(
        P1_U3557) );
  MUX2_X1 U10902 ( .A(n9564), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9563), .Z(
        P1_U3556) );
  OAI21_X1 U10903 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(n9571) );
  INV_X1 U10904 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9568) );
  NOR2_X1 U10905 ( .A1(n10063), .A2(n9568), .ZN(n9569) );
  AOI211_X1 U10906 ( .C1(n10120), .C2(n9571), .A(n9570), .B(n9569), .ZN(n9580)
         );
  INV_X1 U10907 ( .A(n9572), .ZN(n9576) );
  INV_X1 U10908 ( .A(n9573), .ZN(n9575) );
  OAI21_X1 U10909 ( .B1(n9576), .B2(n9575), .A(n9574), .ZN(n9577) );
  AOI22_X1 U10910 ( .A1(n9578), .A2(n10118), .B1(n10124), .B2(n9577), .ZN(
        n9579) );
  NAND3_X1 U10911 ( .A1(n9581), .A2(n9580), .A3(n9579), .ZN(P1_U3245) );
  AOI21_X1 U10912 ( .B1(n9583), .B2(n9587), .A(n9582), .ZN(n9585) );
  XOR2_X1 U10913 ( .A(n9585), .B(n9584), .Z(n9598) );
  OAI21_X1 U10914 ( .B1(n9588), .B2(n9587), .A(n9586), .ZN(n9589) );
  XNOR2_X1 U10915 ( .A(n9589), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9594) );
  OAI22_X1 U10916 ( .A1(n9598), .A2(n10106), .B1(n9594), .B2(n9590), .ZN(n9591) );
  INV_X1 U10917 ( .A(n9591), .ZN(n9600) );
  INV_X1 U10918 ( .A(n9592), .ZN(n9593) );
  NAND2_X1 U10919 ( .A1(n9594), .A2(n9593), .ZN(n9596) );
  NAND2_X1 U10920 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  AOI21_X1 U10921 ( .B1(n9598), .B2(n10120), .A(n9597), .ZN(n9599) );
  MUX2_X1 U10922 ( .A(n9600), .B(n9599), .S(n10148), .Z(n9604) );
  INV_X1 U10923 ( .A(n9601), .ZN(n9602) );
  AOI21_X1 U10924 ( .B1(n10122), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9602), .ZN(
        n9603) );
  NAND2_X1 U10925 ( .A1(n9604), .A2(n9603), .ZN(P1_U3260) );
  OAI21_X1 U10926 ( .B1(n9607), .B2(n9606), .A(n9605), .ZN(n9843) );
  NOR2_X1 U10927 ( .A1(n9607), .A2(n9799), .ZN(n9608) );
  AOI211_X1 U10928 ( .C1(n10157), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9609), .B(
        n9608), .ZN(n9610) );
  OAI21_X1 U10929 ( .B1(n9832), .B2(n9843), .A(n9610), .ZN(P1_U3262) );
  OAI21_X1 U10930 ( .B1(n9612), .B2(n9613), .A(n9611), .ZN(n9853) );
  AND2_X1 U10931 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  OR2_X1 U10932 ( .A1(n4542), .A2(n9615), .ZN(n9618) );
  OAI22_X1 U10933 ( .A1(n9654), .A2(n9818), .B1(n9616), .B2(n9816), .ZN(n9617)
         );
  INV_X1 U10934 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9619) );
  OAI22_X1 U10935 ( .A1(n9620), .A2(n10150), .B1(n9619), .B2(n9810), .ZN(n9621) );
  AOI21_X1 U10936 ( .B1(n9849), .B2(n9830), .A(n9621), .ZN(n9626) );
  OR2_X1 U10937 ( .A1(n9622), .A2(n9631), .ZN(n9624) );
  AND2_X1 U10938 ( .A1(n9624), .A2(n9623), .ZN(n9850) );
  NAND2_X1 U10939 ( .A1(n9850), .A2(n9733), .ZN(n9625) );
  OAI211_X1 U10940 ( .C1(n9852), .C2(n10157), .A(n9626), .B(n9625), .ZN(n9627)
         );
  INV_X1 U10941 ( .A(n9627), .ZN(n9628) );
  OAI21_X1 U10942 ( .B1(n9853), .B2(n9813), .A(n9628), .ZN(P1_U3263) );
  XNOR2_X1 U10943 ( .A(n9630), .B(n9629), .ZN(n9858) );
  AOI21_X1 U10944 ( .B1(n9854), .B2(n9646), .A(n9631), .ZN(n9855) );
  AOI22_X1 U10945 ( .A1(n9632), .A2(n9789), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n10157), .ZN(n9633) );
  OAI21_X1 U10946 ( .B1(n9634), .B2(n9799), .A(n9633), .ZN(n9643) );
  INV_X1 U10947 ( .A(n9635), .ZN(n9637) );
  AOI21_X1 U10948 ( .B1(n9637), .B2(n9636), .A(n9807), .ZN(n9641) );
  OAI22_X1 U10949 ( .A1(n9638), .A2(n9816), .B1(n9671), .B2(n9818), .ZN(n9639)
         );
  AOI21_X1 U10950 ( .B1(n9641), .B2(n9640), .A(n9639), .ZN(n9857) );
  NOR2_X1 U10951 ( .A1(n9857), .A2(n10157), .ZN(n9642) );
  AOI211_X1 U10952 ( .C1(n9733), .C2(n9855), .A(n9643), .B(n9642), .ZN(n9644)
         );
  OAI21_X1 U10953 ( .B1(n9858), .B2(n9813), .A(n9644), .ZN(P1_U3264) );
  XNOR2_X1 U10954 ( .A(n9645), .B(n9651), .ZN(n9863) );
  AOI21_X1 U10955 ( .B1(n9859), .B2(n9675), .A(n4570), .ZN(n9860) );
  AOI22_X1 U10956 ( .A1(n9647), .A2(n9789), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n10157), .ZN(n9648) );
  OAI21_X1 U10957 ( .B1(n9649), .B2(n9799), .A(n9648), .ZN(n9659) );
  INV_X1 U10958 ( .A(n9650), .ZN(n9653) );
  INV_X1 U10959 ( .A(n9651), .ZN(n9652) );
  AOI21_X1 U10960 ( .B1(n9653), .B2(n9652), .A(n9807), .ZN(n9657) );
  OAI22_X1 U10961 ( .A1(n9654), .A2(n9816), .B1(n9687), .B2(n9818), .ZN(n9655)
         );
  AOI21_X1 U10962 ( .B1(n9657), .B2(n9656), .A(n9655), .ZN(n9862) );
  NOR2_X1 U10963 ( .A1(n9862), .A2(n10157), .ZN(n9658) );
  AOI211_X1 U10964 ( .C1(n9860), .C2(n9733), .A(n9659), .B(n9658), .ZN(n9660)
         );
  OAI21_X1 U10965 ( .B1(n9863), .B2(n9813), .A(n9660), .ZN(P1_U3265) );
  OR2_X1 U10966 ( .A1(n9700), .A2(n9661), .ZN(n9663) );
  NAND2_X1 U10967 ( .A1(n9663), .A2(n9662), .ZN(n9666) );
  OAI21_X1 U10968 ( .B1(n9666), .B2(n9665), .A(n9664), .ZN(n9864) );
  INV_X1 U10969 ( .A(n9864), .ZN(n9680) );
  AOI22_X1 U10970 ( .A1(n9667), .A2(n9830), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n10157), .ZN(n9679) );
  XNOR2_X1 U10971 ( .A(n9669), .B(n9668), .ZN(n9670) );
  NAND2_X1 U10972 ( .A1(n9670), .A2(n10135), .ZN(n9674) );
  OAI22_X1 U10973 ( .A1(n9671), .A2(n9816), .B1(n9710), .B2(n9818), .ZN(n9672)
         );
  INV_X1 U10974 ( .A(n9672), .ZN(n9673) );
  NAND2_X1 U10975 ( .A1(n9674), .A2(n9673), .ZN(n9868) );
  OAI211_X1 U10976 ( .C1(n9866), .C2(n9681), .A(n10146), .B(n9675), .ZN(n9865)
         );
  OAI22_X1 U10977 ( .A1(n9865), .A2(n10148), .B1(n10150), .B2(n9676), .ZN(
        n9677) );
  OAI21_X1 U10978 ( .B1(n9868), .B2(n9677), .A(n9810), .ZN(n9678) );
  OAI211_X1 U10979 ( .C1(n9680), .C2(n9813), .A(n9679), .B(n9678), .ZN(
        P1_U3266) );
  AOI211_X1 U10980 ( .C1(n9875), .C2(n9701), .A(n10205), .B(n9681), .ZN(n9874)
         );
  INV_X1 U10981 ( .A(n9682), .ZN(n9683) );
  NOR2_X1 U10982 ( .A1(n9683), .A2(n10150), .ZN(n9689) );
  NAND2_X1 U10983 ( .A1(n9712), .A2(n9684), .ZN(n9685) );
  XNOR2_X1 U10984 ( .A(n9685), .B(n9695), .ZN(n9686) );
  OAI222_X1 U10985 ( .A1(n9818), .A2(n9688), .B1(n9816), .B2(n9687), .C1(n9807), .C2(n9686), .ZN(n9873) );
  AOI211_X1 U10986 ( .C1(n9874), .C2(n9690), .A(n9689), .B(n9873), .ZN(n9699)
         );
  AOI22_X1 U10987 ( .A1(n9875), .A2(n9830), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n10157), .ZN(n9698) );
  OR2_X1 U10988 ( .A1(n9700), .A2(n9691), .ZN(n9694) );
  NAND2_X1 U10989 ( .A1(n9694), .A2(n9692), .ZN(n9872) );
  NAND2_X1 U10990 ( .A1(n9694), .A2(n9693), .ZN(n9696) );
  NAND2_X1 U10991 ( .A1(n9696), .A2(n9695), .ZN(n9871) );
  NAND3_X1 U10992 ( .A1(n9872), .A2(n9871), .A3(n9746), .ZN(n9697) );
  OAI211_X1 U10993 ( .C1(n9699), .C2(n10157), .A(n9698), .B(n9697), .ZN(
        P1_U3267) );
  XOR2_X1 U10994 ( .A(n9708), .B(n9700), .Z(n9882) );
  INV_X1 U10995 ( .A(n9701), .ZN(n9702) );
  AOI21_X1 U10996 ( .B1(n9878), .B2(n9719), .A(n9702), .ZN(n9879) );
  INV_X1 U10997 ( .A(n9703), .ZN(n9704) );
  AOI22_X1 U10998 ( .A1(n9704), .A2(n9789), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n10157), .ZN(n9705) );
  OAI21_X1 U10999 ( .B1(n9706), .B2(n9799), .A(n9705), .ZN(n9715) );
  AOI21_X1 U11000 ( .B1(n4912), .B2(n4917), .A(n9807), .ZN(n9713) );
  OAI22_X1 U11001 ( .A1(n9710), .A2(n9816), .B1(n9709), .B2(n9818), .ZN(n9711)
         );
  AOI21_X1 U11002 ( .B1(n9713), .B2(n9712), .A(n9711), .ZN(n9881) );
  NOR2_X1 U11003 ( .A1(n9881), .A2(n10157), .ZN(n9714) );
  AOI211_X1 U11004 ( .C1(n9879), .C2(n9733), .A(n9715), .B(n9714), .ZN(n9716)
         );
  OAI21_X1 U11005 ( .B1(n9882), .B2(n9813), .A(n9716), .ZN(P1_U3268) );
  XOR2_X1 U11006 ( .A(n9717), .B(n9726), .Z(n9887) );
  INV_X1 U11007 ( .A(n9718), .ZN(n9735) );
  INV_X1 U11008 ( .A(n9719), .ZN(n9720) );
  AOI21_X1 U11009 ( .B1(n9883), .B2(n9735), .A(n9720), .ZN(n9884) );
  INV_X1 U11010 ( .A(n9721), .ZN(n9722) );
  AOI22_X1 U11011 ( .A1(n9722), .A2(n9789), .B1(n10157), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9723) );
  OAI21_X1 U11012 ( .B1(n9724), .B2(n9799), .A(n9723), .ZN(n9732) );
  NAND2_X1 U11013 ( .A1(n9737), .A2(n9725), .ZN(n9727) );
  XNOR2_X1 U11014 ( .A(n9727), .B(n9726), .ZN(n9730) );
  AOI222_X1 U11015 ( .A1(n10135), .A2(n9730), .B1(n9729), .B2(n10140), .C1(
        n9728), .C2(n10137), .ZN(n9886) );
  NOR2_X1 U11016 ( .A1(n9886), .A2(n10157), .ZN(n9731) );
  AOI211_X1 U11017 ( .C1(n9884), .C2(n9733), .A(n9732), .B(n9731), .ZN(n9734)
         );
  OAI21_X1 U11018 ( .B1(n9813), .B2(n9887), .A(n9734), .ZN(P1_U3269) );
  OAI211_X1 U11019 ( .C1(n9736), .C2(n9751), .A(n9735), .B(n10146), .ZN(n9890)
         );
  NOR2_X1 U11020 ( .A1(n9890), .A2(n10148), .ZN(n9741) );
  OAI21_X1 U11021 ( .B1(n4520), .B2(n9744), .A(n9737), .ZN(n9739) );
  AOI222_X1 U11022 ( .A1(n10135), .A2(n9739), .B1(n9738), .B2(n10140), .C1(
        n9773), .C2(n10137), .ZN(n9892) );
  INV_X1 U11023 ( .A(n9892), .ZN(n9740) );
  AOI211_X1 U11024 ( .C1(n9789), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9749)
         );
  AOI22_X1 U11025 ( .A1(n9889), .A2(n9830), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n10157), .ZN(n9748) );
  NAND2_X1 U11026 ( .A1(n9745), .A2(n9744), .ZN(n9888) );
  NAND3_X1 U11027 ( .A1(n9743), .A2(n9888), .A3(n9746), .ZN(n9747) );
  OAI211_X1 U11028 ( .C1(n9749), .C2(n10157), .A(n9748), .B(n9747), .ZN(
        P1_U3270) );
  XNOR2_X1 U11029 ( .A(n9750), .B(n9757), .ZN(n9898) );
  AOI211_X1 U11030 ( .C1(n9896), .C2(n9764), .A(n10205), .B(n9751), .ZN(n9895)
         );
  NOR2_X1 U11031 ( .A1(n9752), .A2(n9799), .ZN(n9756) );
  OAI22_X1 U11032 ( .A1(n9810), .A2(n9754), .B1(n9753), .B2(n10150), .ZN(n9755) );
  AOI211_X1 U11033 ( .C1(n9895), .C2(n9804), .A(n9756), .B(n9755), .ZN(n9762)
         );
  XNOR2_X1 U11034 ( .A(n9758), .B(n9757), .ZN(n9759) );
  OAI222_X1 U11035 ( .A1(n9818), .A2(n9783), .B1(n9816), .B2(n9760), .C1(n9759), .C2(n9807), .ZN(n9894) );
  NAND2_X1 U11036 ( .A1(n9894), .A2(n9810), .ZN(n9761) );
  OAI211_X1 U11037 ( .C1(n9898), .C2(n9813), .A(n9762), .B(n9761), .ZN(
        P1_U3271) );
  XOR2_X1 U11038 ( .A(n9763), .B(n9772), .Z(n9903) );
  INV_X1 U11039 ( .A(n9764), .ZN(n9765) );
  AOI211_X1 U11040 ( .C1(n9900), .C2(n9785), .A(n10205), .B(n9765), .ZN(n9899)
         );
  INV_X1 U11041 ( .A(n9766), .ZN(n9767) );
  AOI22_X1 U11042 ( .A1(n10157), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9767), 
        .B2(n9789), .ZN(n9768) );
  OAI21_X1 U11043 ( .B1(n9769), .B2(n9799), .A(n9768), .ZN(n9777) );
  OAI21_X1 U11044 ( .B1(n9772), .B2(n9771), .A(n9770), .ZN(n9775) );
  AOI222_X1 U11045 ( .A1(n10135), .A2(n9775), .B1(n9774), .B2(n10137), .C1(
        n9773), .C2(n10140), .ZN(n9902) );
  NOR2_X1 U11046 ( .A1(n9902), .A2(n10157), .ZN(n9776) );
  AOI211_X1 U11047 ( .C1(n9804), .C2(n9899), .A(n9777), .B(n9776), .ZN(n9778)
         );
  OAI21_X1 U11048 ( .B1(n9813), .B2(n9903), .A(n9778), .ZN(P1_U3272) );
  XNOR2_X1 U11049 ( .A(n9779), .B(n9781), .ZN(n9908) );
  AOI21_X1 U11050 ( .B1(n9781), .B2(n9780), .A(n4521), .ZN(n9782) );
  OAI222_X1 U11051 ( .A1(n9818), .A2(n9784), .B1(n9816), .B2(n9783), .C1(n9807), .C2(n9782), .ZN(n9904) );
  INV_X1 U11052 ( .A(n9798), .ZN(n9787) );
  INV_X1 U11053 ( .A(n9785), .ZN(n9786) );
  AOI211_X1 U11054 ( .C1(n9906), .C2(n9787), .A(n10205), .B(n9786), .ZN(n9905)
         );
  NAND2_X1 U11055 ( .A1(n9905), .A2(n9804), .ZN(n9792) );
  INV_X1 U11056 ( .A(n9788), .ZN(n9790) );
  AOI22_X1 U11057 ( .A1(n10157), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9790), 
        .B2(n9789), .ZN(n9791) );
  OAI211_X1 U11058 ( .C1(n9793), .C2(n9799), .A(n9792), .B(n9791), .ZN(n9794)
         );
  AOI21_X1 U11059 ( .B1(n9904), .B2(n9810), .A(n9794), .ZN(n9795) );
  OAI21_X1 U11060 ( .B1(n9908), .B2(n9813), .A(n9795), .ZN(P1_U3273) );
  XNOR2_X1 U11061 ( .A(n9796), .B(n9805), .ZN(n9913) );
  AOI211_X1 U11062 ( .C1(n9911), .C2(n4751), .A(n10205), .B(n9798), .ZN(n9910)
         );
  NOR2_X1 U11063 ( .A1(n9800), .A2(n9799), .ZN(n9803) );
  OAI22_X1 U11064 ( .A1(n9810), .A2(n7211), .B1(n9801), .B2(n10150), .ZN(n9802) );
  AOI211_X1 U11065 ( .C1(n9910), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9812)
         );
  XNOR2_X1 U11066 ( .A(n9806), .B(n9805), .ZN(n9808) );
  OAI222_X1 U11067 ( .A1(n9816), .A2(n9809), .B1(n9818), .B2(n9817), .C1(n9808), .C2(n9807), .ZN(n9909) );
  NAND2_X1 U11068 ( .A1(n9909), .A2(n9810), .ZN(n9811) );
  OAI211_X1 U11069 ( .C1(n9913), .C2(n9813), .A(n9812), .B(n9811), .ZN(
        P1_U3274) );
  XNOR2_X1 U11070 ( .A(n9815), .B(n9814), .ZN(n9824) );
  OAI22_X1 U11071 ( .A1(n9819), .A2(n9818), .B1(n9817), .B2(n9816), .ZN(n9823)
         );
  XNOR2_X1 U11072 ( .A(n9821), .B(n9820), .ZN(n9925) );
  NOR2_X1 U11073 ( .A1(n9925), .A2(n10143), .ZN(n9822) );
  AOI211_X1 U11074 ( .C1(n10135), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9924)
         );
  INV_X1 U11075 ( .A(n9925), .ZN(n9835) );
  AND2_X1 U11076 ( .A1(n4560), .A2(n9919), .ZN(n9826) );
  OR2_X1 U11077 ( .A1(n9826), .A2(n9825), .ZN(n9921) );
  OAI22_X1 U11078 ( .A1(n9810), .A2(n9828), .B1(n9827), .B2(n10150), .ZN(n9829) );
  AOI21_X1 U11079 ( .B1(n9919), .B2(n9830), .A(n9829), .ZN(n9831) );
  OAI21_X1 U11080 ( .B1(n9921), .B2(n9832), .A(n9831), .ZN(n9833) );
  AOI21_X1 U11081 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9836) );
  OAI21_X1 U11082 ( .B1(n9924), .B2(n10157), .A(n9836), .ZN(P1_U3276) );
  NAND2_X1 U11083 ( .A1(n9837), .A2(n10146), .ZN(n9838) );
  OAI211_X1 U11084 ( .C1(n9839), .C2(n10204), .A(n9838), .B(n9842), .ZN(n9938)
         );
  MUX2_X1 U11085 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9938), .S(n10223), .Z(
        P1_U3554) );
  NAND2_X1 U11086 ( .A1(n9840), .A2(n10000), .ZN(n9841) );
  OAI211_X1 U11087 ( .C1(n9843), .C2(n10205), .A(n9842), .B(n9841), .ZN(n9939)
         );
  MUX2_X1 U11088 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9939), .S(n10223), .Z(
        P1_U3553) );
  AOI22_X1 U11089 ( .A1(n9850), .A2(n10146), .B1(n10000), .B2(n9849), .ZN(
        n9851) );
  OAI211_X1 U11090 ( .C1(n9853), .C2(n9930), .A(n9852), .B(n9851), .ZN(n9940)
         );
  MUX2_X1 U11091 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9940), .S(n10223), .Z(
        P1_U3551) );
  AOI22_X1 U11092 ( .A1(n9855), .A2(n10146), .B1(n10000), .B2(n9854), .ZN(
        n9856) );
  OAI211_X1 U11093 ( .C1(n9858), .C2(n9930), .A(n9857), .B(n9856), .ZN(n9941)
         );
  MUX2_X1 U11094 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9941), .S(n10223), .Z(
        P1_U3550) );
  AOI22_X1 U11095 ( .A1(n9860), .A2(n10146), .B1(n10000), .B2(n9859), .ZN(
        n9861) );
  OAI211_X1 U11096 ( .C1(n9863), .C2(n9930), .A(n9862), .B(n9861), .ZN(n9942)
         );
  MUX2_X1 U11097 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9942), .S(n10223), .Z(
        P1_U3549) );
  INV_X1 U11098 ( .A(n9930), .ZN(n10194) );
  NAND2_X1 U11099 ( .A1(n9864), .A2(n10194), .ZN(n9870) );
  OAI21_X1 U11100 ( .B1(n9866), .B2(n10204), .A(n9865), .ZN(n9867) );
  NOR2_X1 U11101 ( .A1(n9868), .A2(n9867), .ZN(n9869) );
  NAND2_X1 U11102 ( .A1(n9870), .A2(n9869), .ZN(n9943) );
  MUX2_X1 U11103 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9943), .S(n10223), .Z(
        P1_U3548) );
  NAND3_X1 U11104 ( .A1(n9872), .A2(n10194), .A3(n9871), .ZN(n9877) );
  AOI211_X1 U11105 ( .C1(n10000), .C2(n9875), .A(n9874), .B(n9873), .ZN(n9876)
         );
  NAND2_X1 U11106 ( .A1(n9877), .A2(n9876), .ZN(n9944) );
  INV_X1 U11107 ( .A(n10223), .ZN(n10220) );
  MUX2_X1 U11108 ( .A(n9944), .B(P1_REG1_REG_24__SCAN_IN), .S(n10220), .Z(
        P1_U3547) );
  AOI22_X1 U11109 ( .A1(n9879), .A2(n10146), .B1(n10000), .B2(n9878), .ZN(
        n9880) );
  OAI211_X1 U11110 ( .C1(n9882), .C2(n9930), .A(n9881), .B(n9880), .ZN(n9945)
         );
  MUX2_X1 U11111 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9945), .S(n10223), .Z(
        P1_U3546) );
  AOI22_X1 U11112 ( .A1(n9884), .A2(n10146), .B1(n10000), .B2(n9883), .ZN(
        n9885) );
  OAI211_X1 U11113 ( .C1(n9887), .C2(n9930), .A(n9886), .B(n9885), .ZN(n9946)
         );
  MUX2_X1 U11114 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9946), .S(n10223), .Z(
        P1_U3545) );
  NAND3_X1 U11115 ( .A1(n9743), .A2(n9888), .A3(n10194), .ZN(n9893) );
  NAND2_X1 U11116 ( .A1(n9889), .A2(n10000), .ZN(n9891) );
  NAND4_X1 U11117 ( .A1(n9893), .A2(n9892), .A3(n9891), .A4(n9890), .ZN(n9947)
         );
  MUX2_X1 U11118 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9947), .S(n10223), .Z(
        P1_U3544) );
  AOI211_X1 U11119 ( .C1(n10000), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9897)
         );
  OAI21_X1 U11120 ( .B1(n9898), .B2(n9930), .A(n9897), .ZN(n9948) );
  MUX2_X1 U11121 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9948), .S(n10223), .Z(
        P1_U3543) );
  AOI21_X1 U11122 ( .B1(n10000), .B2(n9900), .A(n9899), .ZN(n9901) );
  OAI211_X1 U11123 ( .C1(n9903), .C2(n9930), .A(n9902), .B(n9901), .ZN(n9949)
         );
  MUX2_X1 U11124 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9949), .S(n10223), .Z(
        P1_U3542) );
  AOI211_X1 U11125 ( .C1(n10000), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9907)
         );
  OAI21_X1 U11126 ( .B1(n9930), .B2(n9908), .A(n9907), .ZN(n9950) );
  MUX2_X1 U11127 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9950), .S(n10223), .Z(
        P1_U3541) );
  AOI211_X1 U11128 ( .C1(n10000), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9912)
         );
  OAI21_X1 U11129 ( .B1(n9913), .B2(n9930), .A(n9912), .ZN(n9951) );
  MUX2_X1 U11130 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9951), .S(n10223), .Z(
        P1_U3540) );
  AOI211_X1 U11131 ( .C1(n10000), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9917)
         );
  OAI21_X1 U11132 ( .B1(n9918), .B2(n9930), .A(n9917), .ZN(n9952) );
  MUX2_X1 U11133 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9952), .S(n10223), .Z(
        P1_U3539) );
  INV_X1 U11134 ( .A(n9919), .ZN(n9920) );
  OAI22_X1 U11135 ( .A1(n9921), .A2(n10205), .B1(n9920), .B2(n10204), .ZN(
        n9922) );
  INV_X1 U11136 ( .A(n9922), .ZN(n9923) );
  OAI211_X1 U11137 ( .C1(n9925), .C2(n9999), .A(n9924), .B(n9923), .ZN(n9953)
         );
  MUX2_X1 U11138 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9953), .S(n10223), .Z(
        P1_U3538) );
  AOI211_X1 U11139 ( .C1(n10000), .C2(n9928), .A(n9927), .B(n9926), .ZN(n9929)
         );
  OAI21_X1 U11140 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(n9954) );
  MUX2_X1 U11141 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9954), .S(n10223), .Z(
        P1_U3537) );
  AOI22_X1 U11142 ( .A1(n9933), .A2(n10146), .B1(n10000), .B2(n9932), .ZN(
        n9934) );
  OAI21_X1 U11143 ( .B1(n9935), .B2(n9999), .A(n9934), .ZN(n9936) );
  MUX2_X1 U11144 ( .A(n9955), .B(P1_REG1_REG_13__SCAN_IN), .S(n10220), .Z(
        P1_U3536) );
  MUX2_X1 U11145 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9938), .S(n10212), .Z(
        P1_U3522) );
  MUX2_X1 U11146 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9939), .S(n10212), .Z(
        P1_U3521) );
  MUX2_X1 U11147 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9940), .S(n10212), .Z(
        P1_U3519) );
  MUX2_X1 U11148 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9941), .S(n10212), .Z(
        P1_U3518) );
  MUX2_X1 U11149 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9942), .S(n10212), .Z(
        P1_U3517) );
  MUX2_X1 U11150 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9943), .S(n10212), .Z(
        P1_U3516) );
  MUX2_X1 U11151 ( .A(n9944), .B(P1_REG0_REG_24__SCAN_IN), .S(n10211), .Z(
        P1_U3515) );
  MUX2_X1 U11152 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9945), .S(n10212), .Z(
        P1_U3514) );
  MUX2_X1 U11153 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9946), .S(n10212), .Z(
        P1_U3513) );
  MUX2_X1 U11154 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9947), .S(n10212), .Z(
        P1_U3512) );
  MUX2_X1 U11155 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9948), .S(n10212), .Z(
        P1_U3511) );
  MUX2_X1 U11156 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9949), .S(n10212), .Z(
        P1_U3510) );
  MUX2_X1 U11157 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9950), .S(n10212), .Z(
        P1_U3508) );
  MUX2_X1 U11158 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9951), .S(n10212), .Z(
        P1_U3505) );
  MUX2_X1 U11159 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9952), .S(n10212), .Z(
        P1_U3502) );
  MUX2_X1 U11160 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9953), .S(n10212), .Z(
        P1_U3499) );
  MUX2_X1 U11161 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9954), .S(n10212), .Z(
        P1_U3496) );
  MUX2_X1 U11162 ( .A(n9955), .B(P1_REG0_REG_13__SCAN_IN), .S(n10211), .Z(
        P1_U3493) );
  MUX2_X1 U11163 ( .A(n9957), .B(P1_D_REG_0__SCAN_IN), .S(n9956), .Z(P1_U3440)
         );
  NAND3_X1 U11164 ( .A1(n8774), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9959) );
  OAI22_X1 U11165 ( .A1(n9958), .A2(n9959), .B1(n5927), .B2(n9968), .ZN(n9960)
         );
  AOI21_X1 U11166 ( .B1(n8092), .B2(n9961), .A(n9960), .ZN(n9962) );
  INV_X1 U11167 ( .A(n9962), .ZN(P1_U3322) );
  OAI222_X1 U11168 ( .A1(n9968), .A2(n9965), .B1(P1_U3084), .B2(n9964), .C1(
        n9971), .C2(n9963), .ZN(P1_U3324) );
  OAI222_X1 U11169 ( .A1(n9968), .A2(n9967), .B1(P1_U3084), .B2(n10065), .C1(
        n9971), .C2(n9966), .ZN(P1_U3326) );
  OAI222_X1 U11170 ( .A1(n9973), .A2(P1_U3084), .B1(n9971), .B2(n9970), .C1(
        n9969), .C2(n9968), .ZN(P1_U3327) );
  MUX2_X1 U11171 ( .A(n9974), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U11172 ( .A1(n10231), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9985) );
  NAND2_X1 U11173 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9977) );
  AOI211_X1 U11174 ( .C1(n9977), .C2(n9976), .A(n9975), .B(n9986), .ZN(n9978)
         );
  AOI21_X1 U11175 ( .B1(n9992), .B2(n9979), .A(n9978), .ZN(n9984) );
  INV_X1 U11176 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10410) );
  NOR2_X1 U11177 ( .A1(n4830), .A2(n10410), .ZN(n9982) );
  OAI211_X1 U11178 ( .C1(n9982), .C2(n9981), .A(n10224), .B(n9980), .ZN(n9983)
         );
  NAND3_X1 U11179 ( .A1(n9985), .A2(n9984), .A3(n9983), .ZN(P2_U3246) );
  AOI22_X1 U11180 ( .A1(n10231), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9998) );
  AOI211_X1 U11181 ( .C1(n9989), .C2(n9988), .A(n9987), .B(n9986), .ZN(n9990)
         );
  AOI21_X1 U11182 ( .B1(n9992), .B2(n9991), .A(n9990), .ZN(n9997) );
  OAI211_X1 U11183 ( .C1(n9995), .C2(n9994), .A(n10224), .B(n9993), .ZN(n9996)
         );
  NAND3_X1 U11184 ( .A1(n9998), .A2(n9997), .A3(n9996), .ZN(P2_U3247) );
  NAND2_X1 U11185 ( .A1(n10001), .A2(n10000), .ZN(n10002) );
  NAND2_X1 U11186 ( .A1(n10003), .A2(n10002), .ZN(n10004) );
  AOI21_X1 U11187 ( .B1(n10005), .B2(n10210), .A(n10004), .ZN(n10006) );
  AND2_X1 U11188 ( .A1(n10007), .A2(n10006), .ZN(n10009) );
  AOI22_X1 U11189 ( .A1(n10212), .A2(n10009), .B1(n10008), .B2(n10211), .ZN(
        P1_U3484) );
  AOI22_X1 U11190 ( .A1(n10223), .A2(n10009), .B1(n6091), .B2(n10220), .ZN(
        P1_U3533) );
  OAI21_X1 U11191 ( .B1(n10011), .B2(n10400), .A(n10010), .ZN(n10012) );
  AOI211_X1 U11192 ( .C1(n10014), .C2(n10407), .A(n10013), .B(n10012), .ZN(
        n10039) );
  AOI22_X1 U11193 ( .A1(n10430), .A2(n10039), .B1(n8070), .B2(n10427), .ZN(
        P2_U3537) );
  INV_X1 U11194 ( .A(n10380), .ZN(n10390) );
  INV_X1 U11195 ( .A(n10015), .ZN(n10016) );
  OAI22_X1 U11196 ( .A1(n10017), .A2(n10402), .B1(n10016), .B2(n10400), .ZN(
        n10019) );
  AOI211_X1 U11197 ( .C1(n10390), .C2(n10020), .A(n10019), .B(n10018), .ZN(
        n10040) );
  AOI22_X1 U11198 ( .A1(n10430), .A2(n10040), .B1(n7238), .B2(n10427), .ZN(
        P2_U3536) );
  OAI22_X1 U11199 ( .A1(n10022), .A2(n10402), .B1(n10021), .B2(n10400), .ZN(
        n10023) );
  AOI211_X1 U11200 ( .C1(n10025), .C2(n10407), .A(n10024), .B(n10023), .ZN(
        n10041) );
  INV_X1 U11201 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10026) );
  AOI22_X1 U11202 ( .A1(n10430), .A2(n10041), .B1(n10026), .B2(n10427), .ZN(
        P2_U3535) );
  OAI22_X1 U11203 ( .A1(n10028), .A2(n10402), .B1(n10027), .B2(n10400), .ZN(
        n10029) );
  AOI211_X1 U11204 ( .C1(n10031), .C2(n10407), .A(n10030), .B(n10029), .ZN(
        n10042) );
  AOI22_X1 U11205 ( .A1(n10430), .A2(n10042), .B1(n10032), .B2(n10427), .ZN(
        P2_U3534) );
  OAI22_X1 U11206 ( .A1(n10034), .A2(n10402), .B1(n10033), .B2(n10400), .ZN(
        n10036) );
  AOI211_X1 U11207 ( .C1(n10390), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        n10043) );
  AOI22_X1 U11208 ( .A1(n10430), .A2(n10043), .B1(n10038), .B2(n10427), .ZN(
        P2_U3533) );
  AOI22_X1 U11209 ( .A1(n10409), .A2(n10039), .B1(n5488), .B2(n10408), .ZN(
        P2_U3502) );
  AOI22_X1 U11210 ( .A1(n10409), .A2(n10040), .B1(n5471), .B2(n10408), .ZN(
        P2_U3499) );
  AOI22_X1 U11211 ( .A1(n10409), .A2(n10041), .B1(n5456), .B2(n10408), .ZN(
        P2_U3496) );
  AOI22_X1 U11212 ( .A1(n10409), .A2(n10042), .B1(n5441), .B2(n10408), .ZN(
        P2_U3493) );
  AOI22_X1 U11213 ( .A1(n10409), .A2(n10043), .B1(n5426), .B2(n10408), .ZN(
        P2_U3490) );
  INV_X1 U11214 ( .A(n10044), .ZN(n10049) );
  OAI21_X1 U11215 ( .B1(n10046), .B2(n10204), .A(n10045), .ZN(n10048) );
  AOI211_X1 U11216 ( .C1(n10210), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        n10059) );
  AOI22_X1 U11217 ( .A1(n10223), .A2(n10059), .B1(n10050), .B2(n10220), .ZN(
        P1_U3535) );
  INV_X1 U11218 ( .A(n10051), .ZN(n10056) );
  OAI21_X1 U11219 ( .B1(n10053), .B2(n10204), .A(n10052), .ZN(n10055) );
  AOI211_X1 U11220 ( .C1(n10210), .C2(n10056), .A(n10055), .B(n10054), .ZN(
        n10061) );
  AOI22_X1 U11221 ( .A1(n10223), .A2(n10061), .B1(n10057), .B2(n10220), .ZN(
        P1_U3534) );
  INV_X1 U11222 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10058) );
  AOI22_X1 U11223 ( .A1(n10212), .A2(n10059), .B1(n10058), .B2(n10211), .ZN(
        P1_U3490) );
  INV_X1 U11224 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10060) );
  AOI22_X1 U11225 ( .A1(n10212), .A2(n10061), .B1(n10060), .B2(n10211), .ZN(
        P1_U3487) );
  XNOR2_X1 U11226 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11227 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI22_X1 U11228 ( .A1(n10063), .A2(n10435), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10062), .ZN(n10064) );
  INV_X1 U11229 ( .A(n10064), .ZN(n10074) );
  INV_X1 U11230 ( .A(P1_U3083), .ZN(n10070) );
  AOI21_X1 U11231 ( .B1(n10065), .B2(n10071), .A(P1_IR_REG_0__SCAN_IN), .ZN(
        n10067) );
  OAI211_X1 U11232 ( .C1(n10068), .C2(n10067), .A(n10066), .B(
        P1_STATE_REG_SCAN_IN), .ZN(n10069) );
  OR2_X1 U11233 ( .A1(n10070), .A2(n10069), .ZN(n10073) );
  NAND3_X1 U11234 ( .A1(n10120), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10071), .ZN(
        n10072) );
  NAND3_X1 U11235 ( .A1(n10074), .A2(n10073), .A3(n10072), .ZN(P1_U3241) );
  AOI211_X1 U11236 ( .C1(n10077), .C2(n10076), .A(n10075), .B(n10106), .ZN(
        n10078) );
  AOI211_X1 U11237 ( .C1(n10118), .C2(n10080), .A(n10079), .B(n10078), .ZN(
        n10086) );
  OAI21_X1 U11238 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(n10084) );
  AOI22_X1 U11239 ( .A1(n10124), .A2(n10084), .B1(n10122), .B2(
        P1_ADDR_REG_5__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U11240 ( .A1(n10086), .A2(n10085), .ZN(P1_U3246) );
  MUX2_X1 U11241 ( .A(n5999), .B(P1_REG1_REG_6__SCAN_IN), .S(n10098), .Z(
        n10087) );
  INV_X1 U11242 ( .A(n10087), .ZN(n10090) );
  OAI21_X1 U11243 ( .B1(n10090), .B2(n10089), .A(n10088), .ZN(n10097) );
  OAI211_X1 U11244 ( .C1(n10093), .C2(n10092), .A(n10124), .B(n10091), .ZN(
        n10094) );
  INV_X1 U11245 ( .A(n10094), .ZN(n10095) );
  AOI211_X1 U11246 ( .C1(n10120), .C2(n10097), .A(n10096), .B(n10095), .ZN(
        n10100) );
  AOI22_X1 U11247 ( .A1(n10118), .A2(n10098), .B1(n10122), .B2(
        P1_ADDR_REG_6__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U11248 ( .A1(n10100), .A2(n10099), .ZN(P1_U3247) );
  AOI22_X1 U11249 ( .A1(n10118), .A2(n10101), .B1(n10122), .B2(
        P1_ADDR_REG_10__SCAN_IN), .ZN(n10114) );
  INV_X1 U11250 ( .A(n10102), .ZN(n10113) );
  AOI21_X1 U11251 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(n10107) );
  OR2_X1 U11252 ( .A1(n10107), .A2(n10106), .ZN(n10112) );
  OAI211_X1 U11253 ( .C1(n10110), .C2(n10109), .A(n10124), .B(n10108), .ZN(
        n10111) );
  NAND4_X1 U11254 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        P1_U3251) );
  INV_X1 U11255 ( .A(n10115), .ZN(n10116) );
  AOI21_X1 U11256 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(n10129) );
  OAI211_X1 U11257 ( .C1(n10121), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10120), 
        .B(n10119), .ZN(n10128) );
  NAND2_X1 U11258 ( .A1(n10122), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n10127) );
  OAI211_X1 U11259 ( .C1(n10125), .C2(P1_REG2_REG_15__SCAN_IN), .A(n10124), 
        .B(n10123), .ZN(n10126) );
  NAND4_X1 U11260 ( .A1(n10129), .A2(n10128), .A3(n10127), .A4(n10126), .ZN(
        P1_U3256) );
  OAI21_X1 U11261 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n10169) );
  XNOR2_X1 U11262 ( .A(n10134), .B(n10133), .ZN(n10136) );
  NAND2_X1 U11263 ( .A1(n10136), .A2(n10135), .ZN(n10142) );
  AOI22_X1 U11264 ( .A1(n10140), .A2(n10139), .B1(n10138), .B2(n10137), .ZN(
        n10141) );
  OAI211_X1 U11265 ( .C1(n10169), .C2(n10143), .A(n10142), .B(n10141), .ZN(
        n10172) );
  NOR2_X1 U11266 ( .A1(n10169), .A2(n10144), .ZN(n10154) );
  OAI211_X1 U11267 ( .C1(n10147), .C2(n10171), .A(n10146), .B(n10145), .ZN(
        n10170) );
  NOR2_X1 U11268 ( .A1(n10170), .A2(n10148), .ZN(n10153) );
  OAI22_X1 U11269 ( .A1(n10171), .A2(n6208), .B1(n10151), .B2(n10150), .ZN(
        n10152) );
  NOR4_X1 U11270 ( .A1(n10172), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10155) );
  AOI22_X1 U11271 ( .A1(n10157), .A2(n10156), .B1(n10155), .B2(n9810), .ZN(
        P1_U3290) );
  AND2_X1 U11272 ( .A1(n10159), .A2(n10158), .ZN(n10168) );
  AND2_X1 U11273 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10165), .ZN(P1_U3292) );
  NOR2_X1 U11274 ( .A1(n10168), .A2(n10160), .ZN(P1_U3293) );
  AND2_X1 U11275 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10165), .ZN(P1_U3294) );
  NOR2_X1 U11276 ( .A1(n10168), .A2(n10161), .ZN(P1_U3295) );
  AND2_X1 U11277 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10165), .ZN(P1_U3296) );
  AND2_X1 U11278 ( .A1(n10165), .A2(P1_D_REG_26__SCAN_IN), .ZN(P1_U3297) );
  AND2_X1 U11279 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10165), .ZN(P1_U3298) );
  AND2_X1 U11280 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10165), .ZN(P1_U3299) );
  NOR2_X1 U11281 ( .A1(n10168), .A2(n10162), .ZN(P1_U3300) );
  AND2_X1 U11282 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10165), .ZN(P1_U3301) );
  NOR2_X1 U11283 ( .A1(n10168), .A2(n10163), .ZN(P1_U3302) );
  AND2_X1 U11284 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10165), .ZN(P1_U3303) );
  AND2_X1 U11285 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10165), .ZN(P1_U3304) );
  AND2_X1 U11286 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10165), .ZN(P1_U3305) );
  AND2_X1 U11287 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10165), .ZN(P1_U3306) );
  NOR2_X1 U11288 ( .A1(n10168), .A2(n10164), .ZN(P1_U3307) );
  AND2_X1 U11289 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10165), .ZN(P1_U3308) );
  AND2_X1 U11290 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10165), .ZN(P1_U3309) );
  AND2_X1 U11291 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10165), .ZN(P1_U3310) );
  AND2_X1 U11292 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10165), .ZN(P1_U3311) );
  AND2_X1 U11293 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10165), .ZN(P1_U3312) );
  AND2_X1 U11294 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10165), .ZN(P1_U3313) );
  AND2_X1 U11295 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10165), .ZN(P1_U3314) );
  AND2_X1 U11296 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10165), .ZN(P1_U3315) );
  AND2_X1 U11297 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10165), .ZN(P1_U3316) );
  AND2_X1 U11298 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10165), .ZN(P1_U3317) );
  AND2_X1 U11299 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10165), .ZN(P1_U3318) );
  AND2_X1 U11300 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10165), .ZN(P1_U3319) );
  NOR2_X1 U11301 ( .A1(n10168), .A2(n10166), .ZN(P1_U3320) );
  NOR2_X1 U11302 ( .A1(n10168), .A2(n10167), .ZN(P1_U3321) );
  INV_X1 U11303 ( .A(n10169), .ZN(n10174) );
  OAI21_X1 U11304 ( .B1(n10171), .B2(n10204), .A(n10170), .ZN(n10173) );
  AOI211_X1 U11305 ( .C1(n10210), .C2(n10174), .A(n10173), .B(n10172), .ZN(
        n10214) );
  INV_X1 U11306 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U11307 ( .A1(n10212), .A2(n10214), .B1(n10175), .B2(n10211), .ZN(
        P1_U3457) );
  OAI22_X1 U11308 ( .A1(n10177), .A2(n10205), .B1(n10176), .B2(n10204), .ZN(
        n10179) );
  AOI211_X1 U11309 ( .C1(n10210), .C2(n10180), .A(n10179), .B(n10178), .ZN(
        n10216) );
  INV_X1 U11310 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U11311 ( .A1(n10212), .A2(n10216), .B1(n10181), .B2(n10211), .ZN(
        P1_U3460) );
  OAI22_X1 U11312 ( .A1(n10183), .A2(n10205), .B1(n10182), .B2(n10204), .ZN(
        n10185) );
  AOI211_X1 U11313 ( .C1(n10210), .C2(n10186), .A(n10185), .B(n10184), .ZN(
        n10217) );
  INV_X1 U11314 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U11315 ( .A1(n10212), .A2(n10217), .B1(n10187), .B2(n10211), .ZN(
        P1_U3466) );
  OAI211_X1 U11316 ( .C1(n10190), .C2(n10204), .A(n10189), .B(n10188), .ZN(
        n10192) );
  AOI211_X1 U11317 ( .C1(n10194), .C2(n10193), .A(n10192), .B(n10191), .ZN(
        n10218) );
  AOI22_X1 U11318 ( .A1(n10212), .A2(n10218), .B1(n6558), .B2(n10211), .ZN(
        P1_U3469) );
  INV_X1 U11319 ( .A(n10195), .ZN(n10200) );
  OAI22_X1 U11320 ( .A1(n10197), .A2(n10205), .B1(n10196), .B2(n10204), .ZN(
        n10199) );
  AOI211_X1 U11321 ( .C1(n10210), .C2(n10200), .A(n10199), .B(n10198), .ZN(
        n10219) );
  INV_X1 U11322 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U11323 ( .A1(n10212), .A2(n10219), .B1(n10201), .B2(n10211), .ZN(
        P1_U3478) );
  INV_X1 U11324 ( .A(n10202), .ZN(n10209) );
  OAI22_X1 U11325 ( .A1(n10206), .A2(n10205), .B1(n4748), .B2(n10204), .ZN(
        n10208) );
  AOI211_X1 U11326 ( .C1(n10210), .C2(n10209), .A(n10208), .B(n10207), .ZN(
        n10222) );
  AOI22_X1 U11327 ( .A1(n10212), .A2(n10222), .B1(n6923), .B2(n10211), .ZN(
        P1_U3481) );
  AOI22_X1 U11328 ( .A1(n10223), .A2(n10214), .B1(n10213), .B2(n10220), .ZN(
        P1_U3524) );
  AOI22_X1 U11329 ( .A1(n10223), .A2(n10216), .B1(n10215), .B2(n10220), .ZN(
        P1_U3525) );
  AOI22_X1 U11330 ( .A1(n10223), .A2(n10217), .B1(n6528), .B2(n10220), .ZN(
        P1_U3527) );
  AOI22_X1 U11331 ( .A1(n10223), .A2(n10218), .B1(n6556), .B2(n10220), .ZN(
        P1_U3528) );
  AOI22_X1 U11332 ( .A1(n10223), .A2(n10219), .B1(n6379), .B2(n10220), .ZN(
        P1_U3531) );
  AOI22_X1 U11333 ( .A1(n10223), .A2(n10222), .B1(n10221), .B2(n10220), .ZN(
        P1_U3532) );
  AOI22_X1 U11334 ( .A1(n10226), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10224), .ZN(n10234) );
  NAND2_X1 U11335 ( .A1(n10226), .A2(n10225), .ZN(n10228) );
  OAI211_X1 U11336 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10229), .A(n10228), .B(
        n10227), .ZN(n10230) );
  INV_X1 U11337 ( .A(n10230), .ZN(n10233) );
  AOI22_X1 U11338 ( .A1(n10231), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10232) );
  OAI221_X1 U11339 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10234), .C1(n4830), .C2(
        n10233), .A(n10232), .ZN(P2_U3245) );
  XNOR2_X1 U11340 ( .A(n10235), .B(n10236), .ZN(n10243) );
  NAND2_X1 U11341 ( .A1(n10237), .A2(n10236), .ZN(n10238) );
  NAND2_X1 U11342 ( .A1(n10239), .A2(n10238), .ZN(n10379) );
  OAI21_X1 U11343 ( .B1(n10379), .B2(n10241), .A(n10240), .ZN(n10242) );
  AOI21_X1 U11344 ( .B1(n10264), .B2(n10243), .A(n10242), .ZN(n10378) );
  AOI222_X1 U11345 ( .A1(n10375), .A2(n10302), .B1(P2_REG2_REG_8__SCAN_IN), 
        .B2(n10308), .C1(n10245), .C2(n10244), .ZN(n10254) );
  INV_X1 U11346 ( .A(n10379), .ZN(n10252) );
  NAND2_X1 U11347 ( .A1(n10246), .A2(n10375), .ZN(n10247) );
  NAND2_X1 U11348 ( .A1(n10247), .A2(n10295), .ZN(n10248) );
  NOR2_X1 U11349 ( .A1(n10249), .A2(n10248), .ZN(n10374) );
  AOI22_X1 U11350 ( .A1(n10252), .A2(n10251), .B1(n10250), .B2(n10374), .ZN(
        n10253) );
  OAI211_X1 U11351 ( .C1(n10308), .C2(n10378), .A(n10254), .B(n10253), .ZN(
        P2_U3288) );
  NAND3_X1 U11352 ( .A1(n10255), .A2(n10265), .A3(n10256), .ZN(n10257) );
  NAND2_X1 U11353 ( .A1(n10258), .A2(n10257), .ZN(n10263) );
  AOI222_X1 U11354 ( .A1(n10264), .A2(n10263), .B1(n10262), .B2(n10261), .C1(
        n10260), .C2(n10259), .ZN(n10363) );
  XNOR2_X1 U11355 ( .A(n10266), .B(n10265), .ZN(n10366) );
  XNOR2_X1 U11356 ( .A(n10267), .B(n10361), .ZN(n10362) );
  INV_X1 U11357 ( .A(n10268), .ZN(n10269) );
  OAI22_X1 U11358 ( .A1(n10299), .A2(n5318), .B1(n10269), .B2(n10297), .ZN(
        n10270) );
  AOI21_X1 U11359 ( .B1(n10302), .B2(n10271), .A(n10270), .ZN(n10272) );
  OAI21_X1 U11360 ( .B1(n10273), .B2(n10362), .A(n10272), .ZN(n10274) );
  AOI21_X1 U11361 ( .B1(n10366), .B2(n10306), .A(n10274), .ZN(n10275) );
  OAI21_X1 U11362 ( .B1(n10308), .B2(n10363), .A(n10275), .ZN(P2_U3290) );
  INV_X1 U11363 ( .A(n10276), .ZN(n10283) );
  INV_X1 U11364 ( .A(n10291), .ZN(n10277) );
  AOI21_X1 U11365 ( .B1(n10279), .B2(n10278), .A(n10277), .ZN(n10280) );
  AOI211_X1 U11366 ( .C1(n10283), .C2(n10282), .A(n10281), .B(n10280), .ZN(
        n10289) );
  OAI22_X1 U11367 ( .A1(n10287), .A2(n10286), .B1(n10285), .B2(n10284), .ZN(
        n10288) );
  NOR2_X1 U11368 ( .A1(n10289), .A2(n10288), .ZN(n10350) );
  XNOR2_X1 U11369 ( .A(n10290), .B(n10291), .ZN(n10353) );
  OAI21_X1 U11370 ( .B1(n10293), .B2(n10292), .A(n10301), .ZN(n10296) );
  NAND3_X1 U11371 ( .A1(n10296), .A2(n10295), .A3(n10294), .ZN(n10349) );
  OAI22_X1 U11372 ( .A1(n10299), .A2(n5285), .B1(n10298), .B2(n10297), .ZN(
        n10300) );
  AOI21_X1 U11373 ( .B1(n10302), .B2(n10301), .A(n10300), .ZN(n10303) );
  OAI21_X1 U11374 ( .B1(n10304), .B2(n10349), .A(n10303), .ZN(n10305) );
  AOI21_X1 U11375 ( .B1(n10306), .B2(n10353), .A(n10305), .ZN(n10307) );
  OAI21_X1 U11376 ( .B1(n10308), .B2(n10350), .A(n10307), .ZN(P2_U3292) );
  AND2_X1 U11377 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10322), .ZN(P2_U3297) );
  AND2_X1 U11378 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10322), .ZN(P2_U3298) );
  AND2_X1 U11379 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10322), .ZN(P2_U3299) );
  AND2_X1 U11380 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10322), .ZN(P2_U3300) );
  NOR2_X1 U11381 ( .A1(n10319), .A2(n10311), .ZN(P2_U3301) );
  AND2_X1 U11382 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10322), .ZN(P2_U3302) );
  AND2_X1 U11383 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10322), .ZN(P2_U3303) );
  AND2_X1 U11384 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10322), .ZN(P2_U3304) );
  NOR2_X1 U11385 ( .A1(n10319), .A2(n10312), .ZN(P2_U3305) );
  AND2_X1 U11386 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10322), .ZN(P2_U3306) );
  AND2_X1 U11387 ( .A1(n10322), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3307) );
  AND2_X1 U11388 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10322), .ZN(P2_U3308) );
  AND2_X1 U11389 ( .A1(n10322), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3309) );
  AND2_X1 U11390 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10322), .ZN(P2_U3310) );
  AND2_X1 U11391 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10322), .ZN(P2_U3311) );
  AND2_X1 U11392 ( .A1(n10322), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3312) );
  AND2_X1 U11393 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10322), .ZN(P2_U3313) );
  AND2_X1 U11394 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10322), .ZN(P2_U3314) );
  NOR2_X1 U11395 ( .A1(n10319), .A2(n10313), .ZN(P2_U3315) );
  NOR2_X1 U11396 ( .A1(n10319), .A2(n10314), .ZN(P2_U3316) );
  AND2_X1 U11397 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10322), .ZN(P2_U3317) );
  NOR2_X1 U11398 ( .A1(n10319), .A2(n10315), .ZN(P2_U3318) );
  AND2_X1 U11399 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10322), .ZN(P2_U3319) );
  AND2_X1 U11400 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10322), .ZN(P2_U3320) );
  AND2_X1 U11401 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10322), .ZN(P2_U3321) );
  AND2_X1 U11402 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10322), .ZN(P2_U3322) );
  NOR2_X1 U11403 ( .A1(n10319), .A2(n10316), .ZN(P2_U3323) );
  NOR2_X1 U11404 ( .A1(n10319), .A2(n10317), .ZN(P2_U3324) );
  AND2_X1 U11405 ( .A1(n10322), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3325) );
  NOR2_X1 U11406 ( .A1(n10319), .A2(n10318), .ZN(P2_U3326) );
  AOI22_X1 U11407 ( .A1(n10321), .A2(n10322), .B1(n10325), .B2(n10320), .ZN(
        P2_U3437) );
  AOI22_X1 U11408 ( .A1(n10325), .A2(n10324), .B1(n10323), .B2(n10322), .ZN(
        P2_U3438) );
  OAI22_X1 U11409 ( .A1(n10328), .A2(n10327), .B1(n4834), .B2(n10326), .ZN(
        n10329) );
  NOR2_X1 U11410 ( .A1(n10330), .A2(n10329), .ZN(n10411) );
  AOI22_X1 U11411 ( .A1(n10409), .A2(n10411), .B1(n5230), .B2(n10408), .ZN(
        P2_U3451) );
  INV_X1 U11412 ( .A(n10331), .ZN(n10337) );
  OAI21_X1 U11413 ( .B1(n10400), .B2(n10333), .A(n10332), .ZN(n10336) );
  INV_X1 U11414 ( .A(n10334), .ZN(n10335) );
  AOI211_X1 U11415 ( .C1(n10407), .C2(n10337), .A(n10336), .B(n10335), .ZN(
        n10413) );
  AOI22_X1 U11416 ( .A1(n10409), .A2(n10413), .B1(n5236), .B2(n10408), .ZN(
        P2_U3454) );
  OAI22_X1 U11417 ( .A1(n10339), .A2(n10402), .B1(n10338), .B2(n10400), .ZN(
        n10341) );
  AOI211_X1 U11418 ( .C1(n10407), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        n10415) );
  AOI22_X1 U11419 ( .A1(n10409), .A2(n10415), .B1(n5255), .B2(n10408), .ZN(
        P2_U3457) );
  OAI21_X1 U11420 ( .B1(n10344), .B2(n10400), .A(n10343), .ZN(n10347) );
  INV_X1 U11421 ( .A(n10345), .ZN(n10346) );
  AOI211_X1 U11422 ( .C1(n10390), .C2(n10348), .A(n10347), .B(n10346), .ZN(
        n10416) );
  AOI22_X1 U11423 ( .A1(n10409), .A2(n10416), .B1(n5270), .B2(n10408), .ZN(
        P2_U3460) );
  OAI211_X1 U11424 ( .C1(n10351), .C2(n10400), .A(n10350), .B(n10349), .ZN(
        n10352) );
  AOI21_X1 U11425 ( .B1(n10407), .B2(n10353), .A(n10352), .ZN(n10417) );
  AOI22_X1 U11426 ( .A1(n10409), .A2(n10417), .B1(n5284), .B2(n10408), .ZN(
        P2_U3463) );
  OAI21_X1 U11427 ( .B1(n10355), .B2(n10400), .A(n10354), .ZN(n10356) );
  INV_X1 U11428 ( .A(n10356), .ZN(n10359) );
  NAND2_X1 U11429 ( .A1(n10357), .A2(n10407), .ZN(n10358) );
  AOI22_X1 U11430 ( .A1(n10409), .A2(n10418), .B1(n5298), .B2(n10408), .ZN(
        P2_U3466) );
  OAI22_X1 U11431 ( .A1(n10362), .A2(n10402), .B1(n10361), .B2(n10400), .ZN(
        n10365) );
  INV_X1 U11432 ( .A(n10363), .ZN(n10364) );
  AOI211_X1 U11433 ( .C1(n10407), .C2(n10366), .A(n10365), .B(n10364), .ZN(
        n10419) );
  AOI22_X1 U11434 ( .A1(n10409), .A2(n10419), .B1(n5317), .B2(n10408), .ZN(
        P2_U3469) );
  OR2_X1 U11435 ( .A1(n10367), .A2(n10400), .ZN(n10368) );
  AND2_X1 U11436 ( .A1(n10369), .A2(n10368), .ZN(n10372) );
  NAND2_X1 U11437 ( .A1(n10370), .A2(n10407), .ZN(n10371) );
  AND3_X1 U11438 ( .A1(n10373), .A2(n10372), .A3(n10371), .ZN(n10420) );
  AOI22_X1 U11439 ( .A1(n10409), .A2(n10420), .B1(n5341), .B2(n10408), .ZN(
        P2_U3472) );
  AOI21_X1 U11440 ( .B1(n10376), .B2(n10375), .A(n10374), .ZN(n10377) );
  OAI211_X1 U11441 ( .C1(n10380), .C2(n10379), .A(n10378), .B(n10377), .ZN(
        n10381) );
  INV_X1 U11442 ( .A(n10381), .ZN(n10422) );
  AOI22_X1 U11443 ( .A1(n10409), .A2(n10422), .B1(n5353), .B2(n10408), .ZN(
        P2_U3475) );
  OAI21_X1 U11444 ( .B1(n10383), .B2(n10400), .A(n10382), .ZN(n10385) );
  AOI211_X1 U11445 ( .C1(n10390), .C2(n10386), .A(n10385), .B(n10384), .ZN(
        n10423) );
  AOI22_X1 U11446 ( .A1(n10409), .A2(n10423), .B1(n5368), .B2(n10408), .ZN(
        P2_U3478) );
  OAI22_X1 U11447 ( .A1(n10388), .A2(n10402), .B1(n10387), .B2(n10400), .ZN(
        n10389) );
  AOI21_X1 U11448 ( .B1(n10391), .B2(n10390), .A(n10389), .ZN(n10392) );
  AOI22_X1 U11449 ( .A1(n10409), .A2(n10424), .B1(n5386), .B2(n10408), .ZN(
        P2_U3481) );
  INV_X1 U11450 ( .A(n10394), .ZN(n10399) );
  OAI22_X1 U11451 ( .A1(n10396), .A2(n10402), .B1(n10395), .B2(n10400), .ZN(
        n10398) );
  AOI211_X1 U11452 ( .C1(n10399), .C2(n10407), .A(n10398), .B(n10397), .ZN(
        n10426) );
  AOI22_X1 U11453 ( .A1(n10409), .A2(n10426), .B1(n5398), .B2(n10408), .ZN(
        P2_U3484) );
  OAI22_X1 U11454 ( .A1(n10403), .A2(n10402), .B1(n10401), .B2(n10400), .ZN(
        n10405) );
  AOI211_X1 U11455 ( .C1(n10407), .C2(n10406), .A(n10405), .B(n10404), .ZN(
        n10429) );
  AOI22_X1 U11456 ( .A1(n10409), .A2(n10429), .B1(n5414), .B2(n10408), .ZN(
        P2_U3487) );
  AOI22_X1 U11457 ( .A1(n10430), .A2(n10411), .B1(n10410), .B2(n10427), .ZN(
        P2_U3520) );
  AOI22_X1 U11458 ( .A1(n10430), .A2(n10413), .B1(n10412), .B2(n10427), .ZN(
        P2_U3521) );
  AOI22_X1 U11459 ( .A1(n10430), .A2(n10415), .B1(n10414), .B2(n10427), .ZN(
        P2_U3522) );
  AOI22_X1 U11460 ( .A1(n10430), .A2(n10416), .B1(n6048), .B2(n10427), .ZN(
        P2_U3523) );
  AOI22_X1 U11461 ( .A1(n10430), .A2(n10417), .B1(n6047), .B2(n10427), .ZN(
        P2_U3524) );
  AOI22_X1 U11462 ( .A1(n10430), .A2(n10418), .B1(n6046), .B2(n10427), .ZN(
        P2_U3525) );
  AOI22_X1 U11463 ( .A1(n10430), .A2(n10419), .B1(n6045), .B2(n10427), .ZN(
        P2_U3526) );
  AOI22_X1 U11464 ( .A1(n10430), .A2(n10420), .B1(n6044), .B2(n10427), .ZN(
        P2_U3527) );
  AOI22_X1 U11465 ( .A1(n10430), .A2(n10422), .B1(n10421), .B2(n10427), .ZN(
        P2_U3528) );
  AOI22_X1 U11466 ( .A1(n10430), .A2(n10423), .B1(n6325), .B2(n10427), .ZN(
        P2_U3529) );
  AOI22_X1 U11467 ( .A1(n10430), .A2(n10424), .B1(n6330), .B2(n10427), .ZN(
        P2_U3530) );
  AOI22_X1 U11468 ( .A1(n10430), .A2(n10426), .B1(n10425), .B2(n10427), .ZN(
        P2_U3531) );
  AOI22_X1 U11469 ( .A1(n10430), .A2(n10429), .B1(n10428), .B2(n10427), .ZN(
        P2_U3532) );
  INV_X1 U11470 ( .A(n10431), .ZN(n10432) );
  NAND2_X1 U11471 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  XNOR2_X1 U11472 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10434), .ZN(ADD_1071_U5)
         );
  INV_X1 U11473 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U11474 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10436), .B2(n10435), .ZN(ADD_1071_U46) );
  OAI21_X1 U11475 ( .B1(n10439), .B2(n10438), .A(n10437), .ZN(ADD_1071_U56) );
  OAI21_X1 U11476 ( .B1(n10442), .B2(n10441), .A(n10440), .ZN(ADD_1071_U57) );
  OAI21_X1 U11477 ( .B1(n10445), .B2(n10444), .A(n10443), .ZN(ADD_1071_U58) );
  OAI21_X1 U11478 ( .B1(n10448), .B2(n10447), .A(n10446), .ZN(ADD_1071_U59) );
  OAI21_X1 U11479 ( .B1(n10451), .B2(n10450), .A(n10449), .ZN(ADD_1071_U60) );
  OAI21_X1 U11480 ( .B1(n10454), .B2(n10453), .A(n10452), .ZN(ADD_1071_U61) );
  AOI21_X1 U11481 ( .B1(n10457), .B2(n10456), .A(n10455), .ZN(ADD_1071_U62) );
  AOI21_X1 U11482 ( .B1(n10460), .B2(n10459), .A(n10458), .ZN(ADD_1071_U63) );
  XOR2_X1 U11483 ( .A(n10461), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U11484 ( .A(n10463), .B(n10462), .Z(ADD_1071_U54) );
  NOR2_X1 U11485 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  XOR2_X1 U11486 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10466), .Z(ADD_1071_U51) );
  OAI21_X1 U11487 ( .B1(n10469), .B2(n10468), .A(n10467), .ZN(n10470) );
  XNOR2_X1 U11488 ( .A(n10470), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11489 ( .B1(n10473), .B2(n10472), .A(n10471), .ZN(ADD_1071_U47) );
  XOR2_X1 U11490 ( .A(n10474), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11491 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10475), .Z(ADD_1071_U48) );
  XOR2_X1 U11492 ( .A(n10477), .B(n10476), .Z(ADD_1071_U53) );
  XNOR2_X1 U11493 ( .A(n10479), .B(n10478), .ZN(ADD_1071_U52) );
  BUF_X1 U4984 ( .A(n6433), .Z(n4476) );
  INV_X1 U4983 ( .A(n4476), .ZN(n7992) );
  CLKBUF_X1 U5202 ( .A(n6506), .Z(n8094) );
  CLKBUF_X1 U5752 ( .A(n5903), .Z(n5915) );
endmodule

