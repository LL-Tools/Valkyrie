

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588;

  NAND2_X1 U4904 ( .A1(n5970), .A2(n5969), .ZN(n8963) );
  OR2_X1 U4905 ( .A1(n7335), .A2(n7334), .ZN(n7374) );
  XNOR2_X1 U4906 ( .A(n4984), .B(n5363), .ZN(n9143) );
  CLKBUF_X2 U4907 ( .A(n8939), .Z(n4840) );
  INV_X1 U4908 ( .A(n5454), .ZN(n8496) );
  OAI21_X1 U4909 ( .B1(n5758), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5779) );
  AND2_X2 U4911 ( .A1(n6151), .A2(n6114), .ZN(n6376) );
  CLKBUF_X1 U4912 ( .A(n9626), .Z(n4839) );
  OAI21_X1 U4913 ( .B1(n7067), .B2(n7065), .A(n10450), .ZN(n9626) );
  AOI21_X2 U4914 ( .B1(n5861), .B2(n5203), .A(n4885), .ZN(n5922) );
  OR2_X2 U4915 ( .A1(n10568), .A2(n9180), .ZN(n7743) );
  INV_X1 U4916 ( .A(n9143), .ZN(n9180) );
  INV_X1 U4917 ( .A(n6659), .ZN(n6642) );
  INV_X1 U4918 ( .A(n8643), .ZN(n8637) );
  INV_X1 U4920 ( .A(n6386), .ZN(n7161) );
  AND2_X1 U4921 ( .A1(n7588), .A2(n7587), .ZN(n7590) );
  INV_X1 U4922 ( .A(n5385), .ZN(n6780) );
  INV_X1 U4923 ( .A(n5452), .ZN(n4845) );
  NAND2_X1 U4924 ( .A1(n5348), .A2(n8423), .ZN(n5452) );
  NAND2_X2 U4925 ( .A1(n6574), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6576) );
  AND2_X2 U4926 ( .A1(n7974), .A2(n8547), .ZN(n7952) );
  OAI22_X2 U4927 ( .A1(n9840), .A2(n9848), .B1(n9867), .B2(n9926), .ZN(n9825)
         );
  OAI22_X2 U4928 ( .A1(n9855), .A2(n8732), .B1(n9624), .B2(n9862), .ZN(n9840)
         );
  NAND4_X2 U4929 ( .A1(n5459), .A2(n5329), .A3(n5330), .A4(n5331), .ZN(n5401)
         );
  NOR2_X2 U4930 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5329) );
  AND2_X1 U4931 ( .A1(n7138), .A2(n7031), .ZN(n8939) );
  INV_X4 U4932 ( .A(n6780), .ZN(n6781) );
  CLKBUF_X2 U4933 ( .A(n7096), .Z(n8949) );
  NAND2_X2 U4934 ( .A1(n7125), .A2(n7687), .ZN(n7041) );
  BUF_X1 U4936 ( .A(n6735), .Z(n4848) );
  AND2_X1 U4937 ( .A1(n6341), .A2(n6184), .ZN(n6287) );
  INV_X4 U4938 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OAI21_X1 U4939 ( .B1(n9764), .B2(n4897), .A(n5234), .ZN(n5233) );
  AND2_X1 U4940 ( .A1(n5146), .A2(n5144), .ZN(n9407) );
  AOI21_X1 U4941 ( .B1(n9233), .B2(n8854), .A(n8853), .ZN(n9222) );
  NAND2_X1 U4942 ( .A1(n9265), .A2(n9273), .ZN(n9264) );
  NAND2_X1 U4943 ( .A1(n8262), .A2(n4865), .ZN(n8273) );
  AND2_X1 U4944 ( .A1(n9312), .A2(n9309), .ZN(n8480) );
  OR2_X1 U4945 ( .A1(n8479), .A2(n9335), .ZN(n9309) );
  OAI21_X1 U4946 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(n8713) );
  AND2_X1 U4947 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  OAI21_X1 U4948 ( .B1(n8113), .B2(n5264), .A(n5262), .ZN(n8340) );
  NOR2_X1 U4949 ( .A1(n8329), .A2(n9952), .ZN(n8361) );
  NOR2_X1 U4950 ( .A1(n7865), .A2(n8083), .ZN(n8052) );
  OAI21_X1 U4951 ( .B1(n7317), .B2(n6409), .A(n6681), .ZN(n7525) );
  OR2_X1 U4952 ( .A1(n7102), .A2(n7101), .ZN(n7103) );
  INV_X2 U4953 ( .A(n10542), .ZN(n4842) );
  INV_X2 U4954 ( .A(n10543), .ZN(n4843) );
  XNOR2_X1 U4955 ( .A(n4942), .B(n5578), .ZN(n6824) );
  NAND2_X1 U4956 ( .A1(n5080), .A2(n5079), .ZN(n5730) );
  NOR2_X1 U4957 ( .A1(n7041), .A2(n6668), .ZN(n7136) );
  INV_X1 U4958 ( .A(n8936), .ZN(n8950) );
  AND4_X1 U4959 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n7972)
         );
  NAND2_X1 U4960 ( .A1(n7024), .A2(n7023), .ZN(n7128) );
  INV_X1 U4961 ( .A(n7392), .ZN(n10481) );
  NAND4_X1 U4962 ( .A1(n6403), .A2(n6402), .A3(n6401), .A4(n6400), .ZN(n9663)
         );
  OAI211_X1 U4963 ( .C1(n6751), .C2(n6934), .A(n5421), .B(n5420), .ZN(n10488)
         );
  NAND2_X1 U4964 ( .A1(n5446), .A2(n5445), .ZN(n7392) );
  NAND2_X1 U4965 ( .A1(n4899), .A2(n4854), .ZN(n7354) );
  INV_X1 U4966 ( .A(n8503), .ZN(n5819) );
  NAND2_X1 U4967 ( .A1(n8874), .A2(n8423), .ZN(n5454) );
  INV_X1 U4968 ( .A(n6151), .ZN(n8470) );
  INV_X1 U4969 ( .A(n5347), .ZN(n8423) );
  INV_X1 U4970 ( .A(n6546), .ZN(n6666) );
  NAND2_X2 U4971 ( .A1(n5364), .A2(n8686), .ZN(n10568) );
  XNOR2_X1 U4972 ( .A(n6109), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6151) );
  OR2_X1 U4973 ( .A1(n9501), .A2(n5343), .ZN(n5344) );
  NAND2_X1 U4974 ( .A1(n6734), .A2(n6735), .ZN(n6405) );
  OR2_X1 U4975 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NAND2_X1 U4976 ( .A1(n9991), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U4977 ( .A1(n6287), .A2(n6185), .ZN(n6198) );
  INV_X2 U4978 ( .A(n9507), .ZN(n7477) );
  INV_X2 U4979 ( .A(n9996), .ZN(n7481) );
  XNOR2_X1 U4980 ( .A(n5498), .B(n10163), .ZN(n5496) );
  NOR2_X1 U4981 ( .A1(n5562), .A2(n5354), .ZN(n5638) );
  NAND2_X2 U4982 ( .A1(n6780), .A2(P1_U3084), .ZN(n8841) );
  INV_X2 U4983 ( .A(n6780), .ZN(n6778) );
  AND2_X1 U4984 ( .A1(n5340), .A2(n4864), .ZN(n5153) );
  AND2_X1 U4985 ( .A1(n6097), .A2(n6105), .ZN(n5006) );
  AND4_X1 U4986 ( .A1(n6096), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n6097)
         );
  AND3_X1 U4987 ( .A1(n6088), .A2(n6087), .A3(n6086), .ZN(n6092) );
  NOR2_X1 U4988 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6083) );
  INV_X1 U4989 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6418) );
  INV_X2 U4990 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4991 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5684) );
  INV_X1 U4992 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5582) );
  NOR2_X2 U4993 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5459) );
  INV_X2 U4994 ( .A(n6183), .ZN(n6099) );
  AOI21_X2 U4995 ( .B1(n5261), .B2(n5259), .A(n4895), .ZN(n9284) );
  NAND2_X1 U4996 ( .A1(n9376), .A2(n9386), .ZN(n5261) );
  OAI21_X2 U4997 ( .B1(n5224), .B2(n5222), .A(n5220), .ZN(n9855) );
  AOI21_X2 U4998 ( .B1(n7952), .B2(n7951), .A(n7950), .ZN(n8113) );
  INV_X1 U4999 ( .A(n7743), .ZN(n4844) );
  INV_X4 U5000 ( .A(n4845), .ZN(n4846) );
  XNOR2_X1 U5001 ( .A(n6103), .B(n6102), .ZN(n6734) );
  AND3_X1 U5002 ( .A1(n6367), .A2(n6366), .A3(n6365), .ZN(n7024) );
  XNOR2_X1 U5003 ( .A(n4956), .B(n6105), .ZN(n6735) );
  NAND2_X2 U5004 ( .A1(n6751), .A2(n6778), .ZN(n8503) );
  INV_X1 U5005 ( .A(n6114), .ZN(n8422) );
  NAND2_X4 U5006 ( .A1(n8470), .A2(n6114), .ZN(n6389) );
  XNOR2_X2 U5007 ( .A(n6112), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6114) );
  AND2_X1 U5008 ( .A1(n9398), .A2(n8646), .ZN(n8513) );
  AND2_X1 U5009 ( .A1(n5598), .A2(n5601), .ZN(n5599) );
  AND2_X1 U5010 ( .A1(n8507), .A2(n8641), .ZN(n8677) );
  OR2_X1 U5011 ( .A1(n9431), .A2(n9186), .ZN(n8624) );
  NOR2_X1 U5012 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  AND2_X1 U5013 ( .A1(n4864), .A2(n5207), .ZN(n4983) );
  INV_X1 U5014 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U5015 ( .A1(n9896), .A2(n9772), .ZN(n5244) );
  OR2_X1 U5016 ( .A1(n9901), .A2(n9783), .ZN(n6644) );
  NAND2_X1 U5017 ( .A1(n9901), .A2(n9783), .ZN(n8721) );
  NAND2_X1 U5018 ( .A1(n9737), .A2(n9715), .ZN(n9729) );
  NAND2_X1 U5019 ( .A1(n5994), .A2(n5993), .ZN(n6068) );
  NAND2_X1 U5020 ( .A1(n5797), .A2(n5796), .ZN(n5818) );
  OAI21_X1 U5021 ( .B1(n5756), .B2(n5104), .A(n5101), .ZN(n5797) );
  AOI21_X1 U5022 ( .B1(n5103), .B2(n5102), .A(n5793), .ZN(n5101) );
  OR2_X1 U5023 ( .A1(n5553), .A2(n5552), .ZN(n5555) );
  INV_X1 U5024 ( .A(n5256), .ZN(n5246) );
  NAND2_X1 U5025 ( .A1(n5252), .A2(n5256), .ZN(n5247) );
  AOI21_X1 U5026 ( .B1(n5251), .B2(n5252), .A(n5250), .ZN(n5249) );
  NAND2_X1 U5027 ( .A1(n8398), .A2(n4870), .ZN(n8845) );
  NAND2_X1 U5028 ( .A1(n6751), .A2(n6780), .ZN(n5520) );
  NAND2_X2 U5029 ( .A1(n8749), .A2(n6053), .ZN(n6751) );
  INV_X1 U5030 ( .A(n9885), .ZN(n9715) );
  NAND2_X1 U5031 ( .A1(n6549), .A2(n9718), .ZN(n8737) );
  INV_X1 U5032 ( .A(n9155), .ZN(n4963) );
  AND2_X1 U5033 ( .A1(n9333), .A2(n9339), .ZN(n8478) );
  OR2_X1 U5034 ( .A1(n9911), .A2(n9819), .ZN(n8733) );
  AND2_X1 U5035 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  OR2_X1 U5036 ( .A1(n5833), .A2(n5832), .ZN(n5835) );
  AND2_X1 U5037 ( .A1(n5182), .A2(n5628), .ZN(n5181) );
  INV_X1 U5038 ( .A(n8145), .ZN(n5182) );
  AND2_X1 U5039 ( .A1(n9422), .A2(n9187), .ZN(n8649) );
  NAND2_X1 U5040 ( .A1(n5956), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5999) );
  OR2_X1 U5041 ( .A1(n9416), .A2(n9069), .ZN(n8633) );
  INV_X1 U5042 ( .A(n9181), .ZN(n9185) );
  NAND2_X1 U5043 ( .A1(n4957), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5912) );
  OR2_X1 U5044 ( .A1(n9437), .A2(n8483), .ZN(n8619) );
  OR2_X1 U5045 ( .A1(n9447), .A2(n9043), .ZN(n8610) );
  AND2_X1 U5046 ( .A1(n8593), .A2(n9336), .ZN(n8476) );
  OR2_X1 U5047 ( .A1(n5565), .A2(n7902), .ZN(n5586) );
  NAND2_X1 U5048 ( .A1(n10481), .A2(n9103), .ZN(n8653) );
  AND2_X1 U5049 ( .A1(n7897), .A2(n8680), .ZN(n8686) );
  NOR2_X1 U5050 ( .A1(n5051), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5048) );
  AND2_X1 U5051 ( .A1(n5356), .A2(n5355), .ZN(n5206) );
  INV_X1 U5052 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5378) );
  INV_X1 U5053 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4949) );
  INV_X1 U5054 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4950) );
  AND2_X1 U5055 ( .A1(n7021), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7022) );
  OR2_X1 U5056 ( .A1(n9922), .A2(n9608), .ZN(n6551) );
  OR2_X1 U5057 ( .A1(n9942), .A2(n8784), .ZN(n8448) );
  OR2_X1 U5058 ( .A1(n9952), .A2(n9569), .ZN(n6623) );
  NAND2_X1 U5059 ( .A1(n9958), .A2(n8765), .ZN(n6621) );
  NAND2_X1 U5060 ( .A1(n7161), .A2(n7072), .ZN(n6676) );
  NAND2_X1 U5061 ( .A1(n6387), .A2(n6386), .ZN(n6674) );
  OR2_X1 U5062 ( .A1(n5818), .A2(n5817), .ZN(n5847) );
  NAND2_X1 U5063 ( .A1(n5730), .A2(n5729), .ZN(n5733) );
  INV_X1 U5064 ( .A(n5728), .ZN(n5729) );
  NAND2_X1 U5065 ( .A1(n5635), .A2(n5634), .ZN(n5656) );
  AND2_X1 U5066 ( .A1(n5603), .A2(n5560), .ZN(n5598) );
  INV_X1 U5067 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U5068 ( .A1(n5554), .A2(n5537), .ZN(n5552) );
  INV_X1 U5069 ( .A(n9055), .ZN(n5192) );
  NAND2_X1 U5070 ( .A1(n5642), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5668) );
  INV_X1 U5071 ( .A(n5643), .ZN(n5642) );
  INV_X1 U5072 ( .A(n5436), .ZN(n5826) );
  INV_X1 U5073 ( .A(n8683), .ZN(n5020) );
  XNOR2_X1 U5074 ( .A(n8685), .B(n8684), .ZN(n4945) );
  INV_X1 U5075 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5331) );
  INV_X1 U5076 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U5077 ( .A1(n8493), .A2(n8492), .ZN(n9405) );
  NOR2_X1 U5078 ( .A1(n8880), .A2(n9405), .ZN(n8883) );
  NAND2_X1 U5079 ( .A1(n9223), .A2(n4919), .ZN(n9198) );
  INV_X1 U5080 ( .A(n9207), .ZN(n8856) );
  OR2_X1 U5081 ( .A1(n9459), .A2(n9058), .ZN(n9272) );
  NAND2_X1 U5082 ( .A1(n5666), .A2(n5665), .ZN(n8396) );
  INV_X1 U5083 ( .A(n5263), .ZN(n5262) );
  OAI21_X1 U5084 ( .B1(n5265), .B2(n5264), .A(n8665), .ZN(n5263) );
  INV_X1 U5085 ( .A(n8114), .ZN(n5264) );
  OR2_X1 U5086 ( .A1(n10527), .A2(n8128), .ZN(n8555) );
  NAND2_X1 U5087 ( .A1(n5996), .A2(n5995), .ZN(n9410) );
  NAND2_X1 U5088 ( .A1(n8419), .A2(n5561), .ZN(n5996) );
  XNOR2_X1 U5089 ( .A(n5346), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5347) );
  AND2_X1 U5090 ( .A1(n5341), .A2(n5269), .ZN(n5268) );
  NOR2_X1 U5091 ( .A1(n5270), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U5092 ( .A1(n6494), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6509) );
  INV_X1 U5093 ( .A(n6507), .ZN(n6494) );
  AND2_X1 U5094 ( .A1(n6652), .A2(n6708), .ZN(n9720) );
  INV_X1 U5095 ( .A(n5233), .ZN(n8738) );
  INV_X1 U5096 ( .A(n5236), .ZN(n5234) );
  NAND2_X1 U5097 ( .A1(n5137), .A2(n4878), .ZN(n9719) );
  OR2_X1 U5098 ( .A1(n8956), .A2(n6535), .ZN(n6528) );
  NAND2_X1 U5099 ( .A1(n8722), .A2(n8721), .ZN(n9758) );
  OR2_X1 U5100 ( .A1(n9901), .A2(n9759), .ZN(n5245) );
  AND2_X1 U5101 ( .A1(n6579), .A2(n8723), .ZN(n9757) );
  NAND2_X1 U5102 ( .A1(n9952), .A2(n9569), .ZN(n8358) );
  INV_X1 U5103 ( .A(n6532), .ZN(n6436) );
  AND2_X1 U5104 ( .A1(n7140), .A2(n4847), .ZN(n9866) );
  AND2_X1 U5105 ( .A1(n7140), .A2(n10402), .ZN(n9864) );
  AND2_X1 U5106 ( .A1(n9729), .A2(n8742), .ZN(n9886) );
  NAND2_X1 U5107 ( .A1(n5890), .A2(n5889), .ZN(n5908) );
  NAND2_X1 U5108 ( .A1(n9758), .A2(n9757), .ZN(n8724) );
  INV_X1 U5109 ( .A(n6405), .ZN(n10265) );
  INV_X1 U5110 ( .A(n9756), .ZN(n9896) );
  OR2_X1 U5111 ( .A1(n8550), .A2(n8551), .ZN(n4979) );
  NAND2_X1 U5112 ( .A1(n4900), .A2(n4977), .ZN(n4976) );
  NAND2_X1 U5113 ( .A1(n8544), .A2(n4978), .ZN(n4977) );
  INV_X1 U5114 ( .A(n8547), .ZN(n4978) );
  NAND2_X1 U5115 ( .A1(n8563), .A2(n8555), .ZN(n4937) );
  AOI21_X1 U5116 ( .B1(n8566), .B2(n8565), .A(n8564), .ZN(n8567) );
  OR3_X1 U5117 ( .A1(n6613), .A2(n6612), .A3(n8259), .ZN(n6615) );
  NAND2_X1 U5118 ( .A1(n6615), .A2(n6614), .ZN(n5009) );
  NOR2_X1 U5119 ( .A1(n8251), .A2(n6659), .ZN(n5008) );
  NAND2_X1 U5120 ( .A1(n6615), .A2(n8249), .ZN(n5012) );
  OAI21_X1 U5121 ( .B1(n5004), .B2(n5002), .A(n5001), .ZN(n5000) );
  AND2_X1 U5122 ( .A1(n6625), .A2(n6624), .ZN(n5001) );
  OAI21_X1 U5123 ( .B1(n6617), .B2(n6659), .A(n5003), .ZN(n5002) );
  NOR2_X1 U5124 ( .A1(n6618), .A2(n6642), .ZN(n5004) );
  NOR2_X1 U5125 ( .A1(n4851), .A2(n4886), .ZN(n4990) );
  INV_X1 U5126 ( .A(n6639), .ZN(n4993) );
  NOR2_X1 U5127 ( .A1(n4851), .A2(n4884), .ZN(n4989) );
  INV_X1 U5128 ( .A(n6643), .ZN(n4988) );
  INV_X1 U5129 ( .A(n8719), .ZN(n4991) );
  OAI21_X1 U5130 ( .B1(n4939), .B2(n4938), .A(n8622), .ZN(n8625) );
  OR2_X1 U5131 ( .A1(n8621), .A2(n8620), .ZN(n4938) );
  AOI21_X1 U5132 ( .B1(n8617), .B2(n8616), .A(n8615), .ZN(n4939) );
  AND2_X1 U5133 ( .A1(n5047), .A2(n4964), .ZN(n5046) );
  NAND2_X1 U5134 ( .A1(n5149), .A2(n9154), .ZN(n5047) );
  AOI21_X1 U5135 ( .B1(n5149), .B2(n5152), .A(n5148), .ZN(n4964) );
  INV_X1 U5136 ( .A(n8639), .ZN(n5148) );
  INV_X1 U5137 ( .A(n5149), .ZN(n5045) );
  AOI21_X1 U5138 ( .B1(n8625), .B2(n9204), .A(n9181), .ZN(n8628) );
  NOR2_X1 U5139 ( .A1(n9422), .A2(n9187), .ZN(n8650) );
  INV_X1 U5140 ( .A(n8065), .ZN(n5287) );
  NOR2_X1 U5141 ( .A1(n5928), .A2(n5113), .ZN(n5112) );
  INV_X1 U5142 ( .A(n5907), .ZN(n5113) );
  OAI21_X1 U5143 ( .B1(n4947), .B2(n4972), .A(n4970), .ZN(n4946) );
  NAND2_X1 U5144 ( .A1(n8634), .A2(n8876), .ZN(n4972) );
  NOR2_X1 U5145 ( .A1(n4872), .A2(n4971), .ZN(n4970) );
  NOR2_X1 U5146 ( .A1(n9154), .A2(n4948), .ZN(n4947) );
  NOR2_X1 U5147 ( .A1(n4969), .A2(n4968), .ZN(n4967) );
  INV_X1 U5148 ( .A(n8640), .ZN(n4969) );
  NAND2_X1 U5149 ( .A1(n8642), .A2(n8641), .ZN(n4968) );
  OR3_X1 U5150 ( .A1(n9143), .A2(n8691), .A3(n8680), .ZN(n8643) );
  NAND2_X1 U5151 ( .A1(n9153), .A2(n9069), .ZN(n5256) );
  OR2_X1 U5152 ( .A1(n9416), .A2(n9422), .ZN(n5177) );
  NOR2_X1 U5153 ( .A1(n8650), .A2(n8649), .ZN(n8859) );
  NOR2_X1 U5154 ( .A1(n9447), .A2(n9452), .ZN(n5173) );
  NAND2_X1 U5155 ( .A1(n8369), .A2(n8575), .ZN(n5026) );
  INV_X1 U5156 ( .A(n8581), .ZN(n5022) );
  INV_X1 U5157 ( .A(n8575), .ZN(n5023) );
  NAND2_X1 U5158 ( .A1(n4896), .A2(n8542), .ZN(n5035) );
  INV_X1 U5159 ( .A(n5035), .ZN(n5028) );
  NAND2_X1 U5160 ( .A1(n5032), .A2(n8543), .ZN(n5030) );
  NOR2_X1 U5161 ( .A1(n5037), .A2(n5033), .ZN(n5032) );
  INV_X1 U5162 ( .A(n7926), .ZN(n5033) );
  NAND2_X1 U5163 ( .A1(n8537), .A2(n8538), .ZN(n8656) );
  OAI21_X1 U5164 ( .B1(n10474), .B2(n7394), .A(n7393), .ZN(n7397) );
  NOR2_X1 U5165 ( .A1(n9103), .A2(n7392), .ZN(n7394) );
  AND2_X1 U5166 ( .A1(n9105), .A2(n7745), .ZN(n7391) );
  OR2_X1 U5167 ( .A1(n8503), .A2(n6785), .ZN(n5442) );
  INV_X1 U5168 ( .A(n10520), .ZN(n8825) );
  NAND2_X1 U5169 ( .A1(n7706), .A2(n8537), .ZN(n7708) );
  NAND2_X1 U5170 ( .A1(n5342), .A2(n5271), .ZN(n5270) );
  INV_X1 U5171 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5271) );
  INV_X1 U5172 ( .A(n9640), .ZN(n5278) );
  NAND2_X1 U5173 ( .A1(n4915), .A2(n9640), .ZN(n5276) );
  AND2_X1 U5174 ( .A1(n5277), .A2(n9522), .ZN(n5275) );
  INV_X1 U5175 ( .A(n9534), .ZN(n5303) );
  NAND2_X1 U5176 ( .A1(n9520), .A2(n9522), .ZN(n5282) );
  OAI211_X1 U5177 ( .C1(n6660), .C2(n6659), .A(n4892), .B(n5076), .ZN(n6665)
         );
  OAI21_X1 U5178 ( .B1(n5017), .B2(n5016), .A(n5013), .ZN(n5076) );
  OR2_X1 U5179 ( .A1(n6658), .A2(n6657), .ZN(n5077) );
  OR2_X1 U5180 ( .A1(n9878), .A2(n9723), .ZN(n6711) );
  NAND2_X1 U5181 ( .A1(n4921), .A2(n8703), .ZN(n5062) );
  OR2_X1 U5182 ( .A1(n9896), .A2(n9744), .ZN(n6579) );
  INV_X1 U5183 ( .A(n9908), .ZN(n8917) );
  INV_X1 U5184 ( .A(n8716), .ZN(n5133) );
  INV_X1 U5185 ( .A(n5132), .ZN(n5131) );
  OAI21_X1 U5186 ( .B1(n9830), .B2(n5133), .A(n9817), .ZN(n5132) );
  AND2_X1 U5187 ( .A1(n9627), .A2(n9865), .ZN(n5224) );
  INV_X1 U5188 ( .A(n6228), .ZN(n6146) );
  AND2_X1 U5189 ( .A1(n5212), .A2(n8279), .ZN(n8276) );
  INV_X1 U5190 ( .A(n8270), .ZN(n5212) );
  NOR2_X1 U5191 ( .A1(n9963), .A2(n8258), .ZN(n5065) );
  AND2_X1 U5192 ( .A1(n7814), .A2(n7812), .ZN(n4951) );
  AND2_X1 U5193 ( .A1(n4913), .A2(n5227), .ZN(n5226) );
  OAI21_X1 U5194 ( .B1(n7131), .B2(n7340), .A(n7130), .ZN(n7132) );
  NAND2_X1 U5195 ( .A1(n6078), .A2(n6077), .ZN(n6125) );
  AND2_X1 U5196 ( .A1(n6100), .A2(n5313), .ZN(n5312) );
  INV_X1 U5197 ( .A(n5096), .ZN(n5095) );
  OAI21_X1 U5198 ( .B1(n5865), .B2(n5848), .A(n5864), .ZN(n5096) );
  NOR2_X1 U5199 ( .A1(n5098), .A2(n5865), .ZN(n5097) );
  INV_X1 U5200 ( .A(n5846), .ZN(n5098) );
  AOI21_X1 U5201 ( .B1(n5082), .B2(n5084), .A(n4887), .ZN(n5079) );
  AND2_X1 U5202 ( .A1(n5326), .A2(n5087), .ZN(n5086) );
  NAND2_X1 U5203 ( .A1(n5657), .A2(n5656), .ZN(n5087) );
  AND2_X1 U5204 ( .A1(n5217), .A2(n5606), .ZN(n5216) );
  NAND2_X1 U5205 ( .A1(n5599), .A2(n5218), .ZN(n5217) );
  INV_X1 U5206 ( .A(n5599), .ZN(n5219) );
  NAND2_X1 U5207 ( .A1(n6370), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4940) );
  INV_X1 U5208 ( .A(n6743), .ZN(n5202) );
  NAND2_X1 U5209 ( .A1(n5187), .A2(n9017), .ZN(n5186) );
  OR2_X1 U5210 ( .A1(n5826), .A2(n6945), .ZN(n5351) );
  NAND2_X1 U5211 ( .A1(n9007), .A2(n9008), .ZN(n9006) );
  INV_X1 U5212 ( .A(n5179), .ZN(n5178) );
  OAI21_X1 U5213 ( .B1(n5181), .B2(n5180), .A(n8219), .ZN(n5179) );
  INV_X1 U5214 ( .A(n5655), .ZN(n5180) );
  NAND2_X1 U5215 ( .A1(n5629), .A2(n5181), .ZN(n8143) );
  NAND2_X1 U5216 ( .A1(n5611), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5643) );
  XNOR2_X1 U5217 ( .A(n5470), .B(n5472), .ZN(n7167) );
  AND4_X1 U5218 ( .A1(n5830), .A2(n5829), .A3(n5828), .A4(n5827), .ZN(n9058)
         );
  OR2_X1 U5219 ( .A1(n5826), .A2(n6977), .ZN(n5547) );
  NOR2_X1 U5220 ( .A1(n5454), .A2(n5435), .ZN(n5267) );
  NAND2_X1 U5221 ( .A1(n8755), .A2(n8883), .ZN(n8836) );
  AND2_X1 U5222 ( .A1(n6046), .A2(n6000), .ZN(n8861) );
  AOI21_X1 U5223 ( .B1(n9167), .B2(n8488), .A(n4889), .ZN(n9155) );
  NOR2_X1 U5224 ( .A1(n8859), .A2(n5254), .ZN(n5253) );
  NOR2_X1 U5225 ( .A1(n8858), .A2(n9181), .ZN(n5254) );
  NAND2_X1 U5226 ( .A1(n8633), .A2(n8632), .ZN(n9154) );
  OR2_X1 U5227 ( .A1(n9195), .A2(n9087), .ZN(n9168) );
  NAND2_X1 U5228 ( .A1(n9168), .A2(n8623), .ZN(n9181) );
  NOR2_X1 U5229 ( .A1(n9195), .A2(n9210), .ZN(n8858) );
  NOR2_X1 U5230 ( .A1(n9431), .A2(n9201), .ZN(n9176) );
  INV_X1 U5231 ( .A(n5912), .ZN(n5911) );
  OR2_X1 U5232 ( .A1(n5936), .A2(n10198), .ZN(n5958) );
  AND2_X1 U5233 ( .A1(n8624), .A2(n8517), .ZN(n9207) );
  NAND2_X1 U5234 ( .A1(n8619), .A2(n9206), .ZN(n9221) );
  AOI21_X1 U5235 ( .B1(n5165), .B2(n5040), .A(n5039), .ZN(n5038) );
  INV_X1 U5236 ( .A(n5165), .ZN(n5041) );
  INV_X1 U5237 ( .A(n8610), .ZN(n5039) );
  NAND2_X1 U5238 ( .A1(n9238), .A2(n9237), .ZN(n9236) );
  INV_X1 U5239 ( .A(n8854), .ZN(n9237) );
  AND2_X1 U5240 ( .A1(n9249), .A2(n8651), .ZN(n5165) );
  NAND2_X1 U5241 ( .A1(n9294), .A2(n8596), .ZN(n8482) );
  AND4_X1 U5242 ( .A1(n5813), .A2(n5812), .A3(n5811), .A4(n5810), .ZN(n9256)
         );
  AND2_X1 U5243 ( .A1(n8610), .A2(n8613), .ZN(n9249) );
  NOR2_X1 U5244 ( .A1(n8847), .A2(n5260), .ZN(n5259) );
  INV_X1 U5245 ( .A(n8846), .ZN(n5260) );
  AND2_X1 U5246 ( .A1(n9378), .A2(n5156), .ZN(n9305) );
  NOR2_X1 U5247 ( .A1(n5157), .A2(n9462), .ZN(n5156) );
  INV_X1 U5248 ( .A(n5158), .ZN(n5157) );
  NAND2_X1 U5249 ( .A1(n5741), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5764) );
  INV_X1 U5250 ( .A(n5742), .ZN(n5741) );
  AND4_X1 U5251 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), .ZN(n8471)
         );
  NOR2_X1 U5252 ( .A1(n8131), .A2(n8136), .ZN(n8132) );
  AND2_X1 U5253 ( .A1(n8663), .A2(n8112), .ZN(n5265) );
  NOR2_X1 U5254 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  AOI21_X1 U5255 ( .B1(n8819), .B2(n8832), .A(n7957), .ZN(n7959) );
  XNOR2_X1 U5256 ( .A(n9096), .B(n10520), .ZN(n8832) );
  NAND2_X1 U5257 ( .A1(n7930), .A2(n8658), .ZN(n5258) );
  NOR2_X1 U5258 ( .A1(n5037), .A2(n5147), .ZN(n5036) );
  OR2_X1 U5259 ( .A1(n7773), .A2(n7718), .ZN(n7977) );
  AND2_X1 U5260 ( .A1(n7388), .A2(n8653), .ZN(n7389) );
  OR2_X1 U5261 ( .A1(n6749), .A2(n6036), .ZN(n8689) );
  AND2_X1 U5262 ( .A1(n6053), .A2(n7398), .ZN(n9390) );
  OR2_X1 U5263 ( .A1(n10568), .A2(n9143), .ZN(n7385) );
  NAND2_X1 U5264 ( .A1(n9405), .A2(n10575), .ZN(n5143) );
  NAND2_X1 U5265 ( .A1(n5740), .A2(n5739), .ZN(n9474) );
  NAND2_X1 U5266 ( .A1(n5688), .A2(n5687), .ZN(n10574) );
  AND2_X1 U5267 ( .A1(n8389), .A2(n8380), .ZN(n5272) );
  AND2_X1 U5268 ( .A1(n8690), .A2(n8686), .ZN(n10575) );
  NAND2_X1 U5269 ( .A1(n7400), .A2(n7399), .ZN(n10564) );
  INV_X1 U5270 ( .A(n5196), .ZN(n5195) );
  OAI21_X1 U5271 ( .B1(n5357), .B2(n5343), .A(n5363), .ZN(n5196) );
  AND2_X1 U5272 ( .A1(n5206), .A2(n5205), .ZN(n5204) );
  INV_X1 U5273 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5205) );
  INV_X1 U5274 ( .A(n9661), .ZN(n7647) );
  XNOR2_X1 U5275 ( .A(n7095), .B(n8947), .ZN(n7247) );
  AND2_X1 U5276 ( .A1(n5301), .A2(n5300), .ZN(n5299) );
  INV_X1 U5277 ( .A(n9590), .ZN(n5300) );
  OR2_X1 U5278 ( .A1(n8914), .A2(n5303), .ZN(n5301) );
  AND2_X1 U5279 ( .A1(n8914), .A2(n5303), .ZN(n5302) );
  OAI21_X1 U5280 ( .B1(n7343), .B2(n7039), .A(n7020), .ZN(n8697) );
  NAND2_X1 U5281 ( .A1(n7026), .A2(n7096), .ZN(n7027) );
  NAND2_X1 U5282 ( .A1(n5294), .A2(n9617), .ZN(n5293) );
  INV_X1 U5283 ( .A(n8811), .ZN(n5292) );
  AND2_X1 U5284 ( .A1(n8796), .A2(n5296), .ZN(n5295) );
  OR2_X1 U5285 ( .A1(n6320), .A2(n6319), .ZN(n6322) );
  AND2_X1 U5286 ( .A1(n9603), .A2(n9599), .ZN(n8907) );
  XNOR2_X1 U5287 ( .A(n7099), .B(n4841), .ZN(n7102) );
  NAND2_X1 U5288 ( .A1(n6140), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U5289 ( .A1(n6482), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U5290 ( .A1(n5280), .A2(n5279), .ZN(n9638) );
  INV_X1 U5291 ( .A(n5281), .ZN(n5280) );
  NAND2_X1 U5292 ( .A1(n5281), .A2(n4915), .ZN(n9637) );
  OAI21_X1 U5293 ( .B1(n6665), .B2(n7110), .A(n6661), .ZN(n5075) );
  AND2_X1 U5294 ( .A1(n6168), .A2(n6167), .ZN(n8813) );
  AND4_X1 U5295 ( .A1(n6262), .A2(n6261), .A3(n6260), .A4(n6259), .ZN(n8765)
         );
  NAND2_X1 U5296 ( .A1(n4904), .A2(n5244), .ZN(n5238) );
  INV_X1 U5297 ( .A(n5245), .ZN(n5239) );
  INV_X1 U5298 ( .A(n9770), .ZN(n5241) );
  AND2_X1 U5299 ( .A1(n6644), .A2(n8721), .ZN(n9770) );
  AOI21_X1 U5300 ( .B1(n8917), .B2(n8916), .A(n8736), .ZN(n9764) );
  NOR2_X1 U5301 ( .A1(n9789), .A2(n8735), .ZN(n8736) );
  AND2_X1 U5302 ( .A1(n9908), .A2(n9806), .ZN(n8735) );
  AND2_X1 U5303 ( .A1(n6550), .A2(n8718), .ZN(n9805) );
  NAND2_X1 U5304 ( .A1(n5228), .A2(n6563), .ZN(n5230) );
  AND2_X1 U5305 ( .A1(n9922), .A2(n9850), .ZN(n5232) );
  NAND2_X1 U5306 ( .A1(n4955), .A2(n8715), .ZN(n9829) );
  OAI21_X1 U5307 ( .B1(n8713), .B2(n5120), .A(n5118), .ZN(n4955) );
  INV_X1 U5308 ( .A(n5121), .ZN(n5120) );
  AOI21_X1 U5309 ( .B1(n5121), .B2(n5125), .A(n5119), .ZN(n5118) );
  NAND2_X1 U5310 ( .A1(n9829), .A2(n9830), .ZN(n9828) );
  INV_X1 U5311 ( .A(n5230), .ZN(n9824) );
  AOI21_X1 U5312 ( .B1(n5124), .B2(n5123), .A(n5122), .ZN(n5121) );
  INV_X1 U5313 ( .A(n8711), .ZN(n5123) );
  OR2_X1 U5314 ( .A1(n9627), .A2(n8794), .ZN(n8712) );
  NAND2_X1 U5315 ( .A1(n5127), .A2(n8711), .ZN(n5126) );
  INV_X1 U5316 ( .A(n8713), .ZN(n5127) );
  NOR2_X1 U5317 ( .A1(n8454), .A2(n5223), .ZN(n5222) );
  INV_X1 U5318 ( .A(n8452), .ZN(n5223) );
  AND2_X1 U5319 ( .A1(n8712), .A2(n8711), .ZN(n8454) );
  OAI21_X1 U5320 ( .B1(n8311), .B2(n4866), .A(n5134), .ZN(n8451) );
  INV_X1 U5321 ( .A(n5135), .ZN(n5134) );
  OAI21_X1 U5322 ( .B1(n4852), .B2(n4866), .A(n8426), .ZN(n5135) );
  NAND2_X1 U5323 ( .A1(n8358), .A2(n6623), .ZN(n8279) );
  INV_X1 U5324 ( .A(n8279), .ZN(n8254) );
  OR2_X1 U5325 ( .A1(n9958), .A2(n8765), .ZN(n8253) );
  NAND2_X1 U5326 ( .A1(n8311), .A2(n4852), .ZN(n8359) );
  NAND2_X1 U5327 ( .A1(n7811), .A2(n7810), .ZN(n7813) );
  NAND2_X1 U5328 ( .A1(n7592), .A2(n7591), .ZN(n7811) );
  AND2_X1 U5329 ( .A1(n6438), .A2(n6437), .ZN(n7665) );
  NAND2_X1 U5330 ( .A1(n7298), .A2(n7297), .ZN(n7315) );
  XNOR2_X1 U5331 ( .A(n7129), .B(n7354), .ZN(n6553) );
  OR3_X1 U5332 ( .A1(n7293), .A2(n9990), .A3(n7292), .ZN(n7542) );
  XNOR2_X1 U5333 ( .A(n9729), .B(n9730), .ZN(n9882) );
  NAND2_X1 U5334 ( .A1(n6173), .A2(n6172), .ZN(n9916) );
  NAND2_X1 U5335 ( .A1(n6215), .A2(n6214), .ZN(n9942) );
  NAND2_X1 U5336 ( .A1(n6266), .A2(n6265), .ZN(n8179) );
  AND2_X1 U5337 ( .A1(n7661), .A2(n8182), .ZN(n10494) );
  INV_X1 U5338 ( .A(n10537), .ZN(n9964) );
  XNOR2_X1 U5339 ( .A(n6125), .B(n6124), .ZN(n8495) );
  XNOR2_X1 U5340 ( .A(n5953), .B(n5952), .ZN(n8351) );
  OAI21_X1 U5341 ( .B1(n5908), .B2(n5111), .A(n5108), .ZN(n5953) );
  INV_X1 U5342 ( .A(n5114), .ZN(n5111) );
  NAND2_X1 U5343 ( .A1(n5908), .A2(n5907), .ZN(n5929) );
  AOI21_X1 U5344 ( .B1(n5847), .B2(n5846), .A(n5099), .ZN(n5866) );
  XNOR2_X1 U5345 ( .A(n5805), .B(n5804), .ZN(n7610) );
  NAND2_X1 U5346 ( .A1(n5100), .A2(n5103), .ZN(n5794) );
  NAND2_X1 U5347 ( .A1(n5756), .A2(n5106), .ZN(n5100) );
  XNOR2_X1 U5348 ( .A(n5730), .B(n5728), .ZN(n6237) );
  NAND2_X1 U5349 ( .A1(n5085), .A2(n5656), .ZN(n5681) );
  OR2_X1 U5350 ( .A1(n5658), .A2(n5657), .ZN(n5085) );
  OR2_X1 U5351 ( .A1(n6198), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U5352 ( .A1(n5574), .A2(n5603), .ZN(n4942) );
  NAND2_X1 U5353 ( .A1(n5893), .A2(n5892), .ZN(n9437) );
  AND4_X1 U5354 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n9063)
         );
  AND4_X1 U5355 ( .A1(n5514), .A2(n5513), .A3(n5512), .A4(n5511), .ZN(n7973)
         );
  OR2_X1 U5356 ( .A1(n4945), .A2(n4927), .ZN(n4944) );
  NAND2_X1 U5357 ( .A1(n5154), .A2(n4864), .ZN(n5538) );
  NAND2_X1 U5358 ( .A1(n8505), .A2(n8504), .ZN(n9398) );
  OAI21_X1 U5359 ( .B1(n8877), .B2(n8876), .A(n5255), .ZN(n8879) );
  INV_X1 U5360 ( .A(n5145), .ZN(n5144) );
  NAND2_X1 U5361 ( .A1(n8888), .A2(n10467), .ZN(n5146) );
  OAI22_X1 U5362 ( .A1(n9156), .A2(n9343), .B1(n8506), .B2(n8890), .ZN(n5145)
         );
  NOR2_X1 U5363 ( .A1(n8883), .A2(n8882), .ZN(n9406) );
  NAND2_X1 U5364 ( .A1(n8864), .A2(n8876), .ZN(n8868) );
  NAND2_X1 U5365 ( .A1(n5372), .A2(n5371), .ZN(n8749) );
  INV_X1 U5366 ( .A(n5367), .ZN(n5371) );
  NAND2_X1 U5367 ( .A1(n6331), .A2(n6330), .ZN(n7854) );
  NAND2_X1 U5368 ( .A1(n8226), .A2(n6340), .ZN(n6481) );
  AND4_X1 U5369 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(n9569)
         );
  AND4_X1 U5370 ( .A1(n6235), .A2(n6234), .A3(n6233), .A4(n6232), .ZN(n9582)
         );
  AND2_X1 U5371 ( .A1(n6157), .A2(n6156), .ZN(n9608) );
  INV_X1 U5372 ( .A(n7125), .ZN(n7030) );
  INV_X1 U5373 ( .A(n9783), .ZN(n9759) );
  AND4_X1 U5374 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n7835)
         );
  AND4_X1 U5375 ( .A1(n6339), .A2(n6338), .A3(n6337), .A4(n6336), .ZN(n7826)
         );
  NAND2_X1 U5376 ( .A1(n6133), .A2(n6132), .ZN(n9874) );
  AOI21_X1 U5377 ( .B1(n9725), .B2(n9869), .A(n9724), .ZN(n9883) );
  AND2_X1 U5378 ( .A1(n8730), .A2(n8729), .ZN(n9888) );
  AOI22_X1 U5379 ( .A1(n9651), .A2(n9866), .B1(n9864), .B2(n5243), .ZN(n8729)
         );
  NAND2_X1 U5380 ( .A1(n6519), .A2(n6518), .ZN(n9885) );
  NAND2_X1 U5381 ( .A1(n8724), .A2(n8723), .ZN(n9743) );
  NAND2_X1 U5382 ( .A1(n4996), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4995) );
  INV_X1 U5383 ( .A(n6532), .ZN(n4996) );
  INV_X1 U5384 ( .A(n7389), .ZN(n8524) );
  NAND2_X1 U5385 ( .A1(n4994), .A2(n6684), .ZN(n6590) );
  NAND2_X1 U5386 ( .A1(n7525), .A2(n7653), .ZN(n4994) );
  INV_X1 U5387 ( .A(n8544), .ZN(n4980) );
  NAND2_X1 U5388 ( .A1(n4974), .A2(n4981), .ZN(n4973) );
  NAND2_X1 U5389 ( .A1(n8545), .A2(n4976), .ZN(n4975) );
  NAND2_X1 U5390 ( .A1(n4979), .A2(n8661), .ZN(n4974) );
  AND3_X1 U5391 ( .A1(n8560), .A2(n4936), .A3(n4935), .ZN(n8566) );
  NAND2_X1 U5392 ( .A1(n8556), .A2(n8643), .ZN(n4935) );
  NAND2_X1 U5393 ( .A1(n4937), .A2(n8637), .ZN(n4936) );
  AND2_X1 U5394 ( .A1(n9368), .A2(n8588), .ZN(n4965) );
  NAND2_X1 U5395 ( .A1(n5012), .A2(n5011), .ZN(n5010) );
  NAND2_X1 U5396 ( .A1(n5009), .A2(n5008), .ZN(n5007) );
  AND2_X1 U5397 ( .A1(n6619), .A2(n6659), .ZN(n5011) );
  AND2_X1 U5398 ( .A1(n6622), .A2(n8254), .ZN(n5003) );
  NOR2_X1 U5399 ( .A1(n4931), .A2(n9342), .ZN(n4930) );
  NAND2_X1 U5400 ( .A1(n5000), .A2(n6626), .ZN(n6627) );
  OAI21_X1 U5401 ( .B1(n4989), .B2(n4991), .A(n4988), .ZN(n4986) );
  NAND2_X1 U5402 ( .A1(n4990), .A2(n4988), .ZN(n4987) );
  AOI21_X1 U5403 ( .B1(n5046), .B2(n5045), .A(n5044), .ZN(n5043) );
  NAND2_X1 U5404 ( .A1(n5046), .A2(n4963), .ZN(n5042) );
  INV_X1 U5405 ( .A(n8638), .ZN(n5044) );
  AOI21_X1 U5406 ( .B1(n8630), .B2(n8631), .A(n8629), .ZN(n4948) );
  NAND2_X1 U5407 ( .A1(n8635), .A2(n8878), .ZN(n4971) );
  OR2_X1 U5408 ( .A1(n9405), .A2(n8866), .ZN(n8638) );
  NOR2_X1 U5409 ( .A1(n5872), .A2(n10212), .ZN(n4957) );
  OR2_X1 U5410 ( .A1(n9467), .A2(n9063), .ZN(n8593) );
  OR2_X1 U5411 ( .A1(n10488), .A2(n7578), .ZN(n8533) );
  NOR2_X1 U5412 ( .A1(n6654), .A2(n6655), .ZN(n5017) );
  AND3_X1 U5413 ( .A1(n8727), .A2(n6651), .A3(n6650), .ZN(n6654) );
  INV_X1 U5414 ( .A(n6653), .ZN(n5016) );
  NOR2_X1 U5415 ( .A1(n5015), .A2(n5014), .ZN(n5013) );
  NOR2_X1 U5416 ( .A1(n6656), .A2(n6711), .ZN(n5015) );
  NAND2_X1 U5417 ( .A1(n6716), .A2(n6657), .ZN(n5014) );
  NAND2_X1 U5418 ( .A1(n9830), .A2(n5231), .ZN(n5227) );
  INV_X1 U5419 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6086) );
  INV_X1 U5420 ( .A(n5106), .ZN(n5102) );
  NAND2_X1 U5421 ( .A1(n5755), .A2(n5757), .ZN(n5105) );
  AOI21_X1 U5422 ( .B1(n5086), .B2(n5083), .A(n4901), .ZN(n5082) );
  INV_X1 U5423 ( .A(n5656), .ZN(n5083) );
  INV_X1 U5424 ( .A(n5682), .ZN(n5209) );
  INV_X1 U5425 ( .A(n5086), .ZN(n5084) );
  INV_X1 U5426 ( .A(n5554), .ZN(n5218) );
  NAND2_X1 U5427 ( .A1(n5535), .A2(n10057), .ZN(n5554) );
  INV_X1 U5428 ( .A(n5496), .ZN(n5072) );
  INV_X1 U5429 ( .A(n5499), .ZN(n5069) );
  NAND2_X1 U5430 ( .A1(n4960), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5852) );
  OR2_X1 U5431 ( .A1(n7972), .A2(n4844), .ZN(n5487) );
  AND2_X1 U5432 ( .A1(n5150), .A2(n8489), .ZN(n5149) );
  NAND2_X1 U5433 ( .A1(n8876), .A2(n5151), .ZN(n5150) );
  INV_X1 U5434 ( .A(n8633), .ZN(n5151) );
  NAND2_X1 U5435 ( .A1(n8638), .A2(n8639), .ZN(n8886) );
  NOR2_X1 U5436 ( .A1(n5177), .A2(n5175), .ZN(n5174) );
  OR2_X1 U5437 ( .A1(n9410), .A2(n9195), .ZN(n5175) );
  INV_X1 U5438 ( .A(n5253), .ZN(n5251) );
  INV_X1 U5439 ( .A(n9154), .ZN(n5250) );
  OR2_X1 U5440 ( .A1(n9442), .A2(n9257), .ZN(n8618) );
  INV_X1 U5441 ( .A(n8596), .ZN(n5040) );
  INV_X1 U5442 ( .A(n4957), .ZN(n5895) );
  OR2_X1 U5443 ( .A1(n9452), .A2(n9256), .ZN(n8652) );
  OR2_X1 U5444 ( .A1(n9281), .A2(n9296), .ZN(n8847) );
  NOR2_X1 U5445 ( .A1(n5764), .A2(n5763), .ZN(n4961) );
  NOR2_X1 U5446 ( .A1(n9467), .A2(n5159), .ZN(n5158) );
  INV_X1 U5447 ( .A(n5160), .ZN(n5159) );
  OR2_X1 U5448 ( .A1(n8472), .A2(n9332), .ZN(n9336) );
  NOR2_X1 U5449 ( .A1(n9474), .A2(n9477), .ZN(n5160) );
  NOR2_X1 U5450 ( .A1(n5170), .A2(n8379), .ZN(n5169) );
  NAND2_X1 U5451 ( .A1(n10554), .A2(n5171), .ZN(n5170) );
  INV_X1 U5452 ( .A(n5509), .ZN(n4958) );
  NAND2_X1 U5453 ( .A1(n7931), .A2(n10504), .ZN(n5164) );
  NAND2_X1 U5454 ( .A1(n7570), .A2(n9102), .ZN(n8528) );
  INV_X1 U5455 ( .A(n7708), .ZN(n7925) );
  AND2_X1 U5456 ( .A1(n5638), .A2(n5355), .ZN(n5664) );
  OAI21_X1 U5457 ( .B1(n5308), .B2(n5318), .A(n5305), .ZN(n7437) );
  NAND2_X1 U5458 ( .A1(n7108), .A2(n5306), .ZN(n5305) );
  AND2_X1 U5459 ( .A1(n5307), .A2(n7109), .ZN(n5306) );
  INV_X1 U5460 ( .A(n7114), .ZN(n7021) );
  AOI21_X1 U5461 ( .B1(n8073), .B2(n5286), .A(n4883), .ZN(n5284) );
  NAND2_X1 U5462 ( .A1(n8073), .A2(n5288), .ZN(n5285) );
  OR2_X1 U5463 ( .A1(n9874), .A2(n8707), .ZN(n6713) );
  OR2_X1 U5464 ( .A1(n8704), .A2(n8959), .ZN(n6652) );
  OR2_X1 U5465 ( .A1(n9885), .A2(n9745), .ZN(n6549) );
  OAI21_X1 U5466 ( .B1(n5238), .B2(n5237), .A(n4898), .ZN(n5236) );
  INV_X1 U5467 ( .A(n9806), .ZN(n8916) );
  NAND2_X1 U5468 ( .A1(n5059), .A2(n9846), .ZN(n5058) );
  INV_X1 U5469 ( .A(n5060), .ZN(n5059) );
  NAND2_X1 U5470 ( .A1(n9862), .A2(n9936), .ZN(n5060) );
  INV_X1 U5471 ( .A(n8358), .ZN(n5136) );
  NOR2_X1 U5472 ( .A1(n8276), .A2(n5210), .ZN(n8272) );
  NAND2_X1 U5473 ( .A1(n8271), .A2(n5211), .ZN(n5210) );
  INV_X1 U5474 ( .A(n8296), .ZN(n5211) );
  NAND2_X1 U5475 ( .A1(n5054), .A2(n5053), .ZN(n7865) );
  NAND2_X1 U5476 ( .A1(n8053), .A2(n4917), .ZN(n8329) );
  NAND2_X1 U5477 ( .A1(n6073), .A2(n6072), .ZN(n6531) );
  NAND2_X1 U5478 ( .A1(n6068), .A2(n6067), .ZN(n6073) );
  AOI21_X1 U5479 ( .B1(n5976), .B2(n5975), .A(n5974), .ZN(n5992) );
  NAND2_X1 U5480 ( .A1(n5116), .A2(n5114), .ZN(n5976) );
  AND2_X1 U5481 ( .A1(n5115), .A2(n5927), .ZN(n5114) );
  INV_X1 U5482 ( .A(n5947), .ZN(n5115) );
  AOI21_X1 U5483 ( .B1(n5110), .B2(n5114), .A(n5109), .ZN(n5108) );
  INV_X1 U5484 ( .A(n5972), .ZN(n5109) );
  INV_X1 U5485 ( .A(n5112), .ZN(n5110) );
  NAND2_X1 U5486 ( .A1(n6726), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U5487 ( .A1(n5908), .A2(n5112), .ZN(n5116) );
  INV_X1 U5488 ( .A(n5884), .ZN(n5093) );
  NOR2_X1 U5489 ( .A1(n5777), .A2(n5107), .ZN(n5106) );
  INV_X1 U5490 ( .A(n5757), .ZN(n5107) );
  XNOR2_X1 U5491 ( .A(n5704), .B(n10024), .ZN(n5703) );
  NAND2_X1 U5492 ( .A1(n5656), .A2(n5637), .ZN(n5657) );
  NAND2_X1 U5493 ( .A1(n5214), .A2(n5213), .ZN(n5658) );
  AOI21_X1 U5494 ( .B1(n4853), .B2(n5219), .A(n4888), .ZN(n5213) );
  NAND2_X1 U5495 ( .A1(n5577), .A2(SI_10_), .ZN(n5601) );
  NAND2_X1 U5496 ( .A1(n5558), .A2(n5557), .ZN(n5603) );
  XNOR2_X1 U5497 ( .A(n5532), .B(SI_7_), .ZN(n5529) );
  INV_X1 U5498 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6084) );
  INV_X1 U5499 ( .A(SI_1_), .ZN(n10169) );
  NAND2_X1 U5500 ( .A1(n5067), .A2(n5066), .ZN(n5385) );
  NAND2_X1 U5501 ( .A1(n5690), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U5502 ( .A1(n4961), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5822) );
  OR2_X1 U5503 ( .A1(n5716), .A2(n5715), .ZN(n5742) );
  AND2_X1 U5504 ( .A1(n4907), .A2(n5860), .ZN(n5203) );
  INV_X1 U5505 ( .A(n7400), .ZN(n5982) );
  INV_X1 U5506 ( .A(n7743), .ZN(n8511) );
  AOI21_X1 U5507 ( .B1(n7900), .B2(n5597), .A(n5328), .ZN(n7987) );
  NOR2_X1 U5508 ( .A1(n5596), .A2(n7908), .ZN(n5328) );
  NAND2_X1 U5509 ( .A1(n5191), .A2(n5190), .ZN(n5189) );
  INV_X1 U5510 ( .A(n9018), .ZN(n5191) );
  AOI21_X1 U5511 ( .B1(n4966), .B2(n8648), .A(n8647), .ZN(n8685) );
  MUX2_X1 U5512 ( .A(n8677), .B(n8678), .S(n8643), .Z(n8648) );
  NAND2_X1 U5513 ( .A1(n4946), .A2(n4967), .ZN(n4966) );
  AND2_X1 U5514 ( .A1(n5902), .A2(n5901), .ZN(n8483) );
  AND2_X1 U5515 ( .A1(n6033), .A2(n6032), .ZN(n6749) );
  NAND2_X1 U5516 ( .A1(n9158), .A2(n8633), .ZN(n8864) );
  AOI21_X1 U5517 ( .B1(n9151), .B2(n6051), .A(n5986), .ZN(n9069) );
  NAND2_X1 U5518 ( .A1(n9437), .A2(n8483), .ZN(n9206) );
  NAND2_X1 U5519 ( .A1(n9287), .A2(n4882), .ZN(n9201) );
  AND2_X1 U5520 ( .A1(n9287), .A2(n4863), .ZN(n9234) );
  NAND2_X1 U5521 ( .A1(n9287), .A2(n5173), .ZN(n5317) );
  NAND2_X1 U5522 ( .A1(n9287), .A2(n9271), .ZN(n9266) );
  AND2_X1 U5523 ( .A1(n9305), .A2(n9289), .ZN(n9287) );
  AND2_X1 U5524 ( .A1(n9272), .A2(n8604), .ZN(n9296) );
  OR2_X1 U5525 ( .A1(n4868), .A2(n8849), .ZN(n9282) );
  INV_X1 U5526 ( .A(n4961), .ZN(n5782) );
  NAND2_X1 U5527 ( .A1(n9378), .A2(n5158), .ZN(n9322) );
  AND2_X1 U5528 ( .A1(n8589), .A2(n9333), .ZN(n9368) );
  NAND2_X1 U5529 ( .A1(n8474), .A2(n9330), .ZN(n9387) );
  NOR2_X1 U5530 ( .A1(n8747), .A2(n10574), .ZN(n9378) );
  NAND2_X1 U5531 ( .A1(n9378), .A2(n9385), .ZN(n9379) );
  INV_X1 U5532 ( .A(n5025), .ZN(n5024) );
  AOI21_X1 U5533 ( .B1(n5025), .B2(n5023), .A(n5022), .ZN(n5021) );
  AND2_X1 U5534 ( .A1(n5026), .A2(n8669), .ZN(n5025) );
  NAND2_X1 U5535 ( .A1(n5168), .A2(n5166), .ZN(n8747) );
  NOR2_X1 U5536 ( .A1(n5167), .A2(n8396), .ZN(n5166) );
  INV_X1 U5537 ( .A(n5169), .ZN(n5167) );
  AND4_X1 U5538 ( .A1(n5649), .A2(n5648), .A3(n5647), .A4(n5646), .ZN(n8372)
         );
  NAND2_X1 U5539 ( .A1(n5168), .A2(n5169), .ZN(n8373) );
  AND4_X1 U5540 ( .A1(n5674), .A2(n5673), .A3(n5672), .A4(n5671), .ZN(n8393)
         );
  NOR2_X1 U5541 ( .A1(n8131), .A2(n5170), .ZN(n8342) );
  OR2_X1 U5542 ( .A1(n7945), .A2(n8829), .ZN(n7949) );
  NAND2_X1 U5543 ( .A1(n4958), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5543) );
  AND2_X1 U5544 ( .A1(n8664), .A2(n8830), .ZN(n8829) );
  NOR2_X1 U5545 ( .A1(n7773), .A2(n5162), .ZN(n8826) );
  NAND2_X1 U5546 ( .A1(n5163), .A2(n10511), .ZN(n5162) );
  INV_X1 U5547 ( .A(n5164), .ZN(n5163) );
  NAND2_X1 U5548 ( .A1(n5029), .A2(n5027), .ZN(n7955) );
  NAND2_X1 U5549 ( .A1(n5030), .A2(n5031), .ZN(n5029) );
  NAND2_X1 U5550 ( .A1(n5035), .A2(n7926), .ZN(n5031) );
  NOR2_X1 U5551 ( .A1(n4850), .A2(n10488), .ZN(n7758) );
  INV_X1 U5552 ( .A(n8657), .ZN(n8530) );
  AND2_X1 U5553 ( .A1(n5442), .A2(n5327), .ZN(n5446) );
  NAND2_X1 U5554 ( .A1(n5821), .A2(n5820), .ZN(n9459) );
  AND2_X1 U5555 ( .A1(n8113), .A2(n8112), .ZN(n8137) );
  INV_X1 U5556 ( .A(n8660), .ZN(n7934) );
  INV_X1 U5557 ( .A(n7778), .ZN(n7703) );
  INV_X1 U5558 ( .A(n5270), .ZN(n5050) );
  NAND2_X1 U5559 ( .A1(n5638), .A2(n5206), .ZN(n5737) );
  AND2_X1 U5560 ( .A1(n5464), .A2(n5463), .ZN(n10385) );
  NAND2_X1 U5561 ( .A1(n4893), .A2(n5067), .ZN(n5432) );
  NAND2_X1 U5562 ( .A1(n6174), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6460) );
  OR2_X1 U5563 ( .A1(n6460), .A2(n9535), .ZN(n6472) );
  OR2_X1 U5564 ( .A1(n6218), .A2(n9620), .ZN(n6209) );
  NOR2_X1 U5565 ( .A1(n9511), .A2(n5311), .ZN(n5310) );
  INV_X1 U5566 ( .A(n8934), .ZN(n5311) );
  NAND2_X1 U5567 ( .A1(n6143), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6320) );
  INV_X1 U5568 ( .A(n6281), .ZN(n6143) );
  AOI21_X1 U5569 ( .B1(n9520), .B2(n5275), .A(n4902), .ZN(n5274) );
  NOR2_X1 U5570 ( .A1(n7253), .A2(n5309), .ZN(n5308) );
  INV_X1 U5571 ( .A(n7250), .ZN(n5309) );
  INV_X1 U5572 ( .A(n8697), .ZN(n5304) );
  OR2_X1 U5573 ( .A1(n6322), .A2(n8241), .ZN(n6310) );
  OR2_X1 U5574 ( .A1(n8906), .A2(n9543), .ZN(n9599) );
  NAND2_X1 U5575 ( .A1(n6144), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6258) );
  INV_X1 U5576 ( .A(n6310), .ZN(n6144) );
  AND4_X1 U5577 ( .A1(n6351), .A2(n6350), .A3(n6349), .A4(n6348), .ZN(n7632)
         );
  NAND2_X1 U5578 ( .A1(n6376), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6380) );
  OR2_X1 U5579 ( .A1(n6389), .A2(n6375), .ZN(n6381) );
  NOR2_X1 U5580 ( .A1(n9729), .A2(n8704), .ZN(n9709) );
  AND2_X1 U5581 ( .A1(n6521), .A2(n6496), .ZN(n9739) );
  NOR3_X1 U5582 ( .A1(n9796), .A2(n9891), .A3(n5062), .ZN(n9737) );
  NOR2_X1 U5583 ( .A1(n9796), .A2(n5062), .ZN(n9752) );
  NAND2_X1 U5584 ( .A1(n5130), .A2(n5128), .ZN(n9804) );
  AOI21_X1 U5585 ( .B1(n5131), .B2(n5133), .A(n5129), .ZN(n5128) );
  INV_X1 U5586 ( .A(n8717), .ZN(n5129) );
  NOR2_X1 U5587 ( .A1(n9916), .A2(n9833), .ZN(n9812) );
  OR2_X1 U5588 ( .A1(n6194), .A2(n6160), .ZN(n6162) );
  NOR2_X1 U5589 ( .A1(n5319), .A2(n5060), .ZN(n9857) );
  INV_X1 U5590 ( .A(n5224), .ZN(n5221) );
  NOR2_X1 U5591 ( .A1(n5319), .A2(n9627), .ZN(n9856) );
  OR2_X1 U5592 ( .A1(n8431), .A2(n9942), .ZN(n5319) );
  AND2_X1 U5593 ( .A1(n8448), .A2(n8449), .ZN(n8444) );
  OR2_X1 U5594 ( .A1(n6244), .A2(n7802), .ZN(n6228) );
  AND3_X1 U5595 ( .A1(n6223), .A2(n6222), .A3(n6221), .ZN(n8784) );
  OR2_X1 U5596 ( .A1(n8322), .A2(n8268), .ZN(n8270) );
  NAND2_X1 U5597 ( .A1(n8253), .A2(n6621), .ZN(n8322) );
  NAND2_X1 U5598 ( .A1(n8248), .A2(n8247), .ZN(n8250) );
  NAND2_X1 U5599 ( .A1(n8053), .A2(n5065), .ZN(n8327) );
  NAND2_X1 U5600 ( .A1(n8053), .A2(n8209), .ZN(n8290) );
  INV_X1 U5601 ( .A(n9658), .ZN(n8089) );
  AND4_X1 U5602 ( .A1(n6315), .A2(n6314), .A3(n6313), .A4(n6312), .ZN(n9524)
         );
  NAND2_X1 U5603 ( .A1(n8040), .A2(n4952), .ZN(n8248) );
  NOR2_X1 U5604 ( .A1(n8041), .A2(n4953), .ZN(n4952) );
  INV_X1 U5605 ( .A(n8039), .ZN(n4953) );
  NAND2_X1 U5606 ( .A1(n8040), .A2(n8039), .ZN(n8173) );
  OR2_X1 U5607 ( .A1(n6295), .A2(n6279), .ZN(n6281) );
  OR2_X1 U5608 ( .A1(n7874), .A2(n9659), .ZN(n7869) );
  NAND2_X1 U5609 ( .A1(n6142), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6295) );
  INV_X1 U5610 ( .A(n6335), .ZN(n6142) );
  NAND2_X1 U5611 ( .A1(n6141), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6347) );
  INV_X1 U5612 ( .A(n6428), .ZN(n6141) );
  OR2_X1 U5613 ( .A1(n6347), .A2(n6333), .ZN(n6335) );
  AND2_X1 U5614 ( .A1(n7664), .A2(n7652), .ZN(n7594) );
  NAND2_X1 U5615 ( .A1(n7526), .A2(n7527), .ZN(n7592) );
  AND2_X1 U5616 ( .A1(n6685), .A2(n6686), .ZN(n7659) );
  NOR2_X1 U5617 ( .A1(n5321), .A2(n7781), .ZN(n7664) );
  NAND2_X1 U5618 ( .A1(n6139), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6426) );
  OR2_X1 U5619 ( .A1(n7323), .A2(n7529), .ZN(n5321) );
  NAND2_X1 U5620 ( .A1(n6683), .A2(n6681), .ZN(n7318) );
  NAND2_X1 U5621 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6411) );
  AND3_X1 U5622 ( .A1(n6408), .A2(n6407), .A3(n6406), .ZN(n7486) );
  NOR2_X1 U5623 ( .A1(n7278), .A2(n7296), .ZN(n7322) );
  NAND2_X1 U5624 ( .A1(n6670), .A2(n7142), .ZN(n7141) );
  NAND2_X1 U5625 ( .A1(n6372), .A2(n5322), .ZN(n7127) );
  NAND2_X1 U5626 ( .A1(n6226), .A2(n6225), .ZN(n9949) );
  AND2_X1 U5627 ( .A1(n6423), .A2(n6422), .ZN(n10497) );
  INV_X1 U5628 ( .A(n7354), .ZN(n10459) );
  INV_X1 U5629 ( .A(n6104), .ZN(n6101) );
  AND2_X1 U5630 ( .A1(n6105), .A2(n6102), .ZN(n5314) );
  XNOR2_X1 U5631 ( .A(n6531), .B(n6530), .ZN(n8490) );
  XNOR2_X1 U5632 ( .A(n6068), .B(n6067), .ZN(n8419) );
  XNOR2_X1 U5633 ( .A(n5992), .B(n5991), .ZN(n8387) );
  XNOR2_X1 U5634 ( .A(n5948), .B(n5947), .ZN(n8226) );
  NAND2_X1 U5635 ( .A1(n5116), .A2(n5927), .ZN(n5948) );
  OAI21_X1 U5636 ( .B1(n5847), .B2(n5092), .A(n5088), .ZN(n5890) );
  AOI21_X1 U5637 ( .B1(n5091), .B2(n5090), .A(n5089), .ZN(n5088) );
  INV_X1 U5638 ( .A(n5883), .ZN(n5089) );
  INV_X1 U5639 ( .A(n5097), .ZN(n5090) );
  NAND2_X1 U5640 ( .A1(n5094), .A2(n5095), .ZN(n5885) );
  NAND2_X1 U5641 ( .A1(n5847), .A2(n5097), .ZN(n5094) );
  INV_X1 U5642 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6667) );
  XNOR2_X1 U5643 ( .A(n5706), .B(n5703), .ZN(n6939) );
  NAND2_X1 U5644 ( .A1(n5683), .A2(n5682), .ZN(n5706) );
  NAND2_X1 U5645 ( .A1(n5081), .A2(n5086), .ZN(n5683) );
  NAND2_X1 U5646 ( .A1(n5658), .A2(n5656), .ZN(n5081) );
  NAND2_X1 U5647 ( .A1(n5215), .A2(n5216), .ZN(n5632) );
  OR2_X1 U5648 ( .A1(n5555), .A2(n5219), .ZN(n5215) );
  AOI21_X1 U5649 ( .B1(n5417), .B2(n5390), .A(n5323), .ZN(n5404) );
  XNOR2_X1 U5650 ( .A(n5405), .B(n10166), .ZN(n5403) );
  XNOR2_X1 U5651 ( .A(n5380), .B(n10169), .ZN(n5444) );
  AND2_X1 U5652 ( .A1(n5385), .A2(SI_0_), .ZN(n6370) );
  INV_X1 U5653 ( .A(n7939), .ZN(n10511) );
  NAND2_X1 U5654 ( .A1(n7516), .A2(n5508), .ZN(n6742) );
  AND2_X1 U5655 ( .A1(n5919), .A2(n5918), .ZN(n9186) );
  AND4_X1 U5656 ( .A1(n5571), .A2(n5570), .A3(n5569), .A4(n5568), .ZN(n8128)
         );
  INV_X1 U5657 ( .A(n10488), .ZN(n7573) );
  AOI21_X1 U5658 ( .B1(n6044), .B2(n6043), .A(n6042), .ZN(n6045) );
  OAI21_X1 U5659 ( .B1(n5504), .B2(n5201), .A(n5197), .ZN(n7731) );
  AOI21_X1 U5660 ( .B1(n5200), .B2(n5199), .A(n5198), .ZN(n5197) );
  INV_X1 U5661 ( .A(n5528), .ZN(n5198) );
  NAND2_X1 U5662 ( .A1(n7731), .A2(n7730), .ZN(n7900) );
  AOI21_X1 U5663 ( .B1(n5184), .B2(n5188), .A(n4856), .ZN(n5183) );
  NAND2_X1 U5664 ( .A1(n5850), .A2(n5849), .ZN(n9447) );
  AND4_X1 U5665 ( .A1(n5619), .A2(n5618), .A3(n5617), .A4(n5616), .ZN(n8337)
         );
  NAND2_X1 U5666 ( .A1(n5629), .A2(n5628), .ZN(n8146) );
  AND4_X1 U5667 ( .A1(n5352), .A2(n5351), .A3(n5350), .A4(n5349), .ZN(n7750)
         );
  AND4_X1 U5668 ( .A1(n5495), .A2(n5494), .A3(n5493), .A4(n5492), .ZN(n7933)
         );
  NAND2_X1 U5669 ( .A1(n9006), .A2(n5754), .ZN(n9018) );
  NAND2_X1 U5670 ( .A1(n5910), .A2(n5909), .ZN(n9431) );
  AND4_X1 U5671 ( .A1(n5591), .A2(n5590), .A3(n5589), .A4(n5588), .ZN(n8106)
         );
  NAND2_X1 U5672 ( .A1(n5564), .A2(n5563), .ZN(n10527) );
  INV_X1 U5673 ( .A(n7745), .ZN(n10470) );
  NAND2_X1 U5674 ( .A1(n8143), .A2(n5655), .ZN(n8218) );
  NAND2_X1 U5675 ( .A1(n5861), .A2(n5860), .ZN(n8970) );
  NAND2_X1 U5676 ( .A1(n5469), .A2(n7167), .ZN(n7172) );
  NAND2_X1 U5677 ( .A1(n5189), .A2(n5773), .ZN(n9056) );
  NAND2_X1 U5678 ( .A1(n5781), .A2(n5780), .ZN(n9462) );
  NAND2_X1 U5679 ( .A1(n5504), .A2(n7513), .ZN(n7516) );
  NAND2_X1 U5680 ( .A1(n8351), .A2(n5561), .ZN(n5955) );
  AND4_X1 U5681 ( .A1(n5748), .A2(n5747), .A3(n5746), .A4(n5745), .ZN(n9344)
         );
  NAND2_X1 U5682 ( .A1(n4959), .A2(n6005), .ZN(n9084) );
  NAND2_X1 U5683 ( .A1(n8861), .A2(n6051), .ZN(n4959) );
  NAND4_X1 U5684 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), .ZN(n9096)
         );
  INV_X1 U5685 ( .A(n7933), .ZN(n9098) );
  INV_X1 U5686 ( .A(n7750), .ZN(n9100) );
  NOR2_X1 U5687 ( .A1(n4879), .A2(n5267), .ZN(n5266) );
  OR2_X1 U5688 ( .A1(n5450), .A2(n5425), .ZN(n5426) );
  XNOR2_X1 U5689 ( .A(n8836), .B(n9398), .ZN(n9400) );
  AOI21_X1 U5690 ( .B1(n8495), .B2(n5561), .A(n8494), .ZN(n8755) );
  NAND2_X1 U5691 ( .A1(n5248), .A2(n5252), .ZN(n9148) );
  AOI21_X1 U5692 ( .B1(n9172), .B2(n10467), .A(n9171), .ZN(n9424) );
  AOI21_X1 U5693 ( .B1(n9182), .B2(n9181), .A(n8858), .ZN(n9163) );
  AND2_X1 U5694 ( .A1(n5958), .A2(n5937), .ZN(n9194) );
  NAND2_X1 U5695 ( .A1(n9223), .A2(n8855), .ZN(n9200) );
  AND2_X1 U5696 ( .A1(n9240), .A2(n9239), .ZN(n9445) );
  NAND2_X1 U5697 ( .A1(n8482), .A2(n5165), .ZN(n9259) );
  NAND2_X1 U5698 ( .A1(n9264), .A2(n8851), .ZN(n9248) );
  AND2_X1 U5699 ( .A1(n9317), .A2(n9316), .ZN(n9465) );
  AND2_X1 U5700 ( .A1(n8398), .A2(n8397), .ZN(n8399) );
  AND2_X1 U5701 ( .A1(n8381), .A2(n8380), .ZN(n8382) );
  NAND2_X1 U5702 ( .A1(n8138), .A2(n8114), .ZN(n8115) );
  NAND2_X1 U5703 ( .A1(n6824), .A2(n5561), .ZN(n4941) );
  NAND2_X1 U5704 ( .A1(n5541), .A2(n5540), .ZN(n10520) );
  NAND2_X1 U5705 ( .A1(n5258), .A2(n7932), .ZN(n7975) );
  NAND2_X1 U5706 ( .A1(n5034), .A2(n8542), .ZN(n7970) );
  NAND2_X1 U5707 ( .A1(n7706), .A2(n5036), .ZN(n5034) );
  OR2_X1 U5708 ( .A1(n8503), .A2(n6790), .ZN(n5408) );
  OR2_X1 U5709 ( .A1(n9393), .A2(n7717), .ZN(n10475) );
  OR2_X1 U5710 ( .A1(n7385), .A2(n8689), .ZN(n10471) );
  INV_X1 U5711 ( .A(n10475), .ZN(n9353) );
  OR2_X1 U5712 ( .A1(n9393), .A2(n10564), .ZN(n10476) );
  NAND2_X1 U5713 ( .A1(n9406), .A2(n10576), .ZN(n5140) );
  INV_X1 U5714 ( .A(n5142), .ZN(n5141) );
  OAI21_X1 U5715 ( .B1(n9408), .B2(n10564), .A(n5143), .ZN(n5142) );
  AND2_X1 U5716 ( .A1(n9413), .A2(n9412), .ZN(n9414) );
  OR2_X1 U5717 ( .A1(n5367), .A2(n5343), .ZN(n5369) );
  XNOR2_X1 U5718 ( .A(n5359), .B(n5358), .ZN(n5364) );
  NAND2_X1 U5719 ( .A1(n5194), .A2(n5193), .ZN(n5359) );
  AOI21_X1 U5720 ( .B1(n5195), .B2(n5343), .A(n5343), .ZN(n5193) );
  NAND2_X1 U5721 ( .A1(n4985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U5722 ( .A1(n5779), .A2(n5357), .ZN(n4985) );
  AND2_X1 U5723 ( .A1(n6515), .A2(n6514), .ZN(n9744) );
  OR2_X1 U5724 ( .A1(n9753), .A2(n6535), .ZN(n6515) );
  NAND2_X1 U5725 ( .A1(n8913), .A2(n8914), .ZN(n9531) );
  OR2_X1 U5726 ( .A1(n8913), .A2(n8914), .ZN(n9532) );
  NAND2_X1 U5727 ( .A1(n6459), .A2(n6458), .ZN(n9911) );
  NAND2_X1 U5728 ( .A1(n7108), .A2(n7109), .ZN(n7251) );
  OR2_X1 U5729 ( .A1(n8795), .A2(n5295), .ZN(n5290) );
  NAND2_X1 U5730 ( .A1(n6191), .A2(n6190), .ZN(n9931) );
  XNOR2_X1 U5731 ( .A(n8952), .B(n8951), .ZN(n8953) );
  AOI21_X1 U5732 ( .B1(n5302), .B2(n5299), .A(n4894), .ZN(n5297) );
  NAND2_X1 U5733 ( .A1(n9638), .A2(n9640), .ZN(n9565) );
  AND2_X1 U5734 ( .A1(n6491), .A2(n6490), .ZN(n9783) );
  OAI21_X1 U5735 ( .B1(n8913), .B2(n5302), .A(n5301), .ZN(n9589) );
  NAND2_X1 U5736 ( .A1(n7251), .A2(n7250), .ZN(n7252) );
  AOI21_X1 U5737 ( .B1(n4862), .B2(n5295), .A(n4922), .ZN(n5291) );
  NAND2_X1 U5738 ( .A1(n6159), .A2(n6158), .ZN(n9926) );
  NAND2_X1 U5739 ( .A1(n6308), .A2(n6307), .ZN(n9963) );
  INV_X1 U5740 ( .A(n9623), .ZN(n9642) );
  INV_X1 U5741 ( .A(n8179), .ZN(n10012) );
  INV_X1 U5742 ( .A(n7665), .ZN(n7781) );
  NAND2_X1 U5743 ( .A1(n6662), .A2(n9834), .ZN(n5078) );
  NAND2_X1 U5744 ( .A1(n5075), .A2(n7541), .ZN(n4999) );
  AND4_X1 U5745 ( .A1(n6326), .A2(n6325), .A3(n6324), .A4(n6323), .ZN(n8196)
         );
  OR3_X1 U5746 ( .A1(n6433), .A2(n6432), .A3(n6431), .ZN(n9661) );
  CLKBUF_X1 U5747 ( .A(n7072), .Z(n9664) );
  OR2_X1 U5748 ( .A1(n6378), .A2(n6354), .ZN(n6355) );
  OR2_X1 U5749 ( .A1(n6389), .A2(n6847), .ZN(n6356) );
  XNOR2_X1 U5750 ( .A(n9708), .B(n9874), .ZN(n9876) );
  NAND2_X1 U5751 ( .A1(n6107), .A2(n6106), .ZN(n9878) );
  NAND2_X1 U5752 ( .A1(n5235), .A2(n5238), .ZN(n9736) );
  NAND2_X1 U5753 ( .A1(n5242), .A2(n4867), .ZN(n5235) );
  AND2_X1 U5754 ( .A1(n6505), .A2(n6504), .ZN(n9756) );
  NAND2_X1 U5755 ( .A1(n8351), .A2(n6340), .ZN(n6505) );
  NAND2_X1 U5756 ( .A1(n5240), .A2(n5245), .ZN(n9751) );
  NAND2_X1 U5757 ( .A1(n5242), .A2(n5241), .ZN(n5240) );
  NAND2_X1 U5758 ( .A1(n6471), .A2(n6470), .ZN(n9908) );
  INV_X1 U5759 ( .A(n9911), .ZN(n9802) );
  NAND2_X1 U5760 ( .A1(n5230), .A2(n5231), .ZN(n5229) );
  NAND2_X1 U5761 ( .A1(n9828), .A2(n8716), .ZN(n9818) );
  NOR2_X1 U5762 ( .A1(n9824), .A2(n5232), .ZN(n9811) );
  NAND2_X1 U5763 ( .A1(n6138), .A2(n6137), .ZN(n9922) );
  NAND2_X1 U5764 ( .A1(n8713), .A2(n5124), .ZN(n5117) );
  INV_X1 U5765 ( .A(n9926), .ZN(n9846) );
  NAND2_X1 U5766 ( .A1(n5126), .A2(n5124), .ZN(n9863) );
  AND2_X1 U5767 ( .A1(n8453), .A2(n5222), .ZN(n8731) );
  NAND2_X1 U5768 ( .A1(n8453), .A2(n8452), .ZN(n8455) );
  NAND2_X1 U5769 ( .A1(n6241), .A2(n6240), .ZN(n9952) );
  NAND2_X1 U5770 ( .A1(n6237), .A2(n6340), .ZN(n6241) );
  AND2_X1 U5771 ( .A1(n8311), .A2(n8253), .ZN(n8255) );
  NAND2_X1 U5772 ( .A1(n6278), .A2(n6277), .ZN(n8083) );
  NAND2_X1 U5773 ( .A1(n7813), .A2(n7812), .ZN(n7815) );
  INV_X1 U5774 ( .A(n10497), .ZN(n7529) );
  AND3_X1 U5775 ( .A1(n6397), .A2(n6396), .A3(n6395), .ZN(n7508) );
  AND2_X1 U5776 ( .A1(n10447), .A2(n7483), .ZN(n10006) );
  AND2_X1 U5777 ( .A1(n10447), .A2(n7311), .ZN(n9827) );
  INV_X1 U5778 ( .A(n7127), .ZN(n10441) );
  NAND2_X1 U5779 ( .A1(n9883), .A2(n4880), .ZN(n9972) );
  AOI21_X1 U5780 ( .B1(n9882), .B2(n9965), .A(n4920), .ZN(n4954) );
  AND2_X1 U5781 ( .A1(n9888), .A2(n9887), .ZN(n9889) );
  XNOR2_X1 U5782 ( .A(n6131), .B(n6130), .ZN(n9997) );
  NAND2_X1 U5783 ( .A1(n6127), .A2(n6126), .ZN(n6131) );
  NAND2_X1 U5784 ( .A1(n6104), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4956) );
  INV_X1 U5785 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6575) );
  NAND2_X1 U5786 ( .A1(n5074), .A2(n5499), .ZN(n5518) );
  NOR2_X1 U5787 ( .A1(n9742), .A2(n5139), .ZN(n5138) );
  NAND2_X1 U5788 ( .A1(n4962), .A2(n5018), .ZN(P2_U3244) );
  OR2_X1 U5789 ( .A1(n8693), .A2(n8692), .ZN(n5018) );
  NAND2_X1 U5790 ( .A1(n4943), .A2(n5019), .ZN(n4962) );
  AND2_X1 U5791 ( .A1(n5137), .A2(n8725), .ZN(n8726) );
  INV_X2 U5792 ( .A(n6378), .ZN(n6424) );
  OR2_X1 U5793 ( .A1(n10469), .A2(n7769), .ZN(n4850) );
  AND2_X1 U5794 ( .A1(n6700), .A2(n6642), .ZN(n4851) );
  NAND2_X1 U5795 ( .A1(n4857), .A2(n8712), .ZN(n5125) );
  AND2_X1 U5796 ( .A1(n8254), .A2(n8253), .ZN(n4852) );
  AND2_X1 U5797 ( .A1(n5216), .A2(n5630), .ZN(n4853) );
  AND2_X1 U5798 ( .A1(n8574), .A2(n8575), .ZN(n8668) );
  NAND2_X1 U5799 ( .A1(n8725), .A2(n6578), .ZN(n9742) );
  INV_X1 U5800 ( .A(n9742), .ZN(n5237) );
  OR2_X1 U5801 ( .A1(n6383), .A2(n6786), .ZN(n4854) );
  AND2_X1 U5802 ( .A1(n4903), .A2(n5312), .ZN(n4855) );
  AND2_X1 U5803 ( .A1(n6600), .A2(n7812), .ZN(n7810) );
  AND2_X1 U5804 ( .A1(n5965), .A2(n5964), .ZN(n9187) );
  OAI21_X1 U5805 ( .B1(n7641), .B2(n7642), .A(n5287), .ZN(n5286) );
  NOR2_X1 U5806 ( .A1(n5843), .A2(n5842), .ZN(n4856) );
  AND2_X1 U5807 ( .A1(n6632), .A2(n8714), .ZN(n4857) );
  AND2_X1 U5808 ( .A1(n6780), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4858) );
  AND2_X1 U5809 ( .A1(n5257), .A2(n9187), .ZN(n4859) );
  AND2_X1 U5810 ( .A1(n7934), .A2(n7932), .ZN(n4860) );
  AND2_X1 U5811 ( .A1(n5314), .A2(n6108), .ZN(n4861) );
  AND2_X1 U5812 ( .A1(n5292), .A2(n5293), .ZN(n4862) );
  NAND2_X1 U5813 ( .A1(n9378), .A2(n5160), .ZN(n5161) );
  AND2_X1 U5814 ( .A1(n5172), .A2(n5173), .ZN(n4863) );
  INV_X1 U5815 ( .A(n7513), .ZN(n5199) );
  NAND2_X1 U5816 ( .A1(n7594), .A2(n7596), .ZN(n7820) );
  INV_X1 U5817 ( .A(n7820), .ZN(n5054) );
  INV_X2 U5818 ( .A(n6383), .ZN(n6340) );
  INV_X1 U5819 ( .A(n7128), .ZN(n7343) );
  NAND2_X1 U5820 ( .A1(n9222), .A2(n9221), .ZN(n9223) );
  AND2_X1 U5821 ( .A1(n5332), .A2(n5155), .ZN(n4864) );
  NOR2_X1 U5822 ( .A1(n8261), .A2(n8266), .ZN(n4865) );
  OR2_X1 U5823 ( .A1(n8427), .A2(n5136), .ZN(n4866) );
  AND2_X1 U5824 ( .A1(n5244), .A2(n5241), .ZN(n4867) );
  NOR2_X1 U5825 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6360) );
  OAI211_X1 U5826 ( .C1(n6803), .C2(n6383), .A(n6385), .B(n4995), .ZN(n6386)
         );
  NOR2_X1 U5827 ( .A1(n9462), .A2(n9089), .ZN(n4868) );
  AND2_X1 U5828 ( .A1(n5360), .A2(n5268), .ZN(n5367) );
  OR2_X1 U5829 ( .A1(n9891), .A2(n8941), .ZN(n8725) );
  NAND2_X1 U5830 ( .A1(n9816), .A2(n9536), .ZN(n4869) );
  AND2_X1 U5831 ( .A1(n8671), .A2(n8397), .ZN(n4870) );
  NAND2_X1 U5832 ( .A1(n5298), .A2(n5297), .ZN(n9554) );
  NAND2_X1 U5833 ( .A1(n5290), .A2(n5293), .ZN(n8810) );
  AND2_X1 U5834 ( .A1(n5229), .A2(n4869), .ZN(n9794) );
  AND2_X1 U5835 ( .A1(n5904), .A2(n5903), .ZN(n4871) );
  NOR3_X1 U5836 ( .A1(n9410), .A2(n9156), .A3(n8637), .ZN(n4872) );
  INV_X1 U5837 ( .A(n7769), .ZN(n7570) );
  OAI211_X1 U5838 ( .C1(n6751), .C2(n6784), .A(n5468), .B(n5467), .ZN(n7769)
         );
  AND2_X1 U5839 ( .A1(n5459), .A2(n5329), .ZN(n5373) );
  NAND2_X1 U5840 ( .A1(n8482), .A2(n8651), .ZN(n9254) );
  OR3_X1 U5841 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4873) );
  INV_X1 U5842 ( .A(n9017), .ZN(n5190) );
  AND2_X1 U5843 ( .A1(n9916), .A2(n9831), .ZN(n4874) );
  AND3_X1 U5844 ( .A1(n6635), .A2(n9848), .A3(n9830), .ZN(n4875) );
  NOR2_X1 U5845 ( .A1(n9178), .A2(n9422), .ZN(n4876) );
  NAND2_X1 U5846 ( .A1(n5153), .A2(n5154), .ZN(n5361) );
  NAND2_X1 U5847 ( .A1(n5807), .A2(n5806), .ZN(n9452) );
  AND2_X1 U5848 ( .A1(n9255), .A2(n8851), .ZN(n4877) );
  AND2_X1 U5849 ( .A1(n8727), .A2(n8725), .ZN(n4878) );
  NAND2_X1 U5850 ( .A1(n8724), .A2(n5138), .ZN(n5137) );
  INV_X1 U5851 ( .A(n5063), .ZN(n9766) );
  NOR3_X1 U5852 ( .A1(n9796), .A2(n9901), .A3(n9908), .ZN(n5063) );
  XNOR2_X1 U5853 ( .A(n5631), .B(n10051), .ZN(n5630) );
  INV_X1 U5854 ( .A(n8543), .ZN(n5147) );
  AND2_X1 U5855 ( .A1(n5436), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4879) );
  AND2_X1 U5856 ( .A1(n9884), .A2(n4954), .ZN(n4880) );
  AND2_X1 U5857 ( .A1(n9756), .A2(n9744), .ZN(n4881) );
  AND2_X1 U5858 ( .A1(n9229), .A2(n4863), .ZN(n4882) );
  AND2_X1 U5859 ( .A1(n8072), .A2(n8071), .ZN(n4883) );
  AND2_X1 U5860 ( .A1(n6503), .A2(n6502), .ZN(n8941) );
  INV_X1 U5861 ( .A(n8941), .ZN(n5243) );
  AND2_X1 U5862 ( .A1(n6641), .A2(n9805), .ZN(n4884) );
  INV_X1 U5863 ( .A(n7641), .ZN(n5288) );
  NOR2_X1 U5864 ( .A1(n4871), .A2(n5906), .ZN(n4885) );
  INV_X1 U5865 ( .A(n5176), .ZN(n9149) );
  NOR2_X1 U5866 ( .A1(n9178), .A2(n5177), .ZN(n5176) );
  INV_X1 U5867 ( .A(n5283), .ZN(n8075) );
  OAI21_X1 U5868 ( .B1(n7640), .B2(n5285), .A(n5284), .ZN(n5283) );
  OR2_X1 U5869 ( .A1(n4993), .A2(n4992), .ZN(n4886) );
  AND2_X1 U5870 ( .A1(n5704), .A2(SI_14_), .ZN(n4887) );
  AND2_X1 U5871 ( .A1(n5631), .A2(SI_11_), .ZN(n4888) );
  AOI21_X1 U5872 ( .B1(n5253), .B2(n8858), .A(n4859), .ZN(n5252) );
  NOR2_X1 U5873 ( .A1(n8649), .A2(n8516), .ZN(n4889) );
  OR2_X1 U5874 ( .A1(n6719), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4890) );
  AND2_X1 U5875 ( .A1(n6669), .A2(n6668), .ZN(n4891) );
  AND2_X1 U5876 ( .A1(n5077), .A2(n6713), .ZN(n4892) );
  AND2_X1 U5877 ( .A1(n6552), .A2(n8715), .ZN(n9848) );
  INV_X1 U5878 ( .A(n9848), .ZN(n5119) );
  INV_X1 U5879 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5049) );
  AND2_X1 U5880 ( .A1(n5066), .A2(n5379), .ZN(n4893) );
  INV_X1 U5881 ( .A(n5201), .ZN(n5200) );
  NAND2_X1 U5882 ( .A1(n5202), .A2(n5508), .ZN(n5201) );
  AND2_X1 U5883 ( .A1(n6551), .A2(n8716), .ZN(n9830) );
  AND2_X1 U5884 ( .A1(n8921), .A2(n8920), .ZN(n4894) );
  INV_X1 U5885 ( .A(n5318), .ZN(n5307) );
  INV_X1 U5886 ( .A(n5185), .ZN(n5184) );
  NAND2_X1 U5887 ( .A1(n5834), .A2(n5186), .ZN(n5185) );
  NOR2_X1 U5888 ( .A1(n9296), .A2(n9282), .ZN(n4895) );
  OR2_X1 U5889 ( .A1(n9098), .A2(n10504), .ZN(n4896) );
  NAND2_X1 U5890 ( .A1(n4867), .A2(n9742), .ZN(n4897) );
  OR2_X1 U5891 ( .A1(n9891), .A2(n5243), .ZN(n4898) );
  AND2_X1 U5892 ( .A1(n5056), .A2(n5055), .ZN(n4899) );
  INV_X1 U5893 ( .A(n4960), .ZN(n5824) );
  NOR2_X1 U5894 ( .A1(n5822), .A2(n10188), .ZN(n4960) );
  OR2_X1 U5895 ( .A1(n8550), .A2(n4980), .ZN(n4900) );
  OR2_X1 U5896 ( .A1(n5705), .A2(n5209), .ZN(n4901) );
  NAND2_X1 U5897 ( .A1(n9564), .A2(n5276), .ZN(n4902) );
  NOR2_X1 U5898 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4903) );
  AOI21_X1 U5899 ( .B1(n7127), .B2(n8936), .A(n7022), .ZN(n7026) );
  OR2_X1 U5900 ( .A1(n4881), .A2(n5239), .ZN(n4904) );
  AND2_X1 U5901 ( .A1(n8509), .A2(n5020), .ZN(n4905) );
  OR2_X1 U5902 ( .A1(n9715), .A2(n9745), .ZN(n4906) );
  NOR2_X1 U5903 ( .A1(n9049), .A2(n4871), .ZN(n4907) );
  NOR2_X1 U5904 ( .A1(n8437), .A2(n8436), .ZN(n4908) );
  AND4_X1 U5905 ( .A1(n5458), .A2(n5457), .A3(n5456), .A4(n5455), .ZN(n7751)
         );
  INV_X1 U5906 ( .A(n7751), .ZN(n9102) );
  NOR2_X1 U5907 ( .A1(n4874), .A2(n5232), .ZN(n5231) );
  AND4_X1 U5908 ( .A1(n5414), .A2(n5413), .A3(n5412), .A4(n5411), .ZN(n7578)
         );
  NOR2_X1 U5909 ( .A1(n8688), .A2(n4905), .ZN(n4909) );
  AND2_X1 U5910 ( .A1(n8440), .A2(n5221), .ZN(n4910) );
  AND2_X1 U5911 ( .A1(n5519), .A2(SI_6_), .ZN(n4911) );
  AND2_X1 U5912 ( .A1(n8587), .A2(n9377), .ZN(n4912) );
  AND2_X1 U5913 ( .A1(n8733), .A2(n4869), .ZN(n4913) );
  AND2_X1 U5914 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n4914) );
  INV_X1 U5915 ( .A(n4982), .ZN(n4981) );
  NAND2_X1 U5916 ( .A1(n8554), .A2(n8832), .ZN(n4982) );
  INV_X2 U5917 ( .A(n6389), .ZN(n6368) );
  NAND2_X1 U5918 ( .A1(n6481), .A2(n6480), .ZN(n9901) );
  NAND2_X1 U5919 ( .A1(n5261), .A2(n8846), .ZN(n9280) );
  XNOR2_X1 U5920 ( .A(n9084), .B(n9410), .ZN(n8876) );
  INV_X1 U5921 ( .A(n8876), .ZN(n5152) );
  NAND2_X1 U5922 ( .A1(n6534), .A2(n6533), .ZN(n8704) );
  AOI21_X1 U5923 ( .B1(n7640), .B2(n7642), .A(n7641), .ZN(n8061) );
  NAND2_X1 U5924 ( .A1(n5274), .A2(n5273), .ZN(n9563) );
  NAND2_X1 U5925 ( .A1(n5189), .A2(n5187), .ZN(n8982) );
  XOR2_X1 U5926 ( .A(n8772), .B(n8947), .Z(n4915) );
  INV_X1 U5927 ( .A(n5092), .ZN(n5091) );
  NAND2_X1 U5928 ( .A1(n5095), .A2(n5093), .ZN(n5092) );
  NAND2_X1 U5929 ( .A1(n8359), .A2(n8358), .ZN(n8428) );
  NAND2_X1 U5930 ( .A1(n5117), .A2(n5121), .ZN(n9847) );
  OAI21_X1 U5931 ( .B1(n9018), .B2(n5185), .A(n5183), .ZN(n8991) );
  NAND2_X1 U5932 ( .A1(n6207), .A2(n6206), .ZN(n9627) );
  INV_X1 U5933 ( .A(n8714), .ZN(n5122) );
  NAND2_X1 U5934 ( .A1(n6254), .A2(n6253), .ZN(n9958) );
  INV_X1 U5935 ( .A(n9958), .ZN(n5064) );
  OAI21_X1 U5936 ( .B1(n8370), .B2(n5024), .A(n5021), .ZN(n8391) );
  NAND2_X1 U5937 ( .A1(n9896), .A2(n9744), .ZN(n8723) );
  INV_X1 U5938 ( .A(n8723), .ZN(n5139) );
  NAND2_X1 U5939 ( .A1(n9176), .A2(n5174), .ZN(n8880) );
  NAND2_X1 U5940 ( .A1(n6493), .A2(n6492), .ZN(n9891) );
  NOR3_X1 U5941 ( .A1(n5319), .A2(n5058), .A3(n9922), .ZN(n5061) );
  AND4_X1 U5942 ( .A1(n5787), .A2(n5786), .A3(n5785), .A4(n5784), .ZN(n9342)
         );
  OR2_X1 U5943 ( .A1(n9802), .A2(n9781), .ZN(n4916) );
  AND2_X1 U5944 ( .A1(n5065), .A2(n5064), .ZN(n4917) );
  NAND2_X1 U5945 ( .A1(n6318), .A2(n6317), .ZN(n8258) );
  INV_X1 U5946 ( .A(n8796), .ZN(n5294) );
  NAND2_X1 U5947 ( .A1(n5713), .A2(n5712), .ZN(n9477) );
  INV_X1 U5948 ( .A(n10504), .ZN(n8549) );
  AND3_X1 U5949 ( .A1(n5503), .A2(n5502), .A3(n5501), .ZN(n10504) );
  INV_X1 U5950 ( .A(n5188), .ZN(n5187) );
  NAND2_X1 U5951 ( .A1(n5192), .A2(n5773), .ZN(n5188) );
  AND2_X1 U5952 ( .A1(n5126), .A2(n8712), .ZN(n4918) );
  AND2_X1 U5953 ( .A1(n8856), .A2(n8855), .ZN(n4919) );
  AND2_X1 U5954 ( .A1(n8704), .A2(n9964), .ZN(n4920) );
  INV_X1 U5955 ( .A(n5125), .ZN(n5124) );
  NAND2_X1 U5956 ( .A1(n9264), .A2(n4877), .ZN(n9246) );
  INV_X1 U5957 ( .A(n5057), .ZN(n9841) );
  NOR2_X1 U5958 ( .A1(n5319), .A2(n5058), .ZN(n5057) );
  NAND2_X1 U5959 ( .A1(n8441), .A2(n8440), .ZN(n8453) );
  INV_X1 U5960 ( .A(n5104), .ZN(n5103) );
  OAI21_X1 U5961 ( .B1(n5777), .B2(n5105), .A(n5776), .ZN(n5104) );
  INV_X1 U5962 ( .A(n5848), .ZN(n5099) );
  NOR2_X1 U5963 ( .A1(n9896), .A2(n9908), .ZN(n4921) );
  NAND2_X1 U5964 ( .A1(n5935), .A2(n5934), .ZN(n9195) );
  INV_X1 U5965 ( .A(n9416), .ZN(n9153) );
  NAND2_X1 U5966 ( .A1(n5981), .A2(n5980), .ZN(n9416) );
  NAND2_X1 U5967 ( .A1(n5279), .A2(n5278), .ZN(n5277) );
  AND2_X1 U5968 ( .A1(n7744), .A2(n10471), .ZN(n9393) );
  XNOR2_X1 U5969 ( .A(n5369), .B(n5368), .ZN(n6053) );
  NAND2_X1 U5970 ( .A1(n4941), .A2(n5585), .ZN(n8136) );
  INV_X1 U5971 ( .A(n8136), .ZN(n5171) );
  NAND2_X1 U5972 ( .A1(n8113), .A2(n5265), .ZN(n8138) );
  AOI21_X1 U5973 ( .B1(n5484), .B2(n7374), .A(n5483), .ZN(n7375) );
  NAND2_X1 U5974 ( .A1(n7813), .A2(n4951), .ZN(n7861) );
  NAND2_X1 U5975 ( .A1(n6398), .A2(n6679), .ZN(n7317) );
  AOI21_X1 U5976 ( .B1(n7525), .B2(n7524), .A(n7523), .ZN(n7526) );
  AND2_X1 U5977 ( .A1(n8802), .A2(n8801), .ZN(n4922) );
  AND2_X1 U5978 ( .A1(n8052), .A2(n10012), .ZN(n8053) );
  NAND2_X1 U5979 ( .A1(n7567), .A2(n7749), .ZN(n7706) );
  NAND2_X1 U5980 ( .A1(n5871), .A2(n5870), .ZN(n9442) );
  INV_X1 U5981 ( .A(n9442), .ZN(n5172) );
  NAND2_X1 U5982 ( .A1(n5955), .A2(n5954), .ZN(n9422) );
  INV_X1 U5983 ( .A(n9422), .ZN(n5257) );
  INV_X1 U5984 ( .A(n4915), .ZN(n5279) );
  OR2_X1 U5985 ( .A1(n6013), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4923) );
  OR2_X1 U5986 ( .A1(n8824), .A2(n10527), .ZN(n8131) );
  INV_X1 U5987 ( .A(n8131), .ZN(n5168) );
  AND2_X1 U5988 ( .A1(n7516), .A2(n5200), .ZN(n4924) );
  NOR2_X1 U5989 ( .A1(n7773), .A2(n5164), .ZN(n4925) );
  AND2_X1 U5990 ( .A1(n5308), .A2(n7251), .ZN(n4926) );
  INV_X1 U5991 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5208) );
  INV_X1 U5992 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U5993 ( .A1(n6292), .A2(n6291), .ZN(n7874) );
  INV_X1 U5994 ( .A(n7874), .ZN(n5053) );
  OAI211_X1 U5995 ( .C1(n6751), .C2(n6968), .A(n5409), .B(n5408), .ZN(n7718)
         );
  OR2_X1 U5996 ( .A1(n8687), .A2(n8686), .ZN(n4927) );
  NOR2_X1 U5997 ( .A1(n5345), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n9501) );
  OR2_X1 U5998 ( .A1(n7151), .A2(n7064), .ZN(n10450) );
  OR2_X1 U5999 ( .A1(n7030), .A2(n9834), .ZN(n6659) );
  XNOR2_X2 U6000 ( .A(n6189), .B(n6188), .ZN(n9834) );
  INV_X2 U6001 ( .A(n7289), .ZN(n9503) );
  NAND2_X1 U6002 ( .A1(n4928), .A2(n8637), .ZN(n8602) );
  NAND2_X1 U6003 ( .A1(n4929), .A2(n8596), .ZN(n4928) );
  NAND2_X1 U6004 ( .A1(n8603), .A2(n4930), .ZN(n4929) );
  INV_X1 U6005 ( .A(n8604), .ZN(n4931) );
  NAND2_X1 U6006 ( .A1(n8598), .A2(n8597), .ZN(n8603) );
  NAND2_X1 U6007 ( .A1(n4932), .A2(n4965), .ZN(n8591) );
  NAND2_X1 U6008 ( .A1(n4933), .A2(n4912), .ZN(n4932) );
  NAND3_X1 U6009 ( .A1(n4934), .A2(n8584), .A3(n8583), .ZN(n4933) );
  NAND3_X1 U6010 ( .A1(n8580), .A2(n8669), .A3(n8579), .ZN(n4934) );
  NAND2_X1 U6011 ( .A1(n4940), .A2(n5432), .ZN(n5380) );
  NAND3_X1 U6012 ( .A1(n4944), .A2(n8682), .A3(n4909), .ZN(n4943) );
  NAND3_X1 U6013 ( .A1(n5378), .A2(n4950), .A3(n4949), .ZN(n5067) );
  INV_X1 U6014 ( .A(n7142), .ZN(n7133) );
  AND2_X1 U6015 ( .A1(n6676), .A2(n6674), .ZN(n7142) );
  NAND2_X1 U6016 ( .A1(n4958), .A2(n4914), .ZN(n5565) );
  OAI211_X1 U6017 ( .C1(n4975), .C2(n4982), .A(n8555), .B(n4973), .ZN(n8557)
         );
  NAND2_X1 U6018 ( .A1(n5154), .A2(n4983), .ZN(n5562) );
  INV_X2 U6019 ( .A(n5401), .ZN(n5154) );
  OAI21_X1 U6020 ( .B1(n4875), .B2(n4987), .A(n4986), .ZN(n6646) );
  INV_X1 U6021 ( .A(n9817), .ZN(n4992) );
  INV_X1 U6022 ( .A(n6590), .ZN(n6589) );
  NAND2_X1 U6023 ( .A1(n4997), .A2(n6738), .ZN(P1_U3240) );
  NAND2_X1 U6024 ( .A1(n4998), .A2(n6725), .ZN(n4997) );
  NAND3_X1 U6025 ( .A1(n4891), .A2(n5078), .A3(n4999), .ZN(n4998) );
  NAND2_X1 U6026 ( .A1(n5005), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6103) );
  NAND4_X1 U6027 ( .A1(n5006), .A2(n6099), .A3(n4855), .A4(n6098), .ZN(n5005)
         );
  NAND4_X1 U6028 ( .A1(n6099), .A2(n4855), .A3(n6098), .A4(n6097), .ZN(n6104)
         );
  NAND3_X1 U6029 ( .A1(n5010), .A2(n5007), .A3(n8312), .ZN(n6616) );
  INV_X1 U6030 ( .A(n8694), .ZN(n5019) );
  NAND2_X1 U6031 ( .A1(n8532), .A2(n8533), .ZN(n8657) );
  OAI21_X1 U6032 ( .B1(n8370), .B2(n8369), .A(n8575), .ZN(n8390) );
  INV_X1 U6033 ( .A(n8391), .ZN(n8392) );
  NAND3_X1 U6034 ( .A1(n7567), .A2(n7749), .A3(n5028), .ZN(n5027) );
  INV_X1 U6035 ( .A(n8537), .ZN(n5037) );
  OAI21_X1 U6036 ( .B1(n9294), .B2(n5041), .A(n5038), .ZN(n9238) );
  NAND2_X1 U6037 ( .A1(n5042), .A2(n5043), .ZN(n8500) );
  OR2_X1 U6038 ( .A1(n9155), .A2(n9154), .ZN(n9158) );
  NAND3_X1 U6039 ( .A1(n5153), .A2(n5048), .A3(n5154), .ZN(n6013) );
  NAND4_X1 U6040 ( .A1(n5153), .A2(n5048), .A3(n5154), .A4(n5050), .ZN(n6017)
         );
  INV_X1 U6041 ( .A(n5341), .ZN(n5051) );
  NAND3_X1 U6042 ( .A1(n5153), .A2(n5154), .A3(n5049), .ZN(n5052) );
  INV_X1 U6043 ( .A(n5052), .ZN(n5360) );
  NAND2_X1 U6044 ( .A1(n6405), .A2(n4858), .ZN(n5056) );
  NAND3_X1 U6045 ( .A1(n4847), .A2(n4848), .A3(n6895), .ZN(n5055) );
  NAND2_X2 U6046 ( .A1(n6405), .A2(n6780), .ZN(n6532) );
  INV_X1 U6047 ( .A(n5061), .ZN(n9833) );
  NOR2_X1 U6048 ( .A1(n9796), .A2(n9908), .ZN(n9765) );
  NAND3_X1 U6049 ( .A1(n5208), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5066) );
  INV_X1 U6050 ( .A(n5517), .ZN(n5073) );
  NAND2_X1 U6051 ( .A1(n5497), .A2(n5496), .ZN(n5074) );
  NAND2_X1 U6052 ( .A1(n5070), .A2(n5068), .ZN(n5531) );
  AOI21_X1 U6053 ( .B1(n5517), .B2(n5069), .A(n4911), .ZN(n5068) );
  NAND2_X1 U6054 ( .A1(n5497), .A2(n5071), .ZN(n5070) );
  NOR2_X1 U6055 ( .A1(n5073), .A2(n5072), .ZN(n5071) );
  NAND2_X1 U6056 ( .A1(n5658), .A2(n5082), .ZN(n5080) );
  OAI21_X1 U6057 ( .B1(n5756), .B2(n5755), .A(n5757), .ZN(n5778) );
  NAND2_X1 U6058 ( .A1(n7135), .A2(n7161), .ZN(n7278) );
  NAND2_X1 U6059 ( .A1(n9802), .A2(n9812), .ZN(n9796) );
  NAND2_X1 U6060 ( .A1(n5992), .A2(n5991), .ZN(n5994) );
  NAND2_X1 U6061 ( .A1(n6405), .A2(n6778), .ZN(n6383) );
  NAND2_X1 U6062 ( .A1(n9829), .A2(n5131), .ZN(n5130) );
  NAND4_X1 U6063 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n5312), .ZN(n6726)
         );
  NAND2_X1 U6064 ( .A1(n7860), .A2(n7861), .ZN(n8040) );
  INV_X1 U6065 ( .A(n8655), .ZN(n7395) );
  NAND2_X1 U6066 ( .A1(n7389), .A2(n8655), .ZN(n7565) );
  AND2_X2 U6067 ( .A1(n8528), .A2(n8527), .ZN(n8655) );
  NAND3_X1 U6068 ( .A1(n9407), .A2(n5141), .A3(n5140), .ZN(n9484) );
  OAI21_X1 U6069 ( .B1(n9158), .B2(n5152), .A(n5149), .ZN(n8887) );
  NOR2_X1 U6070 ( .A1(n5401), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5515) );
  INV_X1 U6071 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6072 ( .A1(n10481), .A2(n10470), .ZN(n10469) );
  INV_X1 U6073 ( .A(n5161), .ZN(n9321) );
  INV_X1 U6074 ( .A(n7773), .ZN(n7713) );
  NAND2_X1 U6075 ( .A1(n9176), .A2(n8748), .ZN(n9178) );
  OAI21_X2 U6076 ( .B1(n5629), .B2(n5180), .A(n5178), .ZN(n8217) );
  NAND2_X1 U6077 ( .A1(n5779), .A2(n5195), .ZN(n5194) );
  NAND2_X1 U6078 ( .A1(n7743), .A2(n9102), .ZN(n5472) );
  XNOR2_X1 U6079 ( .A(n5922), .B(n5920), .ZN(n9028) );
  NAND2_X1 U6080 ( .A1(n5638), .A2(n5204), .ZN(n5758) );
  NAND2_X1 U6081 ( .A1(n5555), .A2(n4853), .ZN(n5214) );
  NAND2_X1 U6082 ( .A1(n5555), .A2(n5554), .ZN(n5600) );
  NAND2_X1 U6083 ( .A1(n8441), .A2(n4910), .ZN(n5220) );
  INV_X1 U6084 ( .A(n9825), .ZN(n5228) );
  NAND2_X1 U6085 ( .A1(n5225), .A2(n5226), .ZN(n8734) );
  NAND2_X1 U6086 ( .A1(n9825), .A2(n5231), .ZN(n5225) );
  INV_X1 U6087 ( .A(n9764), .ZN(n5242) );
  NAND2_X1 U6088 ( .A1(n9182), .A2(n5253), .ZN(n5248) );
  OAI22_X2 U6089 ( .A1(n9182), .A2(n5247), .B1(n5249), .B2(n5246), .ZN(n8877)
         );
  OR2_X1 U6090 ( .A1(n9410), .A2(n9084), .ZN(n5255) );
  NAND2_X1 U6091 ( .A1(n5258), .A2(n4860), .ZN(n7974) );
  NAND3_X2 U6092 ( .A1(n5439), .A2(n5437), .A3(n5266), .ZN(n9103) );
  NAND2_X1 U6093 ( .A1(n8381), .A2(n5272), .ZN(n8398) );
  NAND3_X1 U6094 ( .A1(n5459), .A2(n5329), .A3(n5330), .ZN(n5376) );
  NAND2_X1 U6095 ( .A1(n8771), .A2(n5277), .ZN(n5273) );
  NAND2_X1 U6096 ( .A1(n9519), .A2(n5282), .ZN(n5281) );
  NAND2_X1 U6097 ( .A1(n8795), .A2(n4862), .ZN(n5289) );
  NAND2_X1 U6098 ( .A1(n5289), .A2(n5291), .ZN(n8908) );
  NAND2_X1 U6099 ( .A1(n8795), .A2(n8796), .ZN(n9614) );
  OR2_X1 U6100 ( .A1(n8795), .A2(n8796), .ZN(n9615) );
  INV_X1 U6101 ( .A(n9617), .ZN(n5296) );
  NAND2_X1 U6102 ( .A1(n8913), .A2(n5299), .ZN(n5298) );
  NAND2_X1 U6103 ( .A1(n5304), .A2(n7029), .ZN(n8695) );
  NAND2_X1 U6104 ( .A1(n8935), .A2(n5310), .ZN(n9513) );
  NAND2_X1 U6105 ( .A1(n8935), .A2(n8934), .ZN(n9510) );
  NAND2_X1 U6106 ( .A1(n9513), .A2(n8946), .ZN(n8954) );
  NAND3_X1 U6107 ( .A1(n6099), .A2(n6098), .A3(n6097), .ZN(n6719) );
  AND2_X1 U6108 ( .A1(n6101), .A2(n5314), .ZN(n6111) );
  NAND2_X1 U6109 ( .A1(n6101), .A2(n4861), .ZN(n9991) );
  INV_X1 U6110 ( .A(n9103), .ZN(n7390) );
  NAND2_X1 U6111 ( .A1(n6553), .A2(n7342), .ZN(n7341) );
  NAND2_X1 U6112 ( .A1(n6363), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U6113 ( .A1(n8728), .A2(n9869), .ZN(n8730) );
  AOI21_X1 U6114 ( .B1(n8508), .B2(n8677), .A(n8513), .ZN(n8509) );
  OR2_X1 U6115 ( .A1(n9409), .A2(n10564), .ZN(n9415) );
  XNOR2_X1 U6116 ( .A(n6666), .B(n6667), .ZN(n7018) );
  OAI211_X1 U6117 ( .C1(n9400), .C2(n10568), .A(n9403), .B(n9399), .ZN(n9482)
         );
  NAND2_X1 U6118 ( .A1(n7809), .A2(n7808), .ZN(n7871) );
  INV_X1 U6119 ( .A(n7132), .ZN(n7134) );
  INV_X1 U6120 ( .A(n7041), .ZN(n7063) );
  OR2_X1 U6121 ( .A1(n4846), .A2(n6754), .ZN(n5437) );
  NAND2_X1 U6122 ( .A1(n7128), .A2(n7127), .ZN(n7340) );
  NOR2_X1 U6123 ( .A1(n7129), .A2(n7354), .ZN(n7131) );
  NAND4_X4 U6124 ( .A1(n6393), .A2(n6392), .A3(n6391), .A4(n6390), .ZN(n7092)
         );
  OAI222_X1 U6125 ( .A1(n7477), .A2(n8875), .B1(P2_U3152), .B2(n8874), .C1(
        n8873), .C2(n9503), .ZN(P2_U3328) );
  INV_X1 U6126 ( .A(n8874), .ZN(n5348) );
  OAI22_X2 U6127 ( .A1(n9554), .A2(n8930), .B1(n8929), .B2(n8928), .ZN(n9631)
         );
  AND2_X1 U6128 ( .A1(n6418), .A2(n6084), .ZN(n5315) );
  OR2_X1 U6129 ( .A1(n8903), .A2(n8902), .ZN(n5316) );
  INV_X1 U6130 ( .A(n9249), .ZN(n9255) );
  AND2_X1 U6131 ( .A1(n7434), .A2(n7433), .ZN(n5318) );
  NOR2_X1 U6132 ( .A1(n9467), .A2(n9315), .ZN(n5320) );
  INV_X1 U6133 ( .A(n8444), .ZN(n8440) );
  CLKBUF_X3 U6134 ( .A(n6525), .Z(n6499) );
  AND2_X1 U6135 ( .A1(n6062), .A2(n7398), .ZN(n9388) );
  INV_X1 U6136 ( .A(n9388), .ZN(n9343) );
  INV_X1 U6137 ( .A(n7018), .ZN(n6668) );
  OR2_X1 U6138 ( .A1(n6405), .A2(n6371), .ZN(n5322) );
  NOR2_X1 U6139 ( .A1(n5389), .A2(n5418), .ZN(n5323) );
  AND2_X1 U6140 ( .A1(n9545), .A2(n9543), .ZN(n5324) );
  AND2_X1 U6141 ( .A1(n6064), .A2(n6063), .ZN(n5325) );
  AND2_X1 U6142 ( .A1(n5682), .A2(n5663), .ZN(n5326) );
  INV_X1 U6143 ( .A(n9765), .ZN(n9777) );
  OR2_X1 U6144 ( .A1(n6751), .A2(n6787), .ZN(n5327) );
  INV_X1 U6145 ( .A(n9195), .ZN(n8748) );
  NAND2_X1 U6146 ( .A1(n5946), .A2(n5945), .ZN(n9067) );
  OAI21_X1 U6147 ( .B1(n7871), .B2(n7870), .A(n7869), .ZN(n8046) );
  INV_X1 U6148 ( .A(n7816), .ZN(n7814) );
  NAND2_X1 U6149 ( .A1(n8064), .A2(n8067), .ZN(n8068) );
  INV_X1 U6150 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6371) );
  OR2_X1 U6151 ( .A1(n5852), .A2(n5851), .ZN(n5872) );
  AND2_X1 U6152 ( .A1(n9330), .A2(n8476), .ZN(n8473) );
  INV_X1 U6153 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5579) );
  AND2_X1 U6154 ( .A1(n8069), .A2(n8068), .ZN(n8073) );
  INV_X1 U6155 ( .A(n5613), .ZN(n5611) );
  NOR2_X1 U6156 ( .A1(n5482), .A2(n7370), .ZN(n5483) );
  INV_X1 U6157 ( .A(n5958), .ZN(n5956) );
  INV_X1 U6158 ( .A(n5691), .ZN(n5690) );
  INV_X1 U6159 ( .A(n9327), .ZN(n9339) );
  INV_X1 U6160 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5330) );
  OR2_X1 U6161 ( .A1(n8910), .A2(n8909), .ZN(n8911) );
  INV_X1 U6162 ( .A(n6484), .ZN(n6482) );
  INV_X1 U6163 ( .A(n8188), .ZN(n8189) );
  INV_X1 U6164 ( .A(n6258), .ZN(n6145) );
  INV_X1 U6165 ( .A(n6175), .ZN(n6174) );
  INV_X1 U6166 ( .A(n6209), .ZN(n6147) );
  OR2_X1 U6167 ( .A1(n6509), .A2(n6495), .ZN(n6521) );
  INV_X1 U6168 ( .A(n6162), .ZN(n6148) );
  AND2_X1 U6169 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  INV_X1 U6170 ( .A(n5703), .ZN(n5705) );
  OR2_X1 U6171 ( .A1(n5668), .A2(n5667), .ZN(n5691) );
  INV_X1 U6172 ( .A(n9405), .ZN(n8881) );
  OR2_X1 U6173 ( .A1(n5586), .A2(n10185), .ZN(n5613) );
  INV_X1 U6174 ( .A(n6751), .ZN(n6768) );
  NAND2_X1 U6175 ( .A1(n7758), .A2(n7703), .ZN(n7773) );
  NAND2_X1 U6176 ( .A1(n6146), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6218) );
  INV_X1 U6177 ( .A(n6411), .ZN(n6139) );
  NAND2_X1 U6178 ( .A1(n6145), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6244) );
  OR2_X1 U6179 ( .A1(n6472), .A2(n9591), .ZN(n6484) );
  NAND2_X1 U6180 ( .A1(n6147), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6194) );
  INV_X1 U6181 ( .A(n9901), .ZN(n8703) );
  NAND2_X1 U6182 ( .A1(n6148), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U6183 ( .A1(n7656), .A2(n7534), .ZN(n7536) );
  NAND2_X1 U6184 ( .A1(n8295), .A2(n8296), .ZN(n8314) );
  INV_X1 U6185 ( .A(n7508), .ZN(n7296) );
  NAND2_X1 U6186 ( .A1(n6531), .A2(n6530), .ZN(n6078) );
  INV_X1 U6187 ( .A(n5973), .ZN(n5974) );
  INV_X1 U6188 ( .A(n5774), .ZN(n5777) );
  NAND2_X1 U6189 ( .A1(n5661), .A2(n5660), .ZN(n5682) );
  OR2_X1 U6190 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  NAND2_X1 U6191 ( .A1(n9085), .A2(n9039), .ZN(n6063) );
  AND3_X1 U6192 ( .A1(n5856), .A2(n5855), .A3(n5854), .ZN(n9043) );
  NAND2_X2 U6193 ( .A1(n5348), .A2(n5347), .ZN(n5450) );
  NOR2_X1 U6194 ( .A1(n8881), .A2(n8860), .ZN(n8882) );
  AND3_X1 U6195 ( .A1(n5877), .A2(n5876), .A3(n5875), .ZN(n9257) );
  INV_X1 U6196 ( .A(n8668), .ZN(n8369) );
  INV_X1 U6197 ( .A(n9390), .ZN(n9341) );
  INV_X2 U6198 ( .A(n7096), .ZN(n8943) );
  NAND2_X1 U6199 ( .A1(n8191), .A2(n8190), .ZN(n8234) );
  INV_X1 U6200 ( .A(n6426), .ZN(n6140) );
  OR2_X1 U6201 ( .A1(n9767), .A2(n6535), .ZN(n6491) );
  AND2_X1 U6202 ( .A1(n7213), .A2(n7212), .ZN(n7224) );
  INV_X1 U6203 ( .A(n9819), .ZN(n9781) );
  INV_X1 U6204 ( .A(n9827), .ZN(n10442) );
  INV_X1 U6205 ( .A(n9959), .ZN(n10537) );
  AND4_X1 U6206 ( .A1(n5721), .A2(n5720), .A3(n5719), .A4(n5718), .ZN(n8477)
         );
  INV_X1 U6207 ( .A(n8886), .ZN(n8878) );
  INV_X1 U6208 ( .A(n8848), .ZN(n9312) );
  OR2_X1 U6209 ( .A1(n9280), .A2(n9368), .ZN(n9357) );
  INV_X1 U6210 ( .A(n9393), .ZN(n9373) );
  INV_X1 U6211 ( .A(n6724), .ZN(n6725) );
  AND2_X1 U6212 ( .A1(n6528), .A2(n6527), .ZN(n9745) );
  AND2_X1 U6213 ( .A1(n6619), .A2(n8313), .ZN(n8296) );
  NAND2_X1 U6214 ( .A1(n7300), .A2(n7304), .ZN(n7531) );
  OR3_X1 U6215 ( .A1(n7293), .A2(n7153), .A3(n7152), .ZN(n7181) );
  XNOR2_X1 U6216 ( .A(n5519), .B(n10161), .ZN(n5517) );
  OR3_X1 U6217 ( .A1(n6052), .A2(n7398), .A3(n10575), .ZN(n9081) );
  INV_X1 U6218 ( .A(n9477), .ZN(n9385) );
  INV_X1 U6219 ( .A(n10584), .ZN(n10583) );
  OR2_X1 U6220 ( .A1(n9471), .A2(n9470), .ZN(n9498) );
  INV_X1 U6221 ( .A(n10588), .ZN(n10585) );
  INV_X1 U6222 ( .A(n9891), .ZN(n9741) );
  INV_X1 U6223 ( .A(n9916), .ZN(n9816) );
  INV_X1 U6224 ( .A(n9734), .ZN(n9873) );
  OR2_X1 U6225 ( .A1(n7181), .A2(n7180), .ZN(n10542) );
  OAI21_X1 U6226 ( .B1(n9890), .B2(n10494), .A(n9889), .ZN(n9973) );
  OR2_X1 U6227 ( .A1(n7181), .A2(n9990), .ZN(n10543) );
  NOR2_X1 U6228 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5336) );
  NOR2_X1 U6229 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5335) );
  NOR2_X1 U6230 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5334) );
  NOR2_X1 U6231 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5333) );
  NAND4_X1 U6232 ( .A1(n5336), .A2(n5335), .A3(n5334), .A4(n5333), .ZN(n5339)
         );
  NOR2_X1 U6233 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5337) );
  NAND4_X1 U6234 ( .A1(n5337), .A2(n5684), .A3(n5582), .A4(n5579), .ZN(n5338)
         );
  NOR3_X1 U6235 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5341) );
  INV_X1 U6236 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5342) );
  INV_X1 U6237 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6238 ( .A1(n5367), .A2(n5368), .ZN(n5345) );
  INV_X1 U6239 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5343) );
  INV_X1 U6240 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9502) );
  XNOR2_X2 U6241 ( .A(n5344), .B(n9502), .ZN(n8874) );
  NAND2_X1 U6242 ( .A1(n5345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6243 ( .A1(n8496), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5352) );
  AND2_X2 U6244 ( .A1(n8874), .A2(n5347), .ZN(n5436) );
  INV_X1 U6245 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6945) );
  XNOR2_X1 U6246 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7776) );
  OR2_X1 U6247 ( .A1(n5450), .A2(n7776), .ZN(n5350) );
  INV_X1 U6248 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6952) );
  OR2_X1 U6249 ( .A1(n4846), .A2(n6952), .ZN(n5349) );
  INV_X1 U6250 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5353) );
  NAND3_X1 U6251 ( .A1(n5582), .A2(n5579), .A3(n5353), .ZN(n5354) );
  INV_X1 U6252 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5355) );
  INV_X1 U6253 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5707) );
  INV_X1 U6254 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5710) );
  AND3_X1 U6255 ( .A1(n5684), .A2(n5707), .A3(n5710), .ZN(n5356) );
  INV_X1 U6256 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5357) );
  INV_X1 U6257 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5363) );
  INV_X1 U6258 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6259 ( .A1(n5052), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6008) );
  XNOR2_X1 U6260 ( .A(n6008), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8691) );
  INV_X1 U6261 ( .A(n8691), .ZN(n7897) );
  NAND2_X1 U6262 ( .A1(n5361), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5362) );
  XNOR2_X1 U6263 ( .A(n5362), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8521) );
  INV_X1 U6264 ( .A(n8521), .ZN(n8680) );
  OR2_X1 U6265 ( .A1(n7750), .A2(n4844), .ZN(n5481) );
  NAND2_X1 U6266 ( .A1(n5364), .A2(n8521), .ZN(n5366) );
  NAND2_X1 U6267 ( .A1(n9143), .A2(n8691), .ZN(n5365) );
  NAND2_X4 U6268 ( .A1(n5366), .A2(n5365), .ZN(n7400) );
  NAND2_X1 U6269 ( .A1(n6017), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5370) );
  MUX2_X1 U6270 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5370), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5372) );
  NOR2_X1 U6271 ( .A1(n5373), .A2(n5343), .ZN(n5374) );
  MUX2_X1 U6272 ( .A(n5343), .B(n5374), .S(P2_IR_REG_4__SCAN_IN), .Z(n5375) );
  INV_X1 U6273 ( .A(n5375), .ZN(n5377) );
  NAND2_X1 U6274 ( .A1(n5377), .A2(n5376), .ZN(n6953) );
  AND2_X1 U6275 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5379) );
  MUX2_X1 U6276 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5385), .Z(n5443) );
  NAND2_X1 U6277 ( .A1(n5444), .A2(n5443), .ZN(n5382) );
  NAND2_X1 U6278 ( .A1(n5380), .A2(SI_1_), .ZN(n5381) );
  NAND2_X1 U6279 ( .A1(n5382), .A2(n5381), .ZN(n5465) );
  MUX2_X1 U6280 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5385), .Z(n5384) );
  INV_X1 U6281 ( .A(SI_2_), .ZN(n5383) );
  XNOR2_X1 U6282 ( .A(n5384), .B(n5383), .ZN(n5466) );
  NAND2_X1 U6283 ( .A1(n5465), .A2(n5466), .ZN(n5417) );
  NAND2_X1 U6284 ( .A1(n5384), .A2(SI_2_), .ZN(n5416) );
  INV_X1 U6285 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6779) );
  INV_X1 U6286 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6804) );
  MUX2_X1 U6287 ( .A(n6779), .B(n6804), .S(n5385), .Z(n5388) );
  INV_X1 U6288 ( .A(n5388), .ZN(n5386) );
  NAND2_X1 U6289 ( .A1(n5386), .A2(SI_3_), .ZN(n5387) );
  AND2_X1 U6290 ( .A1(n5416), .A2(n5387), .ZN(n5390) );
  INV_X1 U6291 ( .A(n5387), .ZN(n5389) );
  XNOR2_X1 U6292 ( .A(n5388), .B(SI_3_), .ZN(n5418) );
  MUX2_X1 U6293 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6778), .Z(n5405) );
  INV_X1 U6294 ( .A(SI_4_), .ZN(n10166) );
  XNOR2_X1 U6295 ( .A(n5404), .B(n5403), .ZN(n6808) );
  OR2_X1 U6296 ( .A1(n5520), .A2(n6808), .ZN(n5392) );
  INV_X1 U6297 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6794) );
  OR2_X1 U6298 ( .A1(n8503), .A2(n6794), .ZN(n5391) );
  OAI211_X1 U6299 ( .C1(n6751), .C2(n6953), .A(n5392), .B(n5391), .ZN(n7778)
         );
  XNOR2_X1 U6300 ( .A(n7400), .B(n7778), .ZN(n5479) );
  XNOR2_X1 U6301 ( .A(n5481), .B(n5479), .ZN(n7449) );
  NAND2_X1 U6302 ( .A1(n8496), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5399) );
  INV_X1 U6303 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6946) );
  OR2_X1 U6304 ( .A1(n5826), .A2(n6946), .ZN(n5398) );
  NAND3_X1 U6305 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5489) );
  INV_X1 U6306 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6307 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5393) );
  NAND2_X1 U6308 ( .A1(n5394), .A2(n5393), .ZN(n5395) );
  NAND2_X1 U6309 ( .A1(n5489), .A2(n5395), .ZN(n7714) );
  OR2_X1 U6310 ( .A1(n5450), .A2(n7714), .ZN(n5397) );
  OR2_X1 U6311 ( .A1(n4846), .A2(n7721), .ZN(n5396) );
  NAND2_X1 U6312 ( .A1(n5376), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5400) );
  MUX2_X1 U6313 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5400), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5402) );
  NAND2_X1 U6314 ( .A1(n5402), .A2(n5401), .ZN(n6968) );
  NAND2_X1 U6315 ( .A1(n5404), .A2(n5403), .ZN(n5407) );
  NAND2_X1 U6316 ( .A1(n5405), .A2(SI_4_), .ZN(n5406) );
  NAND2_X1 U6317 ( .A1(n5407), .A2(n5406), .ZN(n5497) );
  MUX2_X1 U6318 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6781), .Z(n5498) );
  INV_X1 U6319 ( .A(SI_5_), .ZN(n10163) );
  XNOR2_X1 U6320 ( .A(n5497), .B(n5496), .ZN(n6789) );
  OR2_X1 U6321 ( .A1(n5520), .A2(n6789), .ZN(n5409) );
  INV_X1 U6322 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6790) );
  XNOR2_X1 U6323 ( .A(n7400), .B(n7718), .ZN(n5485) );
  XNOR2_X1 U6324 ( .A(n5487), .B(n5485), .ZN(n7372) );
  AND2_X1 U6325 ( .A1(n7449), .A2(n7372), .ZN(n5422) );
  NAND2_X1 U6326 ( .A1(n5436), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5414) );
  OR2_X1 U6327 ( .A1(n5450), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5413) );
  INV_X1 U6328 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7761) );
  OR2_X1 U6329 ( .A1(n4846), .A2(n7761), .ZN(n5412) );
  INV_X1 U6330 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5410) );
  OR2_X1 U6331 ( .A1(n5454), .A2(n5410), .ZN(n5411) );
  NOR2_X1 U6332 ( .A1(n7578), .A2(n4844), .ZN(n5474) );
  INV_X1 U6333 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6334 ( .A1(n5461), .A2(n5459), .ZN(n5463) );
  NAND2_X1 U6335 ( .A1(n5463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5415) );
  XNOR2_X1 U6336 ( .A(n5415), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6926) );
  INV_X1 U6337 ( .A(n6926), .ZN(n6934) );
  NAND2_X1 U6338 ( .A1(n5417), .A2(n5416), .ZN(n5419) );
  XNOR2_X1 U6339 ( .A(n5419), .B(n5418), .ZN(n6805) );
  OR2_X1 U6340 ( .A1(n5520), .A2(n6805), .ZN(n5421) );
  OR2_X1 U6341 ( .A1(n8503), .A2(n6779), .ZN(n5420) );
  XNOR2_X1 U6342 ( .A(n7400), .B(n10488), .ZN(n5475) );
  NAND2_X1 U6343 ( .A1(n5474), .A2(n5475), .ZN(n7373) );
  AND2_X1 U6344 ( .A1(n5422), .A2(n7373), .ZN(n5484) );
  NAND2_X1 U6345 ( .A1(n5436), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5429) );
  INV_X1 U6346 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5423) );
  OR2_X1 U6347 ( .A1(n5454), .A2(n5423), .ZN(n5428) );
  INV_X1 U6348 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5424) );
  OR2_X1 U6349 ( .A1(n4846), .A2(n5424), .ZN(n5427) );
  INV_X1 U6350 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5425) );
  NAND4_X2 U6351 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n9105)
         );
  NAND2_X1 U6352 ( .A1(n6780), .A2(SI_0_), .ZN(n5431) );
  INV_X1 U6353 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6354 ( .A1(n5431), .A2(n5430), .ZN(n5433) );
  AND2_X1 U6355 ( .A1(n5433), .A2(n5432), .ZN(n9509) );
  MUX2_X1 U6356 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9509), .S(n6751), .Z(n7745) );
  NAND2_X1 U6357 ( .A1(n7391), .A2(n7743), .ZN(n7261) );
  OR2_X1 U6358 ( .A1(n7745), .A2(n7400), .ZN(n5434) );
  AND2_X1 U6359 ( .A1(n7261), .A2(n5434), .ZN(n7238) );
  INV_X1 U6360 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6754) );
  INV_X1 U6361 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5435) );
  INV_X1 U6362 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5438) );
  OR2_X1 U6363 ( .A1(n5450), .A2(n5438), .ZN(n5439) );
  NAND2_X1 U6364 ( .A1(n9103), .A2(n7743), .ZN(n5448) );
  INV_X1 U6365 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6785) );
  INV_X1 U6366 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6367 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5440) );
  XNOR2_X1 U6368 ( .A(n5441), .B(n5440), .ZN(n6787) );
  XNOR2_X1 U6369 ( .A(n5444), .B(n5443), .ZN(n6786) );
  OR2_X1 U6370 ( .A1(n5520), .A2(n6786), .ZN(n5445) );
  XNOR2_X1 U6371 ( .A(n7400), .B(n7392), .ZN(n5447) );
  XNOR2_X1 U6372 ( .A(n5448), .B(n5447), .ZN(n7237) );
  NAND2_X1 U6373 ( .A1(n7238), .A2(n7237), .ZN(n7168) );
  INV_X1 U6374 ( .A(n5447), .ZN(n5449) );
  NAND2_X1 U6375 ( .A1(n5449), .A2(n5448), .ZN(n7169) );
  NAND2_X1 U6376 ( .A1(n7168), .A2(n7169), .ZN(n5469) );
  NAND2_X1 U6377 ( .A1(n5436), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5458) );
  INV_X1 U6378 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7767) );
  OR2_X1 U6379 ( .A1(n5450), .A2(n7767), .ZN(n5457) );
  INV_X1 U6380 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5451) );
  OR2_X1 U6381 ( .A1(n5452), .A2(n5451), .ZN(n5456) );
  INV_X1 U6382 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5453) );
  OR2_X1 U6383 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  INV_X1 U6384 ( .A(n5459), .ZN(n5460) );
  NAND2_X1 U6385 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5460), .ZN(n5462) );
  MUX2_X1 U6386 ( .A(n5462), .B(P2_IR_REG_31__SCAN_IN), .S(n5461), .Z(n5464)
         );
  INV_X1 U6387 ( .A(n10385), .ZN(n6784) );
  INV_X1 U6388 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6783) );
  OR2_X1 U6389 ( .A1(n8503), .A2(n6783), .ZN(n5468) );
  XNOR2_X1 U6390 ( .A(n5465), .B(n5466), .ZN(n6803) );
  OR2_X1 U6391 ( .A1(n5520), .A2(n6803), .ZN(n5467) );
  XNOR2_X1 U6392 ( .A(n7400), .B(n7769), .ZN(n5470) );
  INV_X1 U6393 ( .A(n5470), .ZN(n5471) );
  NAND2_X1 U6394 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  NAND2_X1 U6395 ( .A1(n7172), .A2(n5473), .ZN(n7335) );
  INV_X1 U6396 ( .A(n5474), .ZN(n5477) );
  INV_X1 U6397 ( .A(n5475), .ZN(n5476) );
  NAND2_X1 U6398 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  NAND2_X1 U6399 ( .A1(n7373), .A2(n5478), .ZN(n7334) );
  INV_X1 U6400 ( .A(n7372), .ZN(n5482) );
  INV_X1 U6401 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U6402 ( .A1(n5481), .A2(n5480), .ZN(n7370) );
  INV_X1 U6403 ( .A(n5485), .ZN(n5486) );
  NAND2_X1 U6404 ( .A1(n5487), .A2(n5486), .ZN(n7514) );
  NAND2_X1 U6405 ( .A1(n7375), .A2(n7514), .ZN(n5504) );
  NAND2_X1 U6406 ( .A1(n8496), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5495) );
  INV_X1 U6407 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6972) );
  OR2_X1 U6408 ( .A1(n5826), .A2(n6972), .ZN(n5494) );
  INV_X1 U6409 ( .A(n5489), .ZN(n5488) );
  NAND2_X1 U6410 ( .A1(n5488), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5509) );
  INV_X1 U6411 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10105) );
  NAND2_X1 U6412 ( .A1(n5489), .A2(n10105), .ZN(n5490) );
  NAND2_X1 U6413 ( .A1(n5509), .A2(n5490), .ZN(n7979) );
  OR2_X1 U6414 ( .A1(n5450), .A2(n7979), .ZN(n5493) );
  INV_X1 U6415 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5491) );
  OR2_X1 U6416 ( .A1(n4846), .A2(n5491), .ZN(n5492) );
  OR2_X1 U6417 ( .A1(n7933), .A2(n8511), .ZN(n5507) );
  NAND2_X1 U6418 ( .A1(n5498), .A2(SI_5_), .ZN(n5499) );
  MUX2_X1 U6419 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6781), .Z(n5519) );
  INV_X1 U6420 ( .A(SI_6_), .ZN(n10161) );
  XNOR2_X1 U6421 ( .A(n5518), .B(n5517), .ZN(n6792) );
  OR2_X1 U6422 ( .A1(n5520), .A2(n6792), .ZN(n5503) );
  INV_X1 U6423 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6793) );
  OR2_X1 U6424 ( .A1(n8503), .A2(n6793), .ZN(n5502) );
  NAND2_X1 U6425 ( .A1(n5401), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5500) );
  XNOR2_X1 U6426 ( .A(n5500), .B(n5155), .ZN(n6983) );
  OR2_X1 U6427 ( .A1(n6751), .A2(n6983), .ZN(n5501) );
  XNOR2_X1 U6428 ( .A(n5982), .B(n10504), .ZN(n5505) );
  XNOR2_X1 U6429 ( .A(n5507), .B(n5505), .ZN(n7513) );
  INV_X1 U6430 ( .A(n5505), .ZN(n5506) );
  NAND2_X1 U6431 ( .A1(n5507), .A2(n5506), .ZN(n5508) );
  NAND2_X1 U6432 ( .A1(n8496), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5514) );
  INV_X1 U6433 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6976) );
  OR2_X1 U6434 ( .A1(n5826), .A2(n6976), .ZN(n5513) );
  NAND2_X1 U6435 ( .A1(n5509), .A2(n6744), .ZN(n5510) );
  NAND2_X1 U6436 ( .A1(n5543), .A2(n5510), .ZN(n7936) );
  OR2_X1 U6437 ( .A1(n5450), .A2(n7936), .ZN(n5512) );
  INV_X1 U6438 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7937) );
  OR2_X1 U6439 ( .A1(n4846), .A2(n7937), .ZN(n5511) );
  NOR2_X1 U6440 ( .A1(n7973), .A2(n8511), .ZN(n5523) );
  OR2_X1 U6441 ( .A1(n5515), .A2(n5343), .ZN(n5516) );
  XNOR2_X1 U6442 ( .A(n5516), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7016) );
  INV_X1 U6443 ( .A(n7016), .ZN(n6975) );
  MUX2_X1 U6444 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6781), .Z(n5532) );
  XNOR2_X1 U6445 ( .A(n5531), .B(n5529), .ZN(n6809) );
  INV_X2 U6446 ( .A(n5520), .ZN(n5561) );
  NAND2_X1 U6447 ( .A1(n6809), .A2(n5561), .ZN(n5522) );
  INV_X1 U6448 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6810) );
  OR2_X1 U6449 ( .A1(n8503), .A2(n6810), .ZN(n5521) );
  OAI211_X1 U6450 ( .C1(n6751), .C2(n6975), .A(n5522), .B(n5521), .ZN(n7939)
         );
  XNOR2_X1 U6451 ( .A(n7939), .B(n7400), .ZN(n5524) );
  NAND2_X1 U6452 ( .A1(n5523), .A2(n5524), .ZN(n5528) );
  INV_X1 U6453 ( .A(n5523), .ZN(n5526) );
  INV_X1 U6454 ( .A(n5524), .ZN(n5525) );
  NAND2_X1 U6455 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  NAND2_X1 U6456 ( .A1(n5528), .A2(n5527), .ZN(n6743) );
  NAND2_X1 U6457 ( .A1(n5531), .A2(n5530), .ZN(n5534) );
  NAND2_X1 U6458 ( .A1(n5532), .A2(SI_7_), .ZN(n5533) );
  NAND2_X1 U6459 ( .A1(n5534), .A2(n5533), .ZN(n5553) );
  INV_X1 U6460 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6828) );
  INV_X1 U6461 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6815) );
  MUX2_X1 U6462 ( .A(n6828), .B(n6815), .S(n6781), .Z(n5535) );
  INV_X1 U6463 ( .A(SI_8_), .ZN(n10057) );
  INV_X1 U6464 ( .A(n5535), .ZN(n5536) );
  NAND2_X1 U6465 ( .A1(n5536), .A2(SI_8_), .ZN(n5537) );
  XNOR2_X1 U6466 ( .A(n5553), .B(n5552), .ZN(n6814) );
  NAND2_X1 U6467 ( .A1(n6814), .A2(n5561), .ZN(n5541) );
  NAND2_X1 U6468 ( .A1(n5538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5539) );
  XNOR2_X1 U6469 ( .A(n5539), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7004) );
  AOI22_X1 U6470 ( .A1(n5819), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6768), .B2(
        n7004), .ZN(n5540) );
  XNOR2_X1 U6471 ( .A(n10520), .B(n7400), .ZN(n5551) );
  NAND2_X1 U6472 ( .A1(n8496), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5548) );
  INV_X1 U6473 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6977) );
  INV_X1 U6474 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U6475 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  NAND2_X1 U6476 ( .A1(n5565), .A2(n5544), .ZN(n8822) );
  OR2_X1 U6477 ( .A1(n5450), .A2(n8822), .ZN(n5546) );
  INV_X1 U6478 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8823) );
  OR2_X1 U6479 ( .A1(n4846), .A2(n8823), .ZN(n5545) );
  NAND2_X1 U6480 ( .A1(n9096), .A2(n7743), .ZN(n5549) );
  XNOR2_X1 U6481 ( .A(n5551), .B(n5549), .ZN(n7730) );
  INV_X1 U6482 ( .A(n5549), .ZN(n5550) );
  NAND2_X1 U6483 ( .A1(n5551), .A2(n5550), .ZN(n7899) );
  INV_X1 U6484 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5556) );
  INV_X1 U6485 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6822) );
  MUX2_X1 U6486 ( .A(n5556), .B(n6822), .S(n6781), .Z(n5558) );
  INV_X1 U6487 ( .A(SI_9_), .ZN(n5557) );
  INV_X1 U6488 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U6489 ( .A1(n5559), .A2(SI_9_), .ZN(n5560) );
  XNOR2_X1 U6490 ( .A(n5600), .B(n5598), .ZN(n6820) );
  NAND2_X1 U6491 ( .A1(n6820), .A2(n5561), .ZN(n5564) );
  NAND2_X1 U6492 ( .A1(n5562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5580) );
  XNOR2_X1 U6493 ( .A(n5580), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7082) );
  AOI22_X1 U6494 ( .A1(n5819), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6768), .B2(
        n7082), .ZN(n5563) );
  XNOR2_X1 U6495 ( .A(n10527), .B(n5982), .ZN(n5595) );
  INV_X1 U6496 ( .A(n5595), .ZN(n5573) );
  NAND2_X1 U6497 ( .A1(n5436), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5571) );
  INV_X1 U6498 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7964) );
  OR2_X1 U6499 ( .A1(n4846), .A2(n7964), .ZN(n5570) );
  INV_X1 U6500 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U6501 ( .A1(n5565), .A2(n7902), .ZN(n5566) );
  NAND2_X1 U6502 ( .A1(n5586), .A2(n5566), .ZN(n7963) );
  OR2_X1 U6503 ( .A1(n5450), .A2(n7963), .ZN(n5569) );
  INV_X1 U6504 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5567) );
  OR2_X1 U6505 ( .A1(n5454), .A2(n5567), .ZN(n5568) );
  OR2_X1 U6506 ( .A1(n8128), .A2(n8511), .ZN(n5594) );
  INV_X1 U6507 ( .A(n5594), .ZN(n5572) );
  NAND2_X1 U6508 ( .A1(n5573), .A2(n5572), .ZN(n7910) );
  NAND2_X1 U6509 ( .A1(n5600), .A2(n5598), .ZN(n5574) );
  INV_X1 U6510 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6826) );
  INV_X1 U6511 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6831) );
  MUX2_X1 U6512 ( .A(n6826), .B(n6831), .S(n6781), .Z(n5576) );
  INV_X1 U6513 ( .A(SI_10_), .ZN(n5575) );
  NAND2_X1 U6514 ( .A1(n5576), .A2(n5575), .ZN(n5602) );
  INV_X1 U6515 ( .A(n5576), .ZN(n5577) );
  AND2_X1 U6516 ( .A1(n5602), .A2(n5601), .ZN(n5578) );
  NAND2_X1 U6517 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  NAND2_X1 U6518 ( .A1(n5581), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5583) );
  OR2_X1 U6519 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  NAND2_X1 U6520 ( .A1(n5583), .A2(n5582), .ZN(n5607) );
  AND2_X1 U6521 ( .A1(n5584), .A2(n5607), .ZN(n7197) );
  AOI22_X1 U6522 ( .A1(n5819), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6768), .B2(
        n7197), .ZN(n5585) );
  XNOR2_X1 U6523 ( .A(n8136), .B(n5982), .ZN(n5622) );
  INV_X1 U6524 ( .A(n5622), .ZN(n5592) );
  NAND2_X1 U6525 ( .A1(n8496), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5591) );
  INV_X1 U6526 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7083) );
  OR2_X1 U6527 ( .A1(n5826), .A2(n7083), .ZN(n5590) );
  INV_X1 U6528 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10185) );
  NAND2_X1 U6529 ( .A1(n5586), .A2(n10185), .ZN(n5587) );
  NAND2_X1 U6530 ( .A1(n5613), .A2(n5587), .ZN(n8129) );
  OR2_X1 U6531 ( .A1(n5450), .A2(n8129), .ZN(n5589) );
  INV_X1 U6532 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8130) );
  OR2_X1 U6533 ( .A1(n4846), .A2(n8130), .ZN(n5588) );
  NOR2_X1 U6534 ( .A1(n8106), .A2(n8511), .ZN(n5621) );
  NAND2_X1 U6535 ( .A1(n5592), .A2(n5621), .ZN(n5620) );
  AND2_X1 U6536 ( .A1(n7910), .A2(n5620), .ZN(n5593) );
  AND2_X1 U6537 ( .A1(n7899), .A2(n5593), .ZN(n5597) );
  INV_X1 U6538 ( .A(n5593), .ZN(n5596) );
  NAND2_X1 U6539 ( .A1(n5595), .A2(n5594), .ZN(n7908) );
  INV_X1 U6540 ( .A(n5601), .ZN(n5605) );
  MUX2_X1 U6541 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6781), .Z(n5631) );
  INV_X1 U6542 ( .A(SI_11_), .ZN(n10051) );
  XNOR2_X1 U6543 ( .A(n5632), .B(n5630), .ZN(n6833) );
  NAND2_X1 U6544 ( .A1(n6833), .A2(n5561), .ZN(n5610) );
  NAND2_X1 U6545 ( .A1(n5607), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5608) );
  XNOR2_X1 U6546 ( .A(n5608), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7364) );
  AOI22_X1 U6547 ( .A1(n5819), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6768), .B2(
        n7364), .ZN(n5609) );
  NAND2_X1 U6548 ( .A1(n5610), .A2(n5609), .ZN(n8338) );
  XNOR2_X1 U6549 ( .A(n8338), .B(n5982), .ZN(n5625) );
  NAND2_X1 U6550 ( .A1(n5436), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5619) );
  INV_X1 U6551 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8119) );
  OR2_X1 U6552 ( .A1(n4846), .A2(n8119), .ZN(n5618) );
  INV_X1 U6553 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U6554 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  NAND2_X1 U6555 ( .A1(n5643), .A2(n5614), .ZN(n8118) );
  OR2_X1 U6556 ( .A1(n5450), .A2(n8118), .ZN(n5617) );
  INV_X1 U6557 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5615) );
  OR2_X1 U6558 ( .A1(n5454), .A2(n5615), .ZN(n5616) );
  NOR2_X1 U6559 ( .A1(n8337), .A2(n8511), .ZN(n5626) );
  XNOR2_X1 U6560 ( .A(n5625), .B(n5626), .ZN(n7988) );
  INV_X1 U6561 ( .A(n5620), .ZN(n5623) );
  XNOR2_X1 U6562 ( .A(n5622), .B(n5621), .ZN(n7912) );
  OR2_X1 U6563 ( .A1(n5623), .A2(n7912), .ZN(n7986) );
  AND2_X1 U6564 ( .A1(n7988), .A2(n7986), .ZN(n5624) );
  NAND2_X1 U6565 ( .A1(n7987), .A2(n5624), .ZN(n5629) );
  INV_X1 U6566 ( .A(n5625), .ZN(n5627) );
  NAND2_X1 U6567 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  INV_X1 U6568 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6844) );
  INV_X1 U6569 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5633) );
  MUX2_X1 U6570 ( .A(n6844), .B(n5633), .S(n6781), .Z(n5635) );
  INV_X1 U6571 ( .A(SI_12_), .ZN(n5634) );
  INV_X1 U6572 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U6573 ( .A1(n5636), .A2(SI_12_), .ZN(n5637) );
  XNOR2_X1 U6574 ( .A(n5658), .B(n5657), .ZN(n6841) );
  NAND2_X1 U6575 ( .A1(n6841), .A2(n5561), .ZN(n5641) );
  OR2_X1 U6576 ( .A1(n5638), .A2(n5343), .ZN(n5639) );
  XNOR2_X1 U6577 ( .A(n5639), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7458) );
  AOI22_X1 U6578 ( .A1(n5819), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6768), .B2(
        n7458), .ZN(n5640) );
  NAND2_X1 U6579 ( .A1(n5641), .A2(n5640), .ZN(n8379) );
  XNOR2_X1 U6580 ( .A(n8379), .B(n5982), .ZN(n5650) );
  INV_X1 U6581 ( .A(n4846), .ZN(n5874) );
  NAND2_X1 U6582 ( .A1(n5874), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5649) );
  INV_X1 U6583 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7464) );
  OR2_X1 U6584 ( .A1(n5826), .A2(n7464), .ZN(n5648) );
  INV_X1 U6585 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10117) );
  NAND2_X1 U6586 ( .A1(n5643), .A2(n10117), .ZN(n5644) );
  NAND2_X1 U6587 ( .A1(n5668), .A2(n5644), .ZN(n8345) );
  OR2_X1 U6588 ( .A1(n5450), .A2(n8345), .ZN(n5647) );
  INV_X1 U6589 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5645) );
  OR2_X1 U6590 ( .A1(n5454), .A2(n5645), .ZN(n5646) );
  OR2_X1 U6591 ( .A1(n8372), .A2(n8511), .ZN(n5651) );
  NAND2_X1 U6592 ( .A1(n5650), .A2(n5651), .ZN(n5655) );
  INV_X1 U6593 ( .A(n5650), .ZN(n5653) );
  INV_X1 U6594 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U6595 ( .A1(n5653), .A2(n5652), .ZN(n5654) );
  NAND2_X1 U6596 ( .A1(n5655), .A2(n5654), .ZN(n8145) );
  INV_X1 U6597 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6924) );
  INV_X1 U6598 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5659) );
  MUX2_X1 U6599 ( .A(n6924), .B(n5659), .S(n6781), .Z(n5661) );
  INV_X1 U6600 ( .A(SI_13_), .ZN(n5660) );
  INV_X1 U6601 ( .A(n5661), .ZN(n5662) );
  NAND2_X1 U6602 ( .A1(n5662), .A2(SI_13_), .ZN(n5663) );
  XNOR2_X1 U6603 ( .A(n5681), .B(n5326), .ZN(n6920) );
  NAND2_X1 U6604 ( .A1(n6920), .A2(n5561), .ZN(n5666) );
  OR2_X1 U6605 ( .A1(n5664), .A2(n5343), .ZN(n5685) );
  XNOR2_X1 U6606 ( .A(n5685), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7618) );
  AOI22_X1 U6607 ( .A1(n5819), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6768), .B2(
        n7618), .ZN(n5665) );
  XNOR2_X1 U6608 ( .A(n8396), .B(n5982), .ZN(n5675) );
  NAND2_X1 U6609 ( .A1(n5874), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5674) );
  INV_X1 U6610 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7463) );
  OR2_X1 U6611 ( .A1(n5826), .A2(n7463), .ZN(n5673) );
  INV_X1 U6612 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U6613 ( .A1(n5668), .A2(n5667), .ZN(n5669) );
  NAND2_X1 U6614 ( .A1(n5691), .A2(n5669), .ZN(n8376) );
  OR2_X1 U6615 ( .A1(n5450), .A2(n8376), .ZN(n5672) );
  INV_X1 U6616 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n5670) );
  OR2_X1 U6617 ( .A1(n5454), .A2(n5670), .ZN(n5671) );
  OR2_X1 U6618 ( .A1(n8393), .A2(n8511), .ZN(n5676) );
  NAND2_X1 U6619 ( .A1(n5675), .A2(n5676), .ZN(n5680) );
  INV_X1 U6620 ( .A(n5675), .ZN(n5678) );
  INV_X1 U6621 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U6622 ( .A1(n5678), .A2(n5677), .ZN(n5679) );
  AND2_X1 U6623 ( .A1(n5680), .A2(n5679), .ZN(n8219) );
  NAND2_X1 U6624 ( .A1(n8217), .A2(n5680), .ZN(n8303) );
  MUX2_X1 U6625 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6781), .Z(n5704) );
  INV_X1 U6626 ( .A(SI_14_), .ZN(n10024) );
  NAND2_X1 U6627 ( .A1(n6939), .A2(n5561), .ZN(n5688) );
  NAND2_X1 U6628 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  NAND2_X1 U6629 ( .A1(n5686), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5708) );
  XNOR2_X1 U6630 ( .A(n5708), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7888) );
  AOI22_X1 U6631 ( .A1(n5819), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6768), .B2(
        n7888), .ZN(n5687) );
  XNOR2_X1 U6632 ( .A(n10574), .B(n5982), .ZN(n5697) );
  NAND2_X1 U6633 ( .A1(n8496), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5696) );
  INV_X1 U6634 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5689) );
  OR2_X1 U6635 ( .A1(n5826), .A2(n5689), .ZN(n5695) );
  INV_X1 U6636 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8402) );
  OR2_X1 U6637 ( .A1(n4846), .A2(n8402), .ZN(n5694) );
  INV_X1 U6638 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U6639 ( .A1(n5691), .A2(n10175), .ZN(n5692) );
  NAND2_X1 U6640 ( .A1(n5716), .A2(n5692), .ZN(n8401) );
  OR2_X1 U6641 ( .A1(n5450), .A2(n8401), .ZN(n5693) );
  OR2_X1 U6642 ( .A1(n8471), .A2(n8511), .ZN(n5698) );
  NAND2_X1 U6643 ( .A1(n5697), .A2(n5698), .ZN(n5702) );
  INV_X1 U6644 ( .A(n5697), .ZN(n5700) );
  INV_X1 U6645 ( .A(n5698), .ZN(n5699) );
  NAND2_X1 U6646 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  AND2_X1 U6647 ( .A1(n5702), .A2(n5701), .ZN(n8304) );
  NAND2_X1 U6648 ( .A1(n8303), .A2(n8304), .ZN(n8302) );
  NAND2_X1 U6649 ( .A1(n8302), .A2(n5702), .ZN(n8408) );
  MUX2_X1 U6650 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6781), .Z(n5731) );
  XNOR2_X1 U6651 ( .A(n5731), .B(SI_15_), .ZN(n5728) );
  NAND2_X1 U6652 ( .A1(n6237), .A2(n5561), .ZN(n5713) );
  NAND2_X1 U6653 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  NAND2_X1 U6654 ( .A1(n5709), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5711) );
  XNOR2_X1 U6655 ( .A(n5711), .B(n5710), .ZN(n8162) );
  INV_X1 U6656 ( .A(n8162), .ZN(n7893) );
  AOI22_X1 U6657 ( .A1(n5819), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6768), .B2(
        n7893), .ZN(n5712) );
  XNOR2_X1 U6658 ( .A(n9477), .B(n5982), .ZN(n5722) );
  NAND2_X1 U6659 ( .A1(n8496), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5721) );
  INV_X1 U6660 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7889) );
  OR2_X1 U6661 ( .A1(n5826), .A2(n7889), .ZN(n5720) );
  INV_X1 U6662 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5714) );
  OR2_X1 U6663 ( .A1(n4846), .A2(n5714), .ZN(n5719) );
  INV_X1 U6664 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U6665 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  NAND2_X1 U6666 ( .A1(n5742), .A2(n5717), .ZN(n8411) );
  OR2_X1 U6667 ( .A1(n5450), .A2(n8411), .ZN(n5718) );
  OR2_X1 U6668 ( .A1(n8477), .A2(n8511), .ZN(n5723) );
  NAND2_X1 U6669 ( .A1(n5722), .A2(n5723), .ZN(n5727) );
  INV_X1 U6670 ( .A(n5722), .ZN(n5725) );
  INV_X1 U6671 ( .A(n5723), .ZN(n5724) );
  NAND2_X1 U6672 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  AND2_X1 U6673 ( .A1(n5727), .A2(n5726), .ZN(n8409) );
  NAND2_X1 U6674 ( .A1(n8408), .A2(n8409), .ZN(n8407) );
  NAND2_X1 U6675 ( .A1(n8407), .A2(n5727), .ZN(n9007) );
  NAND2_X1 U6676 ( .A1(n5731), .A2(SI_15_), .ZN(n5732) );
  NAND2_X2 U6677 ( .A1(n5733), .A2(n5732), .ZN(n5756) );
  INV_X1 U6678 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7232) );
  INV_X1 U6679 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7233) );
  MUX2_X1 U6680 ( .A(n7232), .B(n7233), .S(n6781), .Z(n5734) );
  INV_X1 U6681 ( .A(SI_16_), .ZN(n10147) );
  NAND2_X1 U6682 ( .A1(n5734), .A2(n10147), .ZN(n5757) );
  INV_X1 U6683 ( .A(n5734), .ZN(n5735) );
  NAND2_X1 U6684 ( .A1(n5735), .A2(SI_16_), .ZN(n5736) );
  NAND2_X1 U6685 ( .A1(n5757), .A2(n5736), .ZN(n5755) );
  XNOR2_X1 U6686 ( .A(n5756), .B(n5755), .ZN(n7231) );
  NAND2_X1 U6687 ( .A1(n7231), .A2(n5561), .ZN(n5740) );
  NAND2_X1 U6688 ( .A1(n5737), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5738) );
  XNOR2_X1 U6689 ( .A(n5738), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9110) );
  AOI22_X1 U6690 ( .A1(n5819), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6768), .B2(
        n9110), .ZN(n5739) );
  XNOR2_X1 U6691 ( .A(n9474), .B(n5982), .ZN(n5749) );
  NAND2_X1 U6692 ( .A1(n5874), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5748) );
  INV_X1 U6693 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8156) );
  OR2_X1 U6694 ( .A1(n5826), .A2(n8156), .ZN(n5747) );
  INV_X1 U6695 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U6696 ( .A1(n5742), .A2(n10200), .ZN(n5743) );
  NAND2_X1 U6697 ( .A1(n5764), .A2(n5743), .ZN(n9361) );
  OR2_X1 U6698 ( .A1(n5450), .A2(n9361), .ZN(n5746) );
  INV_X1 U6699 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5744) );
  OR2_X1 U6700 ( .A1(n5454), .A2(n5744), .ZN(n5745) );
  OR2_X1 U6701 ( .A1(n9344), .A2(n8511), .ZN(n5750) );
  NAND2_X1 U6702 ( .A1(n5749), .A2(n5750), .ZN(n5754) );
  INV_X1 U6703 ( .A(n5749), .ZN(n5752) );
  INV_X1 U6704 ( .A(n5750), .ZN(n5751) );
  NAND2_X1 U6705 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  AND2_X1 U6706 ( .A1(n5754), .A2(n5753), .ZN(n9008) );
  MUX2_X1 U6707 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6781), .Z(n5775) );
  INV_X1 U6708 ( .A(SI_17_), .ZN(n10145) );
  XNOR2_X1 U6709 ( .A(n5775), .B(n10145), .ZN(n5774) );
  XNOR2_X1 U6710 ( .A(n5778), .B(n5774), .ZN(n7266) );
  NAND2_X1 U6711 ( .A1(n7266), .A2(n5561), .ZN(n5761) );
  NAND2_X1 U6712 ( .A1(n5758), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5759) );
  XNOR2_X1 U6713 ( .A(n5759), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9124) );
  AOI22_X1 U6714 ( .A1(n5819), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6768), .B2(
        n9124), .ZN(n5760) );
  NAND2_X2 U6715 ( .A1(n5761), .A2(n5760), .ZN(n9467) );
  XNOR2_X1 U6716 ( .A(n9467), .B(n7400), .ZN(n5772) );
  NAND2_X1 U6717 ( .A1(n8496), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5770) );
  INV_X1 U6718 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n5762) );
  OR2_X1 U6719 ( .A1(n5826), .A2(n5762), .ZN(n5769) );
  INV_X1 U6720 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U6721 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  NAND2_X1 U6722 ( .A1(n5782), .A2(n5765), .ZN(n9351) );
  OR2_X1 U6723 ( .A1(n5450), .A2(n9351), .ZN(n5768) );
  INV_X1 U6724 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n5766) );
  OR2_X1 U6725 ( .A1(n4846), .A2(n5766), .ZN(n5767) );
  NOR2_X1 U6726 ( .A1(n9063), .A2(n8511), .ZN(n5771) );
  XNOR2_X1 U6727 ( .A(n5772), .B(n5771), .ZN(n9017) );
  NAND2_X1 U6728 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  NAND2_X1 U6729 ( .A1(n5775), .A2(SI_17_), .ZN(n5776) );
  MUX2_X1 U6730 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6781), .Z(n5795) );
  XNOR2_X1 U6731 ( .A(n5795), .B(SI_18_), .ZN(n5793) );
  XNOR2_X1 U6732 ( .A(n5794), .B(n5793), .ZN(n7286) );
  NAND2_X1 U6733 ( .A1(n7286), .A2(n5561), .ZN(n5781) );
  XNOR2_X1 U6734 ( .A(n5779), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9122) );
  AOI22_X1 U6735 ( .A1(n5819), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6768), .B2(
        n9122), .ZN(n5780) );
  XNOR2_X1 U6736 ( .A(n9462), .B(n5982), .ZN(n5788) );
  NAND2_X1 U6737 ( .A1(n8496), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5787) );
  INV_X1 U6738 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9130) );
  OR2_X1 U6739 ( .A1(n5826), .A2(n9130), .ZN(n5786) );
  INV_X1 U6740 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9135) );
  OR2_X1 U6741 ( .A1(n4846), .A2(n9135), .ZN(n5785) );
  INV_X1 U6742 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10104) );
  NAND2_X1 U6743 ( .A1(n5782), .A2(n10104), .ZN(n5783) );
  NAND2_X1 U6744 ( .A1(n5822), .A2(n5783), .ZN(n9057) );
  OR2_X1 U6745 ( .A1(n5450), .A2(n9057), .ZN(n5784) );
  OR2_X1 U6746 ( .A1(n9342), .A2(n8511), .ZN(n5789) );
  NAND2_X1 U6747 ( .A1(n5788), .A2(n5789), .ZN(n8983) );
  INV_X1 U6748 ( .A(n5788), .ZN(n5791) );
  INV_X1 U6749 ( .A(n5789), .ZN(n5790) );
  NAND2_X1 U6750 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  NAND2_X1 U6751 ( .A1(n8983), .A2(n5792), .ZN(n9055) );
  AND2_X1 U6752 ( .A1(n5982), .A2(n7743), .ZN(n5808) );
  NAND2_X1 U6753 ( .A1(n5795), .A2(SI_18_), .ZN(n5796) );
  INV_X1 U6754 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7478) );
  INV_X1 U6755 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7479) );
  MUX2_X1 U6756 ( .A(n7478), .B(n7479), .S(n6781), .Z(n5798) );
  INV_X1 U6757 ( .A(SI_19_), .ZN(n10122) );
  NAND2_X1 U6758 ( .A1(n5798), .A2(n10122), .ZN(n5845) );
  INV_X1 U6759 ( .A(n5798), .ZN(n5799) );
  NAND2_X1 U6760 ( .A1(n5799), .A2(SI_19_), .ZN(n5800) );
  NAND2_X1 U6761 ( .A1(n5845), .A2(n5800), .ZN(n5817) );
  NAND2_X1 U6762 ( .A1(n5847), .A2(n5845), .ZN(n5805) );
  INV_X1 U6763 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7723) );
  INV_X1 U6764 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7611) );
  MUX2_X1 U6765 ( .A(n7723), .B(n7611), .S(n6781), .Z(n5802) );
  INV_X1 U6766 ( .A(SI_20_), .ZN(n5801) );
  NAND2_X1 U6767 ( .A1(n5802), .A2(n5801), .ZN(n5844) );
  INV_X1 U6768 ( .A(n5802), .ZN(n5803) );
  NAND2_X1 U6769 ( .A1(n5803), .A2(SI_20_), .ZN(n5848) );
  AND2_X1 U6770 ( .A1(n5844), .A2(n5848), .ZN(n5804) );
  NAND2_X1 U6771 ( .A1(n7610), .A2(n5561), .ZN(n5807) );
  OR2_X1 U6772 ( .A1(n8503), .A2(n7723), .ZN(n5806) );
  MUX2_X1 U6773 ( .A(n5808), .B(n7400), .S(n9452), .Z(n5814) );
  INV_X1 U6774 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10188) );
  INV_X1 U6775 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U6776 ( .A1(n5824), .A2(n10210), .ZN(n5809) );
  NAND2_X1 U6777 ( .A1(n5852), .A2(n5809), .ZN(n9040) );
  OR2_X1 U6778 ( .A1(n9040), .A2(n5450), .ZN(n5813) );
  NAND2_X1 U6779 ( .A1(n8496), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U6780 ( .A1(n5436), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U6781 ( .A1(n5874), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5810) );
  INV_X1 U6782 ( .A(n9256), .ZN(n9088) );
  NAND2_X1 U6783 ( .A1(n5814), .A2(n9088), .ZN(n5841) );
  INV_X1 U6784 ( .A(n5841), .ZN(n5833) );
  XNOR2_X1 U6785 ( .A(n9452), .B(n5982), .ZN(n5815) );
  OAI21_X1 U6786 ( .B1(n8511), .B2(n9256), .A(n5815), .ZN(n5816) );
  NAND2_X1 U6787 ( .A1(n5841), .A2(n5816), .ZN(n9037) );
  INV_X1 U6788 ( .A(n9037), .ZN(n5831) );
  XNOR2_X1 U6789 ( .A(n5818), .B(n5817), .ZN(n7476) );
  NAND2_X1 U6790 ( .A1(n7476), .A2(n5561), .ZN(n5821) );
  AOI22_X1 U6791 ( .A1(n5819), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6768), .B2(
        n9180), .ZN(n5820) );
  XNOR2_X1 U6792 ( .A(n9459), .B(n5982), .ZN(n5836) );
  NAND2_X1 U6793 ( .A1(n8496), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U6794 ( .A1(n5822), .A2(n10188), .ZN(n5823) );
  NAND2_X1 U6795 ( .A1(n5824), .A2(n5823), .ZN(n9290) );
  OR2_X1 U6796 ( .A1(n9290), .A2(n5450), .ZN(n5829) );
  INV_X1 U6797 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5825) );
  OR2_X1 U6798 ( .A1(n5826), .A2(n5825), .ZN(n5828) );
  INV_X1 U6799 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9291) );
  OR2_X1 U6800 ( .A1(n4846), .A2(n9291), .ZN(n5827) );
  OR2_X1 U6801 ( .A1(n9058), .A2(n8511), .ZN(n5837) );
  NAND2_X1 U6802 ( .A1(n5836), .A2(n5837), .ZN(n9035) );
  AND2_X1 U6803 ( .A1(n5831), .A2(n9035), .ZN(n5832) );
  AND2_X1 U6804 ( .A1(n8983), .A2(n5835), .ZN(n5834) );
  INV_X1 U6805 ( .A(n5835), .ZN(n5843) );
  INV_X1 U6806 ( .A(n5836), .ZN(n5839) );
  INV_X1 U6807 ( .A(n5837), .ZN(n5838) );
  NAND2_X1 U6808 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  AND2_X1 U6809 ( .A1(n9035), .A2(n5840), .ZN(n8985) );
  AND2_X1 U6810 ( .A1(n8985), .A2(n5841), .ZN(n5842) );
  MUX2_X1 U6811 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6781), .Z(n5863) );
  INV_X1 U6812 ( .A(SI_21_), .ZN(n10044) );
  XNOR2_X1 U6813 ( .A(n5863), .B(n10044), .ZN(n5862) );
  XNOR2_X1 U6814 ( .A(n5866), .B(n5862), .ZN(n7686) );
  NAND2_X1 U6815 ( .A1(n7686), .A2(n5561), .ZN(n5850) );
  INV_X1 U6816 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7689) );
  OR2_X1 U6817 ( .A1(n8503), .A2(n7689), .ZN(n5849) );
  XNOR2_X1 U6818 ( .A(n9447), .B(n7400), .ZN(n5859) );
  INV_X1 U6819 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U6820 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  NAND2_X1 U6821 ( .A1(n5872), .A2(n5853), .ZN(n8993) );
  OR2_X1 U6822 ( .A1(n8993), .A2(n5450), .ZN(n5856) );
  AOI22_X1 U6823 ( .A1(n5436), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n8496), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U6824 ( .A1(n5874), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5854) );
  INV_X1 U6825 ( .A(n9043), .ZN(n9275) );
  NAND2_X1 U6826 ( .A1(n9275), .A2(n7743), .ZN(n5857) );
  XNOR2_X1 U6827 ( .A(n5859), .B(n5857), .ZN(n8992) );
  NAND2_X1 U6828 ( .A1(n8991), .A2(n8992), .ZN(n5861) );
  INV_X1 U6829 ( .A(n5857), .ZN(n5858) );
  NAND2_X1 U6830 ( .A1(n5859), .A2(n5858), .ZN(n5860) );
  INV_X1 U6831 ( .A(n5862), .ZN(n5865) );
  NAND2_X1 U6832 ( .A1(n5863), .A2(SI_21_), .ZN(n5864) );
  INV_X1 U6833 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7898) );
  INV_X1 U6834 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6171) );
  MUX2_X1 U6835 ( .A(n7898), .B(n6171), .S(n6781), .Z(n5867) );
  INV_X1 U6836 ( .A(SI_22_), .ZN(n10137) );
  NAND2_X1 U6837 ( .A1(n5867), .A2(n10137), .ZN(n5883) );
  INV_X1 U6838 ( .A(n5867), .ZN(n5868) );
  NAND2_X1 U6839 ( .A1(n5868), .A2(SI_22_), .ZN(n5869) );
  NAND2_X1 U6840 ( .A1(n5883), .A2(n5869), .ZN(n5884) );
  XNOR2_X1 U6841 ( .A(n5885), .B(n5884), .ZN(n7896) );
  NAND2_X1 U6842 ( .A1(n7896), .A2(n5561), .ZN(n5871) );
  OR2_X1 U6843 ( .A1(n8503), .A2(n7898), .ZN(n5870) );
  XNOR2_X1 U6844 ( .A(n9442), .B(n5982), .ZN(n5878) );
  INV_X1 U6845 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10212) );
  NAND2_X1 U6846 ( .A1(n5872), .A2(n10212), .ZN(n5873) );
  AND2_X1 U6847 ( .A1(n5895), .A2(n5873), .ZN(n9241) );
  INV_X1 U6848 ( .A(n5450), .ZN(n6051) );
  NAND2_X1 U6849 ( .A1(n9241), .A2(n6051), .ZN(n5877) );
  AOI22_X1 U6850 ( .A1(n5436), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n8496), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U6851 ( .A1(n5874), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5875) );
  INV_X1 U6852 ( .A(n9257), .ZN(n9219) );
  NAND2_X1 U6853 ( .A1(n9219), .A2(n7743), .ZN(n5879) );
  NAND2_X1 U6854 ( .A1(n5878), .A2(n5879), .ZN(n8971) );
  INV_X1 U6855 ( .A(n5878), .ZN(n5881) );
  INV_X1 U6856 ( .A(n5879), .ZN(n5880) );
  NAND2_X1 U6857 ( .A1(n5881), .A2(n5880), .ZN(n5882) );
  NAND2_X1 U6858 ( .A1(n8971), .A2(n5882), .ZN(n9049) );
  INV_X1 U6859 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7920) );
  INV_X1 U6860 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7924) );
  MUX2_X1 U6861 ( .A(n7920), .B(n7924), .S(n6778), .Z(n5886) );
  INV_X1 U6862 ( .A(SI_23_), .ZN(n10131) );
  NAND2_X1 U6863 ( .A1(n5886), .A2(n10131), .ZN(n5907) );
  INV_X1 U6864 ( .A(n5886), .ZN(n5887) );
  NAND2_X1 U6865 ( .A1(n5887), .A2(SI_23_), .ZN(n5888) );
  AND2_X1 U6866 ( .A1(n5907), .A2(n5888), .ZN(n5889) );
  OR2_X1 U6867 ( .A1(n5890), .A2(n5889), .ZN(n5891) );
  NAND2_X1 U6868 ( .A1(n5908), .A2(n5891), .ZN(n7921) );
  NAND2_X1 U6869 ( .A1(n7921), .A2(n5561), .ZN(n5893) );
  OR2_X1 U6870 ( .A1(n8503), .A2(n7920), .ZN(n5892) );
  XNOR2_X1 U6871 ( .A(n9437), .B(n5982), .ZN(n8972) );
  INV_X1 U6872 ( .A(n8972), .ZN(n5904) );
  INV_X1 U6873 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6874 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  NAND2_X1 U6875 ( .A1(n5912), .A2(n5896), .ZN(n8976) );
  OR2_X1 U6876 ( .A1(n8976), .A2(n5450), .ZN(n5902) );
  INV_X1 U6877 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U6878 ( .A1(n5436), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U6879 ( .A1(n8496), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5897) );
  OAI211_X1 U6880 ( .C1(n5899), .C2(n4846), .A(n5898), .B(n5897), .ZN(n5900)
         );
  INV_X1 U6881 ( .A(n5900), .ZN(n5901) );
  INV_X1 U6882 ( .A(n8483), .ZN(n9209) );
  NAND2_X1 U6883 ( .A1(n9209), .A2(n7743), .ZN(n8974) );
  INV_X1 U6884 ( .A(n8974), .ZN(n5903) );
  INV_X1 U6885 ( .A(n8971), .ZN(n5905) );
  AOI21_X1 U6886 ( .B1(n8972), .B2(n8974), .A(n5905), .ZN(n5906) );
  MUX2_X1 U6887 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6778), .Z(n5926) );
  INV_X1 U6888 ( .A(SI_24_), .ZN(n10029) );
  XNOR2_X1 U6889 ( .A(n5926), .B(n10029), .ZN(n5925) );
  XNOR2_X1 U6890 ( .A(n5929), .B(n5925), .ZN(n8101) );
  NAND2_X1 U6891 ( .A1(n8101), .A2(n5561), .ZN(n5910) );
  INV_X1 U6892 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8102) );
  OR2_X1 U6893 ( .A1(n8503), .A2(n8102), .ZN(n5909) );
  XNOR2_X1 U6894 ( .A(n9431), .B(n5982), .ZN(n5920) );
  NAND2_X1 U6895 ( .A1(n5911), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5936) );
  INV_X1 U6896 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U6897 ( .A1(n5912), .A2(n10093), .ZN(n5913) );
  NAND2_X1 U6898 ( .A1(n5936), .A2(n5913), .ZN(n9029) );
  OR2_X1 U6899 ( .A1(n9029), .A2(n5450), .ZN(n5919) );
  INV_X1 U6900 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U6901 ( .A1(n5436), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U6902 ( .A1(n8496), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5914) );
  OAI211_X1 U6903 ( .C1(n5916), .C2(n4846), .A(n5915), .B(n5914), .ZN(n5917)
         );
  INV_X1 U6904 ( .A(n5917), .ZN(n5918) );
  NOR2_X1 U6905 ( .A1(n9186), .A2(n8511), .ZN(n9027) );
  NAND2_X1 U6906 ( .A1(n9028), .A2(n9027), .ZN(n5924) );
  INV_X1 U6907 ( .A(n5920), .ZN(n5921) );
  NAND2_X1 U6908 ( .A1(n5922), .A2(n5921), .ZN(n5923) );
  NAND2_X1 U6909 ( .A1(n5924), .A2(n5923), .ZN(n8999) );
  INV_X1 U6910 ( .A(n5925), .ZN(n5928) );
  NAND2_X1 U6911 ( .A1(n5926), .A2(SI_24_), .ZN(n5927) );
  INV_X1 U6912 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8228) );
  INV_X1 U6913 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8229) );
  MUX2_X1 U6914 ( .A(n8228), .B(n8229), .S(n6778), .Z(n5931) );
  INV_X1 U6915 ( .A(SI_25_), .ZN(n5930) );
  NAND2_X1 U6916 ( .A1(n5931), .A2(n5930), .ZN(n5972) );
  INV_X1 U6917 ( .A(n5931), .ZN(n5932) );
  NAND2_X1 U6918 ( .A1(n5932), .A2(SI_25_), .ZN(n5933) );
  NAND2_X1 U6919 ( .A1(n5972), .A2(n5933), .ZN(n5947) );
  NAND2_X1 U6920 ( .A1(n8226), .A2(n5561), .ZN(n5935) );
  OR2_X1 U6921 ( .A1(n8503), .A2(n8228), .ZN(n5934) );
  XNOR2_X1 U6922 ( .A(n9195), .B(n5982), .ZN(n5942) );
  INV_X1 U6923 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10198) );
  NAND2_X1 U6924 ( .A1(n5936), .A2(n10198), .ZN(n5937) );
  INV_X1 U6925 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U6926 ( .A1(n8496), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U6927 ( .A1(n5436), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5938) );
  OAI211_X1 U6928 ( .C1(n5940), .C2(n4846), .A(n5939), .B(n5938), .ZN(n5941)
         );
  AOI21_X1 U6929 ( .B1(n9194), .B2(n6051), .A(n5941), .ZN(n9087) );
  NOR2_X1 U6930 ( .A1(n9087), .A2(n8511), .ZN(n5943) );
  XNOR2_X1 U6931 ( .A(n5942), .B(n5943), .ZN(n9000) );
  NAND2_X1 U6932 ( .A1(n8999), .A2(n9000), .ZN(n5946) );
  INV_X1 U6933 ( .A(n5942), .ZN(n5944) );
  NAND2_X1 U6934 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  INV_X1 U6935 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8352) );
  INV_X1 U6936 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8354) );
  MUX2_X1 U6937 ( .A(n8352), .B(n8354), .S(n6781), .Z(n5950) );
  INV_X1 U6938 ( .A(SI_26_), .ZN(n5949) );
  NAND2_X1 U6939 ( .A1(n5950), .A2(n5949), .ZN(n5971) );
  INV_X1 U6940 ( .A(n5950), .ZN(n5951) );
  NAND2_X1 U6941 ( .A1(n5951), .A2(SI_26_), .ZN(n5973) );
  AND2_X1 U6942 ( .A1(n5971), .A2(n5973), .ZN(n5952) );
  OR2_X1 U6943 ( .A1(n8503), .A2(n8352), .ZN(n5954) );
  XNOR2_X1 U6944 ( .A(n9422), .B(n7400), .ZN(n5968) );
  INV_X1 U6945 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U6946 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  NAND2_X1 U6947 ( .A1(n5999), .A2(n5959), .ZN(n9072) );
  OR2_X1 U6948 ( .A1(n9072), .A2(n5450), .ZN(n5965) );
  INV_X1 U6949 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U6950 ( .A1(n5436), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U6951 ( .A1(n8496), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5960) );
  OAI211_X1 U6952 ( .C1(n5962), .C2(n4846), .A(n5961), .B(n5960), .ZN(n5963)
         );
  INV_X1 U6953 ( .A(n5963), .ZN(n5964) );
  INV_X1 U6954 ( .A(n9187), .ZN(n9086) );
  NAND2_X1 U6955 ( .A1(n9086), .A2(n7743), .ZN(n5966) );
  XNOR2_X1 U6956 ( .A(n5968), .B(n5966), .ZN(n9068) );
  NAND2_X1 U6957 ( .A1(n9067), .A2(n9068), .ZN(n5970) );
  INV_X1 U6958 ( .A(n5966), .ZN(n5967) );
  NAND2_X1 U6959 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  AND2_X1 U6960 ( .A1(n5972), .A2(n5971), .ZN(n5975) );
  INV_X1 U6961 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8418) );
  INV_X1 U6962 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8388) );
  MUX2_X1 U6963 ( .A(n8418), .B(n8388), .S(n6778), .Z(n5977) );
  INV_X1 U6964 ( .A(SI_27_), .ZN(n10032) );
  NAND2_X1 U6965 ( .A1(n5977), .A2(n10032), .ZN(n5993) );
  INV_X1 U6966 ( .A(n5977), .ZN(n5978) );
  NAND2_X1 U6967 ( .A1(n5978), .A2(SI_27_), .ZN(n5979) );
  AND2_X1 U6968 ( .A1(n5993), .A2(n5979), .ZN(n5991) );
  NAND2_X1 U6969 ( .A1(n8387), .A2(n5561), .ZN(n5981) );
  OR2_X1 U6970 ( .A1(n8503), .A2(n8418), .ZN(n5980) );
  XNOR2_X1 U6971 ( .A(n9416), .B(n5982), .ZN(n5987) );
  XNOR2_X1 U6972 ( .A(n5999), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9151) );
  INV_X1 U6973 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U6974 ( .A1(n5436), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U6975 ( .A1(n8496), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5983) );
  OAI211_X1 U6976 ( .C1(n5985), .C2(n4846), .A(n5984), .B(n5983), .ZN(n5986)
         );
  NOR2_X1 U6977 ( .A1(n9069), .A2(n8511), .ZN(n5988) );
  XNOR2_X1 U6978 ( .A(n5987), .B(n5988), .ZN(n8964) );
  INV_X1 U6979 ( .A(n5987), .ZN(n5989) );
  AND2_X1 U6980 ( .A1(n5989), .A2(n5988), .ZN(n5990) );
  AOI21_X1 U6981 ( .B1(n8963), .B2(n8964), .A(n5990), .ZN(n6044) );
  MUX2_X1 U6982 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6778), .Z(n6069) );
  INV_X1 U6983 ( .A(SI_28_), .ZN(n6070) );
  XNOR2_X1 U6984 ( .A(n6069), .B(n6070), .ZN(n6067) );
  INV_X1 U6985 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8420) );
  OR2_X1 U6986 ( .A1(n8503), .A2(n8420), .ZN(n5995) );
  INV_X1 U6987 ( .A(n9410), .ZN(n8863) );
  INV_X1 U6988 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10176) );
  INV_X1 U6989 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5997) );
  OAI21_X1 U6990 ( .B1(n5999), .B2(n10176), .A(n5997), .ZN(n6000) );
  NAND2_X1 U6991 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5998) );
  OR2_X1 U6992 ( .A1(n5999), .A2(n5998), .ZN(n6046) );
  INV_X1 U6993 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U6994 ( .A1(n8496), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U6995 ( .A1(n5436), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6001) );
  OAI211_X1 U6996 ( .C1(n6003), .C2(n4846), .A(n6002), .B(n6001), .ZN(n6004)
         );
  INV_X1 U6997 ( .A(n6004), .ZN(n6005) );
  NAND2_X1 U6998 ( .A1(n9084), .A2(n7743), .ZN(n6006) );
  MUX2_X1 U6999 ( .A(n6006), .B(n9084), .S(n7400), .Z(n6041) );
  INV_X1 U7000 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7001 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  NAND2_X1 U7002 ( .A1(n6009), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6035) );
  INV_X1 U7003 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7004 ( .A1(n6035), .A2(n6034), .ZN(n6010) );
  NAND2_X1 U7005 ( .A1(n6010), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6012) );
  INV_X1 U7006 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6011) );
  XNOR2_X1 U7007 ( .A(n6012), .B(n6011), .ZN(n8103) );
  XNOR2_X1 U7008 ( .A(n8103), .B(P2_B_REG_SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7009 ( .A1(n6013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6014) );
  MUX2_X1 U7010 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6014), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6015) );
  NAND2_X1 U7011 ( .A1(n6015), .A2(n4923), .ZN(n8227) );
  NAND2_X1 U7012 ( .A1(n4923), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6016) );
  MUX2_X1 U7013 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6016), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6018) );
  NAND2_X1 U7014 ( .A1(n6018), .A2(n6017), .ZN(n8353) );
  AOI21_X1 U7015 ( .B1(n6019), .B2(n8227), .A(n8353), .ZN(n6030) );
  INV_X1 U7016 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10353) );
  AND2_X1 U7017 ( .A1(n8103), .A2(n8353), .ZN(n10354) );
  AOI21_X1 U7018 ( .B1(n6030), .B2(n10353), .A(n10354), .ZN(n7699) );
  NOR4_X1 U7019 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6023) );
  NOR4_X1 U7020 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6022) );
  NOR4_X1 U7021 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6021) );
  NOR4_X1 U7022 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6020) );
  NAND4_X1 U7023 ( .A1(n6023), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n6029)
         );
  NOR2_X1 U7024 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6027) );
  NOR4_X1 U7025 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6026) );
  NOR4_X1 U7026 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6025) );
  NOR4_X1 U7027 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6024) );
  NAND4_X1 U7028 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n6028)
         );
  OAI21_X1 U7029 ( .B1(n6029), .B2(n6028), .A(n6030), .ZN(n7383) );
  NAND2_X1 U7030 ( .A1(n7699), .A2(n7383), .ZN(n6031) );
  INV_X1 U7031 ( .A(n6030), .ZN(n10002) );
  NAND2_X1 U7032 ( .A1(n8227), .A2(n8353), .ZN(n10003) );
  OAI21_X1 U7033 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n10002), .A(n10003), .ZN(
        n7698) );
  NOR2_X1 U7034 ( .A1(n6031), .A2(n7698), .ZN(n7173) );
  INV_X1 U7035 ( .A(n8103), .ZN(n6033) );
  NOR2_X1 U7036 ( .A1(n8353), .A2(n8227), .ZN(n6032) );
  XNOR2_X1 U7037 ( .A(n6035), .B(n6034), .ZN(n6056) );
  AND2_X1 U7038 ( .A1(n6056), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10355) );
  INV_X1 U7039 ( .A(n10355), .ZN(n6036) );
  INV_X1 U7040 ( .A(n8689), .ZN(n10001) );
  NAND2_X1 U7041 ( .A1(n7173), .A2(n10001), .ZN(n6052) );
  INV_X1 U7042 ( .A(n8686), .ZN(n10452) );
  OR2_X1 U7043 ( .A1(n5364), .A2(n10452), .ZN(n7717) );
  OR2_X1 U7044 ( .A1(n6052), .A2(n7717), .ZN(n6037) );
  NAND2_X1 U7045 ( .A1(n6037), .A2(n10471), .ZN(n9079) );
  NOR3_X1 U7046 ( .A1(n8863), .A2(n6041), .A3(n9079), .ZN(n6038) );
  AOI21_X1 U7047 ( .B1(n8863), .B2(n6041), .A(n6038), .ZN(n6039) );
  NOR2_X1 U7048 ( .A1(n6044), .A2(n6039), .ZN(n6066) );
  INV_X1 U7049 ( .A(n9079), .ZN(n9016) );
  NAND3_X1 U7050 ( .A1(n9410), .A2(n9016), .A3(n6041), .ZN(n6040) );
  OAI21_X1 U7051 ( .B1(n9410), .B2(n6041), .A(n6040), .ZN(n6043) );
  AND2_X1 U7052 ( .A1(n8691), .A2(n8521), .ZN(n7398) );
  NAND2_X1 U7053 ( .A1(n5364), .A2(n9143), .ZN(n8690) );
  INV_X1 U7054 ( .A(n9081), .ZN(n9009) );
  AOI21_X1 U7055 ( .B1(n9410), .B2(n9079), .A(n9009), .ZN(n6042) );
  INV_X1 U7056 ( .A(n6045), .ZN(n6065) );
  INV_X1 U7057 ( .A(n6046), .ZN(n8884) );
  INV_X1 U7058 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7059 ( .A1(n5436), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7060 ( .A1(n8496), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6047) );
  OAI211_X1 U7061 ( .C1(n6049), .C2(n4846), .A(n6048), .B(n6047), .ZN(n6050)
         );
  AOI21_X1 U7062 ( .B1(n8884), .B2(n6051), .A(n6050), .ZN(n8866) );
  OR2_X1 U7063 ( .A1(n6052), .A2(n8690), .ZN(n9076) );
  OR2_X1 U7064 ( .A1(n9076), .A2(n9341), .ZN(n9059) );
  INV_X1 U7065 ( .A(n7173), .ZN(n6055) );
  OAI22_X1 U7066 ( .A1(n10575), .A2(P2_U3152), .B1(n8689), .B2(n7717), .ZN(
        n6054) );
  NAND2_X1 U7067 ( .A1(n6055), .A2(n6054), .ZN(n6059) );
  AOI21_X1 U7068 ( .B1(n8690), .B2(n7398), .A(n6749), .ZN(n7384) );
  OR2_X1 U7069 ( .A1(n6056), .A2(P2_U3152), .ZN(n8694) );
  OAI21_X1 U7070 ( .B1(n7384), .B2(P2_U3152), .A(n8694), .ZN(n6057) );
  INV_X1 U7071 ( .A(n6057), .ZN(n6058) );
  NAND2_X1 U7072 ( .A1(n6059), .A2(n6058), .ZN(n9074) );
  AOI22_X1 U7073 ( .A1(n8861), .A2(n9074), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6060) );
  OAI21_X1 U7074 ( .B1(n8866), .B2(n9059), .A(n6060), .ZN(n6061) );
  INV_X1 U7075 ( .A(n6061), .ZN(n6064) );
  INV_X1 U7076 ( .A(n9069), .ZN(n9085) );
  INV_X1 U7077 ( .A(n6053), .ZN(n6062) );
  OR2_X1 U7078 ( .A1(n9076), .A2(n9343), .ZN(n9062) );
  INV_X1 U7079 ( .A(n9062), .ZN(n9039) );
  OAI21_X1 U7080 ( .B1(n6066), .B2(n6065), .A(n5325), .ZN(P2_U3222) );
  INV_X1 U7081 ( .A(n6069), .ZN(n6071) );
  NAND2_X1 U7082 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  MUX2_X1 U7083 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6778), .Z(n6074) );
  INV_X1 U7084 ( .A(SI_29_), .ZN(n6075) );
  XNOR2_X1 U7085 ( .A(n6074), .B(n6075), .ZN(n6530) );
  INV_X1 U7086 ( .A(n6074), .ZN(n6076) );
  NAND2_X1 U7087 ( .A1(n6076), .A2(n6075), .ZN(n6077) );
  INV_X1 U7088 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8873) );
  INV_X1 U7089 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8469) );
  MUX2_X1 U7090 ( .A(n8873), .B(n8469), .S(n6778), .Z(n6080) );
  INV_X1 U7091 ( .A(SI_30_), .ZN(n6079) );
  NAND2_X1 U7092 ( .A1(n6080), .A2(n6079), .ZN(n6126) );
  INV_X1 U7093 ( .A(n6080), .ZN(n6081) );
  NAND2_X1 U7094 ( .A1(n6081), .A2(SI_30_), .ZN(n6082) );
  AND2_X1 U7095 ( .A1(n6126), .A2(n6082), .ZN(n6124) );
  NAND2_X1 U7096 ( .A1(n6360), .A2(n6083), .ZN(n6404) );
  INV_X1 U7097 ( .A(n6404), .ZN(n6085) );
  NAND2_X1 U7098 ( .A1(n6085), .A2(n5315), .ZN(n6183) );
  INV_X1 U7099 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6088) );
  INV_X1 U7100 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6087) );
  NOR2_X1 U7101 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6091) );
  NOR2_X1 U7102 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6090) );
  NOR2_X1 U7103 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6089) );
  NAND4_X1 U7104 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n6186)
         );
  INV_X1 U7105 ( .A(n6186), .ZN(n6098) );
  NOR2_X1 U7106 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6096) );
  NOR2_X1 U7107 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6095) );
  NOR2_X1 U7108 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6094) );
  NOR2_X1 U7109 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6093) );
  INV_X1 U7110 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6100) );
  INV_X1 U7111 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6102) );
  INV_X1 U7112 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7113 ( .A1(n8495), .A2(n6340), .ZN(n6107) );
  OR2_X1 U7114 ( .A1(n6532), .A2(n8469), .ZN(n6106) );
  INV_X1 U7115 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6108) );
  INV_X1 U7116 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6110) );
  INV_X1 U7117 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6113) );
  OR2_X1 U7118 ( .A1(n6389), .A2(n6113), .ZN(n6118) );
  NAND2_X4 U7119 ( .A1(n6151), .A2(n8422), .ZN(n6525) );
  INV_X1 U7120 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9712) );
  OR2_X1 U7121 ( .A1(n6525), .A2(n9712), .ZN(n6117) );
  NAND2_X2 U7122 ( .A1(n8470), .A2(n8422), .ZN(n6378) );
  INV_X1 U7123 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6115) );
  OR2_X1 U7124 ( .A1(n6378), .A2(n6115), .ZN(n6116) );
  AND3_X1 U7125 ( .A1(n6118), .A2(n6117), .A3(n6116), .ZN(n9723) );
  INV_X1 U7126 ( .A(n6711), .ZN(n6135) );
  INV_X1 U7127 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6119) );
  OR2_X1 U7128 ( .A1(n6389), .A2(n6119), .ZN(n6123) );
  INV_X1 U7129 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8708) );
  OR2_X1 U7130 ( .A1(n6525), .A2(n8708), .ZN(n6122) );
  INV_X1 U7131 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6120) );
  OR2_X1 U7132 ( .A1(n6378), .A2(n6120), .ZN(n6121) );
  AND3_X1 U7133 ( .A1(n6123), .A2(n6122), .A3(n6121), .ZN(n8707) );
  INV_X1 U7134 ( .A(n8707), .ZN(n6817) );
  NAND2_X1 U7135 ( .A1(n6125), .A2(n6124), .ZN(n6127) );
  MUX2_X1 U7136 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6778), .Z(n6129) );
  INV_X1 U7137 ( .A(SI_31_), .ZN(n6128) );
  XNOR2_X1 U7138 ( .A(n6129), .B(n6128), .ZN(n6130) );
  NAND2_X1 U7139 ( .A1(n9997), .A2(n6340), .ZN(n6133) );
  INV_X1 U7140 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9993) );
  OR2_X1 U7141 ( .A1(n6532), .A2(n9993), .ZN(n6132) );
  NAND2_X1 U7142 ( .A1(n9874), .A2(n8707), .ZN(n6716) );
  INV_X1 U7143 ( .A(n6716), .ZN(n6134) );
  AOI21_X1 U7144 ( .B1(n6135), .B2(n6817), .A(n6134), .ZN(n6660) );
  NAND2_X1 U7145 ( .A1(n7686), .A2(n6340), .ZN(n6138) );
  INV_X1 U7146 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6136) );
  OR2_X1 U7147 ( .A1(n6532), .A2(n6136), .ZN(n6137) );
  INV_X1 U7148 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6333) );
  INV_X1 U7149 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6279) );
  INV_X1 U7150 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6319) );
  INV_X1 U7151 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8241) );
  INV_X1 U7152 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7802) );
  INV_X1 U7153 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9620) );
  INV_X1 U7154 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6160) );
  INV_X1 U7155 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7156 ( .A1(n6162), .A2(n6149), .ZN(n6150) );
  NAND2_X1 U7157 ( .A1(n6175), .A2(n6150), .ZN(n9836) );
  OR2_X1 U7158 ( .A1(n9836), .A2(n6535), .ZN(n6157) );
  INV_X1 U7159 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7160 ( .A1(n6368), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7161 ( .A1(n6424), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6152) );
  OAI211_X1 U7162 ( .C1(n6154), .C2(n6525), .A(n6153), .B(n6152), .ZN(n6155)
         );
  INV_X1 U7163 ( .A(n6155), .ZN(n6156) );
  NAND2_X1 U7164 ( .A1(n7610), .A2(n6340), .ZN(n6159) );
  OR2_X1 U7165 ( .A1(n6532), .A2(n7611), .ZN(n6158) );
  NAND2_X1 U7166 ( .A1(n6194), .A2(n6160), .ZN(n6161) );
  AND2_X1 U7167 ( .A1(n6162), .A2(n6161), .ZN(n9844) );
  NAND2_X1 U7168 ( .A1(n9844), .A2(n6376), .ZN(n6168) );
  INV_X1 U7169 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7170 ( .A1(n6424), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7171 ( .A1(n6368), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6163) );
  OAI211_X1 U7172 ( .C1(n6165), .C2(n6499), .A(n6164), .B(n6163), .ZN(n6166)
         );
  INV_X1 U7173 ( .A(n6166), .ZN(n6167) );
  NAND2_X1 U7174 ( .A1(n9926), .A2(n8813), .ZN(n8715) );
  INV_X1 U7175 ( .A(n8715), .ZN(n6169) );
  NAND2_X1 U7176 ( .A1(n6551), .A2(n6169), .ZN(n6170) );
  NAND2_X1 U7177 ( .A1(n9922), .A2(n9608), .ZN(n8716) );
  AND2_X1 U7178 ( .A1(n6170), .A2(n8716), .ZN(n6637) );
  NAND2_X1 U7179 ( .A1(n7896), .A2(n6340), .ZN(n6173) );
  OR2_X1 U7180 ( .A1(n6532), .A2(n6171), .ZN(n6172) );
  INV_X1 U7181 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U7182 ( .A1(n6175), .A2(n9606), .ZN(n6176) );
  NAND2_X1 U7183 ( .A1(n6460), .A2(n6176), .ZN(n9813) );
  OR2_X1 U7184 ( .A1(n9813), .A2(n6535), .ZN(n6182) );
  INV_X1 U7185 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7186 ( .A1(n6368), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7187 ( .A1(n6424), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6177) );
  OAI211_X1 U7188 ( .C1(n6499), .C2(n6179), .A(n6178), .B(n6177), .ZN(n6180)
         );
  INV_X1 U7189 ( .A(n6180), .ZN(n6181) );
  NAND2_X1 U7190 ( .A1(n6182), .A2(n6181), .ZN(n9831) );
  INV_X1 U7191 ( .A(n9831), .ZN(n9536) );
  NAND2_X1 U7192 ( .A1(n9916), .A2(n9536), .ZN(n8717) );
  NAND2_X1 U7193 ( .A1(n6637), .A2(n8717), .ZN(n6456) );
  NAND2_X1 U7194 ( .A1(n7476), .A2(n6340), .ZN(n6191) );
  BUF_X1 U7195 ( .A(n6183), .Z(n6434) );
  NOR2_X2 U7196 ( .A1(n6434), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6341) );
  INV_X1 U7197 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6184) );
  NOR2_X1 U7198 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6185) );
  NOR2_X2 U7199 ( .A1(n6198), .A2(n6186), .ZN(n6545) );
  INV_X1 U7200 ( .A(n6545), .ZN(n6187) );
  NAND2_X1 U7201 ( .A1(n6187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6189) );
  INV_X1 U7202 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6188) );
  INV_X1 U7203 ( .A(n9834), .ZN(n7541) );
  AOI22_X1 U7204 ( .A1(n6436), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7541), .B2(
        n10265), .ZN(n6190) );
  INV_X1 U7205 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6197) );
  INV_X1 U7206 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7207 ( .A1(n6209), .A2(n6192), .ZN(n6193) );
  NAND2_X1 U7208 ( .A1(n6194), .A2(n6193), .ZN(n9859) );
  OR2_X1 U7209 ( .A1(n9859), .A2(n6535), .ZN(n6196) );
  AOI22_X1 U7210 ( .A1(n6424), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n6368), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n6195) );
  OAI211_X1 U7211 ( .C1(n6525), .C2(n6197), .A(n6196), .B(n6195), .ZN(n9849)
         );
  INV_X1 U7212 ( .A(n9849), .ZN(n9624) );
  NAND2_X1 U7213 ( .A1(n9931), .A2(n9624), .ZN(n8714) );
  NOR2_X1 U7214 ( .A1(n6456), .A2(n5122), .ZN(n6696) );
  NAND2_X1 U7215 ( .A1(n7286), .A2(n6340), .ZN(n6207) );
  NOR2_X1 U7216 ( .A1(n6274), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6303) );
  NOR2_X1 U7217 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6199) );
  NAND2_X1 U7218 ( .A1(n6303), .A2(n6199), .ZN(n6249) );
  OR2_X1 U7219 ( .A1(n6249), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6251) );
  OR2_X1 U7220 ( .A1(n6251), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7221 ( .A1(n6200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6224) );
  INV_X1 U7222 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7223 ( .A1(n6224), .A2(n6201), .ZN(n6202) );
  NAND2_X1 U7224 ( .A1(n6202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6213) );
  INV_X1 U7225 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7226 ( .A1(n6213), .A2(n6203), .ZN(n6204) );
  NAND2_X1 U7227 ( .A1(n6204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6205) );
  XNOR2_X1 U7228 ( .A(n6205), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U7229 ( .A1(n9699), .A2(n10265), .B1(n6436), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7230 ( .A1(n6218), .A2(n9620), .ZN(n6208) );
  AND2_X1 U7231 ( .A1(n6209), .A2(n6208), .ZN(n9618) );
  NAND2_X1 U7232 ( .A1(n9618), .A2(n6376), .ZN(n6212) );
  AOI22_X1 U7233 ( .A1(n6363), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n6368), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7234 ( .A1(n6424), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6210) );
  AND3_X1 U7235 ( .A1(n6212), .A2(n6211), .A3(n6210), .ZN(n8794) );
  NAND2_X1 U7236 ( .A1(n9627), .A2(n8794), .ZN(n8711) );
  NAND2_X1 U7237 ( .A1(n7266), .A2(n6340), .ZN(n6215) );
  XNOR2_X1 U7238 ( .A(n6213), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9687) );
  AOI22_X1 U7239 ( .A1(n9687), .A2(n10265), .B1(n6436), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n6214) );
  INV_X1 U7240 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7241 ( .A1(n6228), .A2(n6216), .ZN(n6217) );
  NAND2_X1 U7242 ( .A1(n6218), .A2(n6217), .ZN(n9583) );
  OR2_X1 U7243 ( .A1(n9583), .A2(n6535), .ZN(n6223) );
  NAND2_X1 U7244 ( .A1(n6424), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7245 ( .A1(n6368), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6219) );
  AND2_X1 U7246 ( .A1(n6220), .A2(n6219), .ZN(n6222) );
  NAND2_X1 U7247 ( .A1(n6374), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7248 ( .A1(n9942), .A2(n8784), .ZN(n8449) );
  NAND2_X1 U7249 ( .A1(n7231), .A2(n6340), .ZN(n6226) );
  XNOR2_X1 U7250 ( .A(n6224), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9675) );
  AOI22_X1 U7251 ( .A1(n9675), .A2(n10265), .B1(n6436), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7252 ( .A1(n6244), .A2(n7802), .ZN(n6227) );
  AND2_X1 U7253 ( .A1(n6228), .A2(n6227), .ZN(n9571) );
  NAND2_X1 U7254 ( .A1(n9571), .A2(n6376), .ZN(n6235) );
  INV_X1 U7255 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n6229) );
  OR2_X1 U7256 ( .A1(n6389), .A2(n6229), .ZN(n6234) );
  INV_X1 U7257 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6230) );
  OR2_X1 U7258 ( .A1(n6378), .A2(n6230), .ZN(n6233) );
  INV_X1 U7259 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6231) );
  OR2_X1 U7260 ( .A1(n6499), .A2(n6231), .ZN(n6232) );
  NAND2_X1 U7261 ( .A1(n9949), .A2(n9582), .ZN(n8425) );
  AND2_X1 U7262 ( .A1(n8449), .A2(n8425), .ZN(n6236) );
  NAND2_X1 U7263 ( .A1(n8711), .A2(n6236), .ZN(n6449) );
  NAND2_X1 U7264 ( .A1(n6251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6238) );
  XNOR2_X1 U7265 ( .A(n6238), .B(n6088), .ZN(n7797) );
  INV_X1 U7266 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7155) );
  OAI22_X1 U7267 ( .A1(n7797), .A2(n6405), .B1(n6532), .B2(n7155), .ZN(n6239)
         );
  INV_X1 U7268 ( .A(n6239), .ZN(n6240) );
  NAND2_X1 U7269 ( .A1(n6424), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6248) );
  INV_X1 U7270 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7679) );
  OR2_X1 U7271 ( .A1(n6389), .A2(n7679), .ZN(n6247) );
  INV_X1 U7272 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7273 ( .A1(n6258), .A2(n6242), .ZN(n6243) );
  NAND2_X1 U7274 ( .A1(n6244), .A2(n6243), .ZN(n9645) );
  OR2_X1 U7275 ( .A1(n6535), .A2(n9645), .ZN(n6246) );
  INV_X1 U7276 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8281) );
  OR2_X1 U7277 ( .A1(n6525), .A2(n8281), .ZN(n6245) );
  NAND2_X1 U7278 ( .A1(n6939), .A2(n6340), .ZN(n6254) );
  NAND2_X1 U7279 ( .A1(n6249), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6250) );
  MUX2_X1 U7280 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6250), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6252) );
  AND2_X1 U7281 ( .A1(n6252), .A2(n6251), .ZN(n7676) );
  AOI22_X1 U7282 ( .A1(n6436), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7676), .B2(
        n10265), .ZN(n6253) );
  NAND2_X1 U7283 ( .A1(n6424), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6262) );
  INV_X1 U7284 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6255) );
  OR2_X1 U7285 ( .A1(n6389), .A2(n6255), .ZN(n6261) );
  INV_X1 U7286 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7287 ( .A1(n6310), .A2(n6256), .ZN(n6257) );
  NAND2_X1 U7288 ( .A1(n6258), .A2(n6257), .ZN(n9527) );
  OR2_X1 U7289 ( .A1(n6535), .A2(n9527), .ZN(n6260) );
  INV_X1 U7290 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8325) );
  OR2_X1 U7291 ( .A1(n6499), .A2(n8325), .ZN(n6259) );
  NAND2_X1 U7292 ( .A1(n6833), .A2(n6340), .ZN(n6266) );
  NAND2_X1 U7293 ( .A1(n6274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6264) );
  INV_X1 U7294 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6263) );
  XNOR2_X1 U7295 ( .A(n6264), .B(n6263), .ZN(n7215) );
  INV_X1 U7296 ( .A(n7215), .ZN(n7423) );
  AOI22_X1 U7297 ( .A1(n6436), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10265), 
        .B2(n7423), .ZN(n6265) );
  NAND2_X1 U7298 ( .A1(n6424), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6272) );
  INV_X1 U7299 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6267) );
  OR2_X1 U7300 ( .A1(n6389), .A2(n6267), .ZN(n6271) );
  INV_X1 U7301 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7218) );
  NAND2_X1 U7302 ( .A1(n6281), .A2(n7218), .ZN(n6268) );
  NAND2_X1 U7303 ( .A1(n6320), .A2(n6268), .ZN(n8095) );
  OR2_X1 U7304 ( .A1(n6535), .A2(n8095), .ZN(n6270) );
  INV_X1 U7305 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7214) );
  OR2_X1 U7306 ( .A1(n6525), .A2(n7214), .ZN(n6269) );
  NAND4_X1 U7307 ( .A1(n6272), .A2(n6271), .A3(n6270), .A4(n6269), .ZN(n9658)
         );
  AND2_X1 U7308 ( .A1(n8179), .A2(n8089), .ZN(n8041) );
  NAND2_X1 U7309 ( .A1(n6824), .A2(n6340), .ZN(n6278) );
  NAND2_X1 U7310 ( .A1(n6198), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6273) );
  MUX2_X1 U7311 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6273), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n6275) );
  NAND2_X1 U7312 ( .A1(n6275), .A2(n6274), .ZN(n10290) );
  INV_X1 U7313 ( .A(n10290), .ZN(n6276) );
  AOI22_X1 U7314 ( .A1(n6436), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10265), 
        .B2(n6276), .ZN(n6277) );
  NAND2_X1 U7315 ( .A1(n6374), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6286) );
  INV_X1 U7316 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7208) );
  OR2_X1 U7317 ( .A1(n6389), .A2(n7208), .ZN(n6285) );
  NAND2_X1 U7318 ( .A1(n6295), .A2(n6279), .ZN(n6280) );
  NAND2_X1 U7319 ( .A1(n6281), .A2(n6280), .ZN(n8081) );
  OR2_X1 U7320 ( .A1(n6535), .A2(n8081), .ZN(n6284) );
  INV_X1 U7321 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6282) );
  OR2_X1 U7322 ( .A1(n6378), .A2(n6282), .ZN(n6283) );
  OR2_X1 U7323 ( .A1(n8083), .A2(n7835), .ZN(n6606) );
  NAND2_X1 U7324 ( .A1(n6820), .A2(n6340), .ZN(n6292) );
  OR2_X1 U7325 ( .A1(n6287), .A2(n6110), .ZN(n6329) );
  INV_X1 U7326 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7327 ( .A1(n6329), .A2(n6288), .ZN(n6289) );
  NAND2_X1 U7328 ( .A1(n6289), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6290) );
  XNOR2_X1 U7329 ( .A(n6290), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7211) );
  AOI22_X1 U7330 ( .A1(n6436), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10265), .B2(
        n7211), .ZN(n6291) );
  NAND2_X1 U7331 ( .A1(n6424), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6299) );
  INV_X1 U7332 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6293) );
  OR2_X1 U7333 ( .A1(n6389), .A2(n6293), .ZN(n6298) );
  INV_X1 U7334 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6908) );
  NAND2_X1 U7335 ( .A1(n6335), .A2(n6908), .ZN(n6294) );
  NAND2_X1 U7336 ( .A1(n6295), .A2(n6294), .ZN(n7840) );
  OR2_X1 U7337 ( .A1(n6535), .A2(n7840), .ZN(n6297) );
  INV_X1 U7338 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7821) );
  OR2_X1 U7339 ( .A1(n6525), .A2(n7821), .ZN(n6296) );
  NAND4_X1 U7340 ( .A1(n6299), .A2(n6298), .A3(n6297), .A4(n6296), .ZN(n9659)
         );
  INV_X1 U7341 ( .A(n9659), .ZN(n6440) );
  NAND2_X1 U7342 ( .A1(n7874), .A2(n6440), .ZN(n6603) );
  INV_X1 U7343 ( .A(n6603), .ZN(n6300) );
  NAND2_X1 U7344 ( .A1(n6606), .A2(n6300), .ZN(n6301) );
  NAND2_X1 U7345 ( .A1(n8083), .A2(n7835), .ZN(n8039) );
  NAND2_X1 U7346 ( .A1(n6301), .A2(n8039), .ZN(n6302) );
  NOR2_X1 U7347 ( .A1(n8041), .A2(n6302), .ZN(n6327) );
  NAND2_X1 U7348 ( .A1(n6920), .A2(n6340), .ZN(n6308) );
  OR2_X1 U7349 ( .A1(n6303), .A2(n6110), .ZN(n6316) );
  INV_X1 U7350 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7351 ( .A1(n6316), .A2(n6304), .ZN(n6305) );
  NAND2_X1 U7352 ( .A1(n6305), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6306) );
  XNOR2_X1 U7353 ( .A(n6306), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U7354 ( .A1(n6436), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10316), 
        .B2(n10265), .ZN(n6307) );
  NAND2_X1 U7355 ( .A1(n6424), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6315) );
  INV_X1 U7356 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7419) );
  OR2_X1 U7357 ( .A1(n6389), .A2(n7419), .ZN(n6314) );
  NAND2_X1 U7358 ( .A1(n6322), .A2(n8241), .ZN(n6309) );
  NAND2_X1 U7359 ( .A1(n6310), .A2(n6309), .ZN(n8291) );
  OR2_X1 U7360 ( .A1(n6535), .A2(n8291), .ZN(n6313) );
  INV_X1 U7361 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6311) );
  OR2_X1 U7362 ( .A1(n6525), .A2(n6311), .ZN(n6312) );
  NAND2_X1 U7363 ( .A1(n9963), .A2(n9524), .ZN(n8313) );
  NAND2_X1 U7364 ( .A1(n6841), .A2(n6340), .ZN(n6318) );
  XNOR2_X1 U7365 ( .A(n6316), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U7366 ( .A1(n6436), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10265), 
        .B2(n10302), .ZN(n6317) );
  NAND2_X1 U7367 ( .A1(n6424), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6326) );
  INV_X1 U7368 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7420) );
  OR2_X1 U7369 ( .A1(n6389), .A2(n7420), .ZN(n6325) );
  NAND2_X1 U7370 ( .A1(n6320), .A2(n6319), .ZN(n6321) );
  NAND2_X1 U7371 ( .A1(n6322), .A2(n6321), .ZN(n8204) );
  OR2_X1 U7372 ( .A1(n6535), .A2(n8204), .ZN(n6324) );
  INV_X1 U7373 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8054) );
  OR2_X1 U7374 ( .A1(n6499), .A2(n8054), .ZN(n6323) );
  NAND2_X1 U7375 ( .A1(n8258), .A2(n8196), .ZN(n8249) );
  AND4_X1 U7376 ( .A1(n6621), .A2(n6327), .A3(n8313), .A4(n8249), .ZN(n6328)
         );
  AND2_X1 U7377 ( .A1(n8358), .A2(n6328), .ZN(n6442) );
  INV_X1 U7378 ( .A(n6442), .ZN(n6353) );
  NAND2_X1 U7379 ( .A1(n6814), .A2(n6340), .ZN(n6331) );
  XNOR2_X1 U7380 ( .A(n6329), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6912) );
  AOI22_X1 U7381 ( .A1(n6436), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10265), .B2(
        n6912), .ZN(n6330) );
  NAND2_X1 U7382 ( .A1(n6424), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6339) );
  INV_X1 U7383 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6332) );
  OR2_X1 U7384 ( .A1(n6389), .A2(n6332), .ZN(n6338) );
  NAND2_X1 U7385 ( .A1(n6347), .A2(n6333), .ZN(n6334) );
  NAND2_X1 U7386 ( .A1(n6335), .A2(n6334), .ZN(n7852) );
  OR2_X1 U7387 ( .A1(n6535), .A2(n7852), .ZN(n6337) );
  INV_X1 U7388 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7597) );
  OR2_X1 U7389 ( .A1(n6499), .A2(n7597), .ZN(n6336) );
  NAND2_X1 U7390 ( .A1(n7854), .A2(n7826), .ZN(n7812) );
  NAND2_X1 U7391 ( .A1(n6809), .A2(n6340), .ZN(n6344) );
  OR2_X1 U7392 ( .A1(n6341), .A2(n6110), .ZN(n6342) );
  XNOR2_X1 U7393 ( .A(n6342), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6888) );
  AOI22_X1 U7394 ( .A1(n6436), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10265), .B2(
        n6888), .ZN(n6343) );
  NAND2_X1 U7395 ( .A1(n6344), .A2(n6343), .ZN(n7631) );
  NAND2_X1 U7396 ( .A1(n6424), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6351) );
  INV_X1 U7397 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6345) );
  OR2_X1 U7398 ( .A1(n6389), .A2(n6345), .ZN(n6350) );
  INV_X1 U7399 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7538) );
  OR2_X1 U7400 ( .A1(n6525), .A2(n7538), .ZN(n6349) );
  INV_X1 U7401 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U7402 ( .A1(n6428), .A2(n6885), .ZN(n6346) );
  NAND2_X1 U7403 ( .A1(n6347), .A2(n6346), .ZN(n7644) );
  OR2_X1 U7404 ( .A1(n6535), .A2(n7644), .ZN(n6348) );
  NAND2_X1 U7405 ( .A1(n7631), .A2(n7632), .ZN(n7591) );
  NAND2_X1 U7406 ( .A1(n7812), .A2(n7591), .ZN(n6352) );
  OR3_X1 U7407 ( .A1(n6449), .A2(n6353), .A3(n6352), .ZN(n6694) );
  NAND2_X1 U7408 ( .A1(n6376), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6357) );
  INV_X1 U7409 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6847) );
  INV_X1 U7410 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6354) );
  NAND4_X2 U7411 ( .A1(n6358), .A2(n6357), .A3(n6356), .A4(n6355), .ZN(n7129)
         );
  NAND2_X1 U7412 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6359) );
  MUX2_X1 U7413 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6359), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n6362) );
  INV_X1 U7414 ( .A(n6360), .ZN(n6361) );
  NAND2_X1 U7415 ( .A1(n6362), .A2(n6361), .ZN(n6864) );
  INV_X1 U7416 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6782) );
  INV_X1 U7417 ( .A(n6525), .ZN(n6363) );
  NAND2_X1 U7418 ( .A1(n6363), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6367) );
  INV_X1 U7419 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6364) );
  OR2_X1 U7420 ( .A1(n6378), .A2(n6364), .ZN(n6366) );
  NAND2_X1 U7421 ( .A1(n6376), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U7422 ( .A1(n6368), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7023) );
  INV_X1 U7423 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6369) );
  XNOR2_X1 U7424 ( .A(n6370), .B(n6369), .ZN(n9999) );
  NAND2_X1 U7425 ( .A1(n6405), .A2(n9999), .ZN(n6372) );
  NOR2_X1 U7426 ( .A1(n7128), .A2(n10441), .ZN(n7342) );
  OR2_X1 U7427 ( .A1(n7129), .A2(n10459), .ZN(n6373) );
  NAND2_X1 U7428 ( .A1(n7341), .A2(n6373), .ZN(n6670) );
  INV_X1 U7429 ( .A(n6525), .ZN(n6374) );
  NAND2_X1 U7430 ( .A1(n6374), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6382) );
  INV_X1 U7431 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6375) );
  INV_X1 U7432 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6377) );
  OR2_X1 U7433 ( .A1(n6378), .A2(n6377), .ZN(n6379) );
  NAND4_X1 U7434 ( .A1(n6382), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(n7072)
         );
  INV_X1 U7435 ( .A(n7072), .ZN(n6387) );
  INV_X1 U7436 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6802) );
  OR2_X1 U7437 ( .A1(n6360), .A2(n6110), .ZN(n6384) );
  XNOR2_X1 U7438 ( .A(n6384), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10417) );
  INV_X1 U7439 ( .A(n10417), .ZN(n6848) );
  OR2_X1 U7440 ( .A1(n6405), .A2(n6848), .ZN(n6385) );
  NAND2_X1 U7441 ( .A1(n7141), .A2(n6674), .ZN(n7274) );
  NAND2_X1 U7442 ( .A1(n6424), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6393) );
  OR2_X1 U7443 ( .A1(n6535), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6392) );
  INV_X1 U7444 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6388) );
  OR2_X1 U7445 ( .A1(n6499), .A2(n6388), .ZN(n6391) );
  INV_X1 U7446 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6846) );
  OR2_X1 U7447 ( .A1(n6389), .A2(n6846), .ZN(n6390) );
  OR2_X1 U7448 ( .A1(n6383), .A2(n6805), .ZN(n6397) );
  OR2_X1 U7449 ( .A1(n6532), .A2(n6804), .ZN(n6396) );
  NAND2_X1 U7450 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4873), .ZN(n6394) );
  XNOR2_X1 U7451 ( .A(n6394), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10340) );
  INV_X1 U7452 ( .A(n10340), .ZN(n6806) );
  OR2_X1 U7453 ( .A1(n6405), .A2(n6806), .ZN(n6395) );
  NAND2_X1 U7454 ( .A1(n7092), .A2(n7508), .ZN(n6677) );
  NAND2_X1 U7455 ( .A1(n7274), .A2(n6677), .ZN(n6398) );
  OR2_X1 U7456 ( .A1(n7092), .A2(n7508), .ZN(n6679) );
  NAND2_X1 U7457 ( .A1(n6424), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6403) );
  INV_X1 U7458 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6399) );
  OR2_X1 U7459 ( .A1(n6389), .A2(n6399), .ZN(n6402) );
  OAI21_X1 U7460 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6411), .ZN(n7484) );
  OR2_X1 U7461 ( .A1(n6535), .A2(n7484), .ZN(n6401) );
  INV_X1 U7462 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7485) );
  OR2_X1 U7463 ( .A1(n6525), .A2(n7485), .ZN(n6400) );
  OR2_X1 U7464 ( .A1(n6808), .A2(n6383), .ZN(n6408) );
  NAND2_X1 U7465 ( .A1(n6404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6419) );
  XNOR2_X1 U7466 ( .A(n6419), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10428) );
  INV_X1 U7467 ( .A(n10428), .ZN(n6850) );
  OR2_X1 U7468 ( .A1(n6405), .A2(n6850), .ZN(n6407) );
  INV_X1 U7469 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6807) );
  OR2_X1 U7470 ( .A1(n6532), .A2(n6807), .ZN(n6406) );
  OR2_X1 U7471 ( .A1(n9663), .A2(n7486), .ZN(n6683) );
  INV_X1 U7472 ( .A(n6683), .ZN(n6409) );
  NAND2_X1 U7473 ( .A1(n9663), .A2(n7486), .ZN(n6681) );
  NAND2_X1 U7474 ( .A1(n6424), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6417) );
  INV_X1 U7475 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6852) );
  OR2_X1 U7476 ( .A1(n6389), .A2(n6852), .ZN(n6416) );
  INV_X1 U7477 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U7478 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  NAND2_X1 U7479 ( .A1(n6426), .A2(n6412), .ZN(n7443) );
  OR2_X1 U7480 ( .A1(n6535), .A2(n7443), .ZN(n6415) );
  INV_X1 U7481 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6413) );
  OR2_X1 U7482 ( .A1(n6499), .A2(n6413), .ZN(n6414) );
  NAND4_X1 U7483 ( .A1(n6417), .A2(n6416), .A3(n6415), .A4(n6414), .ZN(n9662)
         );
  OR2_X1 U7484 ( .A1(n6789), .A2(n6383), .ZN(n6423) );
  NAND2_X1 U7485 ( .A1(n6419), .A2(n6418), .ZN(n6420) );
  NAND2_X1 U7486 ( .A1(n6420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6421) );
  XNOR2_X1 U7487 ( .A(n6421), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U7488 ( .A1(n6436), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10265), .B2(
        n10328), .ZN(n6422) );
  NAND2_X1 U7489 ( .A1(n9662), .A2(n10497), .ZN(n6684) );
  INV_X1 U7490 ( .A(n6684), .ZN(n6581) );
  OR2_X1 U7491 ( .A1(n7525), .A2(n6581), .ZN(n7654) );
  NAND2_X1 U7492 ( .A1(n6424), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6430) );
  INV_X1 U7493 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U7494 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  NAND2_X1 U7495 ( .A1(n6428), .A2(n6427), .ZN(n7666) );
  OR2_X1 U7496 ( .A1(n6535), .A2(n7666), .ZN(n6429) );
  NAND2_X1 U7497 ( .A1(n6430), .A2(n6429), .ZN(n6433) );
  INV_X1 U7498 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6845) );
  NOR2_X1 U7499 ( .A1(n6389), .A2(n6845), .ZN(n6432) );
  INV_X1 U7500 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7667) );
  NOR2_X1 U7501 ( .A1(n6499), .A2(n7667), .ZN(n6431) );
  OR2_X1 U7502 ( .A1(n6792), .A2(n6383), .ZN(n6438) );
  NAND2_X1 U7503 ( .A1(n6434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6435) );
  XNOR2_X1 U7504 ( .A(n6435), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U7505 ( .A1(n6436), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10265), .B2(
        n10271), .ZN(n6437) );
  NAND2_X1 U7506 ( .A1(n7647), .A2(n7781), .ZN(n6686) );
  OR2_X1 U7507 ( .A1(n9662), .A2(n10497), .ZN(n7653) );
  AND2_X1 U7508 ( .A1(n6686), .A2(n7653), .ZN(n7524) );
  OR2_X1 U7509 ( .A1(n7631), .A2(n7632), .ZN(n6688) );
  NAND2_X1 U7510 ( .A1(n7665), .A2(n9661), .ZN(n6685) );
  NAND2_X1 U7511 ( .A1(n6688), .A2(n6685), .ZN(n6439) );
  AOI21_X1 U7512 ( .B1(n7654), .B2(n7524), .A(n6439), .ZN(n6450) );
  OR2_X1 U7513 ( .A1(n7874), .A2(n6440), .ZN(n7857) );
  OR2_X1 U7514 ( .A1(n7854), .A2(n7826), .ZN(n6600) );
  NAND3_X1 U7515 ( .A1(n6606), .A2(n7857), .A3(n6600), .ZN(n6441) );
  NAND2_X1 U7516 ( .A1(n6442), .A2(n6441), .ZN(n6447) );
  OR2_X1 U7517 ( .A1(n9949), .A2(n9582), .ZN(n8426) );
  OR2_X1 U7518 ( .A1(n9963), .A2(n9524), .ZN(n6619) );
  OR2_X1 U7519 ( .A1(n8258), .A2(n8196), .ZN(n6614) );
  OR2_X1 U7520 ( .A1(n8179), .A2(n8089), .ZN(n8042) );
  AND2_X1 U7521 ( .A1(n6614), .A2(n8042), .ZN(n8247) );
  INV_X1 U7522 ( .A(n8247), .ZN(n6443) );
  NAND3_X1 U7523 ( .A1(n6443), .A2(n8313), .A3(n8249), .ZN(n6444) );
  NAND3_X1 U7524 ( .A1(n8253), .A2(n6619), .A3(n6444), .ZN(n6445) );
  NAND3_X1 U7525 ( .A1(n8358), .A2(n6621), .A3(n6445), .ZN(n6446) );
  AND4_X1 U7526 ( .A1(n6447), .A2(n8426), .A3(n6623), .A4(n6446), .ZN(n6448)
         );
  OR2_X1 U7527 ( .A1(n6449), .A2(n6448), .ZN(n6692) );
  OAI21_X1 U7528 ( .B1(n6694), .B2(n6450), .A(n6692), .ZN(n6451) );
  NAND2_X1 U7529 ( .A1(n6696), .A2(n6451), .ZN(n6468) );
  OR2_X1 U7530 ( .A1(n9926), .A2(n8813), .ZN(n6552) );
  NAND2_X1 U7531 ( .A1(n6551), .A2(n6552), .ZN(n6636) );
  NAND2_X1 U7532 ( .A1(n8712), .A2(n8448), .ZN(n6452) );
  NAND3_X1 U7533 ( .A1(n8714), .A2(n8711), .A3(n6452), .ZN(n6453) );
  OR2_X1 U7534 ( .A1(n9931), .A2(n9624), .ZN(n6632) );
  NAND2_X1 U7535 ( .A1(n6453), .A2(n6632), .ZN(n6454) );
  NOR2_X1 U7536 ( .A1(n6636), .A2(n6454), .ZN(n6455) );
  OR2_X1 U7537 ( .A1(n6456), .A2(n6455), .ZN(n6457) );
  OR2_X1 U7538 ( .A1(n9916), .A2(n9536), .ZN(n6640) );
  AND2_X1 U7539 ( .A1(n6457), .A2(n6640), .ZN(n6698) );
  NAND2_X1 U7540 ( .A1(n7921), .A2(n6340), .ZN(n6459) );
  OR2_X1 U7541 ( .A1(n6532), .A2(n7924), .ZN(n6458) );
  INV_X1 U7542 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U7543 ( .A1(n6460), .A2(n9535), .ZN(n6461) );
  NAND2_X1 U7544 ( .A1(n6472), .A2(n6461), .ZN(n9799) );
  OR2_X1 U7545 ( .A1(n9799), .A2(n6535), .ZN(n6467) );
  INV_X1 U7546 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U7547 ( .A1(n6424), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U7548 ( .A1(n6368), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6462) );
  OAI211_X1 U7549 ( .C1(n6464), .C2(n6499), .A(n6463), .B(n6462), .ZN(n6465)
         );
  INV_X1 U7550 ( .A(n6465), .ZN(n6466) );
  NAND2_X1 U7551 ( .A1(n6467), .A2(n6466), .ZN(n9819) );
  NAND2_X1 U7552 ( .A1(n9911), .A2(n9781), .ZN(n8718) );
  INV_X1 U7553 ( .A(n8718), .ZN(n6697) );
  AOI21_X1 U7554 ( .B1(n6468), .B2(n6698), .A(n6697), .ZN(n6479) );
  NAND2_X1 U7555 ( .A1(n8101), .A2(n6340), .ZN(n6471) );
  INV_X1 U7556 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n6469) );
  OR2_X1 U7557 ( .A1(n6532), .A2(n6469), .ZN(n6470) );
  INV_X1 U7558 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U7559 ( .A1(n6472), .A2(n9591), .ZN(n6473) );
  AND2_X1 U7560 ( .A1(n6484), .A2(n6473), .ZN(n9785) );
  NAND2_X1 U7561 ( .A1(n9785), .A2(n6376), .ZN(n6478) );
  INV_X1 U7562 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9786) );
  NAND2_X1 U7563 ( .A1(n6424), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U7564 ( .A1(n6368), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6474) );
  OAI211_X1 U7565 ( .C1(n9786), .C2(n6499), .A(n6475), .B(n6474), .ZN(n6476)
         );
  INV_X1 U7566 ( .A(n6476), .ZN(n6477) );
  NAND2_X1 U7567 ( .A1(n6478), .A2(n6477), .ZN(n9806) );
  OR2_X1 U7568 ( .A1(n9908), .A2(n8916), .ZN(n6580) );
  OR2_X1 U7569 ( .A1(n9911), .A2(n9781), .ZN(n6550) );
  NAND2_X1 U7570 ( .A1(n6580), .A2(n6550), .ZN(n6700) );
  NOR2_X1 U7571 ( .A1(n6479), .A2(n6700), .ZN(n6516) );
  OR2_X1 U7572 ( .A1(n6532), .A2(n8229), .ZN(n6480) );
  INV_X1 U7573 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U7574 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  NAND2_X1 U7575 ( .A1(n6507), .A2(n6485), .ZN(n9767) );
  INV_X1 U7576 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7577 ( .A1(n6368), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7578 ( .A1(n6424), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6486) );
  OAI211_X1 U7579 ( .C1(n6488), .C2(n6499), .A(n6487), .B(n6486), .ZN(n6489)
         );
  INV_X1 U7580 ( .A(n6489), .ZN(n6490) );
  NAND2_X1 U7581 ( .A1(n9908), .A2(n8916), .ZN(n8719) );
  NAND2_X1 U7582 ( .A1(n8721), .A2(n8719), .ZN(n6703) );
  NAND2_X1 U7583 ( .A1(n8387), .A2(n6340), .ZN(n6493) );
  OR2_X1 U7584 ( .A1(n6532), .A2(n8388), .ZN(n6492) );
  INV_X1 U7585 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U7586 ( .A1(n6509), .A2(n6495), .ZN(n6496) );
  NAND2_X1 U7587 ( .A1(n9739), .A2(n6376), .ZN(n6503) );
  INV_X1 U7588 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U7589 ( .A1(n6368), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U7590 ( .A1(n6424), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6497) );
  OAI211_X1 U7591 ( .C1(n6500), .C2(n6499), .A(n6498), .B(n6497), .ZN(n6501)
         );
  INV_X1 U7592 ( .A(n6501), .ZN(n6502) );
  OR2_X1 U7593 ( .A1(n6532), .A2(n8354), .ZN(n6504) );
  INV_X1 U7594 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U7595 ( .A1(n6507), .A2(n6506), .ZN(n6508) );
  NAND2_X1 U7596 ( .A1(n6509), .A2(n6508), .ZN(n9753) );
  INV_X1 U7597 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U7598 ( .A1(n6368), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U7599 ( .A1(n6424), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6510) );
  OAI211_X1 U7600 ( .C1(n6512), .C2(n6525), .A(n6511), .B(n6510), .ZN(n6513)
         );
  INV_X1 U7601 ( .A(n6513), .ZN(n6514) );
  AND2_X1 U7602 ( .A1(n6579), .A2(n6644), .ZN(n6702) );
  OAI211_X1 U7603 ( .C1(n6516), .C2(n6703), .A(n8725), .B(n6702), .ZN(n6517)
         );
  INV_X1 U7604 ( .A(n6517), .ZN(n6542) );
  NAND2_X1 U7605 ( .A1(n8419), .A2(n6340), .ZN(n6519) );
  INV_X1 U7606 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8467) );
  OR2_X1 U7607 ( .A1(n6532), .A2(n8467), .ZN(n6518) );
  INV_X1 U7608 ( .A(n6521), .ZN(n6520) );
  NAND2_X1 U7609 ( .A1(n6520), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9727) );
  INV_X1 U7610 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U7611 ( .A1(n6521), .A2(n8955), .ZN(n6522) );
  NAND2_X1 U7612 ( .A1(n9727), .A2(n6522), .ZN(n8956) );
  INV_X1 U7613 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U7614 ( .A1(n6424), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U7615 ( .A1(n6368), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6523) );
  OAI211_X1 U7616 ( .C1(n8739), .C2(n6525), .A(n6524), .B(n6523), .ZN(n6526)
         );
  INV_X1 U7617 ( .A(n6526), .ZN(n6527) );
  NAND2_X1 U7618 ( .A1(n9885), .A2(n9745), .ZN(n9718) );
  NAND2_X1 U7619 ( .A1(n9891), .A2(n8941), .ZN(n6578) );
  NAND2_X1 U7620 ( .A1(n8725), .A2(n5139), .ZN(n6529) );
  NAND3_X1 U7621 ( .A1(n9718), .A2(n6578), .A3(n6529), .ZN(n6707) );
  NAND2_X1 U7622 ( .A1(n8490), .A2(n6340), .ZN(n6534) );
  INV_X1 U7623 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8421) );
  OR2_X1 U7624 ( .A1(n6532), .A2(n8421), .ZN(n6533) );
  OR2_X1 U7625 ( .A1(n9727), .A2(n6535), .ZN(n6540) );
  INV_X1 U7626 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U7627 ( .A1(n6424), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U7628 ( .A1(n6368), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6536) );
  OAI211_X1 U7629 ( .C1(n9726), .C2(n6499), .A(n6537), .B(n6536), .ZN(n6538)
         );
  INV_X1 U7630 ( .A(n6538), .ZN(n6539) );
  NAND2_X1 U7631 ( .A1(n6540), .A2(n6539), .ZN(n9651) );
  INV_X1 U7632 ( .A(n9651), .ZN(n8959) );
  NAND2_X1 U7633 ( .A1(n6652), .A2(n6549), .ZN(n6709) );
  INV_X1 U7634 ( .A(n6709), .ZN(n6541) );
  OAI21_X1 U7635 ( .B1(n6542), .B2(n6707), .A(n6541), .ZN(n6544) );
  NAND2_X1 U7636 ( .A1(n8704), .A2(n8959), .ZN(n6708) );
  OR2_X1 U7637 ( .A1(n9723), .A2(n8707), .ZN(n6543) );
  NAND2_X1 U7638 ( .A1(n9878), .A2(n6543), .ZN(n6657) );
  NAND3_X1 U7639 ( .A1(n6544), .A2(n6708), .A3(n6657), .ZN(n6548) );
  INV_X1 U7640 ( .A(n6713), .ZN(n6663) );
  AOI21_X1 U7641 ( .B1(n6545), .B2(n6188), .A(n6110), .ZN(n6546) );
  NAND2_X1 U7642 ( .A1(n6666), .A2(n6667), .ZN(n6547) );
  NAND2_X2 U7643 ( .A1(n6547), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6573) );
  XNOR2_X2 U7644 ( .A(n6573), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7019) );
  INV_X1 U7645 ( .A(n7019), .ZN(n7687) );
  AOI211_X1 U7646 ( .C1(n6660), .C2(n6548), .A(n6663), .B(n7687), .ZN(n6571)
         );
  NAND2_X1 U7647 ( .A1(n6713), .A2(n6716), .ZN(n6569) );
  INV_X1 U7648 ( .A(n9757), .ZN(n6566) );
  INV_X1 U7649 ( .A(n9805), .ZN(n9795) );
  INV_X1 U7650 ( .A(n9830), .ZN(n6563) );
  NAND2_X1 U7651 ( .A1(n8426), .A2(n8425), .ZN(n8436) );
  NAND2_X1 U7652 ( .A1(n6614), .A2(n8249), .ZN(n8259) );
  INV_X1 U7653 ( .A(n8259), .ZN(n8050) );
  NAND2_X1 U7654 ( .A1(n6606), .A2(n8039), .ZN(n8045) );
  NAND2_X1 U7655 ( .A1(n7857), .A2(n6603), .ZN(n7816) );
  AND2_X1 U7656 ( .A1(n7128), .A2(n10441), .ZN(n6671) );
  NOR2_X1 U7657 ( .A1(n7342), .A2(n6671), .ZN(n7184) );
  NAND2_X1 U7658 ( .A1(n6679), .A2(n6677), .ZN(n7273) );
  INV_X1 U7659 ( .A(n7273), .ZN(n6554) );
  NAND4_X1 U7660 ( .A1(n7184), .A2(n6554), .A3(n7142), .A4(n6553), .ZN(n6555)
         );
  NOR2_X1 U7661 ( .A1(n6555), .A2(n7318), .ZN(n6556) );
  NAND2_X1 U7662 ( .A1(n6688), .A2(n7591), .ZN(n7535) );
  INV_X1 U7663 ( .A(n7535), .ZN(n7527) );
  AND2_X1 U7664 ( .A1(n7653), .A2(n6684), .ZN(n7301) );
  NAND4_X1 U7665 ( .A1(n6556), .A2(n7527), .A3(n7659), .A4(n7301), .ZN(n6557)
         );
  NOR4_X1 U7666 ( .A1(n8045), .A2(n7816), .A3(n7589), .A4(n6557), .ZN(n6559)
         );
  NOR2_X1 U7667 ( .A1(n8179), .A2(n9658), .ZN(n8261) );
  NAND2_X1 U7668 ( .A1(n8179), .A2(n9658), .ZN(n8264) );
  INV_X1 U7669 ( .A(n8264), .ZN(n6558) );
  OR2_X1 U7670 ( .A1(n8261), .A2(n6558), .ZN(n8172) );
  NAND4_X1 U7671 ( .A1(n8296), .A2(n8050), .A3(n6559), .A4(n8172), .ZN(n6560)
         );
  NOR4_X1 U7672 ( .A1(n8436), .A2(n8279), .A3(n8322), .A4(n6560), .ZN(n6561)
         );
  NAND4_X1 U7673 ( .A1(n4857), .A2(n8454), .A3(n8444), .A4(n6561), .ZN(n6562)
         );
  NOR4_X1 U7674 ( .A1(n9795), .A2(n6563), .A3(n5119), .A4(n6562), .ZN(n6564)
         );
  XNOR2_X1 U7675 ( .A(n9908), .B(n9806), .ZN(n9788) );
  XNOR2_X1 U7676 ( .A(n9916), .B(n9831), .ZN(n9817) );
  NAND4_X1 U7677 ( .A1(n9770), .A2(n6564), .A3(n9788), .A4(n9817), .ZN(n6565)
         );
  NOR4_X1 U7678 ( .A1(n8737), .A2(n9742), .A3(n6566), .A4(n6565), .ZN(n6567)
         );
  NAND2_X1 U7679 ( .A1(n9878), .A2(n9723), .ZN(n6714) );
  NAND4_X1 U7680 ( .A1(n6567), .A2(n9720), .A3(n6714), .A4(n6711), .ZN(n6568)
         );
  OAI21_X1 U7681 ( .B1(n6569), .B2(n6568), .A(n7687), .ZN(n6661) );
  INV_X1 U7682 ( .A(n6661), .ZN(n6570) );
  NOR2_X1 U7683 ( .A1(n6571), .A2(n6570), .ZN(n6662) );
  INV_X1 U7684 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U7685 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  XNOR2_X2 U7686 ( .A(n6576), .B(n6575), .ZN(n7125) );
  NAND2_X1 U7687 ( .A1(n6716), .A2(n6659), .ZN(n6658) );
  INV_X1 U7688 ( .A(n9874), .ZN(n6656) );
  NAND2_X1 U7689 ( .A1(n6708), .A2(n9718), .ZN(n6577) );
  MUX2_X1 U7690 ( .A(n6577), .B(n6709), .S(n6659), .Z(n6655) );
  INV_X1 U7691 ( .A(n8737), .ZN(n8727) );
  MUX2_X1 U7692 ( .A(n8725), .B(n6578), .S(n6659), .Z(n6651) );
  MUX2_X1 U7693 ( .A(n8723), .B(n6579), .S(n6659), .Z(n6649) );
  OAI21_X1 U7694 ( .B1(n6642), .B2(n6580), .A(n9770), .ZN(n6647) );
  NAND4_X1 U7695 ( .A1(n6589), .A2(n6642), .A3(n6688), .A4(n6685), .ZN(n6598)
         );
  NAND2_X1 U7696 ( .A1(n7647), .A2(n6642), .ZN(n6583) );
  NAND2_X1 U7697 ( .A1(n7632), .A2(n6642), .ZN(n6582) );
  OAI21_X1 U7698 ( .B1(n6583), .B2(n7665), .A(n6582), .ZN(n6588) );
  INV_X1 U7699 ( .A(n6583), .ZN(n6584) );
  NAND2_X1 U7700 ( .A1(n6584), .A2(n7632), .ZN(n6585) );
  NAND2_X1 U7701 ( .A1(n6585), .A2(n7781), .ZN(n6587) );
  NAND2_X1 U7702 ( .A1(n9661), .A2(n6659), .ZN(n6591) );
  OAI21_X1 U7703 ( .B1(n7632), .B2(n6591), .A(n7665), .ZN(n6586) );
  AOI22_X1 U7704 ( .A1(n7631), .A2(n6588), .B1(n6587), .B2(n6586), .ZN(n6597)
         );
  NAND4_X1 U7705 ( .A1(n6590), .A2(n7591), .A3(n6686), .A4(n6659), .ZN(n6596)
         );
  INV_X1 U7706 ( .A(n6591), .ZN(n6592) );
  NAND2_X1 U7707 ( .A1(n6592), .A2(n7665), .ZN(n6593) );
  OAI21_X1 U7708 ( .B1(n7632), .B2(n6642), .A(n6593), .ZN(n6594) );
  INV_X1 U7709 ( .A(n7631), .ZN(n7652) );
  NAND2_X1 U7710 ( .A1(n6594), .A2(n7652), .ZN(n6595) );
  NAND4_X1 U7711 ( .A1(n6598), .A2(n6597), .A3(n6596), .A4(n6595), .ZN(n6599)
         );
  NAND2_X1 U7712 ( .A1(n6599), .A2(n7810), .ZN(n6602) );
  MUX2_X1 U7713 ( .A(n7812), .B(n6600), .S(n6659), .Z(n6601) );
  NAND3_X1 U7714 ( .A1(n6602), .A2(n7814), .A3(n6601), .ZN(n6605) );
  MUX2_X1 U7715 ( .A(n6603), .B(n7857), .S(n6642), .Z(n6604) );
  NAND2_X1 U7716 ( .A1(n6605), .A2(n6604), .ZN(n6610) );
  INV_X1 U7717 ( .A(n8045), .ZN(n6609) );
  MUX2_X1 U7718 ( .A(n8039), .B(n6606), .S(n6642), .Z(n6607) );
  NAND2_X1 U7719 ( .A1(n8172), .A2(n6607), .ZN(n6608) );
  AOI21_X1 U7720 ( .B1(n6610), .B2(n6609), .A(n6608), .ZN(n6613) );
  INV_X1 U7721 ( .A(n8042), .ZN(n6611) );
  MUX2_X1 U7722 ( .A(n8041), .B(n6611), .S(n6659), .Z(n6612) );
  INV_X1 U7723 ( .A(n8322), .ZN(n8312) );
  INV_X1 U7724 ( .A(n8313), .ZN(n8251) );
  OAI21_X1 U7725 ( .B1(n6616), .B2(n8251), .A(n8253), .ZN(n6618) );
  NAND2_X1 U7726 ( .A1(n6616), .A2(n6621), .ZN(n6617) );
  INV_X1 U7727 ( .A(n6619), .ZN(n6620) );
  NAND3_X1 U7728 ( .A1(n6621), .A2(n6620), .A3(n6642), .ZN(n6622) );
  INV_X1 U7729 ( .A(n8436), .ZN(n6625) );
  MUX2_X1 U7730 ( .A(n6623), .B(n8358), .S(n6642), .Z(n6624) );
  MUX2_X1 U7731 ( .A(n8426), .B(n8425), .S(n6659), .Z(n6626) );
  NAND2_X1 U7732 ( .A1(n6627), .A2(n8444), .ZN(n6629) );
  MUX2_X1 U7733 ( .A(n8448), .B(n8449), .S(n6659), .Z(n6628) );
  NAND3_X1 U7734 ( .A1(n6629), .A2(n8454), .A3(n6628), .ZN(n6631) );
  MUX2_X1 U7735 ( .A(n8711), .B(n8712), .S(n6659), .Z(n6630) );
  NAND3_X1 U7736 ( .A1(n6631), .A2(n4857), .A3(n6630), .ZN(n6634) );
  MUX2_X1 U7737 ( .A(n8714), .B(n6632), .S(n6642), .Z(n6633) );
  NAND2_X1 U7738 ( .A1(n6634), .A2(n6633), .ZN(n6635) );
  NAND2_X1 U7739 ( .A1(n6636), .A2(n8716), .ZN(n6638) );
  MUX2_X1 U7740 ( .A(n6638), .B(n6637), .S(n6659), .Z(n6639) );
  MUX2_X1 U7741 ( .A(n6640), .B(n8717), .S(n6642), .Z(n6641) );
  AOI21_X1 U7742 ( .B1(n8719), .B2(n8718), .A(n6642), .ZN(n6643) );
  MUX2_X1 U7743 ( .A(n6644), .B(n8721), .S(n6659), .Z(n6645) );
  OAI211_X1 U7744 ( .C1(n6647), .C2(n6646), .A(n9757), .B(n6645), .ZN(n6648)
         );
  NAND3_X1 U7745 ( .A1(n5237), .A2(n6649), .A3(n6648), .ZN(n6650) );
  MUX2_X1 U7746 ( .A(n6652), .B(n6708), .S(n6659), .Z(n6653) );
  NAND2_X1 U7747 ( .A1(n7030), .A2(n7019), .ZN(n7110) );
  NOR3_X1 U7748 ( .A1(n6663), .A2(n7030), .A3(n7687), .ZN(n6664) );
  NAND2_X1 U7749 ( .A1(n6665), .A2(n6664), .ZN(n6669) );
  INV_X1 U7750 ( .A(n6671), .ZN(n6673) );
  NAND2_X1 U7751 ( .A1(n7129), .A2(n10459), .ZN(n6672) );
  NAND3_X1 U7752 ( .A1(n6673), .A2(n7019), .A3(n6672), .ZN(n6675) );
  NAND2_X1 U7753 ( .A1(n6675), .A2(n6674), .ZN(n6678) );
  OAI211_X1 U7754 ( .C1(n6670), .C2(n6678), .A(n6677), .B(n6676), .ZN(n6680)
         );
  NAND2_X1 U7755 ( .A1(n6680), .A2(n6679), .ZN(n6682) );
  NAND2_X1 U7756 ( .A1(n6682), .A2(n6681), .ZN(n6691) );
  AND2_X1 U7757 ( .A1(n7524), .A2(n6683), .ZN(n6690) );
  NAND2_X1 U7758 ( .A1(n6685), .A2(n6684), .ZN(n6687) );
  NAND2_X1 U7759 ( .A1(n6687), .A2(n6686), .ZN(n7522) );
  NAND2_X1 U7760 ( .A1(n7522), .A2(n6688), .ZN(n6689) );
  AOI21_X1 U7761 ( .B1(n6691), .B2(n6690), .A(n6689), .ZN(n6693) );
  OAI21_X1 U7762 ( .B1(n6694), .B2(n6693), .A(n6692), .ZN(n6695) );
  NAND2_X1 U7763 ( .A1(n6696), .A2(n6695), .ZN(n6699) );
  AOI21_X1 U7764 ( .B1(n6699), .B2(n6698), .A(n6697), .ZN(n6701) );
  NOR2_X1 U7765 ( .A1(n6701), .A2(n6700), .ZN(n6704) );
  OAI21_X1 U7766 ( .B1(n6704), .B2(n6703), .A(n6702), .ZN(n6705) );
  NOR2_X1 U7767 ( .A1(n9742), .A2(n6705), .ZN(n6706) );
  NOR2_X1 U7768 ( .A1(n6707), .A2(n6706), .ZN(n6710) );
  OAI21_X1 U7769 ( .B1(n6710), .B2(n6709), .A(n6708), .ZN(n6712) );
  NAND2_X1 U7770 ( .A1(n6712), .A2(n6711), .ZN(n6715) );
  NAND3_X1 U7771 ( .A1(n6715), .A2(n6714), .A3(n6713), .ZN(n6717) );
  NAND2_X1 U7772 ( .A1(n6717), .A2(n6716), .ZN(n6723) );
  NAND2_X1 U7773 ( .A1(n7018), .A2(n7541), .ZN(n7126) );
  NAND2_X1 U7774 ( .A1(n7018), .A2(n9834), .ZN(n7042) );
  INV_X1 U7775 ( .A(n7042), .ZN(n6718) );
  NAND2_X1 U7776 ( .A1(n6723), .A2(n6718), .ZN(n6722) );
  NAND2_X1 U7777 ( .A1(n6719), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6720) );
  XNOR2_X1 U7778 ( .A(n6720), .B(n5313), .ZN(n7113) );
  OR2_X1 U7779 ( .A1(n7113), .A2(P1_U3084), .ZN(n7922) );
  INV_X1 U7780 ( .A(n7922), .ZN(n6721) );
  OAI211_X1 U7781 ( .C1(n6723), .C2(n7126), .A(n6722), .B(n6721), .ZN(n6724)
         );
  OR2_X1 U7782 ( .A1(n7110), .A2(n7042), .ZN(n7182) );
  INV_X1 U7783 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U7784 ( .A1(n6730), .A2(n6727), .ZN(n6728) );
  NAND2_X1 U7785 ( .A1(n6728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6729) );
  XNOR2_X1 U7786 ( .A(n6729), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6800) );
  XNOR2_X1 U7787 ( .A(n6730), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U7788 ( .A1(n4890), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6731) );
  XNOR2_X1 U7789 ( .A(n6731), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6796) );
  AND2_X1 U7790 ( .A1(n6795), .A2(n6796), .ZN(n6732) );
  NAND2_X1 U7791 ( .A1(n6800), .A2(n6732), .ZN(n7114) );
  AND2_X1 U7792 ( .A1(n7113), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6733) );
  AND2_X1 U7793 ( .A1(n7114), .A2(n6733), .ZN(n9989) );
  INV_X1 U7794 ( .A(n9989), .ZN(n7064) );
  OR2_X1 U7795 ( .A1(n7182), .A2(n7064), .ZN(n7062) );
  NOR3_X1 U7796 ( .A1(n7062), .A2(n4847), .A3(n4848), .ZN(n6737) );
  OAI21_X1 U7797 ( .B1(n7030), .B2(n7922), .A(P1_B_REG_SCAN_IN), .ZN(n6736) );
  OR2_X1 U7798 ( .A1(n6737), .A2(n6736), .ZN(n6738) );
  INV_X1 U7799 ( .A(n7113), .ZN(n6739) );
  OR2_X1 U7800 ( .A1(n7110), .A2(n6739), .ZN(n6740) );
  OR2_X1 U7801 ( .A1(n7114), .A2(n6739), .ZN(n6872) );
  NAND2_X1 U7802 ( .A1(n6740), .A2(n6872), .ZN(n6859) );
  OR2_X1 U7803 ( .A1(n6859), .A2(n10265), .ZN(n6741) );
  NAND2_X1 U7804 ( .A1(n6741), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U7805 ( .A1(n6749), .A2(n10355), .ZN(n9104) );
  INV_X2 U7806 ( .A(n9104), .ZN(P2_U3966) );
  OR2_X1 U7807 ( .A1(n6872), .A2(P1_U3084), .ZN(n9665) );
  INV_X2 U7808 ( .A(n9665), .ZN(P1_U4006) );
  AOI211_X1 U7809 ( .C1(n6743), .C2(n6742), .A(n9081), .B(n4924), .ZN(n6748)
         );
  NOR2_X1 U7810 ( .A1(n9016), .A2(n10511), .ZN(n6747) );
  INV_X1 U7811 ( .A(n9074), .ZN(n9019) );
  INV_X1 U7812 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6744) );
  OAI22_X1 U7813 ( .A1(n9019), .A2(n7936), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6744), .ZN(n6746) );
  INV_X1 U7814 ( .A(n9096), .ZN(n7956) );
  OAI22_X1 U7815 ( .A1(n7956), .A2(n9059), .B1(n9062), .B2(n7933), .ZN(n6745)
         );
  OR4_X1 U7816 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(P2_U3215)
         );
  NAND2_X1 U7817 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6749), .ZN(n6750) );
  OAI211_X1 U7818 ( .C1(n8689), .C2(n7398), .A(n6750), .B(n8694), .ZN(n6752)
         );
  AND2_X1 U7819 ( .A1(n6752), .A2(n6751), .ZN(n6765) );
  INV_X1 U7820 ( .A(n6765), .ZN(n6753) );
  NAND2_X1 U7821 ( .A1(n6753), .A2(n9104), .ZN(n6759) );
  AND2_X1 U7822 ( .A1(n6759), .A2(n6053), .ZN(n10386) );
  INV_X1 U7823 ( .A(n10386), .ZN(n10356) );
  NOR2_X1 U7824 ( .A1(n10356), .A2(n6934), .ZN(n6777) );
  OR2_X1 U7825 ( .A1(n6787), .A2(n6754), .ZN(n6755) );
  MUX2_X1 U7826 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6754), .S(n6787), .Z(n10365)
         );
  NAND2_X1 U7827 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10364) );
  OR2_X1 U7828 ( .A1(n10365), .A2(n10364), .ZN(n10366) );
  AND2_X1 U7829 ( .A1(n6755), .A2(n10366), .ZN(n10380) );
  NAND2_X1 U7830 ( .A1(n10385), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6756) );
  OAI21_X1 U7831 ( .B1(n10385), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6756), .ZN(
        n10381) );
  NOR2_X1 U7832 ( .A1(n10380), .A2(n10381), .ZN(n10382) );
  AOI21_X1 U7833 ( .B1(n10385), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10382), .ZN(
        n6761) );
  NAND2_X1 U7834 ( .A1(n6926), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6757) );
  OAI21_X1 U7835 ( .B1(n6926), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6757), .ZN(
        n6760) );
  NOR2_X1 U7836 ( .A1(n6761), .A2(n6760), .ZN(n6932) );
  NOR2_X1 U7837 ( .A1(n6053), .A2(n8749), .ZN(n6758) );
  NAND2_X1 U7838 ( .A1(n6759), .A2(n6758), .ZN(n10394) );
  AOI211_X1 U7839 ( .C1(n6761), .C2(n6760), .A(n6932), .B(n10394), .ZN(n6776)
         );
  INV_X1 U7840 ( .A(n6787), .ZN(n10368) );
  INV_X1 U7841 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6762) );
  MUX2_X1 U7842 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6762), .S(n6787), .Z(n10371)
         );
  NAND2_X1 U7843 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10370) );
  NOR2_X1 U7844 ( .A1(n10371), .A2(n10370), .ZN(n10369) );
  AOI21_X1 U7845 ( .B1(n10368), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10369), .ZN(
        n10388) );
  NAND2_X1 U7846 ( .A1(n10385), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6763) );
  OAI21_X1 U7847 ( .B1(n10385), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6763), .ZN(
        n10389) );
  NOR2_X1 U7848 ( .A1(n10388), .A2(n10389), .ZN(n10387) );
  AOI21_X1 U7849 ( .B1(n10385), .B2(P2_REG1_REG_2__SCAN_IN), .A(n10387), .ZN(
        n6767) );
  NAND2_X1 U7850 ( .A1(n6926), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6764) );
  OAI21_X1 U7851 ( .B1(n6926), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6764), .ZN(
        n6766) );
  NOR2_X1 U7852 ( .A1(n6767), .A2(n6766), .ZN(n6925) );
  NAND2_X1 U7853 ( .A1(n6765), .A2(n8749), .ZN(n10357) );
  AOI211_X1 U7854 ( .C1(n6767), .C2(n6766), .A(n6925), .B(n10357), .ZN(n6775)
         );
  NAND2_X1 U7855 ( .A1(n10001), .A2(n7398), .ZN(n6771) );
  NAND2_X1 U7856 ( .A1(n8689), .A2(n8694), .ZN(n6769) );
  NAND2_X1 U7857 ( .A1(n6769), .A2(n6768), .ZN(n6770) );
  AND2_X1 U7858 ( .A1(n6771), .A2(n6770), .ZN(n9116) );
  INV_X1 U7859 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U7860 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n6772) );
  OAI21_X1 U7861 ( .B1(n9116), .B2(n6773), .A(n6772), .ZN(n6774) );
  OR4_X1 U7862 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(P2_U3248)
         );
  AND2_X1 U7863 ( .A1(n6778), .A2(P2_U3152), .ZN(n7289) );
  NOR2_X1 U7864 ( .A1(n6778), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9507) );
  OAI222_X1 U7865 ( .A1(n9503), .A2(n6779), .B1(n7477), .B2(n6805), .C1(
        P2_U3152), .C2(n6934), .ZN(P2_U3355) );
  AND2_X1 U7866 ( .A1(n6781), .A2(P1_U3084), .ZN(n9996) );
  OAI222_X1 U7867 ( .A1(n8841), .A2(n6782), .B1(n7481), .B2(n6786), .C1(n6864), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  OAI222_X1 U7868 ( .A1(P2_U3152), .A2(n6784), .B1(n7477), .B2(n6803), .C1(
        n6783), .C2(n9503), .ZN(P2_U3356) );
  OAI222_X1 U7869 ( .A1(P2_U3152), .A2(n6787), .B1(n7477), .B2(n6786), .C1(
        n6785), .C2(n9503), .ZN(P2_U3357) );
  INV_X1 U7870 ( .A(n10328), .ZN(n6863) );
  INV_X1 U7871 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6788) );
  OAI222_X1 U7872 ( .A1(n6863), .A2(P1_U3084), .B1(n7481), .B2(n6789), .C1(
        n6788), .C2(n8841), .ZN(P1_U3348) );
  OAI222_X1 U7873 ( .A1(n9503), .A2(n6790), .B1(n7477), .B2(n6789), .C1(
        P2_U3152), .C2(n6968), .ZN(P2_U3353) );
  INV_X1 U7874 ( .A(n8841), .ZN(n7287) );
  AOI22_X1 U7875 ( .A1(n10271), .A2(P1_STATE_REG_SCAN_IN), .B1(n7287), .B2(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n6791) );
  OAI21_X1 U7876 ( .B1(n6792), .B2(n7481), .A(n6791), .ZN(P1_U3347) );
  OAI222_X1 U7877 ( .A1(n9503), .A2(n6793), .B1(n7477), .B2(n6792), .C1(
        P2_U3152), .C2(n6983), .ZN(P2_U3352) );
  OAI222_X1 U7878 ( .A1(n9503), .A2(n6794), .B1(n7477), .B2(n6808), .C1(
        P2_U3152), .C2(n6953), .ZN(P2_U3354) );
  INV_X1 U7879 ( .A(n6795), .ZN(n8231) );
  NAND2_X1 U7880 ( .A1(n8231), .A2(P1_B_REG_SCAN_IN), .ZN(n6797) );
  INV_X1 U7881 ( .A(n6796), .ZN(n8105) );
  MUX2_X1 U7882 ( .A(P1_B_REG_SCAN_IN), .B(n6797), .S(n8105), .Z(n6798) );
  AND2_X1 U7883 ( .A1(n6798), .A2(n6800), .ZN(n7057) );
  INV_X1 U7884 ( .A(n7057), .ZN(n6799) );
  NAND2_X1 U7885 ( .A1(n6799), .A2(n9989), .ZN(n10000) );
  INV_X1 U7886 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7045) );
  AND2_X1 U7887 ( .A1(n10000), .A2(n7045), .ZN(n6801) );
  INV_X1 U7888 ( .A(n6800), .ZN(n8356) );
  AND2_X1 U7889 ( .A1(n8356), .A2(n8231), .ZN(n7044) );
  OAI22_X1 U7890 ( .A1(n6801), .A2(n7044), .B1(n9989), .B2(n7045), .ZN(
        P1_U3441) );
  OAI222_X1 U7891 ( .A1(n6848), .A2(P1_U3084), .B1(n7481), .B2(n6803), .C1(
        n6802), .C2(n8841), .ZN(P1_U3351) );
  OAI222_X1 U7892 ( .A1(n6806), .A2(P1_U3084), .B1(n7481), .B2(n6805), .C1(
        n6804), .C2(n8841), .ZN(P1_U3350) );
  OAI222_X1 U7893 ( .A1(n6850), .A2(P1_U3084), .B1(n7481), .B2(n6808), .C1(
        n6807), .C2(n8841), .ZN(P1_U3349) );
  INV_X1 U7894 ( .A(n6809), .ZN(n6812) );
  OAI222_X1 U7895 ( .A1(n9503), .A2(n6810), .B1(n7477), .B2(n6812), .C1(
        P2_U3152), .C2(n6975), .ZN(P2_U3351) );
  INV_X1 U7896 ( .A(n6888), .ZN(n6854) );
  INV_X1 U7897 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6811) );
  OAI222_X1 U7898 ( .A1(n6854), .A2(P1_U3084), .B1(n7481), .B2(n6812), .C1(
        n6811), .C2(n8841), .ZN(P1_U3346) );
  NAND2_X1 U7899 ( .A1(n9665), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6813) );
  OAI21_X1 U7900 ( .B1(n9723), .B2(n9665), .A(n6813), .ZN(P1_U3585) );
  INV_X1 U7901 ( .A(n6912), .ZN(n6856) );
  INV_X1 U7902 ( .A(n6814), .ZN(n6816) );
  OAI222_X1 U7903 ( .A1(n6856), .A2(P1_U3084), .B1(n7481), .B2(n6816), .C1(
        n6815), .C2(n8841), .ZN(P1_U3345) );
  INV_X1 U7904 ( .A(n7004), .ZN(n6978) );
  OAI222_X1 U7905 ( .A1(n9503), .A2(n6828), .B1(n7477), .B2(n6816), .C1(
        P2_U3152), .C2(n6978), .ZN(P2_U3350) );
  INV_X1 U7906 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U7907 ( .A1(n6817), .A2(P1_U4006), .ZN(n6818) );
  OAI21_X1 U7908 ( .B1(P1_U4006), .B2(n6819), .A(n6818), .ZN(P1_U3586) );
  INV_X1 U7909 ( .A(n6820), .ZN(n6823) );
  AOI22_X1 U7910 ( .A1(n7082), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n7289), .ZN(n6821) );
  OAI21_X1 U7911 ( .B1(n6823), .B2(n7477), .A(n6821), .ZN(P2_U3349) );
  INV_X1 U7912 ( .A(n7211), .ZN(n6905) );
  OAI222_X1 U7913 ( .A1(P1_U3084), .A2(n6905), .B1(n7481), .B2(n6823), .C1(
        n6822), .C2(n8841), .ZN(P1_U3344) );
  INV_X1 U7914 ( .A(n6824), .ZN(n6832) );
  AOI22_X1 U7915 ( .A1(n7197), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n7289), .ZN(n6825) );
  OAI21_X1 U7916 ( .B1(n6832), .B2(n7477), .A(n6825), .ZN(P2_U3348) );
  MUX2_X1 U7917 ( .A(n6826), .B(n7835), .S(P1_U4006), .Z(n6827) );
  INV_X1 U7918 ( .A(n6827), .ZN(P1_U3565) );
  MUX2_X1 U7919 ( .A(n6828), .B(n7826), .S(P1_U4006), .Z(n6829) );
  INV_X1 U7920 ( .A(n6829), .ZN(P1_U3563) );
  MUX2_X1 U7921 ( .A(n6844), .B(n8196), .S(P1_U4006), .Z(n6830) );
  INV_X1 U7922 ( .A(n6830), .ZN(P1_U3567) );
  OAI222_X1 U7923 ( .A1(P1_U3084), .A2(n10290), .B1(n7481), .B2(n6832), .C1(
        n6831), .C2(n8841), .ZN(P1_U3343) );
  INV_X1 U7924 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6834) );
  INV_X1 U7925 ( .A(n6833), .ZN(n6835) );
  OAI222_X1 U7926 ( .A1(n8841), .A2(n6834), .B1(n7481), .B2(n6835), .C1(
        P1_U3084), .C2(n7215), .ZN(P1_U3342) );
  INV_X1 U7927 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6836) );
  INV_X1 U7928 ( .A(n7364), .ZN(n7205) );
  OAI222_X1 U7929 ( .A1(n9503), .A2(n6836), .B1(n7477), .B2(n6835), .C1(n7205), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7930 ( .A(n9116), .ZN(n10379) );
  NOR2_X1 U7931 ( .A1(n10379), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7932 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U7933 ( .A1(n5436), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6839) );
  INV_X1 U7934 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6837) );
  OR2_X1 U7935 ( .A1(n5454), .A2(n6837), .ZN(n6838) );
  OAI211_X1 U7936 ( .C1(n4846), .C2(n8837), .A(n6839), .B(n6838), .ZN(n8752)
         );
  NAND2_X1 U7937 ( .A1(n8752), .A2(P2_U3966), .ZN(n6840) );
  OAI21_X1 U7938 ( .B1(n9993), .B2(P2_U3966), .A(n6840), .ZN(P2_U3583) );
  INV_X1 U7939 ( .A(n6841), .ZN(n6843) );
  AOI22_X1 U7940 ( .A1(n10302), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7287), .ZN(n6842) );
  OAI21_X1 U7941 ( .B1(n6843), .B2(n7481), .A(n6842), .ZN(P1_U3341) );
  INV_X1 U7942 ( .A(n7458), .ZN(n7465) );
  OAI222_X1 U7943 ( .A1(n9503), .A2(n6844), .B1(n7477), .B2(n6843), .C1(
        P2_U3152), .C2(n7465), .ZN(P2_U3346) );
  NOR2_X1 U7944 ( .A1(n6888), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U7945 ( .A1(n10271), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6853) );
  MUX2_X1 U7946 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6845), .S(n10271), .Z(n10277) );
  NOR2_X1 U7947 ( .A1(n10428), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U7948 ( .A1(n10340), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6849) );
  MUX2_X1 U7949 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6846), .S(n10340), .Z(n10346) );
  XNOR2_X1 U7950 ( .A(n6848), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10409) );
  INV_X1 U7951 ( .A(n6864), .ZN(n6895) );
  MUX2_X1 U7952 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6847), .S(n6895), .Z(n6897)
         );
  NAND3_X1 U7953 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n6897), .ZN(n6896) );
  OAI21_X1 U7954 ( .B1(n6864), .B2(n6847), .A(n6896), .ZN(n10408) );
  NAND2_X1 U7955 ( .A1(n10409), .A2(n10408), .ZN(n10406) );
  OAI21_X1 U7956 ( .B1(n6848), .B2(n6375), .A(n10406), .ZN(n10347) );
  NAND2_X1 U7957 ( .A1(n10346), .A2(n10347), .ZN(n10345) );
  NAND2_X1 U7958 ( .A1(n6849), .A2(n10345), .ZN(n10431) );
  AOI22_X1 U7959 ( .A1(n10428), .A2(n6399), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n6850), .ZN(n10430) );
  NOR2_X1 U7960 ( .A1(n10431), .A2(n10430), .ZN(n10429) );
  NOR2_X1 U7961 ( .A1(n6851), .A2(n10429), .ZN(n10335) );
  MUX2_X1 U7962 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6852), .S(n10328), .Z(n10334) );
  NAND2_X1 U7963 ( .A1(n10335), .A2(n10334), .ZN(n10333) );
  OAI21_X1 U7964 ( .B1(n6863), .B2(n6852), .A(n10333), .ZN(n10278) );
  NAND2_X1 U7965 ( .A1(n10277), .A2(n10278), .ZN(n10276) );
  NAND2_X1 U7966 ( .A1(n6853), .A2(n10276), .ZN(n6880) );
  AOI22_X1 U7967 ( .A1(n6888), .A2(n6345), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n6854), .ZN(n6879) );
  NOR2_X1 U7968 ( .A1(n6880), .A2(n6879), .ZN(n6878) );
  NOR2_X1 U7969 ( .A1(n6855), .A2(n6878), .ZN(n6858) );
  AOI22_X1 U7970 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6856), .B1(n6912), .B2(
        n6332), .ZN(n6857) );
  NOR2_X1 U7971 ( .A1(n6858), .A2(n6857), .ZN(n6903) );
  AOI21_X1 U7972 ( .B1(n6858), .B2(n6857), .A(n6903), .ZN(n6877) );
  OR2_X1 U7973 ( .A1(n6859), .A2(P1_U3084), .ZN(n10264) );
  INV_X1 U7974 ( .A(n4848), .ZN(n10263) );
  OR2_X1 U7975 ( .A1(n4847), .A2(n10263), .ZN(n6860) );
  OR2_X1 U7976 ( .A1(n10264), .A2(n6860), .ZN(n10433) );
  NOR2_X1 U7977 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6912), .ZN(n6861) );
  AOI21_X1 U7978 ( .B1(n6912), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6861), .ZN(
        n6870) );
  NAND2_X1 U7979 ( .A1(n10271), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6862) );
  OAI21_X1 U7980 ( .B1(n10271), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6862), .ZN(
        n10274) );
  AOI22_X1 U7981 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10328), .B1(n6863), .B2(
        n6413), .ZN(n10330) );
  NAND2_X1 U7982 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10399) );
  INV_X1 U7983 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7351) );
  MUX2_X1 U7984 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7351), .S(n6864), .Z(n6893)
         );
  NOR2_X1 U7985 ( .A1(n10399), .A2(n6893), .ZN(n6892) );
  AOI21_X1 U7986 ( .B1(n6895), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6892), .ZN(
        n10414) );
  NAND2_X1 U7987 ( .A1(n10417), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6865) );
  OAI21_X1 U7988 ( .B1(n10417), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6865), .ZN(
        n10413) );
  NOR2_X1 U7989 ( .A1(n10414), .A2(n10413), .ZN(n10412) );
  AOI21_X1 U7990 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n10417), .A(n10412), .ZN(
        n10342) );
  NAND2_X1 U7991 ( .A1(n10340), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6866) );
  OAI21_X1 U7992 ( .B1(n10340), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6866), .ZN(
        n10343) );
  NOR2_X1 U7993 ( .A1(n10342), .A2(n10343), .ZN(n10341) );
  AOI21_X1 U7994 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n10340), .A(n10341), .ZN(
        n10424) );
  NOR2_X1 U7995 ( .A1(n10428), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6867) );
  AOI21_X1 U7996 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n10428), .A(n6867), .ZN(
        n10423) );
  NAND2_X1 U7997 ( .A1(n10424), .A2(n10423), .ZN(n10422) );
  OAI21_X1 U7998 ( .B1(n10428), .B2(P1_REG2_REG_4__SCAN_IN), .A(n10422), .ZN(
        n10331) );
  NAND2_X1 U7999 ( .A1(n10330), .A2(n10331), .ZN(n10329) );
  OAI21_X1 U8000 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n10328), .A(n10329), .ZN(
        n10273) );
  NOR2_X1 U8001 ( .A1(n10274), .A2(n10273), .ZN(n10272) );
  AOI21_X1 U8002 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n10271), .A(n10272), .ZN(
        n6883) );
  NOR2_X1 U8003 ( .A1(n6888), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6868) );
  AOI21_X1 U8004 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6888), .A(n6868), .ZN(
        n6882) );
  NAND2_X1 U8005 ( .A1(n6883), .A2(n6882), .ZN(n6881) );
  OAI21_X1 U8006 ( .B1(n6888), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6881), .ZN(
        n6869) );
  NAND2_X1 U8007 ( .A1(n6870), .A2(n6869), .ZN(n6911) );
  OAI21_X1 U8008 ( .B1(n6870), .B2(n6869), .A(n6911), .ZN(n6871) );
  NOR2_X1 U8009 ( .A1(n10264), .A2(n4848), .ZN(n7217) );
  INV_X1 U8010 ( .A(n4847), .ZN(n10402) );
  NAND2_X1 U8011 ( .A1(n7217), .A2(n10402), .ZN(n10411) );
  INV_X1 U8012 ( .A(n10411), .ZN(n10426) );
  NAND2_X1 U8013 ( .A1(n6871), .A2(n10426), .ZN(n6876) );
  NAND2_X1 U8014 ( .A1(n7217), .A2(n4847), .ZN(n10318) );
  INV_X1 U8015 ( .A(n10318), .ZN(n10427) );
  INV_X1 U8016 ( .A(n6872), .ZN(n6873) );
  OR2_X1 U8017 ( .A1(P1_U3083), .A2(n6873), .ZN(n10420) );
  INV_X1 U8018 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U8019 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7848) );
  OAI21_X1 U8020 ( .B1(n10420), .B2(n8013), .A(n7848), .ZN(n6874) );
  AOI21_X1 U8021 ( .B1(n10427), .B2(n6912), .A(n6874), .ZN(n6875) );
  OAI211_X1 U8022 ( .C1(n6877), .C2(n10433), .A(n6876), .B(n6875), .ZN(
        P1_U3249) );
  AOI21_X1 U8023 ( .B1(n6880), .B2(n6879), .A(n6878), .ZN(n6891) );
  OAI21_X1 U8024 ( .B1(n6883), .B2(n6882), .A(n6881), .ZN(n6884) );
  NAND2_X1 U8025 ( .A1(n6884), .A2(n10426), .ZN(n6890) );
  INV_X1 U8026 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8009) );
  NOR2_X1 U8027 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6885), .ZN(n7645) );
  INV_X1 U8028 ( .A(n7645), .ZN(n6886) );
  OAI21_X1 U8029 ( .B1(n10420), .B2(n8009), .A(n6886), .ZN(n6887) );
  AOI21_X1 U8030 ( .B1(n10427), .B2(n6888), .A(n6887), .ZN(n6889) );
  OAI211_X1 U8031 ( .C1(n6891), .C2(n10433), .A(n6890), .B(n6889), .ZN(
        P1_U3248) );
  AOI211_X1 U8032 ( .C1(n10399), .C2(n6893), .A(n6892), .B(n10411), .ZN(n6894)
         );
  AOI21_X1 U8033 ( .B1(n10427), .B2(n6895), .A(n6894), .ZN(n6902) );
  INV_X1 U8034 ( .A(n10420), .ZN(n10436) );
  INV_X1 U8035 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7348) );
  INV_X1 U8036 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7189) );
  NOR2_X1 U8037 ( .A1(n6371), .A2(n7189), .ZN(n6898) );
  INV_X1 U8038 ( .A(n10433), .ZN(n10407) );
  OAI211_X1 U8039 ( .C1(n6898), .C2(n6897), .A(n6896), .B(n10407), .ZN(n6899)
         );
  OAI21_X1 U8040 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7348), .A(n6899), .ZN(n6900) );
  AOI21_X1 U8041 ( .B1(n10436), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n6900), .ZN(
        n6901) );
  NAND2_X1 U8042 ( .A1(n6902), .A2(n6901), .ZN(P1_U3242) );
  NOR2_X1 U8043 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6912), .ZN(n6904) );
  NOR2_X1 U8044 ( .A1(n6904), .A2(n6903), .ZN(n6907) );
  AOI22_X1 U8045 ( .A1(n7211), .A2(n6293), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6905), .ZN(n6906) );
  NOR2_X1 U8046 ( .A1(n6907), .A2(n6906), .ZN(n7207) );
  AOI21_X1 U8047 ( .B1(n6907), .B2(n6906), .A(n7207), .ZN(n6919) );
  INV_X1 U8048 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6910) );
  NOR2_X1 U8049 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6908), .ZN(n7836) );
  INV_X1 U8050 ( .A(n7836), .ZN(n6909) );
  OAI21_X1 U8051 ( .B1(n10420), .B2(n6910), .A(n6909), .ZN(n6917) );
  OAI21_X1 U8052 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6912), .A(n6911), .ZN(
        n6915) );
  NAND2_X1 U8053 ( .A1(n7211), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6913) );
  OAI21_X1 U8054 ( .B1(n7211), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6913), .ZN(
        n6914) );
  NOR2_X1 U8055 ( .A1(n6914), .A2(n6915), .ZN(n7210) );
  AOI211_X1 U8056 ( .C1(n6915), .C2(n6914), .A(n7210), .B(n10411), .ZN(n6916)
         );
  AOI211_X1 U8057 ( .C1(n10427), .C2(n7211), .A(n6917), .B(n6916), .ZN(n6918)
         );
  OAI21_X1 U8058 ( .B1(n6919), .B2(n10433), .A(n6918), .ZN(P1_U3250) );
  INV_X1 U8059 ( .A(n6920), .ZN(n6923) );
  AOI22_X1 U8060 ( .A1(n10316), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7287), .ZN(n6921) );
  OAI21_X1 U8061 ( .B1(n6923), .B2(n7481), .A(n6921), .ZN(P1_U3340) );
  NAND2_X1 U8062 ( .A1(n9275), .A2(P2_U3966), .ZN(n6922) );
  OAI21_X1 U8063 ( .B1(n6136), .B2(P2_U3966), .A(n6922), .ZN(P2_U3573) );
  INV_X1 U8064 ( .A(n7618), .ZN(n7475) );
  OAI222_X1 U8065 ( .A1(n9503), .A2(n6924), .B1(n7477), .B2(n6923), .C1(n7475), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  AOI21_X1 U8066 ( .B1(n6926), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6925), .ZN(
        n6928) );
  XOR2_X1 U8067 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6953), .Z(n6927) );
  NOR2_X1 U8068 ( .A1(n6927), .A2(n6928), .ZN(n6943) );
  AOI211_X1 U8069 ( .C1(n6928), .C2(n6927), .A(n6943), .B(n10357), .ZN(n6931)
         );
  INV_X1 U8070 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U8071 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7451) );
  OAI21_X1 U8072 ( .B1(n9116), .B2(n6929), .A(n7451), .ZN(n6930) );
  NOR2_X1 U8073 ( .A1(n6931), .A2(n6930), .ZN(n6938) );
  XNOR2_X1 U8074 ( .A(n6953), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6936) );
  INV_X1 U8075 ( .A(n6932), .ZN(n6933) );
  OAI21_X1 U8076 ( .B1(n6934), .B2(n7761), .A(n6933), .ZN(n6935) );
  INV_X1 U8077 ( .A(n10394), .ZN(n10359) );
  NAND2_X1 U8078 ( .A1(n6936), .A2(n6935), .ZN(n6951) );
  OAI211_X1 U8079 ( .C1(n6936), .C2(n6935), .A(n10359), .B(n6951), .ZN(n6937)
         );
  OAI211_X1 U8080 ( .C1(n10356), .C2(n6953), .A(n6938), .B(n6937), .ZN(
        P2_U3249) );
  INV_X1 U8081 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6940) );
  INV_X1 U8082 ( .A(n6939), .ZN(n6941) );
  INV_X1 U8083 ( .A(n7676), .ZN(n7418) );
  OAI222_X1 U8084 ( .A1(n8841), .A2(n6940), .B1(n7481), .B2(n6941), .C1(
        P1_U3084), .C2(n7418), .ZN(P1_U3339) );
  INV_X1 U8085 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6942) );
  INV_X1 U8086 ( .A(n7888), .ZN(n7622) );
  OAI222_X1 U8087 ( .A1(n9503), .A2(n6942), .B1(n7477), .B2(n6941), .C1(n7622), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8088 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10236) );
  XNOR2_X1 U8089 ( .A(n6983), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n6948) );
  INV_X1 U8090 ( .A(n6943), .ZN(n6944) );
  OAI21_X1 U8091 ( .B1(n6953), .B2(n6945), .A(n6944), .ZN(n6959) );
  MUX2_X1 U8092 ( .A(n6946), .B(P2_REG1_REG_5__SCAN_IN), .S(n6968), .Z(n6960)
         );
  NAND2_X1 U8093 ( .A1(n6959), .A2(n6960), .ZN(n6958) );
  OAI21_X1 U8094 ( .B1(n6968), .B2(n6946), .A(n6958), .ZN(n6947) );
  INV_X1 U8095 ( .A(n10357), .ZN(n10391) );
  NAND2_X1 U8096 ( .A1(n6947), .A2(n6948), .ZN(n6971) );
  OAI211_X1 U8097 ( .C1(n6948), .C2(n6947), .A(n10391), .B(n6971), .ZN(n6949)
         );
  NAND2_X1 U8098 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7517) );
  OAI211_X1 U8099 ( .C1(n9116), .C2(n10236), .A(n6949), .B(n7517), .ZN(n6950)
         );
  INV_X1 U8100 ( .A(n6950), .ZN(n6957) );
  XNOR2_X1 U8101 ( .A(n6983), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6955) );
  OAI21_X1 U8102 ( .B1(n6953), .B2(n6952), .A(n6951), .ZN(n6964) );
  INV_X1 U8103 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7721) );
  MUX2_X1 U8104 ( .A(n7721), .B(P2_REG2_REG_5__SCAN_IN), .S(n6968), .Z(n6965)
         );
  NAND2_X1 U8105 ( .A1(n6964), .A2(n6965), .ZN(n6963) );
  OAI21_X1 U8106 ( .B1(n6968), .B2(n7721), .A(n6963), .ZN(n6954) );
  NAND2_X1 U8107 ( .A1(n6954), .A2(n6955), .ZN(n6984) );
  OAI211_X1 U8108 ( .C1(n6955), .C2(n6954), .A(n10359), .B(n6984), .ZN(n6956)
         );
  OAI211_X1 U8109 ( .C1(n10356), .C2(n6983), .A(n6957), .B(n6956), .ZN(
        P2_U3251) );
  INV_X1 U8110 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10234) );
  OAI211_X1 U8111 ( .C1(n6960), .C2(n6959), .A(n10391), .B(n6958), .ZN(n6961)
         );
  NAND2_X1 U8112 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7378) );
  OAI211_X1 U8113 ( .C1(n9116), .C2(n10234), .A(n6961), .B(n7378), .ZN(n6962)
         );
  INV_X1 U8114 ( .A(n6962), .ZN(n6967) );
  OAI211_X1 U8115 ( .C1(n6965), .C2(n6964), .A(n10359), .B(n6963), .ZN(n6966)
         );
  OAI211_X1 U8116 ( .C1(n10356), .C2(n6968), .A(n6967), .B(n6966), .ZN(
        P2_U3250) );
  NAND2_X1 U8117 ( .A1(n9219), .A2(P2_U3966), .ZN(n6969) );
  OAI21_X1 U8118 ( .B1(n6171), .B2(P2_U3966), .A(n6969), .ZN(P2_U3574) );
  NAND2_X1 U8119 ( .A1(n9819), .A2(P1_U4006), .ZN(n6970) );
  OAI21_X1 U8120 ( .B1(P1_U4006), .B2(n7920), .A(n6970), .ZN(P1_U3578) );
  INV_X1 U8121 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10242) );
  INV_X1 U8122 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10533) );
  MUX2_X1 U8123 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10533), .S(n7082), .Z(n6980)
         );
  OAI21_X1 U8124 ( .B1(n6972), .B2(n6983), .A(n6971), .ZN(n7007) );
  NAND2_X1 U8125 ( .A1(n7016), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6973) );
  OAI21_X1 U8126 ( .B1(n7016), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6973), .ZN(
        n6974) );
  INV_X1 U8127 ( .A(n6974), .ZN(n7008) );
  NAND2_X1 U8128 ( .A1(n7007), .A2(n7008), .ZN(n7006) );
  OAI21_X1 U8129 ( .B1(n6976), .B2(n6975), .A(n7006), .ZN(n6995) );
  MUX2_X1 U8130 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6977), .S(n7004), .Z(n6996)
         );
  NAND2_X1 U8131 ( .A1(n6995), .A2(n6996), .ZN(n6994) );
  OAI21_X1 U8132 ( .B1(n6978), .B2(n6977), .A(n6994), .ZN(n6979) );
  NAND2_X1 U8133 ( .A1(n6979), .A2(n6980), .ZN(n7080) );
  OAI211_X1 U8134 ( .C1(n6980), .C2(n6979), .A(n10391), .B(n7080), .ZN(n6982)
         );
  NAND2_X1 U8135 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6981) );
  OAI211_X1 U8136 ( .C1(n9116), .C2(n10242), .A(n6982), .B(n6981), .ZN(n6992)
         );
  INV_X1 U8137 ( .A(n6983), .ZN(n6986) );
  INV_X1 U8138 ( .A(n6984), .ZN(n6985) );
  AOI21_X1 U8139 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6986), .A(n6985), .ZN(
        n7013) );
  NAND2_X1 U8140 ( .A1(n7016), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6987) );
  OAI21_X1 U8141 ( .B1(n7016), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6987), .ZN(
        n7012) );
  NOR2_X1 U8142 ( .A1(n7013), .A2(n7012), .ZN(n7011) );
  AOI21_X1 U8143 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7016), .A(n7011), .ZN(
        n7001) );
  XNOR2_X1 U8144 ( .A(n7004), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7000) );
  NOR2_X1 U8145 ( .A1(n7001), .A2(n7000), .ZN(n6999) );
  AOI21_X1 U8146 ( .B1(n7004), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6999), .ZN(
        n6990) );
  NAND2_X1 U8147 ( .A1(n7082), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6988) );
  OAI21_X1 U8148 ( .B1(n7082), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6988), .ZN(
        n6989) );
  NOR2_X1 U8149 ( .A1(n6990), .A2(n6989), .ZN(n7076) );
  AOI211_X1 U8150 ( .C1(n6990), .C2(n6989), .A(n10394), .B(n7076), .ZN(n6991)
         );
  AOI211_X1 U8151 ( .C1(n10386), .C2(n7082), .A(n6992), .B(n6991), .ZN(n6993)
         );
  INV_X1 U8152 ( .A(n6993), .ZN(P2_U3254) );
  INV_X1 U8153 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10240) );
  OAI211_X1 U8154 ( .C1(n6996), .C2(n6995), .A(n10391), .B(n6994), .ZN(n6998)
         );
  NAND2_X1 U8155 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6997) );
  OAI211_X1 U8156 ( .C1(n9116), .C2(n10240), .A(n6998), .B(n6997), .ZN(n7003)
         );
  AOI211_X1 U8157 ( .C1(n7001), .C2(n7000), .A(n6999), .B(n10394), .ZN(n7002)
         );
  AOI211_X1 U8158 ( .C1(n10386), .C2(n7004), .A(n7003), .B(n7002), .ZN(n7005)
         );
  INV_X1 U8159 ( .A(n7005), .ZN(P2_U3253) );
  INV_X1 U8160 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10238) );
  OAI211_X1 U8161 ( .C1(n7008), .C2(n7007), .A(n10391), .B(n7006), .ZN(n7010)
         );
  NAND2_X1 U8162 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n7009) );
  OAI211_X1 U8163 ( .C1(n9116), .C2(n10238), .A(n7010), .B(n7009), .ZN(n7015)
         );
  AOI211_X1 U8164 ( .C1(n7013), .C2(n7012), .A(n7011), .B(n10394), .ZN(n7014)
         );
  AOI211_X1 U8165 ( .C1(n10386), .C2(n7016), .A(n7015), .B(n7014), .ZN(n7017)
         );
  INV_X1 U8166 ( .A(n7017), .ZN(P2_U3252) );
  NAND2_X1 U8167 ( .A1(n7136), .A2(n9834), .ZN(n7482) );
  NAND2_X2 U8168 ( .A1(n7019), .A2(n7018), .ZN(n7138) );
  AND2_X4 U8169 ( .A1(n7138), .A2(n7114), .ZN(n8936) );
  NAND2_X1 U8170 ( .A1(n7482), .A2(n8936), .ZN(n7039) );
  OR2_X2 U8171 ( .A1(n7138), .A2(n7021), .ZN(n7096) );
  INV_X4 U8172 ( .A(n7096), .ZN(n8898) );
  AOI22_X1 U8173 ( .A1(n8898), .A2(n7127), .B1(n7021), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n7020) );
  AND2_X1 U8174 ( .A1(n7026), .A2(n7023), .ZN(n7025) );
  NAND2_X1 U8175 ( .A1(n7025), .A2(n7024), .ZN(n7028) );
  NAND2_X2 U8176 ( .A1(n7028), .A2(n7027), .ZN(n8698) );
  INV_X1 U8177 ( .A(n8698), .ZN(n7029) );
  NAND2_X1 U8178 ( .A1(n7030), .A2(n9834), .ZN(n7031) );
  INV_X4 U8179 ( .A(n8939), .ZN(n8947) );
  NAND2_X1 U8180 ( .A1(n8698), .A2(n8947), .ZN(n7032) );
  NAND2_X1 U8181 ( .A1(n8695), .A2(n7032), .ZN(n7037) );
  NAND2_X1 U8182 ( .A1(n7129), .A2(n8898), .ZN(n7034) );
  NAND2_X1 U8183 ( .A1(n7354), .A2(n8936), .ZN(n7033) );
  NAND2_X1 U8184 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  XNOR2_X1 U8185 ( .A(n7035), .B(n4840), .ZN(n7036) );
  NOR2_X2 U8186 ( .A1(n7037), .A2(n7036), .ZN(n7106) );
  NAND2_X1 U8187 ( .A1(n7037), .A2(n7036), .ZN(n7104) );
  INV_X1 U8188 ( .A(n7104), .ZN(n7038) );
  NOR2_X1 U8189 ( .A1(n7106), .A2(n7038), .ZN(n7040) );
  INV_X1 U8190 ( .A(n7129), .ZN(n8699) );
  INV_X1 U8191 ( .A(n7039), .ZN(n7243) );
  INV_X1 U8192 ( .A(n7243), .ZN(n8195) );
  OAI22_X1 U8193 ( .A1(n8699), .A2(n8195), .B1(n10459), .B2(n8949), .ZN(n7105)
         );
  XNOR2_X1 U8194 ( .A(n7040), .B(n7105), .ZN(n7075) );
  AND2_X1 U8195 ( .A1(n7063), .A2(n7042), .ZN(n9959) );
  NAND2_X1 U8196 ( .A1(n7110), .A2(n9989), .ZN(n7043) );
  NOR2_X1 U8197 ( .A1(n9964), .A2(n7043), .ZN(n7061) );
  AOI21_X1 U8198 ( .B1(n7057), .B2(n7045), .A(n7044), .ZN(n7153) );
  NOR2_X1 U8199 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n7049) );
  NOR4_X1 U8200 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n7048) );
  NOR4_X1 U8201 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n7047) );
  NOR4_X1 U8202 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n7046) );
  NAND4_X1 U8203 ( .A1(n7049), .A2(n7048), .A3(n7047), .A4(n7046), .ZN(n7055)
         );
  NOR4_X1 U8204 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n7053) );
  NOR4_X1 U8205 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n7052) );
  NOR4_X1 U8206 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n7051) );
  NOR4_X1 U8207 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n7050) );
  NAND4_X1 U8208 ( .A1(n7053), .A2(n7052), .A3(n7051), .A4(n7050), .ZN(n7054)
         );
  OAI21_X1 U8209 ( .B1(n7055), .B2(n7054), .A(n7057), .ZN(n7150) );
  NAND2_X1 U8210 ( .A1(n7153), .A2(n7150), .ZN(n7292) );
  INV_X1 U8211 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7056) );
  NAND2_X1 U8212 ( .A1(n7057), .A2(n7056), .ZN(n7059) );
  NAND2_X1 U8213 ( .A1(n8356), .A2(n8105), .ZN(n7058) );
  NAND2_X1 U8214 ( .A1(n7059), .A2(n7058), .ZN(n7180) );
  OR2_X1 U8215 ( .A1(n7292), .A2(n7180), .ZN(n7067) );
  INV_X1 U8216 ( .A(n7067), .ZN(n7060) );
  NAND2_X1 U8217 ( .A1(n7061), .A2(n7060), .ZN(n9649) );
  NOR2_X1 U8218 ( .A1(n7067), .A2(n7062), .ZN(n7070) );
  AND2_X1 U8219 ( .A1(n7070), .A2(n10402), .ZN(n9641) );
  OR2_X1 U8220 ( .A1(n7041), .A2(n7018), .ZN(n7310) );
  OR2_X1 U8221 ( .A1(n7310), .A2(n7064), .ZN(n7065) );
  OR2_X1 U8222 ( .A1(n7041), .A2(n7126), .ZN(n7151) );
  AOI22_X1 U8223 ( .A1(n9641), .A2(n7128), .B1(n7354), .B2(n4839), .ZN(n7074)
         );
  NAND2_X1 U8224 ( .A1(n10537), .A2(n7067), .ZN(n7111) );
  INV_X1 U8225 ( .A(n7111), .ZN(n7069) );
  NAND2_X1 U8226 ( .A1(n7182), .A2(n7310), .ZN(n7066) );
  AND3_X1 U8227 ( .A1(n7067), .A2(n9989), .A3(n7066), .ZN(n7117) );
  INV_X1 U8228 ( .A(n7110), .ZN(n7140) );
  NAND2_X1 U8229 ( .A1(n7182), .A2(n7140), .ZN(n7068) );
  NAND2_X1 U8230 ( .A1(n7068), .A2(n9989), .ZN(n7293) );
  NOR3_X1 U8231 ( .A1(n7069), .A2(n7117), .A3(n7293), .ZN(n7162) );
  INV_X1 U8232 ( .A(n7162), .ZN(n8701) );
  INV_X1 U8233 ( .A(n7070), .ZN(n7071) );
  OR2_X1 U8234 ( .A1(n7071), .A2(n10402), .ZN(n9623) );
  AOI22_X1 U8235 ( .A1(n8701), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9642), .B2(
        n9664), .ZN(n7073) );
  OAI211_X1 U8236 ( .C1(n7075), .C2(n9649), .A(n7074), .B(n7073), .ZN(P1_U3220) );
  AOI21_X1 U8237 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7082), .A(n7076), .ZN(
        n7079) );
  MUX2_X1 U8238 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8130), .S(n7197), .Z(n7077)
         );
  INV_X1 U8239 ( .A(n7077), .ZN(n7078) );
  NOR2_X1 U8240 ( .A1(n7079), .A2(n7078), .ZN(n7190) );
  AOI211_X1 U8241 ( .C1(n7079), .C2(n7078), .A(n7190), .B(n10394), .ZN(n7091)
         );
  INV_X1 U8242 ( .A(n7080), .ZN(n7081) );
  AOI21_X1 U8243 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7082), .A(n7081), .ZN(
        n7085) );
  MUX2_X1 U8244 ( .A(n7083), .B(P2_REG1_REG_10__SCAN_IN), .S(n7197), .Z(n7084)
         );
  NOR2_X1 U8245 ( .A1(n7085), .A2(n7084), .ZN(n7196) );
  AOI211_X1 U8246 ( .C1(n7085), .C2(n7084), .A(n7196), .B(n10357), .ZN(n7090)
         );
  INV_X1 U8247 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7088) );
  NAND2_X1 U8248 ( .A1(n10386), .A2(n7197), .ZN(n7087) );
  NAND2_X1 U8249 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7086) );
  OAI211_X1 U8250 ( .C1(n9116), .C2(n7088), .A(n7087), .B(n7086), .ZN(n7089)
         );
  OR3_X1 U8251 ( .A1(n7091), .A2(n7090), .A3(n7089), .ZN(P2_U3255) );
  AOI22_X1 U8252 ( .A1(n7243), .A2(n7092), .B1(n8898), .B2(n7296), .ZN(n7248)
         );
  NAND2_X1 U8253 ( .A1(n7092), .A2(n8898), .ZN(n7094) );
  OR2_X1 U8254 ( .A1(n7508), .A2(n8950), .ZN(n7093) );
  NAND2_X1 U8255 ( .A1(n7094), .A2(n7093), .ZN(n7095) );
  XNOR2_X1 U8256 ( .A(n7248), .B(n7247), .ZN(n7109) );
  OR2_X1 U8257 ( .A1(n7161), .A2(n8950), .ZN(n7098) );
  NAND2_X1 U8258 ( .A1(n9664), .A2(n8943), .ZN(n7097) );
  NAND2_X1 U8259 ( .A1(n7098), .A2(n7097), .ZN(n7099) );
  NOR2_X1 U8260 ( .A1(n7161), .A2(n7096), .ZN(n7100) );
  AOI21_X1 U8261 ( .B1(n7243), .B2(n9664), .A(n7100), .ZN(n7101) );
  NAND2_X1 U8262 ( .A1(n7102), .A2(n7101), .ZN(n7107) );
  AND2_X1 U8263 ( .A1(n7103), .A2(n7107), .ZN(n7160) );
  OAI21_X1 U8264 ( .B1(n7106), .B2(n7105), .A(n7104), .ZN(n7159) );
  NAND2_X1 U8265 ( .A1(n7160), .A2(n7159), .ZN(n7158) );
  NAND2_X1 U8266 ( .A1(n7158), .A2(n7107), .ZN(n7108) );
  OAI21_X1 U8267 ( .B1(n7109), .B2(n7108), .A(n7251), .ZN(n7123) );
  INV_X1 U8268 ( .A(n9649), .ZN(n9604) );
  NAND2_X1 U8269 ( .A1(n7111), .A2(n7110), .ZN(n7112) );
  NAND2_X1 U8270 ( .A1(n7112), .A2(n7182), .ZN(n7116) );
  AND2_X1 U8271 ( .A1(n7114), .A2(n7113), .ZN(n7115) );
  NAND2_X1 U8272 ( .A1(n7116), .A2(n7115), .ZN(n7118) );
  AOI21_X2 U8273 ( .B1(n7118), .B2(P1_STATE_REG_SCAN_IN), .A(n7117), .ZN(n9646) );
  NAND2_X1 U8274 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10350) );
  INV_X1 U8275 ( .A(n10350), .ZN(n7119) );
  AOI21_X1 U8276 ( .B1(n4839), .B2(n7296), .A(n7119), .ZN(n7121) );
  AOI22_X1 U8277 ( .A1(n9642), .A2(n9663), .B1(n9641), .B2(n9664), .ZN(n7120)
         );
  OAI211_X1 U8278 ( .C1(n9646), .C2(P1_REG3_REG_3__SCAN_IN), .A(n7121), .B(
        n7120), .ZN(n7122) );
  AOI21_X1 U8279 ( .B1(n7123), .B2(n9604), .A(n7122), .ZN(n7124) );
  INV_X1 U8280 ( .A(n7124), .ZN(P1_U3216) );
  INV_X1 U8281 ( .A(n7126), .ZN(n7294) );
  NAND2_X1 U8282 ( .A1(n7125), .A2(n7294), .ZN(n8182) );
  INV_X1 U8283 ( .A(n8182), .ZN(n10463) );
  NAND2_X1 U8284 ( .A1(n7129), .A2(n7354), .ZN(n7130) );
  NAND2_X1 U8285 ( .A1(n7134), .A2(n7133), .ZN(n7271) );
  OAI21_X1 U8286 ( .B1(n7134), .B2(n7133), .A(n7271), .ZN(n7149) );
  NAND2_X1 U8287 ( .A1(n10459), .A2(n10441), .ZN(n7347) );
  INV_X1 U8288 ( .A(n7347), .ZN(n7135) );
  OAI21_X1 U8289 ( .B1(n7135), .B2(n7161), .A(n7278), .ZN(n7497) );
  INV_X1 U8290 ( .A(n7136), .ZN(n7137) );
  INV_X1 U8291 ( .A(n7137), .ZN(n9965) );
  OAI22_X1 U8292 ( .A1(n7497), .A2(n7137), .B1(n7161), .B2(n10537), .ZN(n7148)
         );
  INV_X1 U8293 ( .A(n7149), .ZN(n7499) );
  AOI21_X1 U8294 ( .B1(n7125), .B2(n7138), .A(n7541), .ZN(n7139) );
  NAND2_X1 U8295 ( .A1(n7182), .A2(n7139), .ZN(n7661) );
  AOI22_X1 U8296 ( .A1(n9866), .A2(n7092), .B1(n7129), .B2(n9864), .ZN(n7147)
         );
  OAI21_X1 U8297 ( .B1(n7142), .B2(n6670), .A(n7141), .ZN(n7145) );
  NAND2_X1 U8298 ( .A1(n7030), .A2(n7541), .ZN(n7144) );
  NAND2_X1 U8299 ( .A1(n7019), .A2(n6668), .ZN(n7143) );
  NAND2_X1 U8300 ( .A1(n7144), .A2(n7143), .ZN(n9869) );
  NAND2_X1 U8301 ( .A1(n7145), .A2(n9869), .ZN(n7146) );
  OAI211_X1 U8302 ( .C1(n7499), .C2(n7661), .A(n7147), .B(n7146), .ZN(n7494)
         );
  AOI211_X1 U8303 ( .C1(n10463), .C2(n7149), .A(n7148), .B(n7494), .ZN(n7229)
         );
  NAND2_X1 U8304 ( .A1(n7151), .A2(n7150), .ZN(n7152) );
  NAND2_X1 U8305 ( .A1(n10542), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7154) );
  OAI21_X1 U8306 ( .B1(n7229), .B2(n10542), .A(n7154), .ZN(P1_U3525) );
  INV_X1 U8307 ( .A(n6237), .ZN(n7156) );
  OAI222_X1 U8308 ( .A1(n8841), .A2(n7155), .B1(n7481), .B2(n7156), .C1(n7797), 
        .C2(P1_U3084), .ZN(P1_U3338) );
  INV_X1 U8309 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7157) );
  OAI222_X1 U8310 ( .A1(n9503), .A2(n7157), .B1(n7477), .B2(n7156), .C1(
        P2_U3152), .C2(n8162), .ZN(P2_U3343) );
  OAI21_X1 U8311 ( .B1(n7160), .B2(n7159), .A(n7158), .ZN(n7165) );
  INV_X1 U8312 ( .A(n9641), .ZN(n9607) );
  INV_X1 U8313 ( .A(n4839), .ZN(n9613) );
  OAI22_X1 U8314 ( .A1(n9607), .A2(n8699), .B1(n7161), .B2(n9613), .ZN(n7164)
         );
  INV_X1 U8315 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7495) );
  INV_X1 U8316 ( .A(n7092), .ZN(n7316) );
  OAI22_X1 U8317 ( .A1(n7162), .A2(n7495), .B1(n7316), .B2(n9623), .ZN(n7163)
         );
  AOI211_X1 U8318 ( .C1(n7165), .C2(n9604), .A(n7164), .B(n7163), .ZN(n7166)
         );
  INV_X1 U8319 ( .A(n7166), .ZN(P1_U3235) );
  INV_X1 U8320 ( .A(n7167), .ZN(n7170) );
  NAND3_X1 U8321 ( .A1(n7170), .A2(n7168), .A3(n7169), .ZN(n7171) );
  AND2_X1 U8322 ( .A1(n7172), .A2(n7171), .ZN(n7178) );
  INV_X1 U8323 ( .A(n9059), .ZN(n9022) );
  INV_X1 U8324 ( .A(n7578), .ZN(n9101) );
  AOI22_X1 U8325 ( .A1(n9039), .A2(n9103), .B1(n9022), .B2(n9101), .ZN(n7177)
         );
  INV_X1 U8326 ( .A(n7385), .ZN(n7408) );
  OR2_X1 U8327 ( .A1(n7173), .A2(n7408), .ZN(n7175) );
  AND2_X1 U8328 ( .A1(n7384), .A2(n10355), .ZN(n7174) );
  NAND2_X1 U8329 ( .A1(n7175), .A2(n7174), .ZN(n7258) );
  AOI22_X1 U8330 ( .A1(n9079), .A2(n7769), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n7258), .ZN(n7176) );
  OAI211_X1 U8331 ( .C1(n7178), .C2(n9081), .A(n7177), .B(n7176), .ZN(P2_U3239) );
  INV_X1 U8332 ( .A(n9186), .ZN(n9218) );
  NAND2_X1 U8333 ( .A1(n9218), .A2(P2_U3966), .ZN(n7179) );
  OAI21_X1 U8334 ( .B1(n6469), .B2(P2_U3966), .A(n7179), .ZN(P2_U3576) );
  INV_X1 U8335 ( .A(n7180), .ZN(n9990) );
  NAND2_X1 U8336 ( .A1(n7182), .A2(n7041), .ZN(n7183) );
  INV_X1 U8337 ( .A(n9866), .ZN(n9784) );
  OAI22_X1 U8338 ( .A1(n7184), .A2(n7183), .B1(n8699), .B2(n9784), .ZN(n10446)
         );
  INV_X1 U8339 ( .A(n10446), .ZN(n7185) );
  OAI21_X1 U8340 ( .B1(n10441), .B2(n7041), .A(n7185), .ZN(n7187) );
  NAND2_X1 U8341 ( .A1(n7187), .A2(n4843), .ZN(n7186) );
  OAI21_X1 U8342 ( .B1(n4843), .B2(n6364), .A(n7186), .ZN(P1_U3454) );
  NAND2_X1 U8343 ( .A1(n7187), .A2(n4842), .ZN(n7188) );
  OAI21_X1 U8344 ( .B1(n4842), .B2(n7189), .A(n7188), .ZN(P1_U3523) );
  AOI21_X1 U8345 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7197), .A(n7190), .ZN(
        n7193) );
  NOR2_X1 U8346 ( .A1(n7364), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7191) );
  AOI21_X1 U8347 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7364), .A(n7191), .ZN(
        n7192) );
  NAND2_X1 U8348 ( .A1(n7193), .A2(n7192), .ZN(n7363) );
  OAI21_X1 U8349 ( .B1(n7193), .B2(n7192), .A(n7363), .ZN(n7194) );
  NAND2_X1 U8350 ( .A1(n7194), .A2(n10359), .ZN(n7204) );
  INV_X1 U8351 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7195) );
  MUX2_X1 U8352 ( .A(n7195), .B(P2_REG1_REG_11__SCAN_IN), .S(n7364), .Z(n7199)
         );
  AOI21_X1 U8353 ( .B1(n7197), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7196), .ZN(
        n7198) );
  NOR2_X1 U8354 ( .A1(n7198), .A2(n7199), .ZN(n7357) );
  AOI21_X1 U8355 ( .B1(n7199), .B2(n7198), .A(n7357), .ZN(n7202) );
  INV_X1 U8356 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7200) );
  NAND2_X1 U8357 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7991) );
  OAI21_X1 U8358 ( .B1(n9116), .B2(n7200), .A(n7991), .ZN(n7201) );
  AOI21_X1 U8359 ( .B1(n10391), .B2(n7202), .A(n7201), .ZN(n7203) );
  OAI211_X1 U8360 ( .C1(n10356), .C2(n7205), .A(n7204), .B(n7203), .ZN(
        P2_U3256) );
  NOR2_X1 U8361 ( .A1(n7211), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7206) );
  NOR2_X1 U8362 ( .A1(n7207), .A2(n7206), .ZN(n10294) );
  MUX2_X1 U8363 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7208), .S(n10290), .Z(
        n10293) );
  NOR2_X1 U8364 ( .A1(n10294), .A2(n10293), .ZN(n10292) );
  AOI21_X1 U8365 ( .B1(n10290), .B2(n7208), .A(n10292), .ZN(n7421) );
  NOR2_X1 U8366 ( .A1(n7215), .A2(n6267), .ZN(n7422) );
  AOI21_X1 U8367 ( .B1(n7215), .B2(n6267), .A(n7422), .ZN(n7209) );
  XNOR2_X1 U8368 ( .A(n7421), .B(n7209), .ZN(n7228) );
  INV_X1 U8369 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7221) );
  INV_X1 U8370 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7864) );
  OR2_X1 U8371 ( .A1(n10290), .A2(n7864), .ZN(n7213) );
  AOI21_X1 U8372 ( .B1(n7211), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7210), .ZN(
        n10283) );
  MUX2_X1 U8373 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7864), .S(n10290), .Z(
        n10284) );
  NOR2_X1 U8374 ( .A1(n10283), .A2(n10284), .ZN(n10286) );
  INV_X1 U8375 ( .A(n10286), .ZN(n7212) );
  OR2_X1 U8376 ( .A1(n7215), .A2(n7214), .ZN(n7222) );
  NOR2_X1 U8377 ( .A1(n7224), .A2(n7222), .ZN(n7216) );
  NAND2_X1 U8378 ( .A1(n7217), .A2(n7216), .ZN(n7220) );
  NOR2_X1 U8379 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7218), .ZN(n8096) );
  INV_X1 U8380 ( .A(n8096), .ZN(n7219) );
  OAI211_X1 U8381 ( .C1(n10420), .C2(n7221), .A(n7220), .B(n7219), .ZN(n7226)
         );
  NOR2_X1 U8382 ( .A1(n7423), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7223) );
  OAI21_X1 U8383 ( .B1(n7223), .B2(n7224), .A(n7222), .ZN(n10309) );
  AOI211_X1 U8384 ( .C1(n7224), .C2(n7223), .A(n10309), .B(n10411), .ZN(n7225)
         );
  AOI211_X1 U8385 ( .C1(n10427), .C2(n7423), .A(n7226), .B(n7225), .ZN(n7227)
         );
  OAI21_X1 U8386 ( .B1(n7228), .B2(n10433), .A(n7227), .ZN(P1_U3252) );
  OR2_X1 U8387 ( .A1(n7229), .A2(n10543), .ZN(n7230) );
  OAI21_X1 U8388 ( .B1(n4843), .B2(n6377), .A(n7230), .ZN(P1_U3460) );
  INV_X1 U8389 ( .A(n7231), .ZN(n7234) );
  INV_X1 U8390 ( .A(n9110), .ZN(n8160) );
  OAI222_X1 U8391 ( .A1(n9503), .A2(n7232), .B1(n7477), .B2(n7234), .C1(
        P2_U3152), .C2(n8160), .ZN(P2_U3342) );
  INV_X1 U8392 ( .A(n9675), .ZN(n7804) );
  OAI222_X1 U8393 ( .A1(n7804), .A2(P1_U3084), .B1(n7481), .B2(n7234), .C1(
        n7233), .C2(n8841), .ZN(P1_U3337) );
  INV_X1 U8394 ( .A(n9076), .ZN(n7990) );
  OR2_X1 U8395 ( .A1(n7751), .A2(n9341), .ZN(n7236) );
  NAND2_X1 U8396 ( .A1(n9105), .A2(n9388), .ZN(n7235) );
  NAND2_X1 U8397 ( .A1(n7236), .A2(n7235), .ZN(n10466) );
  AOI22_X1 U8398 ( .A1(n7990), .A2(n10466), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n7258), .ZN(n7241) );
  OAI21_X1 U8399 ( .B1(n7238), .B2(n7237), .A(n7168), .ZN(n7239) );
  NAND2_X1 U8400 ( .A1(n9009), .A2(n7239), .ZN(n7240) );
  OAI211_X1 U8401 ( .C1(n10481), .C2(n9016), .A(n7241), .B(n7240), .ZN(
        P2_U3224) );
  NOR2_X1 U8402 ( .A1(n7486), .A2(n8949), .ZN(n7242) );
  AOI21_X1 U8403 ( .B1(n7243), .B2(n9663), .A(n7242), .ZN(n7432) );
  NAND2_X1 U8404 ( .A1(n9663), .A2(n8943), .ZN(n7245) );
  INV_X1 U8405 ( .A(n7486), .ZN(n7326) );
  NAND2_X1 U8406 ( .A1(n7326), .A2(n8936), .ZN(n7244) );
  NAND2_X1 U8407 ( .A1(n7245), .A2(n7244), .ZN(n7246) );
  XNOR2_X1 U8408 ( .A(n7246), .B(n8947), .ZN(n7434) );
  XOR2_X1 U8409 ( .A(n7432), .B(n7434), .Z(n7253) );
  INV_X1 U8410 ( .A(n7247), .ZN(n7249) );
  NAND2_X1 U8411 ( .A1(n7249), .A2(n7248), .ZN(n7250) );
  AOI211_X1 U8412 ( .C1(n7253), .C2(n7252), .A(n9649), .B(n4926), .ZN(n7257)
         );
  AND2_X1 U8413 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10435) );
  AOI21_X1 U8414 ( .B1(n4839), .B2(n7326), .A(n10435), .ZN(n7255) );
  AOI22_X1 U8415 ( .A1(n9642), .A2(n9662), .B1(n9641), .B2(n7092), .ZN(n7254)
         );
  OAI211_X1 U8416 ( .C1(n9646), .C2(n7484), .A(n7255), .B(n7254), .ZN(n7256)
         );
  OR2_X1 U8417 ( .A1(n7257), .A2(n7256), .ZN(P1_U3228) );
  NAND2_X1 U8418 ( .A1(n7258), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7263) );
  NAND2_X1 U8419 ( .A1(n9105), .A2(n7743), .ZN(n7259) );
  NAND2_X1 U8420 ( .A1(n7259), .A2(n10470), .ZN(n7260) );
  NAND3_X1 U8421 ( .A1(n9009), .A2(n7261), .A3(n7260), .ZN(n7262) );
  OAI211_X1 U8422 ( .C1(n9016), .C2(n10470), .A(n7263), .B(n7262), .ZN(n7264)
         );
  AOI21_X1 U8423 ( .B1(n9022), .B2(n9103), .A(n7264), .ZN(n7265) );
  INV_X1 U8424 ( .A(n7265), .ZN(P2_U3234) );
  INV_X1 U8425 ( .A(n7266), .ZN(n7269) );
  AOI22_X1 U8426 ( .A1(n9124), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n7289), .ZN(n7267) );
  OAI21_X1 U8427 ( .B1(n7269), .B2(n7477), .A(n7267), .ZN(P2_U3341) );
  AOI22_X1 U8428 ( .A1(n9687), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7287), .ZN(n7268) );
  OAI21_X1 U8429 ( .B1(n7269), .B2(n7481), .A(n7268), .ZN(P1_U3336) );
  INV_X1 U8430 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7282) );
  OR2_X1 U8431 ( .A1(n7072), .A2(n6386), .ZN(n7270) );
  NAND2_X1 U8432 ( .A1(n7271), .A2(n7270), .ZN(n7272) );
  NAND2_X1 U8433 ( .A1(n7272), .A2(n7273), .ZN(n7298) );
  OAI21_X1 U8434 ( .B1(n7272), .B2(n7273), .A(n7298), .ZN(n7510) );
  INV_X1 U8435 ( .A(n7510), .ZN(n7280) );
  INV_X1 U8436 ( .A(n7661), .ZN(n8457) );
  INV_X1 U8437 ( .A(n9864), .ZN(n9782) );
  INV_X1 U8438 ( .A(n9663), .ZN(n7442) );
  OAI22_X1 U8439 ( .A1(n6387), .A2(n9782), .B1(n7442), .B2(n9784), .ZN(n7277)
         );
  XNOR2_X1 U8440 ( .A(n7274), .B(n7273), .ZN(n7275) );
  INV_X1 U8441 ( .A(n9869), .ZN(n9780) );
  NOR2_X1 U8442 ( .A1(n7275), .A2(n9780), .ZN(n7276) );
  AOI211_X1 U8443 ( .C1(n8457), .C2(n7510), .A(n7277), .B(n7276), .ZN(n7512)
         );
  AOI21_X1 U8444 ( .B1(n7296), .B2(n7278), .A(n7322), .ZN(n7504) );
  AOI22_X1 U8445 ( .A1(n7504), .A2(n9965), .B1(n9964), .B2(n7296), .ZN(n7279)
         );
  OAI211_X1 U8446 ( .C1(n7280), .C2(n8182), .A(n7512), .B(n7279), .ZN(n7283)
         );
  NAND2_X1 U8447 ( .A1(n7283), .A2(n4843), .ZN(n7281) );
  OAI21_X1 U8448 ( .B1(n4843), .B2(n7282), .A(n7281), .ZN(P1_U3463) );
  NAND2_X1 U8449 ( .A1(n7283), .A2(n4842), .ZN(n7284) );
  OAI21_X1 U8450 ( .B1(n4842), .B2(n6846), .A(n7284), .ZN(P1_U3526) );
  NAND2_X1 U8451 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n9104), .ZN(n7285) );
  OAI21_X1 U8452 ( .B1(n8866), .B2(n9104), .A(n7285), .ZN(P2_U3581) );
  INV_X1 U8453 ( .A(n7286), .ZN(n7291) );
  AOI22_X1 U8454 ( .A1(n9699), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7287), .ZN(n7288) );
  OAI21_X1 U8455 ( .B1(n7291), .B2(n7481), .A(n7288), .ZN(P1_U3335) );
  AOI22_X1 U8456 ( .A1(n9122), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7289), .ZN(n7290) );
  OAI21_X1 U8457 ( .B1(n7291), .B2(n7477), .A(n7290), .ZN(P2_U3340) );
  NAND2_X2 U8458 ( .A1(n7542), .A2(n10450), .ZN(n10447) );
  NAND2_X1 U8459 ( .A1(n7294), .A2(n7019), .ZN(n7353) );
  NAND2_X1 U8460 ( .A1(n7661), .A2(n7353), .ZN(n7295) );
  AND2_X1 U8461 ( .A1(n10447), .A2(n7295), .ZN(n9734) );
  OR2_X1 U8462 ( .A1(n7092), .A2(n7296), .ZN(n7297) );
  NAND2_X1 U8463 ( .A1(n7315), .A2(n7318), .ZN(n7314) );
  OR2_X1 U8464 ( .A1(n9663), .A2(n7326), .ZN(n7299) );
  NAND2_X1 U8465 ( .A1(n7314), .A2(n7299), .ZN(n7302) );
  INV_X1 U8466 ( .A(n7302), .ZN(n7300) );
  INV_X1 U8467 ( .A(n7301), .ZN(n7304) );
  NAND2_X1 U8468 ( .A1(n7302), .A2(n7301), .ZN(n7303) );
  NAND2_X1 U8469 ( .A1(n7531), .A2(n7303), .ZN(n10495) );
  XNOR2_X1 U8470 ( .A(n7525), .B(n7304), .ZN(n7305) );
  NAND2_X1 U8471 ( .A1(n7305), .A2(n9869), .ZN(n7307) );
  AOI22_X1 U8472 ( .A1(n9864), .A2(n9663), .B1(n9661), .B2(n9866), .ZN(n7306)
         );
  NAND2_X1 U8473 ( .A1(n7307), .A2(n7306), .ZN(n10500) );
  NAND2_X1 U8474 ( .A1(n7322), .A2(n7486), .ZN(n7323) );
  AOI21_X1 U8475 ( .B1(n7323), .B2(n7529), .A(n7137), .ZN(n7308) );
  NAND2_X1 U8476 ( .A1(n7308), .A2(n5321), .ZN(n10496) );
  OAI22_X1 U8477 ( .A1(n10496), .A2(n7541), .B1(n10450), .B2(n7443), .ZN(n7309) );
  OAI21_X1 U8478 ( .B1(n10500), .B2(n7309), .A(n10447), .ZN(n7313) );
  INV_X1 U8479 ( .A(n7310), .ZN(n7311) );
  INV_X2 U8480 ( .A(n10447), .ZN(n9843) );
  AOI22_X1 U8481 ( .A1(n9827), .A2(n7529), .B1(n9843), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n7312) );
  OAI211_X1 U8482 ( .C1(n9873), .C2(n10495), .A(n7313), .B(n7312), .ZN(
        P1_U3286) );
  INV_X1 U8483 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7330) );
  OAI21_X1 U8484 ( .B1(n7315), .B2(n7318), .A(n7314), .ZN(n7490) );
  INV_X1 U8485 ( .A(n7490), .ZN(n7328) );
  INV_X1 U8486 ( .A(n9662), .ZN(n7561) );
  OAI22_X1 U8487 ( .A1(n7316), .A2(n9782), .B1(n7561), .B2(n9784), .ZN(n7321)
         );
  XNOR2_X1 U8488 ( .A(n7317), .B(n7318), .ZN(n7319) );
  NOR2_X1 U8489 ( .A1(n7319), .A2(n9780), .ZN(n7320) );
  AOI211_X1 U8490 ( .C1(n8457), .C2(n7490), .A(n7321), .B(n7320), .ZN(n7493)
         );
  INV_X1 U8491 ( .A(n7322), .ZN(n7325) );
  INV_X1 U8492 ( .A(n7323), .ZN(n7324) );
  AOI21_X1 U8493 ( .B1(n7326), .B2(n7325), .A(n7324), .ZN(n7489) );
  AOI22_X1 U8494 ( .A1(n7489), .A2(n9965), .B1(n9964), .B2(n7326), .ZN(n7327)
         );
  OAI211_X1 U8495 ( .C1(n7328), .C2(n8182), .A(n7493), .B(n7327), .ZN(n7331)
         );
  NAND2_X1 U8496 ( .A1(n7331), .A2(n4843), .ZN(n7329) );
  OAI21_X1 U8497 ( .B1(n4843), .B2(n7330), .A(n7329), .ZN(P1_U3466) );
  NAND2_X1 U8498 ( .A1(n7331), .A2(n4842), .ZN(n7332) );
  OAI21_X1 U8499 ( .B1(n4842), .B2(n6399), .A(n7332), .ZN(P1_U3527) );
  INV_X1 U8500 ( .A(n7374), .ZN(n7333) );
  AOI211_X1 U8501 ( .C1(n7335), .C2(n7334), .A(n9081), .B(n7333), .ZN(n7339)
         );
  AOI22_X1 U8502 ( .A1(n9039), .A2(n9102), .B1(n9022), .B2(n9100), .ZN(n7337)
         );
  INV_X1 U8503 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7759) );
  MUX2_X1 U8504 ( .A(P2_STATE_REG_SCAN_IN), .B(n9019), .S(n7759), .Z(n7336) );
  OAI211_X1 U8505 ( .C1(n7573), .C2(n9016), .A(n7337), .B(n7336), .ZN(n7338)
         );
  OR2_X1 U8506 ( .A1(n7339), .A2(n7338), .ZN(P2_U3220) );
  XNOR2_X1 U8507 ( .A(n7340), .B(n6553), .ZN(n7352) );
  OAI21_X1 U8508 ( .B1(n7342), .B2(n6553), .A(n7341), .ZN(n7345) );
  OAI22_X1 U8509 ( .A1(n7343), .A2(n9782), .B1(n6387), .B2(n9784), .ZN(n7344)
         );
  AOI21_X1 U8510 ( .B1(n7345), .B2(n9869), .A(n7344), .ZN(n7346) );
  OAI21_X1 U8511 ( .B1(n7352), .B2(n7661), .A(n7346), .ZN(n10460) );
  OAI211_X1 U8512 ( .C1(n10459), .C2(n10441), .A(n9965), .B(n7347), .ZN(n10458) );
  OAI22_X1 U8513 ( .A1(n10458), .A2(n7541), .B1(n7348), .B2(n10450), .ZN(n7349) );
  NOR2_X1 U8514 ( .A1(n10460), .A2(n7349), .ZN(n7350) );
  MUX2_X1 U8515 ( .A(n7351), .B(n7350), .S(n10447), .Z(n7356) );
  INV_X1 U8516 ( .A(n7352), .ZN(n10462) );
  NOR2_X1 U8517 ( .A1(n9843), .A2(n7353), .ZN(n10014) );
  AOI22_X1 U8518 ( .A1(n10462), .A2(n10014), .B1(n9827), .B2(n7354), .ZN(n7355) );
  NAND2_X1 U8519 ( .A1(n7356), .A2(n7355), .ZN(P1_U3290) );
  INV_X1 U8520 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7362) );
  AOI21_X1 U8521 ( .B1(n7364), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7357), .ZN(
        n7359) );
  MUX2_X1 U8522 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7464), .S(n7458), .Z(n7358)
         );
  NAND2_X1 U8523 ( .A1(n7359), .A2(n7358), .ZN(n7467) );
  OAI21_X1 U8524 ( .B1(n7359), .B2(n7358), .A(n7467), .ZN(n7360) );
  NAND2_X1 U8525 ( .A1(n10391), .A2(n7360), .ZN(n7361) );
  NAND2_X1 U8526 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8147) );
  OAI211_X1 U8527 ( .C1(n9116), .C2(n7362), .A(n7361), .B(n8147), .ZN(n7368)
         );
  OAI21_X1 U8528 ( .B1(n7364), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7363), .ZN(
        n7366) );
  XNOR2_X1 U8529 ( .A(n7458), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7365) );
  NOR2_X1 U8530 ( .A1(n7366), .A2(n7365), .ZN(n7457) );
  AOI211_X1 U8531 ( .C1(n7366), .C2(n7365), .A(n10394), .B(n7457), .ZN(n7367)
         );
  AOI211_X1 U8532 ( .C1(n10386), .C2(n7458), .A(n7368), .B(n7367), .ZN(n7369)
         );
  INV_X1 U8533 ( .A(n7369), .ZN(P2_U3257) );
  INV_X1 U8534 ( .A(n7370), .ZN(n7371) );
  NOR2_X1 U8535 ( .A1(n7372), .A2(n7371), .ZN(n7377) );
  AND2_X1 U8536 ( .A1(n7374), .A2(n7373), .ZN(n7450) );
  NAND2_X1 U8537 ( .A1(n7450), .A2(n7449), .ZN(n7448) );
  INV_X1 U8538 ( .A(n7375), .ZN(n7376) );
  AOI21_X1 U8539 ( .B1(n7377), .B2(n7448), .A(n7376), .ZN(n7382) );
  OAI21_X1 U8540 ( .B1(n9019), .B2(n7714), .A(n7378), .ZN(n7380) );
  OAI22_X1 U8541 ( .A1(n7750), .A2(n9062), .B1(n9059), .B2(n7933), .ZN(n7379)
         );
  AOI211_X1 U8542 ( .C1(n7718), .C2(n9079), .A(n7380), .B(n7379), .ZN(n7381)
         );
  OAI21_X1 U8543 ( .B1(n7382), .B2(n9081), .A(n7381), .ZN(P2_U3229) );
  AND3_X1 U8544 ( .A1(n7384), .A2(n10355), .A3(n7383), .ZN(n7701) );
  AND2_X1 U8545 ( .A1(n7701), .A2(n7698), .ZN(n7410) );
  AND2_X1 U8546 ( .A1(n7699), .A2(n7385), .ZN(n7386) );
  AND2_X2 U8547 ( .A1(n7410), .A2(n7386), .ZN(n10584) );
  INV_X1 U8548 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7407) );
  INV_X1 U8549 ( .A(n10575), .ZN(n10566) );
  INV_X1 U8550 ( .A(n5364), .ZN(n8687) );
  NAND2_X1 U8551 ( .A1(n8687), .A2(n8521), .ZN(n8510) );
  NAND2_X1 U8552 ( .A1(n9180), .A2(n8691), .ZN(n8684) );
  NAND2_X1 U8553 ( .A1(n8510), .A2(n8684), .ZN(n10467) );
  NAND2_X1 U8554 ( .A1(n7390), .A2(n7392), .ZN(n8654) );
  INV_X1 U8555 ( .A(n9105), .ZN(n7387) );
  NAND2_X1 U8556 ( .A1(n7387), .A2(n7745), .ZN(n10465) );
  NAND2_X1 U8557 ( .A1(n8654), .A2(n10465), .ZN(n7388) );
  NAND2_X1 U8558 ( .A1(n7751), .A2(n7769), .ZN(n8527) );
  OAI21_X1 U8559 ( .B1(n7389), .B2(n8655), .A(n7565), .ZN(n7404) );
  OAI22_X1 U8560 ( .A1(n7390), .A2(n9343), .B1(n7578), .B2(n9341), .ZN(n7403)
         );
  INV_X1 U8561 ( .A(n7391), .ZN(n10474) );
  NAND2_X1 U8562 ( .A1(n9103), .A2(n7392), .ZN(n7393) );
  INV_X1 U8563 ( .A(n7397), .ZN(n7396) );
  NAND2_X1 U8564 ( .A1(n7396), .A2(n7395), .ZN(n7571) );
  NAND2_X1 U8565 ( .A1(n8655), .A2(n7397), .ZN(n7401) );
  INV_X1 U8566 ( .A(n7398), .ZN(n7399) );
  AOI21_X1 U8567 ( .B1(n7571), .B2(n7401), .A(n10564), .ZN(n7402) );
  AOI211_X1 U8568 ( .C1(n10467), .C2(n7404), .A(n7403), .B(n7402), .ZN(n7771)
         );
  INV_X1 U8569 ( .A(n10568), .ZN(n10576) );
  NAND2_X1 U8570 ( .A1(n10469), .A2(n7769), .ZN(n7764) );
  NAND3_X1 U8571 ( .A1(n4850), .A2(n10576), .A3(n7764), .ZN(n7405) );
  OAI211_X1 U8572 ( .C1(n7570), .C2(n10566), .A(n7771), .B(n7405), .ZN(n7411)
         );
  NAND2_X1 U8573 ( .A1(n7411), .A2(n10584), .ZN(n7406) );
  OAI21_X1 U8574 ( .B1(n10584), .B2(n7407), .A(n7406), .ZN(P2_U3522) );
  NOR2_X1 U8575 ( .A1(n7699), .A2(n7408), .ZN(n7409) );
  AND2_X2 U8576 ( .A1(n7410), .A2(n7409), .ZN(n10588) );
  NAND2_X1 U8577 ( .A1(n7411), .A2(n10588), .ZN(n7412) );
  OAI21_X1 U8578 ( .B1(n10588), .B2(n5453), .A(n7412), .ZN(P2_U3457) );
  NOR2_X1 U8579 ( .A1(n7418), .A2(n8325), .ZN(n7673) );
  AOI21_X1 U8580 ( .B1(n8325), .B2(n7418), .A(n7673), .ZN(n7417) );
  NAND2_X1 U8581 ( .A1(n10316), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7416) );
  MUX2_X1 U8582 ( .A(n6311), .B(P1_REG2_REG_13__SCAN_IN), .S(n10316), .Z(n7413) );
  INV_X1 U8583 ( .A(n7413), .ZN(n10323) );
  NAND2_X1 U8584 ( .A1(n10302), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7415) );
  MUX2_X1 U8585 ( .A(n8054), .B(P1_REG2_REG_12__SCAN_IN), .S(n10302), .Z(n7414) );
  INV_X1 U8586 ( .A(n7414), .ZN(n10308) );
  NAND2_X1 U8587 ( .A1(n10308), .A2(n10309), .ZN(n10307) );
  NAND2_X1 U8588 ( .A1(n7415), .A2(n10307), .ZN(n10324) );
  NAND2_X1 U8589 ( .A1(n10323), .A2(n10324), .ZN(n10322) );
  NAND2_X1 U8590 ( .A1(n7416), .A2(n10322), .ZN(n7674) );
  XOR2_X1 U8591 ( .A(n7417), .B(n7674), .Z(n7430) );
  NOR2_X1 U8592 ( .A1(n10318), .A2(n7418), .ZN(n7429) );
  INV_X1 U8593 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7427) );
  XNOR2_X1 U8594 ( .A(n7676), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7678) );
  XNOR2_X1 U8595 ( .A(n10316), .B(n7419), .ZN(n10315) );
  MUX2_X1 U8596 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7420), .S(n10302), .Z(
        n10301) );
  OAI22_X1 U8597 ( .A1(n7423), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n7422), .B2(
        n7421), .ZN(n10300) );
  NAND2_X1 U8598 ( .A1(n10301), .A2(n10300), .ZN(n10299) );
  OAI21_X1 U8599 ( .B1(n10302), .B2(P1_REG1_REG_12__SCAN_IN), .A(n10299), .ZN(
        n10314) );
  NAND2_X1 U8600 ( .A1(n10315), .A2(n10314), .ZN(n10313) );
  OAI21_X1 U8601 ( .B1(n10316), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10313), .ZN(
        n7424) );
  INV_X1 U8602 ( .A(n7424), .ZN(n7677) );
  XNOR2_X1 U8603 ( .A(n7678), .B(n7677), .ZN(n7425) );
  NAND2_X1 U8604 ( .A1(n10407), .A2(n7425), .ZN(n7426) );
  NAND2_X1 U8605 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9523) );
  OAI211_X1 U8606 ( .C1(n10420), .C2(n7427), .A(n7426), .B(n9523), .ZN(n7428)
         );
  AOI211_X1 U8607 ( .C1(n7430), .C2(n10426), .A(n7429), .B(n7428), .ZN(n7431)
         );
  INV_X1 U8608 ( .A(n7431), .ZN(P1_U3255) );
  INV_X1 U8609 ( .A(n7432), .ZN(n7433) );
  AOI22_X1 U8610 ( .A1(n7529), .A2(n8936), .B1(n9662), .B2(n8898), .ZN(n7435)
         );
  XNOR2_X1 U8611 ( .A(n7435), .B(n8947), .ZN(n7436) );
  NOR2_X1 U8612 ( .A1(n7437), .A2(n7436), .ZN(n7555) );
  NAND2_X1 U8613 ( .A1(n7437), .A2(n7436), .ZN(n7553) );
  INV_X1 U8614 ( .A(n7553), .ZN(n7438) );
  NOR2_X1 U8615 ( .A1(n7555), .A2(n7438), .ZN(n7439) );
  INV_X1 U8616 ( .A(n7243), .ZN(n8236) );
  OAI22_X1 U8617 ( .A1(n7561), .A2(n8236), .B1(n10497), .B2(n7096), .ZN(n7554)
         );
  XNOR2_X1 U8618 ( .A(n7439), .B(n7554), .ZN(n7447) );
  NAND2_X1 U8619 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10338) );
  INV_X1 U8620 ( .A(n10338), .ZN(n7440) );
  AOI21_X1 U8621 ( .B1(n9642), .B2(n9661), .A(n7440), .ZN(n7441) );
  OAI21_X1 U8622 ( .B1(n7442), .B2(n9607), .A(n7441), .ZN(n7445) );
  NOR2_X1 U8623 ( .A1(n9646), .A2(n7443), .ZN(n7444) );
  AOI211_X1 U8624 ( .C1(n7529), .C2(n4839), .A(n7445), .B(n7444), .ZN(n7446)
         );
  OAI21_X1 U8625 ( .B1(n7447), .B2(n9649), .A(n7446), .ZN(P1_U3225) );
  OAI21_X1 U8626 ( .B1(n7450), .B2(n7449), .A(n7448), .ZN(n7455) );
  NAND2_X1 U8627 ( .A1(n9079), .A2(n7778), .ZN(n7452) );
  OAI211_X1 U8628 ( .C1(n9019), .C2(n7776), .A(n7452), .B(n7451), .ZN(n7454)
         );
  OAI22_X1 U8629 ( .A1(n7972), .A2(n9059), .B1(n9062), .B2(n7578), .ZN(n7453)
         );
  AOI211_X1 U8630 ( .C1(n7455), .C2(n9009), .A(n7454), .B(n7453), .ZN(n7456)
         );
  INV_X1 U8631 ( .A(n7456), .ZN(P2_U3232) );
  AOI21_X1 U8632 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7458), .A(n7457), .ZN(
        n7461) );
  NOR2_X1 U8633 ( .A1(n7618), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7459) );
  AOI21_X1 U8634 ( .B1(n7618), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7459), .ZN(
        n7460) );
  NAND2_X1 U8635 ( .A1(n7461), .A2(n7460), .ZN(n7613) );
  OAI21_X1 U8636 ( .B1(n7461), .B2(n7460), .A(n7613), .ZN(n7462) );
  NAND2_X1 U8637 ( .A1(n7462), .A2(n10359), .ZN(n7474) );
  MUX2_X1 U8638 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n7463), .S(n7618), .Z(n7469)
         );
  NAND2_X1 U8639 ( .A1(n7465), .A2(n7464), .ZN(n7466) );
  NAND2_X1 U8640 ( .A1(n7467), .A2(n7466), .ZN(n7468) );
  NAND2_X1 U8641 ( .A1(n7468), .A2(n7469), .ZN(n7617) );
  OAI21_X1 U8642 ( .B1(n7469), .B2(n7468), .A(n7617), .ZN(n7472) );
  INV_X1 U8643 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7470) );
  NAND2_X1 U8644 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8221) );
  OAI21_X1 U8645 ( .B1(n9116), .B2(n7470), .A(n8221), .ZN(n7471) );
  AOI21_X1 U8646 ( .B1(n10391), .B2(n7472), .A(n7471), .ZN(n7473) );
  OAI211_X1 U8647 ( .C1(n10356), .C2(n7475), .A(n7474), .B(n7473), .ZN(
        P2_U3258) );
  INV_X1 U8648 ( .A(n7476), .ZN(n7480) );
  OAI222_X1 U8649 ( .A1(n9503), .A2(n7478), .B1(n7477), .B2(n7480), .C1(n9143), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8650 ( .A1(n9834), .A2(P1_U3084), .B1(n7481), .B2(n7480), .C1(
        n7479), .C2(n8841), .ZN(P1_U3334) );
  INV_X1 U8651 ( .A(n7482), .ZN(n7483) );
  OAI22_X1 U8652 ( .A1(n10447), .A2(n7485), .B1(n7484), .B2(n10450), .ZN(n7488) );
  NOR2_X1 U8653 ( .A1(n10442), .A2(n7486), .ZN(n7487) );
  AOI211_X1 U8654 ( .C1(n7489), .C2(n10006), .A(n7488), .B(n7487), .ZN(n7492)
         );
  NAND2_X1 U8655 ( .A1(n7490), .A2(n10014), .ZN(n7491) );
  OAI211_X1 U8656 ( .C1(n7493), .C2(n9843), .A(n7492), .B(n7491), .ZN(P1_U3287) );
  INV_X1 U8657 ( .A(n7494), .ZN(n7503) );
  INV_X1 U8658 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7496) );
  OAI22_X1 U8659 ( .A1(n10447), .A2(n7496), .B1(n7495), .B2(n10450), .ZN(n7501) );
  INV_X1 U8660 ( .A(n10014), .ZN(n7498) );
  INV_X1 U8661 ( .A(n10006), .ZN(n10443) );
  OAI22_X1 U8662 ( .A1(n7499), .A2(n7498), .B1(n10443), .B2(n7497), .ZN(n7500)
         );
  AOI211_X1 U8663 ( .C1(n9827), .C2(n6386), .A(n7501), .B(n7500), .ZN(n7502)
         );
  OAI21_X1 U8664 ( .B1(n9843), .B2(n7503), .A(n7502), .ZN(P1_U3289) );
  NAND2_X1 U8665 ( .A1(n7504), .A2(n10006), .ZN(n7507) );
  NOR2_X1 U8666 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(n10450), .ZN(n7505) );
  AOI21_X1 U8667 ( .B1(n9843), .B2(P1_REG2_REG_3__SCAN_IN), .A(n7505), .ZN(
        n7506) );
  OAI211_X1 U8668 ( .C1(n7508), .C2(n10442), .A(n7507), .B(n7506), .ZN(n7509)
         );
  AOI21_X1 U8669 ( .B1(n7510), .B2(n10014), .A(n7509), .ZN(n7511) );
  OAI21_X1 U8670 ( .B1(n7512), .B2(n9843), .A(n7511), .ZN(P1_U3288) );
  NAND3_X1 U8671 ( .A1(n7375), .A2(n5199), .A3(n7514), .ZN(n7515) );
  AOI21_X1 U8672 ( .B1(n7516), .B2(n7515), .A(n9081), .ZN(n7521) );
  NAND2_X1 U8673 ( .A1(n9079), .A2(n8549), .ZN(n7518) );
  OAI211_X1 U8674 ( .C1(n9019), .C2(n7979), .A(n7518), .B(n7517), .ZN(n7520)
         );
  OAI22_X1 U8675 ( .A1(n7972), .A2(n9062), .B1(n9059), .B2(n7973), .ZN(n7519)
         );
  OR3_X1 U8676 ( .A1(n7521), .A2(n7520), .A3(n7519), .ZN(P2_U3241) );
  INV_X1 U8677 ( .A(n7522), .ZN(n7523) );
  OAI21_X1 U8678 ( .B1(n7526), .B2(n7527), .A(n7592), .ZN(n7528) );
  INV_X1 U8679 ( .A(n7826), .ZN(n7837) );
  AOI222_X1 U8680 ( .A1(n9869), .A2(n7528), .B1(n7837), .B2(n9866), .C1(n9661), 
        .C2(n9864), .ZN(n7604) );
  NAND2_X1 U8681 ( .A1(n9662), .A2(n7529), .ZN(n7530) );
  NAND2_X1 U8682 ( .A1(n7531), .A2(n7530), .ZN(n7658) );
  INV_X1 U8683 ( .A(n7658), .ZN(n7533) );
  INV_X1 U8684 ( .A(n7659), .ZN(n7532) );
  NAND2_X1 U8685 ( .A1(n7533), .A2(n7532), .ZN(n7656) );
  NAND2_X1 U8686 ( .A1(n7665), .A2(n7647), .ZN(n7534) );
  NAND2_X1 U8687 ( .A1(n7536), .A2(n7535), .ZN(n7588) );
  OAI21_X1 U8688 ( .B1(n7536), .B2(n7535), .A(n7588), .ZN(n7537) );
  INV_X1 U8689 ( .A(n7537), .ZN(n7605) );
  OAI22_X1 U8690 ( .A1(n10447), .A2(n7538), .B1(n7644), .B2(n10450), .ZN(n7539) );
  AOI21_X1 U8691 ( .B1(n9827), .B2(n7631), .A(n7539), .ZN(n7544) );
  OAI21_X1 U8692 ( .B1(n7664), .B2(n7652), .A(n9965), .ZN(n7540) );
  NOR2_X1 U8693 ( .A1(n7540), .A2(n7594), .ZN(n7602) );
  NOR2_X1 U8694 ( .A1(n7542), .A2(n7541), .ZN(n8364) );
  NAND2_X1 U8695 ( .A1(n7602), .A2(n8364), .ZN(n7543) );
  OAI211_X1 U8696 ( .C1(n7605), .C2(n9873), .A(n7544), .B(n7543), .ZN(n7545)
         );
  INV_X1 U8697 ( .A(n7545), .ZN(n7546) );
  OAI21_X1 U8698 ( .B1(n7604), .B2(n9843), .A(n7546), .ZN(P1_U3284) );
  NAND2_X1 U8699 ( .A1(n9661), .A2(n8943), .ZN(n7547) );
  OAI21_X1 U8700 ( .B1(n7665), .B2(n8950), .A(n7547), .ZN(n7548) );
  XNOR2_X1 U8701 ( .A(n7548), .B(n8947), .ZN(n7552) );
  NAND2_X1 U8702 ( .A1(n8925), .A2(n9661), .ZN(n7550) );
  OR2_X1 U8703 ( .A1(n7665), .A2(n8949), .ZN(n7549) );
  NAND2_X1 U8704 ( .A1(n7550), .A2(n7549), .ZN(n7551) );
  NOR2_X1 U8705 ( .A1(n7552), .A2(n7551), .ZN(n7627) );
  AOI21_X1 U8706 ( .B1(n7552), .B2(n7551), .A(n7627), .ZN(n7557) );
  OAI21_X1 U8707 ( .B1(n7555), .B2(n7554), .A(n7553), .ZN(n7556) );
  NAND2_X1 U8708 ( .A1(n7556), .A2(n7557), .ZN(n7640) );
  OAI21_X1 U8709 ( .B1(n7557), .B2(n7556), .A(n7640), .ZN(n7558) );
  NAND2_X1 U8710 ( .A1(n7558), .A2(n9604), .ZN(n7564) );
  INV_X1 U8711 ( .A(n7632), .ZN(n9660) );
  NAND2_X1 U8712 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10281) );
  INV_X1 U8713 ( .A(n10281), .ZN(n7559) );
  AOI21_X1 U8714 ( .B1(n9642), .B2(n9660), .A(n7559), .ZN(n7560) );
  OAI21_X1 U8715 ( .B1(n7561), .B2(n9607), .A(n7560), .ZN(n7562) );
  AOI21_X1 U8716 ( .B1(n7781), .B2(n4839), .A(n7562), .ZN(n7563) );
  OAI211_X1 U8717 ( .C1(n9646), .C2(n7666), .A(n7564), .B(n7563), .ZN(P1_U3237) );
  INV_X1 U8718 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U8719 ( .A1(n7565), .A2(n8527), .ZN(n7748) );
  NAND2_X1 U8720 ( .A1(n7578), .A2(n10488), .ZN(n8532) );
  NAND2_X1 U8721 ( .A1(n7748), .A2(n8530), .ZN(n7749) );
  NAND2_X1 U8722 ( .A1(n9100), .A2(n7703), .ZN(n8537) );
  NAND2_X1 U8723 ( .A1(n7750), .A2(n7778), .ZN(n8538) );
  INV_X1 U8724 ( .A(n8532), .ZN(n7566) );
  NOR2_X1 U8725 ( .A1(n8656), .A2(n7566), .ZN(n7567) );
  INV_X1 U8726 ( .A(n7706), .ZN(n7569) );
  INV_X1 U8727 ( .A(n8656), .ZN(n8535) );
  AOI21_X1 U8728 ( .B1(n7749), .B2(n8532), .A(n8535), .ZN(n7568) );
  INV_X1 U8729 ( .A(n10467), .ZN(n9371) );
  NOR3_X1 U8730 ( .A1(n7569), .A2(n7568), .A3(n9371), .ZN(n7581) );
  NAND2_X1 U8731 ( .A1(n7751), .A2(n7570), .ZN(n7752) );
  NAND2_X1 U8732 ( .A1(n7571), .A2(n7752), .ZN(n7572) );
  NAND2_X1 U8733 ( .A1(n7572), .A2(n8657), .ZN(n7575) );
  NAND2_X1 U8734 ( .A1(n7578), .A2(n7573), .ZN(n7576) );
  NAND2_X1 U8735 ( .A1(n7575), .A2(n7576), .ZN(n7574) );
  NAND2_X1 U8736 ( .A1(n7574), .A2(n8656), .ZN(n7705) );
  NAND3_X1 U8737 ( .A1(n7575), .A2(n8535), .A3(n7576), .ZN(n7577) );
  AOI21_X1 U8738 ( .B1(n7705), .B2(n7577), .A(n10564), .ZN(n7580) );
  OAI22_X1 U8739 ( .A1(n7972), .A2(n9341), .B1(n7578), .B2(n9343), .ZN(n7579)
         );
  NOR3_X1 U8740 ( .A1(n7581), .A2(n7580), .A3(n7579), .ZN(n7780) );
  OR2_X1 U8741 ( .A1(n7758), .A2(n7703), .ZN(n7772) );
  NAND3_X1 U8742 ( .A1(n7772), .A2(n10576), .A3(n7773), .ZN(n7582) );
  OAI211_X1 U8743 ( .C1(n7703), .C2(n10566), .A(n7780), .B(n7582), .ZN(n7585)
         );
  NAND2_X1 U8744 ( .A1(n7585), .A2(n10588), .ZN(n7583) );
  OAI21_X1 U8745 ( .B1(n10588), .B2(n7584), .A(n7583), .ZN(P2_U3463) );
  NAND2_X1 U8746 ( .A1(n7585), .A2(n10584), .ZN(n7586) );
  OAI21_X1 U8747 ( .B1(n10584), .B2(n6945), .A(n7586), .ZN(P2_U3524) );
  OR2_X1 U8748 ( .A1(n7631), .A2(n9660), .ZN(n7587) );
  INV_X1 U8749 ( .A(n7810), .ZN(n7589) );
  NAND2_X1 U8750 ( .A1(n7590), .A2(n7589), .ZN(n7809) );
  OAI21_X1 U8751 ( .B1(n7590), .B2(n7589), .A(n7809), .ZN(n7693) );
  XNOR2_X1 U8752 ( .A(n7811), .B(n7810), .ZN(n7593) );
  AOI222_X1 U8753 ( .A1(n9869), .A2(n7593), .B1(n9659), .B2(n9866), .C1(n9660), 
        .C2(n9864), .ZN(n7692) );
  OR2_X1 U8754 ( .A1(n7692), .A2(n9843), .ZN(n7601) );
  INV_X1 U8755 ( .A(n7594), .ZN(n7595) );
  INV_X1 U8756 ( .A(n7854), .ZN(n7596) );
  AOI21_X1 U8757 ( .B1(n7854), .B2(n7595), .A(n5054), .ZN(n7690) );
  NOR2_X1 U8758 ( .A1(n7596), .A2(n10442), .ZN(n7599) );
  OAI22_X1 U8759 ( .A1(n10447), .A2(n7597), .B1(n7852), .B2(n10450), .ZN(n7598) );
  AOI211_X1 U8760 ( .C1(n7690), .C2(n10006), .A(n7599), .B(n7598), .ZN(n7600)
         );
  OAI211_X1 U8761 ( .C1(n7693), .C2(n9873), .A(n7601), .B(n7600), .ZN(P1_U3283) );
  AOI21_X1 U8762 ( .B1(n9959), .B2(n7631), .A(n7602), .ZN(n7603) );
  OAI211_X1 U8763 ( .C1(n10494), .C2(n7605), .A(n7604), .B(n7603), .ZN(n7607)
         );
  NAND2_X1 U8764 ( .A1(n7607), .A2(n4842), .ZN(n7606) );
  OAI21_X1 U8765 ( .B1(n4842), .B2(n6345), .A(n7606), .ZN(P1_U3530) );
  INV_X1 U8766 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U8767 ( .A1(n7607), .A2(n4843), .ZN(n7608) );
  OAI21_X1 U8768 ( .B1(n4843), .B2(n7609), .A(n7608), .ZN(P1_U3475) );
  INV_X1 U8769 ( .A(n7610), .ZN(n7722) );
  OAI222_X1 U8770 ( .A1(P1_U3084), .A2(n7018), .B1(n7481), .B2(n7722), .C1(
        n7611), .C2(n8841), .ZN(P1_U3333) );
  NOR2_X1 U8771 ( .A1(n7888), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7612) );
  AOI21_X1 U8772 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7888), .A(n7612), .ZN(
        n7615) );
  OAI21_X1 U8773 ( .B1(n7618), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7613), .ZN(
        n7614) );
  NAND2_X1 U8774 ( .A1(n7615), .A2(n7614), .ZN(n7883) );
  OAI21_X1 U8775 ( .B1(n7615), .B2(n7614), .A(n7883), .ZN(n7616) );
  INV_X1 U8776 ( .A(n7616), .ZN(n7626) );
  AOI22_X1 U8777 ( .A1(n7888), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n5689), .B2(
        n7622), .ZN(n7620) );
  OAI21_X1 U8778 ( .B1(n7618), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7617), .ZN(
        n7619) );
  NAND2_X1 U8779 ( .A1(n7620), .A2(n7619), .ZN(n7887) );
  OAI21_X1 U8780 ( .B1(n7620), .B2(n7619), .A(n7887), .ZN(n7624) );
  NAND2_X1 U8781 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U8782 ( .A1(n10379), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7621) );
  OAI211_X1 U8783 ( .C1(n10356), .C2(n7622), .A(n8306), .B(n7621), .ZN(n7623)
         );
  AOI21_X1 U8784 ( .B1(n7624), .B2(n10391), .A(n7623), .ZN(n7625) );
  OAI21_X1 U8785 ( .B1(n7626), .B2(n10394), .A(n7625), .ZN(P2_U3259) );
  INV_X1 U8786 ( .A(n7627), .ZN(n7642) );
  NAND2_X1 U8787 ( .A1(n7631), .A2(n8936), .ZN(n7629) );
  OR2_X1 U8788 ( .A1(n7632), .A2(n8949), .ZN(n7628) );
  NAND2_X1 U8789 ( .A1(n7629), .A2(n7628), .ZN(n7630) );
  XNOR2_X1 U8790 ( .A(n7630), .B(n4840), .ZN(n7635) );
  NAND2_X1 U8791 ( .A1(n7631), .A2(n8898), .ZN(n7634) );
  OR2_X1 U8792 ( .A1(n7632), .A2(n8236), .ZN(n7633) );
  AND2_X1 U8793 ( .A1(n7634), .A2(n7633), .ZN(n7636) );
  NAND2_X1 U8794 ( .A1(n7635), .A2(n7636), .ZN(n8063) );
  INV_X1 U8795 ( .A(n7635), .ZN(n7638) );
  INV_X1 U8796 ( .A(n7636), .ZN(n7637) );
  NAND2_X1 U8797 ( .A1(n7638), .A2(n7637), .ZN(n7639) );
  NAND2_X1 U8798 ( .A1(n8063), .A2(n7639), .ZN(n7641) );
  AND3_X1 U8799 ( .A1(n7640), .A2(n7642), .A3(n7641), .ZN(n7643) );
  OAI21_X1 U8800 ( .B1(n8061), .B2(n7643), .A(n9604), .ZN(n7651) );
  INV_X1 U8801 ( .A(n7644), .ZN(n7649) );
  INV_X1 U8802 ( .A(n9646), .ZN(n9619) );
  AOI21_X1 U8803 ( .B1(n9642), .B2(n7837), .A(n7645), .ZN(n7646) );
  OAI21_X1 U8804 ( .B1(n7647), .B2(n9607), .A(n7646), .ZN(n7648) );
  AOI21_X1 U8805 ( .B1(n7649), .B2(n9619), .A(n7648), .ZN(n7650) );
  OAI211_X1 U8806 ( .C1(n7652), .C2(n9613), .A(n7651), .B(n7650), .ZN(P1_U3211) );
  NAND2_X1 U8807 ( .A1(n7654), .A2(n7653), .ZN(n7655) );
  XNOR2_X1 U8808 ( .A(n7655), .B(n7659), .ZN(n7663) );
  INV_X1 U8809 ( .A(n7656), .ZN(n7657) );
  AOI21_X1 U8810 ( .B1(n7659), .B2(n7658), .A(n7657), .ZN(n7785) );
  AOI22_X1 U8811 ( .A1(n9660), .A2(n9866), .B1(n9864), .B2(n9662), .ZN(n7660)
         );
  OAI21_X1 U8812 ( .B1(n7785), .B2(n7661), .A(n7660), .ZN(n7662) );
  AOI21_X1 U8813 ( .B1(n7663), .B2(n9869), .A(n7662), .ZN(n7784) );
  AOI21_X1 U8814 ( .B1(n7781), .B2(n5321), .A(n7664), .ZN(n7782) );
  NOR2_X1 U8815 ( .A1(n10442), .A2(n7665), .ZN(n7669) );
  OAI22_X1 U8816 ( .A1(n10447), .A2(n7667), .B1(n7666), .B2(n10450), .ZN(n7668) );
  AOI211_X1 U8817 ( .C1(n7782), .C2(n10006), .A(n7669), .B(n7668), .ZN(n7672)
         );
  INV_X1 U8818 ( .A(n7785), .ZN(n7670) );
  NAND2_X1 U8819 ( .A1(n7670), .A2(n10014), .ZN(n7671) );
  OAI211_X1 U8820 ( .C1(n7784), .C2(n9843), .A(n7672), .B(n7671), .ZN(P1_U3285) );
  OAI22_X1 U8821 ( .A1(n7674), .A2(n7673), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n7676), .ZN(n7790) );
  XNOR2_X1 U8822 ( .A(n7790), .B(n7797), .ZN(n7675) );
  NOR2_X1 U8823 ( .A1(n8281), .A2(n7675), .ZN(n7791) );
  AOI211_X1 U8824 ( .C1(n7675), .C2(n8281), .A(n7791), .B(n10411), .ZN(n7685)
         );
  OAI22_X1 U8825 ( .A1(n7678), .A2(n7677), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n7676), .ZN(n7796) );
  XNOR2_X1 U8826 ( .A(n7796), .B(n7797), .ZN(n7680) );
  NOR2_X1 U8827 ( .A1(n7679), .A2(n7680), .ZN(n7798) );
  AOI211_X1 U8828 ( .C1(n7680), .C2(n7679), .A(n7798), .B(n10433), .ZN(n7684)
         );
  NAND2_X1 U8829 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3084), .ZN(n7682) );
  NAND2_X1 U8830 ( .A1(n10436), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7681) );
  OAI211_X1 U8831 ( .C1(n10318), .C2(n7797), .A(n7682), .B(n7681), .ZN(n7683)
         );
  OR3_X1 U8832 ( .A1(n7685), .A2(n7684), .A3(n7683), .ZN(P1_U3256) );
  INV_X1 U8833 ( .A(n7686), .ZN(n7688) );
  OAI222_X1 U8834 ( .A1(n7687), .A2(P1_U3084), .B1(n8841), .B2(n6136), .C1(
        n7688), .C2(n7481), .ZN(P1_U3332) );
  OAI222_X1 U8835 ( .A1(n9503), .A2(n7689), .B1(P2_U3152), .B2(n8680), .C1(
        n7477), .C2(n7688), .ZN(P2_U3337) );
  INV_X1 U8836 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7695) );
  AOI22_X1 U8837 ( .A1(n7690), .A2(n9965), .B1(n9964), .B2(n7854), .ZN(n7691)
         );
  OAI211_X1 U8838 ( .C1(n10494), .C2(n7693), .A(n7692), .B(n7691), .ZN(n7696)
         );
  NAND2_X1 U8839 ( .A1(n7696), .A2(n4843), .ZN(n7694) );
  OAI21_X1 U8840 ( .B1(n4843), .B2(n7695), .A(n7694), .ZN(P1_U3478) );
  NAND2_X1 U8841 ( .A1(n7696), .A2(n4842), .ZN(n7697) );
  OAI21_X1 U8842 ( .B1(n4842), .B2(n6332), .A(n7697), .ZN(P1_U3531) );
  INV_X1 U8843 ( .A(n7698), .ZN(n7702) );
  INV_X1 U8844 ( .A(n7699), .ZN(n7700) );
  NAND3_X1 U8845 ( .A1(n7702), .A2(n7701), .A3(n7700), .ZN(n7744) );
  NAND2_X1 U8846 ( .A1(n7750), .A2(n7703), .ZN(n7704) );
  NAND2_X1 U8847 ( .A1(n7705), .A2(n7704), .ZN(n7930) );
  INV_X1 U8848 ( .A(n7930), .ZN(n7707) );
  OAI22_X1 U8849 ( .A1(n7707), .A2(n10564), .B1(n7925), .B2(n9371), .ZN(n7710)
         );
  OAI22_X1 U8850 ( .A1(n7930), .A2(n10564), .B1(n7708), .B2(n9371), .ZN(n7709)
         );
  NAND2_X1 U8851 ( .A1(n7972), .A2(n7718), .ZN(n8542) );
  INV_X1 U8852 ( .A(n7972), .ZN(n9099) );
  INV_X1 U8853 ( .A(n7718), .ZN(n7931) );
  NAND2_X1 U8854 ( .A1(n9099), .A2(n7931), .ZN(n8543) );
  NAND2_X1 U8855 ( .A1(n8542), .A2(n8543), .ZN(n8658) );
  INV_X1 U8856 ( .A(n8658), .ZN(n8540) );
  MUX2_X1 U8857 ( .A(n7710), .B(n7709), .S(n8540), .Z(n7712) );
  OAI22_X1 U8858 ( .A1(n7750), .A2(n9343), .B1(n7933), .B2(n9341), .ZN(n7711)
         );
  NOR2_X1 U8859 ( .A1(n7712), .A2(n7711), .ZN(n7725) );
  INV_X1 U8860 ( .A(n7725), .ZN(n7716) );
  OAI211_X1 U8861 ( .C1(n7931), .C2(n7713), .A(n7977), .B(n10576), .ZN(n7724)
         );
  OAI22_X1 U8862 ( .A1(n7724), .A2(n9180), .B1(n10471), .B2(n7714), .ZN(n7715)
         );
  OAI21_X1 U8863 ( .B1(n7716), .B2(n7715), .A(n9373), .ZN(n7720) );
  NAND2_X1 U8864 ( .A1(n9353), .A2(n7718), .ZN(n7719) );
  OAI211_X1 U8865 ( .C1(n7721), .C2(n9373), .A(n7720), .B(n7719), .ZN(P2_U3291) );
  OAI222_X1 U8866 ( .A1(n9503), .A2(n7723), .B1(P2_U3152), .B2(n5364), .C1(
        n7477), .C2(n7722), .ZN(P2_U3338) );
  INV_X1 U8867 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7727) );
  OAI211_X1 U8868 ( .C1(n7931), .C2(n10566), .A(n7725), .B(n7724), .ZN(n7728)
         );
  NAND2_X1 U8869 ( .A1(n7728), .A2(n10588), .ZN(n7726) );
  OAI21_X1 U8870 ( .B1(n10588), .B2(n7727), .A(n7726), .ZN(P2_U3466) );
  NAND2_X1 U8871 ( .A1(n7728), .A2(n10584), .ZN(n7729) );
  OAI21_X1 U8872 ( .B1(n10584), .B2(n6946), .A(n7729), .ZN(P2_U3525) );
  OAI211_X1 U8873 ( .C1(n7731), .C2(n7730), .A(n7900), .B(n9009), .ZN(n7739)
         );
  OR2_X1 U8874 ( .A1(n8128), .A2(n9341), .ZN(n7733) );
  OR2_X1 U8875 ( .A1(n7973), .A2(n9343), .ZN(n7732) );
  NAND2_X1 U8876 ( .A1(n7733), .A2(n7732), .ZN(n8820) );
  INV_X1 U8877 ( .A(n8820), .ZN(n7736) );
  INV_X1 U8878 ( .A(n8822), .ZN(n7734) );
  AOI22_X1 U8879 ( .A1(n9074), .A2(n7734), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n7735) );
  OAI21_X1 U8880 ( .B1(n7736), .B2(n9076), .A(n7735), .ZN(n7737) );
  AOI21_X1 U8881 ( .B1(n10520), .B2(n9079), .A(n7737), .ZN(n7738) );
  NAND2_X1 U8882 ( .A1(n7739), .A2(n7738), .ZN(P2_U3223) );
  NAND2_X1 U8883 ( .A1(n9105), .A2(n10470), .ZN(n8522) );
  AND2_X1 U8884 ( .A1(n10465), .A2(n8522), .ZN(n10453) );
  OR2_X1 U8885 ( .A1(n10453), .A2(n9371), .ZN(n7741) );
  NAND2_X1 U8886 ( .A1(n9103), .A2(n9390), .ZN(n7740) );
  AND2_X1 U8887 ( .A1(n7741), .A2(n7740), .ZN(n10451) );
  INV_X1 U8888 ( .A(n9373), .ZN(n9164) );
  OAI22_X1 U8889 ( .A1(n10451), .A2(n9164), .B1(n5425), .B2(n10471), .ZN(n7742) );
  AOI21_X1 U8890 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9393), .A(n7742), .ZN(
        n7747) );
  OR2_X1 U8891 ( .A1(n7744), .A2(n7743), .ZN(n10472) );
  INV_X1 U8892 ( .A(n10472), .ZN(n9396) );
  OAI21_X1 U8893 ( .B1(n9353), .B2(n9396), .A(n7745), .ZN(n7746) );
  OAI211_X1 U8894 ( .C1(n10453), .C2(n10476), .A(n7747), .B(n7746), .ZN(
        P2_U3296) );
  OAI21_X1 U8895 ( .B1(n8530), .B2(n7748), .A(n7749), .ZN(n7756) );
  OAI22_X1 U8896 ( .A1(n7751), .A2(n9343), .B1(n7750), .B2(n9341), .ZN(n7755)
         );
  NAND3_X1 U8897 ( .A1(n7571), .A2(n8530), .A3(n7752), .ZN(n7753) );
  AOI21_X1 U8898 ( .B1(n7575), .B2(n7753), .A(n10564), .ZN(n7754) );
  AOI211_X1 U8899 ( .C1(n10467), .C2(n7756), .A(n7755), .B(n7754), .ZN(n10491)
         );
  AND2_X1 U8900 ( .A1(n4850), .A2(n10488), .ZN(n7757) );
  NOR2_X1 U8901 ( .A1(n7758), .A2(n7757), .ZN(n10489) );
  INV_X1 U8902 ( .A(n10471), .ZN(n9382) );
  AOI22_X1 U8903 ( .A1(n9396), .A2(n10489), .B1(n9382), .B2(n7759), .ZN(n7760)
         );
  OAI21_X1 U8904 ( .B1(n7761), .B2(n9373), .A(n7760), .ZN(n7762) );
  AOI21_X1 U8905 ( .B1(n9353), .B2(n10488), .A(n7762), .ZN(n7763) );
  OAI21_X1 U8906 ( .B1(n10491), .B2(n9164), .A(n7763), .ZN(P2_U3293) );
  NAND3_X1 U8907 ( .A1(n9396), .A2(n4850), .A3(n7764), .ZN(n7766) );
  NAND2_X1 U8908 ( .A1(n9393), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7765) );
  OAI211_X1 U8909 ( .C1(n10471), .C2(n7767), .A(n7766), .B(n7765), .ZN(n7768)
         );
  AOI21_X1 U8910 ( .B1(n9353), .B2(n7769), .A(n7768), .ZN(n7770) );
  OAI21_X1 U8911 ( .B1(n7771), .B2(n9164), .A(n7770), .ZN(P2_U3294) );
  NAND3_X1 U8912 ( .A1(n9396), .A2(n7773), .A3(n7772), .ZN(n7775) );
  NAND2_X1 U8913 ( .A1(n9393), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7774) );
  OAI211_X1 U8914 ( .C1(n10471), .C2(n7776), .A(n7775), .B(n7774), .ZN(n7777)
         );
  AOI21_X1 U8915 ( .B1(n9353), .B2(n7778), .A(n7777), .ZN(n7779) );
  OAI21_X1 U8916 ( .B1(n7780), .B2(n9164), .A(n7779), .ZN(P2_U3292) );
  INV_X1 U8917 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7787) );
  AOI22_X1 U8918 ( .A1(n7782), .A2(n9965), .B1(n9964), .B2(n7781), .ZN(n7783)
         );
  OAI211_X1 U8919 ( .C1(n7785), .C2(n8182), .A(n7784), .B(n7783), .ZN(n7788)
         );
  NAND2_X1 U8920 ( .A1(n7788), .A2(n4843), .ZN(n7786) );
  OAI21_X1 U8921 ( .B1(n4843), .B2(n7787), .A(n7786), .ZN(P1_U3472) );
  NAND2_X1 U8922 ( .A1(n7788), .A2(n4842), .ZN(n7789) );
  OAI21_X1 U8923 ( .B1(n4842), .B2(n6845), .A(n7789), .ZN(P1_U3529) );
  NOR2_X1 U8924 ( .A1(n7797), .A2(n7790), .ZN(n7792) );
  NOR2_X1 U8925 ( .A1(n7792), .A2(n7791), .ZN(n7795) );
  NAND2_X1 U8926 ( .A1(n9675), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7793) );
  OAI21_X1 U8927 ( .B1(n9675), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7793), .ZN(
        n7794) );
  NOR2_X1 U8928 ( .A1(n7795), .A2(n7794), .ZN(n9666) );
  AOI211_X1 U8929 ( .C1(n7795), .C2(n7794), .A(n9666), .B(n10411), .ZN(n7807)
         );
  NOR2_X1 U8930 ( .A1(n7797), .A2(n7796), .ZN(n7799) );
  NOR2_X1 U8931 ( .A1(n7799), .A2(n7798), .ZN(n7801) );
  XNOR2_X1 U8932 ( .A(n9675), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7800) );
  NOR2_X1 U8933 ( .A1(n7801), .A2(n7800), .ZN(n9674) );
  AOI211_X1 U8934 ( .C1(n7801), .C2(n7800), .A(n9674), .B(n10433), .ZN(n7806)
         );
  NOR2_X1 U8935 ( .A1(n7802), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9567) );
  AOI21_X1 U8936 ( .B1(n10436), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9567), .ZN(
        n7803) );
  OAI21_X1 U8937 ( .B1(n7804), .B2(n10318), .A(n7803), .ZN(n7805) );
  OR3_X1 U8938 ( .A1(n7807), .A2(n7806), .A3(n7805), .ZN(P1_U3257) );
  NAND2_X1 U8939 ( .A1(n7854), .A2(n7837), .ZN(n7808) );
  XNOR2_X1 U8940 ( .A(n7871), .B(n7816), .ZN(n7878) );
  INV_X1 U8941 ( .A(n7861), .ZN(n7858) );
  AOI211_X1 U8942 ( .C1(n7816), .C2(n7815), .A(n9780), .B(n7858), .ZN(n7818)
         );
  OAI22_X1 U8943 ( .A1(n7826), .A2(n9782), .B1(n7835), .B2(n9784), .ZN(n7817)
         );
  NOR2_X1 U8944 ( .A1(n7818), .A2(n7817), .ZN(n7877) );
  OAI21_X1 U8945 ( .B1(n7840), .B2(n10450), .A(n7877), .ZN(n7819) );
  NAND2_X1 U8946 ( .A1(n7819), .A2(n10447), .ZN(n7824) );
  INV_X1 U8947 ( .A(n7865), .ZN(n7866) );
  AOI21_X1 U8948 ( .B1(n7874), .B2(n7820), .A(n7866), .ZN(n7875) );
  OAI22_X1 U8949 ( .A1(n5053), .A2(n10442), .B1(n7821), .B2(n10447), .ZN(n7822) );
  AOI21_X1 U8950 ( .B1(n7875), .B2(n10006), .A(n7822), .ZN(n7823) );
  OAI211_X1 U8951 ( .C1(n7878), .C2(n9873), .A(n7824), .B(n7823), .ZN(P1_U3282) );
  INV_X1 U8952 ( .A(n8063), .ZN(n7825) );
  NOR2_X1 U8953 ( .A1(n8061), .A2(n7825), .ZN(n7830) );
  INV_X1 U8954 ( .A(n8236), .ZN(n8925) );
  AOI22_X1 U8955 ( .A1(n7854), .A2(n8943), .B1(n8925), .B2(n7837), .ZN(n8062)
         );
  INV_X1 U8956 ( .A(n8062), .ZN(n8067) );
  NOR2_X1 U8957 ( .A1(n7830), .A2(n8067), .ZN(n7844) );
  NAND2_X1 U8958 ( .A1(n7854), .A2(n8936), .ZN(n7828) );
  OR2_X1 U8959 ( .A1(n7826), .A2(n8949), .ZN(n7827) );
  NAND2_X1 U8960 ( .A1(n7828), .A2(n7827), .ZN(n7829) );
  XNOR2_X1 U8961 ( .A(n7829), .B(n4841), .ZN(n8066) );
  NAND2_X1 U8962 ( .A1(n7830), .A2(n8067), .ZN(n7845) );
  OAI21_X1 U8963 ( .B1(n7844), .B2(n8066), .A(n7845), .ZN(n7834) );
  NAND2_X1 U8964 ( .A1(n7874), .A2(n8936), .ZN(n7832) );
  NAND2_X1 U8965 ( .A1(n9659), .A2(n8943), .ZN(n7831) );
  NAND2_X1 U8966 ( .A1(n7832), .A2(n7831), .ZN(n7833) );
  XNOR2_X1 U8967 ( .A(n7833), .B(n8947), .ZN(n8070) );
  AOI22_X1 U8968 ( .A1(n7874), .A2(n8943), .B1(n8925), .B2(n9659), .ZN(n8071)
         );
  XNOR2_X1 U8969 ( .A(n8070), .B(n8071), .ZN(n8069) );
  XNOR2_X1 U8970 ( .A(n7834), .B(n8069), .ZN(n7843) );
  INV_X1 U8971 ( .A(n7835), .ZN(n8174) );
  AOI21_X1 U8972 ( .B1(n9642), .B2(n8174), .A(n7836), .ZN(n7839) );
  NAND2_X1 U8973 ( .A1(n9641), .A2(n7837), .ZN(n7838) );
  OAI211_X1 U8974 ( .C1(n9646), .C2(n7840), .A(n7839), .B(n7838), .ZN(n7841)
         );
  AOI21_X1 U8975 ( .B1(n7874), .B2(n4839), .A(n7841), .ZN(n7842) );
  OAI21_X1 U8976 ( .B1(n7843), .B2(n9649), .A(n7842), .ZN(P1_U3229) );
  INV_X1 U8977 ( .A(n7844), .ZN(n7846) );
  NAND2_X1 U8978 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  XNOR2_X1 U8979 ( .A(n7847), .B(n8066), .ZN(n7856) );
  INV_X1 U8980 ( .A(n7848), .ZN(n7849) );
  AOI21_X1 U8981 ( .B1(n9642), .B2(n9659), .A(n7849), .ZN(n7851) );
  NAND2_X1 U8982 ( .A1(n9641), .A2(n9660), .ZN(n7850) );
  OAI211_X1 U8983 ( .C1(n9646), .C2(n7852), .A(n7851), .B(n7850), .ZN(n7853)
         );
  AOI21_X1 U8984 ( .B1(n7854), .B2(n4839), .A(n7853), .ZN(n7855) );
  OAI21_X1 U8985 ( .B1(n7856), .B2(n9649), .A(n7855), .ZN(P1_U3219) );
  INV_X1 U8986 ( .A(n7857), .ZN(n7859) );
  OAI21_X1 U8987 ( .B1(n7858), .B2(n7859), .A(n8045), .ZN(n7862) );
  NOR2_X1 U8988 ( .A1(n8045), .A2(n7859), .ZN(n7860) );
  NAND2_X1 U8989 ( .A1(n7862), .A2(n8040), .ZN(n7863) );
  AOI222_X1 U8990 ( .A1(n9869), .A2(n7863), .B1(n9658), .B2(n9866), .C1(n9659), 
        .C2(n9864), .ZN(n10536) );
  OAI22_X1 U8991 ( .A1(n10447), .A2(n7864), .B1(n8081), .B2(n10450), .ZN(n7868) );
  INV_X1 U8992 ( .A(n8083), .ZN(n10538) );
  INV_X1 U8993 ( .A(n8052), .ZN(n8178) );
  OAI211_X1 U8994 ( .C1(n10538), .C2(n7866), .A(n8178), .B(n9965), .ZN(n10535)
         );
  INV_X1 U8995 ( .A(n8364), .ZN(n8057) );
  NOR2_X1 U8996 ( .A1(n10535), .A2(n8057), .ZN(n7867) );
  AOI211_X1 U8997 ( .C1(n9827), .C2(n8083), .A(n7868), .B(n7867), .ZN(n7873)
         );
  AND2_X1 U8998 ( .A1(n7874), .A2(n9659), .ZN(n7870) );
  XNOR2_X1 U8999 ( .A(n8046), .B(n8045), .ZN(n10540) );
  NAND2_X1 U9000 ( .A1(n10540), .A2(n9734), .ZN(n7872) );
  OAI211_X1 U9001 ( .C1(n10536), .C2(n9843), .A(n7873), .B(n7872), .ZN(
        P1_U3281) );
  AOI22_X1 U9002 ( .A1(n7875), .A2(n9965), .B1(n9964), .B2(n7874), .ZN(n7876)
         );
  OAI211_X1 U9003 ( .C1(n10494), .C2(n7878), .A(n7877), .B(n7876), .ZN(n7880)
         );
  NAND2_X1 U9004 ( .A1(n7880), .A2(n4842), .ZN(n7879) );
  OAI21_X1 U9005 ( .B1(n4842), .B2(n6293), .A(n7879), .ZN(P1_U3532) );
  INV_X1 U9006 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U9007 ( .A1(n7880), .A2(n4843), .ZN(n7881) );
  OAI21_X1 U9008 ( .B1(n4843), .B2(n7882), .A(n7881), .ZN(P1_U3481) );
  OAI21_X1 U9009 ( .B1(n7888), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7883), .ZN(
        n8161) );
  XNOR2_X1 U9010 ( .A(n8161), .B(n7893), .ZN(n7884) );
  NAND2_X1 U9011 ( .A1(n7884), .A2(n5714), .ZN(n8163) );
  OAI21_X1 U9012 ( .B1(n7884), .B2(n5714), .A(n8163), .ZN(n7885) );
  INV_X1 U9013 ( .A(n7885), .ZN(n7895) );
  INV_X1 U9014 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U9015 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8413) );
  OAI21_X1 U9016 ( .B1(n9116), .B2(n7886), .A(n8413), .ZN(n7892) );
  OAI21_X1 U9017 ( .B1(n7888), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7887), .ZN(
        n8153) );
  XNOR2_X1 U9018 ( .A(n8153), .B(n8162), .ZN(n7890) );
  NOR2_X1 U9019 ( .A1(n7889), .A2(n7890), .ZN(n8154) );
  AOI211_X1 U9020 ( .C1(n7890), .C2(n7889), .A(n8154), .B(n10357), .ZN(n7891)
         );
  AOI211_X1 U9021 ( .C1(n10386), .C2(n7893), .A(n7892), .B(n7891), .ZN(n7894)
         );
  OAI21_X1 U9022 ( .B1(n7895), .B2(n10394), .A(n7894), .ZN(P2_U3260) );
  INV_X1 U9023 ( .A(n7896), .ZN(n8842) );
  OAI222_X1 U9024 ( .A1(n9503), .A2(n7898), .B1(n7477), .B2(n8842), .C1(n7897), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U9025 ( .A1(n7908), .A2(n7910), .ZN(n7901) );
  NAND2_X1 U9026 ( .A1(n7900), .A2(n7899), .ZN(n7909) );
  XOR2_X1 U9027 ( .A(n7901), .B(n7909), .Z(n7907) );
  OAI22_X1 U9028 ( .A1(n9019), .A2(n7963), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7902), .ZN(n7903) );
  AOI21_X1 U9029 ( .B1(n9039), .B2(n9096), .A(n7903), .ZN(n7904) );
  OAI21_X1 U9030 ( .B1(n8106), .B2(n9059), .A(n7904), .ZN(n7905) );
  AOI21_X1 U9031 ( .B1(n10527), .B2(n9079), .A(n7905), .ZN(n7906) );
  OAI21_X1 U9032 ( .B1(n7907), .B2(n9081), .A(n7906), .ZN(P2_U3233) );
  NAND2_X1 U9033 ( .A1(n7909), .A2(n7908), .ZN(n7911) );
  NAND2_X1 U9034 ( .A1(n7911), .A2(n7910), .ZN(n7913) );
  XNOR2_X1 U9035 ( .A(n7913), .B(n7912), .ZN(n7918) );
  INV_X1 U9036 ( .A(n8337), .ZN(n9093) );
  OAI22_X1 U9037 ( .A1(n9019), .A2(n8129), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10185), .ZN(n7914) );
  AOI21_X1 U9038 ( .B1(n9022), .B2(n9093), .A(n7914), .ZN(n7915) );
  OAI21_X1 U9039 ( .B1(n8128), .B2(n9062), .A(n7915), .ZN(n7916) );
  AOI21_X1 U9040 ( .B1(n8136), .B2(n9079), .A(n7916), .ZN(n7917) );
  OAI21_X1 U9041 ( .B1(n7918), .B2(n9081), .A(n7917), .ZN(P2_U3219) );
  NAND2_X1 U9042 ( .A1(n7921), .A2(n9507), .ZN(n7919) );
  OAI211_X1 U9043 ( .C1(n7920), .C2(n9503), .A(n7919), .B(n8694), .ZN(P2_U3335) );
  NAND2_X1 U9044 ( .A1(n7921), .A2(n9996), .ZN(n7923) );
  OAI211_X1 U9045 ( .C1(n7924), .C2(n8841), .A(n7923), .B(n7922), .ZN(P1_U3330) );
  NAND2_X1 U9046 ( .A1(n9098), .A2(n10504), .ZN(n7926) );
  NAND2_X1 U9047 ( .A1(n7973), .A2(n7939), .ZN(n8552) );
  INV_X1 U9048 ( .A(n7973), .ZN(n9097) );
  NAND2_X1 U9049 ( .A1(n9097), .A2(n10511), .ZN(n8553) );
  NAND2_X1 U9050 ( .A1(n8552), .A2(n8553), .ZN(n8546) );
  XNOR2_X1 U9051 ( .A(n7955), .B(n8546), .ZN(n7927) );
  NAND2_X1 U9052 ( .A1(n7927), .A2(n10467), .ZN(n7929) );
  AOI22_X1 U9053 ( .A1(n9098), .A2(n9388), .B1(n9390), .B2(n9096), .ZN(n7928)
         );
  NAND2_X1 U9054 ( .A1(n7929), .A2(n7928), .ZN(n10513) );
  INV_X1 U9055 ( .A(n10513), .ZN(n7943) );
  NAND2_X1 U9056 ( .A1(n7972), .A2(n7931), .ZN(n7932) );
  NAND2_X1 U9057 ( .A1(n7933), .A2(n10504), .ZN(n8548) );
  NAND2_X1 U9058 ( .A1(n9098), .A2(n8549), .ZN(n8547) );
  NAND2_X1 U9059 ( .A1(n8548), .A2(n8547), .ZN(n8660) );
  NAND2_X1 U9060 ( .A1(n7952), .A2(n8546), .ZN(n8831) );
  OAI21_X1 U9061 ( .B1(n7952), .B2(n8546), .A(n8831), .ZN(n10515) );
  INV_X1 U9062 ( .A(n10476), .ZN(n9224) );
  INV_X1 U9063 ( .A(n8826), .ZN(n7935) );
  OAI21_X1 U9064 ( .B1(n10511), .B2(n4925), .A(n7935), .ZN(n10512) );
  OAI22_X1 U9065 ( .A1(n9373), .A2(n7937), .B1(n7936), .B2(n10471), .ZN(n7938)
         );
  AOI21_X1 U9066 ( .B1(n9353), .B2(n7939), .A(n7938), .ZN(n7940) );
  OAI21_X1 U9067 ( .B1(n10512), .B2(n10472), .A(n7940), .ZN(n7941) );
  AOI21_X1 U9068 ( .B1(n10515), .B2(n9224), .A(n7941), .ZN(n7942) );
  OAI21_X1 U9069 ( .B1(n7943), .B2(n9164), .A(n7942), .ZN(P2_U3289) );
  NAND2_X1 U9070 ( .A1(n9096), .A2(n10520), .ZN(n7944) );
  AND2_X1 U9071 ( .A1(n8546), .A2(n7944), .ZN(n7947) );
  NAND2_X1 U9072 ( .A1(n7952), .A2(n7947), .ZN(n7946) );
  INV_X1 U9073 ( .A(n7944), .ZN(n7945) );
  INV_X1 U9074 ( .A(n8832), .ZN(n8664) );
  NAND2_X1 U9075 ( .A1(n7973), .A2(n10511), .ZN(n8830) );
  NAND2_X1 U9076 ( .A1(n7946), .A2(n7949), .ZN(n7953) );
  NAND2_X1 U9077 ( .A1(n10527), .A2(n8128), .ZN(n8559) );
  NAND2_X1 U9078 ( .A1(n8555), .A2(n8559), .ZN(n7958) );
  AND2_X1 U9079 ( .A1(n7947), .A2(n7958), .ZN(n7951) );
  INV_X1 U9080 ( .A(n7958), .ZN(n7948) );
  OAI21_X1 U9081 ( .B1(n7953), .B2(n7958), .A(n8113), .ZN(n10532) );
  INV_X1 U9082 ( .A(n10532), .ZN(n7969) );
  INV_X1 U9083 ( .A(n8553), .ZN(n7954) );
  OAI21_X1 U9084 ( .B1(n7955), .B2(n7954), .A(n8552), .ZN(n8819) );
  NAND2_X1 U9085 ( .A1(n7956), .A2(n10520), .ZN(n8558) );
  INV_X1 U9086 ( .A(n8558), .ZN(n7957) );
  NAND2_X1 U9087 ( .A1(n7959), .A2(n7948), .ZN(n8109) );
  OAI211_X1 U9088 ( .C1(n7959), .C2(n7948), .A(n8109), .B(n10467), .ZN(n7961)
         );
  INV_X1 U9089 ( .A(n8106), .ZN(n9094) );
  AOI22_X1 U9090 ( .A1(n9094), .A2(n9390), .B1(n9388), .B2(n9096), .ZN(n7960)
         );
  NAND2_X1 U9091 ( .A1(n7961), .A2(n7960), .ZN(n10530) );
  NAND2_X1 U9092 ( .A1(n8826), .A2(n8825), .ZN(n8824) );
  NAND2_X1 U9093 ( .A1(n8824), .A2(n10527), .ZN(n7962) );
  NAND2_X1 U9094 ( .A1(n8131), .A2(n7962), .ZN(n10529) );
  OAI22_X1 U9095 ( .A1(n9373), .A2(n7964), .B1(n7963), .B2(n10471), .ZN(n7965)
         );
  AOI21_X1 U9096 ( .B1(n9353), .B2(n10527), .A(n7965), .ZN(n7966) );
  OAI21_X1 U9097 ( .B1(n10529), .B2(n10472), .A(n7966), .ZN(n7967) );
  AOI21_X1 U9098 ( .B1(n10530), .B2(n9373), .A(n7967), .ZN(n7968) );
  OAI21_X1 U9099 ( .B1(n7969), .B2(n10476), .A(n7968), .ZN(P2_U3287) );
  XOR2_X1 U9100 ( .A(n8660), .B(n7970), .Z(n7971) );
  OAI222_X1 U9101 ( .A1(n9341), .A2(n7973), .B1(n9343), .B2(n7972), .C1(n9371), 
        .C2(n7971), .ZN(n10506) );
  INV_X1 U9102 ( .A(n7974), .ZN(n7976) );
  AND2_X1 U9103 ( .A1(n7975), .A2(n8660), .ZN(n10503) );
  NOR3_X1 U9104 ( .A1(n7976), .A2(n10503), .A3(n10476), .ZN(n7984) );
  AND2_X1 U9105 ( .A1(n7977), .A2(n8549), .ZN(n7978) );
  OR2_X1 U9106 ( .A1(n7978), .A2(n4925), .ZN(n10505) );
  NOR2_X1 U9107 ( .A1(n10471), .A2(n7979), .ZN(n7980) );
  AOI21_X1 U9108 ( .B1(n9164), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7980), .ZN(
        n7982) );
  NAND2_X1 U9109 ( .A1(n9353), .A2(n8549), .ZN(n7981) );
  OAI211_X1 U9110 ( .C1(n10505), .C2(n10472), .A(n7982), .B(n7981), .ZN(n7983)
         );
  AOI211_X1 U9111 ( .C1(n10506), .C2(n9373), .A(n7984), .B(n7983), .ZN(n7985)
         );
  INV_X1 U9112 ( .A(n7985), .ZN(P2_U3290) );
  AND2_X1 U9113 ( .A1(n7987), .A2(n7986), .ZN(n7989) );
  XNOR2_X1 U9114 ( .A(n7989), .B(n7988), .ZN(n7995) );
  OAI22_X1 U9115 ( .A1(n8106), .A2(n9343), .B1(n8372), .B2(n9341), .ZN(n8110)
         );
  NAND2_X1 U9116 ( .A1(n7990), .A2(n8110), .ZN(n7992) );
  OAI211_X1 U9117 ( .C1(n9019), .C2(n8118), .A(n7992), .B(n7991), .ZN(n7993)
         );
  AOI21_X1 U9118 ( .B1(n8338), .B2(n9079), .A(n7993), .ZN(n7994) );
  OAI21_X1 U9119 ( .B1(n7995), .B2(n9081), .A(n7994), .ZN(P2_U3238) );
  NOR2_X1 U9120 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8034) );
  NOR2_X1 U9121 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8032) );
  NOR2_X1 U9122 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8030) );
  NOR2_X1 U9123 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8028) );
  NOR2_X1 U9124 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8026) );
  NOR2_X1 U9125 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8024) );
  NAND2_X1 U9126 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8022) );
  XOR2_X1 U9127 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10247) );
  NAND2_X1 U9128 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8020) );
  XOR2_X1 U9129 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10245) );
  NOR2_X1 U9130 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8002) );
  XNOR2_X1 U9131 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10231) );
  NAND2_X1 U9132 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8000) );
  XOR2_X1 U9133 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10229) );
  NAND2_X1 U9134 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7998) );
  XOR2_X1 U9135 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10227) );
  AOI21_X1 U9136 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10222) );
  INV_X1 U9137 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7996) );
  NAND3_X1 U9138 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10224) );
  OAI21_X1 U9139 ( .B1(n10222), .B2(n7996), .A(n10224), .ZN(n10226) );
  NAND2_X1 U9140 ( .A1(n10227), .A2(n10226), .ZN(n7997) );
  NAND2_X1 U9141 ( .A1(n7998), .A2(n7997), .ZN(n10228) );
  NAND2_X1 U9142 ( .A1(n10229), .A2(n10228), .ZN(n7999) );
  NAND2_X1 U9143 ( .A1(n8000), .A2(n7999), .ZN(n10230) );
  NOR2_X1 U9144 ( .A1(n10231), .A2(n10230), .ZN(n8001) );
  NOR2_X1 U9145 ( .A1(n8002), .A2(n8001), .ZN(n8003) );
  NOR2_X1 U9146 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8003), .ZN(n10232) );
  AND2_X1 U9147 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8003), .ZN(n10233) );
  NOR2_X1 U9148 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10233), .ZN(n8004) );
  NOR2_X1 U9149 ( .A1(n10232), .A2(n8004), .ZN(n8005) );
  NAND2_X1 U9150 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n8005), .ZN(n8007) );
  XOR2_X1 U9151 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n8005), .Z(n10237) );
  NAND2_X1 U9152 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10237), .ZN(n8006) );
  NAND2_X1 U9153 ( .A1(n8007), .A2(n8006), .ZN(n8008) );
  NAND2_X1 U9154 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8008), .ZN(n8011) );
  XNOR2_X1 U9155 ( .A(n8009), .B(n8008), .ZN(n10239) );
  NAND2_X1 U9156 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10239), .ZN(n8010) );
  NAND2_X1 U9157 ( .A1(n8011), .A2(n8010), .ZN(n8012) );
  NAND2_X1 U9158 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8012), .ZN(n8015) );
  XNOR2_X1 U9159 ( .A(n8013), .B(n8012), .ZN(n10241) );
  NAND2_X1 U9160 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10241), .ZN(n8014) );
  NAND2_X1 U9161 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  NAND2_X1 U9162 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n8016), .ZN(n8018) );
  XOR2_X1 U9163 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n8016), .Z(n10243) );
  NAND2_X1 U9164 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10243), .ZN(n8017) );
  NAND2_X1 U9165 ( .A1(n8018), .A2(n8017), .ZN(n10244) );
  NAND2_X1 U9166 ( .A1(n10245), .A2(n10244), .ZN(n8019) );
  NAND2_X1 U9167 ( .A1(n8020), .A2(n8019), .ZN(n10246) );
  NAND2_X1 U9168 ( .A1(n10247), .A2(n10246), .ZN(n8021) );
  NAND2_X1 U9169 ( .A1(n8022), .A2(n8021), .ZN(n10249) );
  XNOR2_X1 U9170 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10248) );
  NOR2_X1 U9171 ( .A1(n10249), .A2(n10248), .ZN(n8023) );
  NOR2_X1 U9172 ( .A1(n8024), .A2(n8023), .ZN(n10251) );
  XNOR2_X1 U9173 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10250) );
  NOR2_X1 U9174 ( .A1(n10251), .A2(n10250), .ZN(n8025) );
  NOR2_X1 U9175 ( .A1(n8026), .A2(n8025), .ZN(n10253) );
  XNOR2_X1 U9176 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10252) );
  NOR2_X1 U9177 ( .A1(n10253), .A2(n10252), .ZN(n8027) );
  NOR2_X1 U9178 ( .A1(n8028), .A2(n8027), .ZN(n10255) );
  XNOR2_X1 U9179 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10254) );
  NOR2_X1 U9180 ( .A1(n10255), .A2(n10254), .ZN(n8029) );
  NOR2_X1 U9181 ( .A1(n8030), .A2(n8029), .ZN(n10257) );
  XNOR2_X1 U9182 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10256) );
  NOR2_X1 U9183 ( .A1(n10257), .A2(n10256), .ZN(n8031) );
  NOR2_X1 U9184 ( .A1(n8032), .A2(n8031), .ZN(n10259) );
  XNOR2_X1 U9185 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10258) );
  NOR2_X1 U9186 ( .A1(n10259), .A2(n10258), .ZN(n8033) );
  NOR2_X1 U9187 ( .A1(n8034), .A2(n8033), .ZN(n8035) );
  AND2_X1 U9188 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8035), .ZN(n10260) );
  NOR2_X1 U9189 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10260), .ZN(n8036) );
  NOR2_X1 U9190 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8035), .ZN(n10261) );
  NOR2_X1 U9191 ( .A1(n8036), .A2(n10261), .ZN(n8038) );
  XNOR2_X1 U9192 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8037) );
  XNOR2_X1 U9193 ( .A(n8038), .B(n8037), .ZN(ADD_1071_U4) );
  NAND2_X1 U9194 ( .A1(n8248), .A2(n8042), .ZN(n8043) );
  XNOR2_X1 U9195 ( .A(n8043), .B(n8050), .ZN(n8044) );
  OAI222_X1 U9196 ( .A1(n9784), .A2(n9524), .B1(n9782), .B2(n8089), .C1(n9780), 
        .C2(n8044), .ZN(n8210) );
  INV_X1 U9197 ( .A(n8210), .ZN(n8060) );
  NAND2_X1 U9198 ( .A1(n8046), .A2(n8045), .ZN(n8048) );
  OR2_X1 U9199 ( .A1(n8083), .A2(n8174), .ZN(n8047) );
  NAND2_X1 U9200 ( .A1(n8048), .A2(n8047), .ZN(n8257) );
  OR2_X1 U9201 ( .A1(n8257), .A2(n8261), .ZN(n8049) );
  NAND2_X1 U9202 ( .A1(n8049), .A2(n8264), .ZN(n8051) );
  XNOR2_X1 U9203 ( .A(n8051), .B(n8050), .ZN(n8212) );
  INV_X1 U9204 ( .A(n8258), .ZN(n8209) );
  OAI211_X1 U9205 ( .C1(n8053), .C2(n8209), .A(n9965), .B(n8290), .ZN(n8208)
         );
  OAI22_X1 U9206 ( .A1(n10447), .A2(n8054), .B1(n8204), .B2(n10450), .ZN(n8055) );
  AOI21_X1 U9207 ( .B1(n8258), .B2(n9827), .A(n8055), .ZN(n8056) );
  OAI21_X1 U9208 ( .B1(n8208), .B2(n8057), .A(n8056), .ZN(n8058) );
  AOI21_X1 U9209 ( .B1(n8212), .B2(n9734), .A(n8058), .ZN(n8059) );
  OAI21_X1 U9210 ( .B1(n8060), .B2(n9843), .A(n8059), .ZN(P1_U3279) );
  INV_X1 U9211 ( .A(n8066), .ZN(n8064) );
  OAI21_X1 U9212 ( .B1(n8064), .B2(n8067), .A(n8063), .ZN(n8065) );
  INV_X1 U9213 ( .A(n8070), .ZN(n8072) );
  AOI22_X1 U9214 ( .A1(n8083), .A2(n8936), .B1(n8898), .B2(n8174), .ZN(n8074)
         );
  XOR2_X1 U9215 ( .A(n8947), .B(n8074), .Z(n8076) );
  NAND2_X1 U9216 ( .A1(n8075), .A2(n8076), .ZN(n8087) );
  INV_X1 U9217 ( .A(n8076), .ZN(n8077) );
  NAND2_X1 U9218 ( .A1(n5283), .A2(n8077), .ZN(n8091) );
  NAND2_X1 U9219 ( .A1(n8087), .A2(n8091), .ZN(n8078) );
  AOI22_X1 U9220 ( .A1(n8083), .A2(n8943), .B1(n8925), .B2(n8174), .ZN(n8086)
         );
  XNOR2_X1 U9221 ( .A(n8078), .B(n8086), .ZN(n8085) );
  AND2_X1 U9222 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10287) );
  NOR2_X1 U9223 ( .A1(n9623), .A2(n8089), .ZN(n8079) );
  AOI211_X1 U9224 ( .C1(n9641), .C2(n9659), .A(n10287), .B(n8079), .ZN(n8080)
         );
  OAI21_X1 U9225 ( .B1(n9646), .B2(n8081), .A(n8080), .ZN(n8082) );
  AOI21_X1 U9226 ( .B1(n8083), .B2(n4839), .A(n8082), .ZN(n8084) );
  OAI21_X1 U9227 ( .B1(n8085), .B2(n9649), .A(n8084), .ZN(P1_U3215) );
  NAND2_X1 U9228 ( .A1(n8087), .A2(n8086), .ZN(n8092) );
  AND2_X1 U9229 ( .A1(n8092), .A2(n8091), .ZN(n8094) );
  OAI22_X1 U9230 ( .A1(n10012), .A2(n8950), .B1(n8089), .B2(n8949), .ZN(n8088)
         );
  XNOR2_X1 U9231 ( .A(n8088), .B(n8947), .ZN(n8187) );
  NOR2_X1 U9232 ( .A1(n8089), .A2(n8236), .ZN(n8090) );
  AOI21_X1 U9233 ( .B1(n8179), .B2(n8943), .A(n8090), .ZN(n8188) );
  XNOR2_X1 U9234 ( .A(n8187), .B(n8188), .ZN(n8093) );
  NAND3_X1 U9235 ( .A1(n8092), .A2(n8091), .A3(n8093), .ZN(n8191) );
  OAI211_X1 U9236 ( .C1(n8094), .C2(n8093), .A(n9604), .B(n8191), .ZN(n8100)
         );
  INV_X1 U9237 ( .A(n8095), .ZN(n10009) );
  AOI21_X1 U9238 ( .B1(n9641), .B2(n8174), .A(n8096), .ZN(n8097) );
  OAI21_X1 U9239 ( .B1(n8196), .B2(n9623), .A(n8097), .ZN(n8098) );
  AOI21_X1 U9240 ( .B1(n9619), .B2(n10009), .A(n8098), .ZN(n8099) );
  OAI211_X1 U9241 ( .C1(n10012), .C2(n9613), .A(n8100), .B(n8099), .ZN(
        P1_U3234) );
  INV_X1 U9242 ( .A(n8101), .ZN(n8104) );
  OAI222_X1 U9243 ( .A1(P2_U3152), .A2(n8103), .B1(n7477), .B2(n8104), .C1(
        n8102), .C2(n9503), .ZN(P2_U3334) );
  OAI222_X1 U9244 ( .A1(P1_U3084), .A2(n8105), .B1(n8841), .B2(n6469), .C1(
        n8104), .C2(n7481), .ZN(P1_U3329) );
  OR2_X1 U9245 ( .A1(n8136), .A2(n8106), .ZN(n8563) );
  NAND2_X1 U9246 ( .A1(n8136), .A2(n8106), .ZN(n8560) );
  NAND2_X1 U9247 ( .A1(n8563), .A2(n8560), .ZN(n8663) );
  INV_X1 U9248 ( .A(n8555), .ZN(n8107) );
  NOR2_X1 U9249 ( .A1(n8663), .A2(n8107), .ZN(n8108) );
  NAND2_X1 U9250 ( .A1(n8109), .A2(n8108), .ZN(n8124) );
  NAND2_X1 U9251 ( .A1(n8124), .A2(n8560), .ZN(n8335) );
  OR2_X1 U9252 ( .A1(n8338), .A2(n8337), .ZN(n8573) );
  NAND2_X1 U9253 ( .A1(n8338), .A2(n8337), .ZN(n8571) );
  NAND2_X1 U9254 ( .A1(n8573), .A2(n8571), .ZN(n8665) );
  XOR2_X1 U9255 ( .A(n8335), .B(n8665), .Z(n8111) );
  AOI21_X1 U9256 ( .B1(n8111), .B2(n10467), .A(n8110), .ZN(n10553) );
  INV_X1 U9257 ( .A(n8128), .ZN(n9095) );
  OR2_X1 U9258 ( .A1(n10527), .A2(n9095), .ZN(n8112) );
  NAND2_X1 U9259 ( .A1(n8136), .A2(n9094), .ZN(n8114) );
  OAI21_X1 U9260 ( .B1(n8115), .B2(n8665), .A(n8340), .ZN(n8116) );
  INV_X1 U9261 ( .A(n8116), .ZN(n10556) );
  INV_X1 U9262 ( .A(n8338), .ZN(n10554) );
  OAI21_X1 U9263 ( .B1(n8132), .B2(n10554), .A(n10576), .ZN(n8117) );
  OR2_X1 U9264 ( .A1(n8117), .A2(n8342), .ZN(n10552) );
  NOR2_X1 U9265 ( .A1(n9164), .A2(n9180), .ZN(n9365) );
  INV_X1 U9266 ( .A(n9365), .ZN(n9356) );
  OAI22_X1 U9267 ( .A1(n9373), .A2(n8119), .B1(n8118), .B2(n10471), .ZN(n8120)
         );
  AOI21_X1 U9268 ( .B1(n9353), .B2(n8338), .A(n8120), .ZN(n8121) );
  OAI21_X1 U9269 ( .B1(n10552), .B2(n9356), .A(n8121), .ZN(n8122) );
  AOI21_X1 U9270 ( .B1(n10556), .B2(n9224), .A(n8122), .ZN(n8123) );
  OAI21_X1 U9271 ( .B1(n9164), .B2(n10553), .A(n8123), .ZN(P2_U3285) );
  NAND2_X1 U9272 ( .A1(n8109), .A2(n8555), .ZN(n8126) );
  INV_X1 U9273 ( .A(n8124), .ZN(n8125) );
  AOI21_X1 U9274 ( .B1(n8663), .B2(n8126), .A(n8125), .ZN(n8127) );
  OAI222_X1 U9275 ( .A1(n9341), .A2(n8337), .B1(n9343), .B2(n8128), .C1(n9371), 
        .C2(n8127), .ZN(n10547) );
  INV_X1 U9276 ( .A(n10547), .ZN(n8142) );
  OAI22_X1 U9277 ( .A1(n9373), .A2(n8130), .B1(n8129), .B2(n10471), .ZN(n8135)
         );
  INV_X1 U9278 ( .A(n8132), .ZN(n8133) );
  OAI21_X1 U9279 ( .B1(n5171), .B2(n5168), .A(n8133), .ZN(n10546) );
  NOR2_X1 U9280 ( .A1(n10546), .A2(n10472), .ZN(n8134) );
  AOI211_X1 U9281 ( .C1(n9353), .C2(n8136), .A(n8135), .B(n8134), .ZN(n8141)
         );
  NOR2_X1 U9282 ( .A1(n8137), .A2(n8663), .ZN(n10545) );
  INV_X1 U9283 ( .A(n10545), .ZN(n8139) );
  NAND3_X1 U9284 ( .A1(n8139), .A2(n9224), .A3(n8138), .ZN(n8140) );
  OAI211_X1 U9285 ( .C1(n8142), .C2(n9164), .A(n8141), .B(n8140), .ZN(P2_U3286) );
  INV_X1 U9286 ( .A(n8143), .ZN(n8144) );
  AOI21_X1 U9287 ( .B1(n8146), .B2(n8145), .A(n8144), .ZN(n8152) );
  INV_X1 U9288 ( .A(n8393), .ZN(n9091) );
  OAI21_X1 U9289 ( .B1(n9019), .B2(n8345), .A(n8147), .ZN(n8148) );
  AOI21_X1 U9290 ( .B1(n9022), .B2(n9091), .A(n8148), .ZN(n8149) );
  OAI21_X1 U9291 ( .B1(n8337), .B2(n9062), .A(n8149), .ZN(n8150) );
  AOI21_X1 U9292 ( .B1(n8379), .B2(n9079), .A(n8150), .ZN(n8151) );
  OAI21_X1 U9293 ( .B1(n8152), .B2(n9081), .A(n8151), .ZN(P2_U3226) );
  NOR2_X1 U9294 ( .A1(n8162), .A2(n8153), .ZN(n8155) );
  NOR2_X1 U9295 ( .A1(n8155), .A2(n8154), .ZN(n8158) );
  AOI22_X1 U9296 ( .A1(n9110), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8156), .B2(
        n8160), .ZN(n8157) );
  NAND2_X1 U9297 ( .A1(n8158), .A2(n8157), .ZN(n9106) );
  OAI21_X1 U9298 ( .B1(n8158), .B2(n8157), .A(n9106), .ZN(n8170) );
  NOR2_X1 U9299 ( .A1(n10200), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9012) );
  AOI21_X1 U9300 ( .B1(n10379), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n9012), .ZN(
        n8159) );
  OAI21_X1 U9301 ( .B1(n10356), .B2(n8160), .A(n8159), .ZN(n8169) );
  NAND2_X1 U9302 ( .A1(n8162), .A2(n8161), .ZN(n8164) );
  NAND2_X1 U9303 ( .A1(n8164), .A2(n8163), .ZN(n8167) );
  NAND2_X1 U9304 ( .A1(n9110), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8165) );
  OAI21_X1 U9305 ( .B1(n9110), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8165), .ZN(
        n8166) );
  NOR2_X1 U9306 ( .A1(n8167), .A2(n8166), .ZN(n9109) );
  AOI211_X1 U9307 ( .C1(n8167), .C2(n8166), .A(n9109), .B(n10394), .ZN(n8168)
         );
  AOI211_X1 U9308 ( .C1(n8170), .C2(n10391), .A(n8169), .B(n8168), .ZN(n8171)
         );
  INV_X1 U9309 ( .A(n8171), .ZN(P2_U3261) );
  INV_X1 U9310 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8184) );
  XOR2_X1 U9311 ( .A(n8257), .B(n8172), .Z(n10015) );
  INV_X1 U9312 ( .A(n10015), .ZN(n8181) );
  XOR2_X1 U9313 ( .A(n8173), .B(n8172), .Z(n8176) );
  INV_X1 U9314 ( .A(n8196), .ZN(n8297) );
  AOI22_X1 U9315 ( .A1(n9864), .A2(n8174), .B1(n8297), .B2(n9866), .ZN(n8175)
         );
  OAI21_X1 U9316 ( .B1(n8176), .B2(n9780), .A(n8175), .ZN(n8177) );
  AOI21_X1 U9317 ( .B1(n10015), .B2(n8457), .A(n8177), .ZN(n10017) );
  AOI21_X1 U9318 ( .B1(n8179), .B2(n8178), .A(n8053), .ZN(n10007) );
  AOI22_X1 U9319 ( .A1(n10007), .A2(n9965), .B1(n9964), .B2(n8179), .ZN(n8180)
         );
  OAI211_X1 U9320 ( .C1(n8182), .C2(n8181), .A(n10017), .B(n8180), .ZN(n8185)
         );
  NAND2_X1 U9321 ( .A1(n8185), .A2(n4843), .ZN(n8183) );
  OAI21_X1 U9322 ( .B1(n4843), .B2(n8184), .A(n8183), .ZN(P1_U3487) );
  NAND2_X1 U9323 ( .A1(n8185), .A2(n4842), .ZN(n8186) );
  OAI21_X1 U9324 ( .B1(n4842), .B2(n6267), .A(n8186), .ZN(P1_U3534) );
  NAND2_X1 U9325 ( .A1(n8187), .A2(n8189), .ZN(n8190) );
  NAND2_X1 U9326 ( .A1(n8258), .A2(n8936), .ZN(n8193) );
  OR2_X1 U9327 ( .A1(n8196), .A2(n8949), .ZN(n8192) );
  NAND2_X1 U9328 ( .A1(n8193), .A2(n8192), .ZN(n8194) );
  XNOR2_X1 U9329 ( .A(n8194), .B(n4840), .ZN(n8199) );
  NOR2_X1 U9330 ( .A1(n8196), .A2(n8195), .ZN(n8197) );
  AOI21_X1 U9331 ( .B1(n8258), .B2(n8898), .A(n8197), .ZN(n8198) );
  NOR2_X1 U9332 ( .A1(n8199), .A2(n8198), .ZN(n8232) );
  NAND2_X1 U9333 ( .A1(n8199), .A2(n8198), .ZN(n8233) );
  INV_X1 U9334 ( .A(n8233), .ZN(n8200) );
  NOR2_X1 U9335 ( .A1(n8232), .A2(n8200), .ZN(n8201) );
  XNOR2_X1 U9336 ( .A(n8234), .B(n8201), .ZN(n8207) );
  AND2_X1 U9337 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10305) );
  NOR2_X1 U9338 ( .A1(n9623), .A2(n9524), .ZN(n8202) );
  AOI211_X1 U9339 ( .C1(n9641), .C2(n9658), .A(n10305), .B(n8202), .ZN(n8203)
         );
  OAI21_X1 U9340 ( .B1(n9646), .B2(n8204), .A(n8203), .ZN(n8205) );
  AOI21_X1 U9341 ( .B1(n8258), .B2(n4839), .A(n8205), .ZN(n8206) );
  OAI21_X1 U9342 ( .B1(n8207), .B2(n9649), .A(n8206), .ZN(P1_U3222) );
  INV_X1 U9343 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8214) );
  INV_X1 U9344 ( .A(n10494), .ZN(n10541) );
  OAI21_X1 U9345 ( .B1(n8209), .B2(n10537), .A(n8208), .ZN(n8211) );
  AOI211_X1 U9346 ( .C1(n8212), .C2(n10541), .A(n8211), .B(n8210), .ZN(n8215)
         );
  OR2_X1 U9347 ( .A1(n8215), .A2(n10543), .ZN(n8213) );
  OAI21_X1 U9348 ( .B1(n4843), .B2(n8214), .A(n8213), .ZN(P1_U3490) );
  OR2_X1 U9349 ( .A1(n8215), .A2(n10542), .ZN(n8216) );
  OAI21_X1 U9350 ( .B1(n4842), .B2(n7420), .A(n8216), .ZN(P1_U3535) );
  INV_X1 U9351 ( .A(n8396), .ZN(n10567) );
  OAI21_X1 U9352 ( .B1(n8219), .B2(n8218), .A(n8217), .ZN(n8220) );
  NAND2_X1 U9353 ( .A1(n8220), .A2(n9009), .ZN(n8225) );
  INV_X1 U9354 ( .A(n8372), .ZN(n9092) );
  INV_X1 U9355 ( .A(n8471), .ZN(n9389) );
  NAND2_X1 U9356 ( .A1(n9022), .A2(n9389), .ZN(n8222) );
  OAI211_X1 U9357 ( .C1(n9019), .C2(n8376), .A(n8222), .B(n8221), .ZN(n8223)
         );
  AOI21_X1 U9358 ( .B1(n9039), .B2(n9092), .A(n8223), .ZN(n8224) );
  OAI211_X1 U9359 ( .C1(n10567), .C2(n9016), .A(n8225), .B(n8224), .ZN(
        P2_U3236) );
  INV_X1 U9360 ( .A(n8226), .ZN(n8230) );
  OAI222_X1 U9361 ( .A1(n9503), .A2(n8228), .B1(n7477), .B2(n8230), .C1(
        P2_U3152), .C2(n8227), .ZN(P2_U3333) );
  OAI222_X1 U9362 ( .A1(P1_U3084), .A2(n8231), .B1(n7481), .B2(n8230), .C1(
        n8229), .C2(n8841), .ZN(P1_U3328) );
  AOI21_X2 U9363 ( .B1(n8234), .B2(n8233), .A(n8232), .ZN(n8762) );
  INV_X1 U9364 ( .A(n9524), .ZN(n9657) );
  AOI22_X1 U9365 ( .A1(n9963), .A2(n8936), .B1(n8898), .B2(n9657), .ZN(n8235)
         );
  XNOR2_X1 U9366 ( .A(n8235), .B(n8947), .ZN(n8761) );
  INV_X1 U9367 ( .A(n8761), .ZN(n8239) );
  NAND2_X1 U9368 ( .A1(n9963), .A2(n8943), .ZN(n8238) );
  OR2_X1 U9369 ( .A1(n9524), .A2(n8236), .ZN(n8237) );
  NAND2_X1 U9370 ( .A1(n8238), .A2(n8237), .ZN(n8769) );
  XNOR2_X1 U9371 ( .A(n8239), .B(n8769), .ZN(n8240) );
  XNOR2_X1 U9372 ( .A(n8762), .B(n8240), .ZN(n8246) );
  NOR2_X1 U9373 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8241), .ZN(n10320) );
  NOR2_X1 U9374 ( .A1(n9623), .A2(n8765), .ZN(n8242) );
  AOI211_X1 U9375 ( .C1(n9641), .C2(n8297), .A(n10320), .B(n8242), .ZN(n8243)
         );
  OAI21_X1 U9376 ( .B1(n9646), .B2(n8291), .A(n8243), .ZN(n8244) );
  AOI21_X1 U9377 ( .B1(n9963), .B2(n4839), .A(n8244), .ZN(n8245) );
  OAI21_X1 U9378 ( .B1(n8246), .B2(n9649), .A(n8245), .ZN(P1_U3232) );
  NAND2_X1 U9379 ( .A1(n8250), .A2(n8249), .ZN(n8295) );
  NOR2_X1 U9380 ( .A1(n8322), .A2(n8251), .ZN(n8252) );
  NAND2_X1 U9381 ( .A1(n8314), .A2(n8252), .ZN(n8311) );
  OAI21_X1 U9382 ( .B1(n8255), .B2(n8254), .A(n8359), .ZN(n8256) );
  INV_X1 U9383 ( .A(n9582), .ZN(n9654) );
  INV_X1 U9384 ( .A(n8765), .ZN(n9656) );
  AOI222_X1 U9385 ( .A1(n9869), .A2(n8256), .B1(n9654), .B2(n9866), .C1(n9656), 
        .C2(n9864), .ZN(n9955) );
  INV_X1 U9386 ( .A(n8257), .ZN(n8262) );
  NAND2_X1 U9387 ( .A1(n8258), .A2(n8297), .ZN(n8263) );
  INV_X1 U9388 ( .A(n8263), .ZN(n8260) );
  NOR2_X1 U9389 ( .A1(n8260), .A2(n8259), .ZN(n8266) );
  AND2_X1 U9390 ( .A1(n8264), .A2(n8263), .ZN(n8265) );
  OR2_X1 U9391 ( .A1(n8266), .A2(n8265), .ZN(n8271) );
  NAND2_X1 U9392 ( .A1(n8273), .A2(n8271), .ZN(n8288) );
  OR2_X1 U9393 ( .A1(n8288), .A2(n8296), .ZN(n8320) );
  OR2_X1 U9394 ( .A1(n9963), .A2(n9657), .ZN(n8319) );
  OR2_X1 U9395 ( .A1(n9958), .A2(n9656), .ZN(n8267) );
  AND2_X1 U9396 ( .A1(n8319), .A2(n8267), .ZN(n8274) );
  NAND2_X1 U9397 ( .A1(n8320), .A2(n8274), .ZN(n8269) );
  INV_X1 U9398 ( .A(n8267), .ZN(n8268) );
  NAND2_X1 U9399 ( .A1(n8269), .A2(n8270), .ZN(n8280) );
  NAND2_X1 U9400 ( .A1(n8273), .A2(n8272), .ZN(n8278) );
  AND2_X1 U9401 ( .A1(n8274), .A2(n8279), .ZN(n8275) );
  OR2_X1 U9402 ( .A1(n8276), .A2(n8275), .ZN(n8277) );
  NAND2_X1 U9403 ( .A1(n8278), .A2(n8277), .ZN(n8439) );
  OAI21_X1 U9404 ( .B1(n8280), .B2(n8279), .A(n8439), .ZN(n9956) );
  OAI22_X1 U9405 ( .A1(n10447), .A2(n8281), .B1(n9645), .B2(n10450), .ZN(n8282) );
  AOI21_X1 U9406 ( .B1(n9952), .B2(n9827), .A(n8282), .ZN(n8285) );
  AND2_X1 U9407 ( .A1(n8329), .A2(n9952), .ZN(n8283) );
  NOR2_X1 U9408 ( .A1(n8361), .A2(n8283), .ZN(n9953) );
  NAND2_X1 U9409 ( .A1(n9953), .A2(n10006), .ZN(n8284) );
  OAI211_X1 U9410 ( .C1(n9956), .C2(n9873), .A(n8285), .B(n8284), .ZN(n8286)
         );
  INV_X1 U9411 ( .A(n8286), .ZN(n8287) );
  OAI21_X1 U9412 ( .B1(n9843), .B2(n9955), .A(n8287), .ZN(P1_U3276) );
  XOR2_X1 U9413 ( .A(n8296), .B(n8288), .Z(n9969) );
  INV_X1 U9414 ( .A(n8327), .ZN(n8289) );
  AOI21_X1 U9415 ( .B1(n9963), .B2(n8290), .A(n8289), .ZN(n9966) );
  INV_X1 U9416 ( .A(n9963), .ZN(n8294) );
  INV_X1 U9417 ( .A(n8291), .ZN(n8292) );
  INV_X1 U9418 ( .A(n10450), .ZN(n10008) );
  AOI22_X1 U9419 ( .A1(n9843), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8292), .B2(
        n10008), .ZN(n8293) );
  OAI21_X1 U9420 ( .B1(n8294), .B2(n10442), .A(n8293), .ZN(n8300) );
  OAI21_X1 U9421 ( .B1(n8296), .B2(n8295), .A(n8314), .ZN(n8298) );
  AOI222_X1 U9422 ( .A1(n9869), .A2(n8298), .B1(n9656), .B2(n9866), .C1(n8297), 
        .C2(n9864), .ZN(n9968) );
  NOR2_X1 U9423 ( .A1(n9968), .A2(n9843), .ZN(n8299) );
  AOI211_X1 U9424 ( .C1(n9966), .C2(n10006), .A(n8300), .B(n8299), .ZN(n8301)
         );
  OAI21_X1 U9425 ( .B1(n9873), .B2(n9969), .A(n8301), .ZN(P1_U3278) );
  INV_X1 U9426 ( .A(n10574), .ZN(n8400) );
  OAI21_X1 U9427 ( .B1(n8304), .B2(n8303), .A(n8302), .ZN(n8305) );
  NAND2_X1 U9428 ( .A1(n8305), .A2(n9009), .ZN(n8310) );
  INV_X1 U9429 ( .A(n8477), .ZN(n9090) );
  NAND2_X1 U9430 ( .A1(n9022), .A2(n9090), .ZN(n8307) );
  OAI211_X1 U9431 ( .C1(n9019), .C2(n8401), .A(n8307), .B(n8306), .ZN(n8308)
         );
  AOI21_X1 U9432 ( .B1(n9039), .B2(n9091), .A(n8308), .ZN(n8309) );
  OAI211_X1 U9433 ( .C1(n8400), .C2(n9016), .A(n8310), .B(n8309), .ZN(P2_U3217) );
  INV_X1 U9434 ( .A(n8311), .ZN(n8316) );
  AOI21_X1 U9435 ( .B1(n8314), .B2(n8313), .A(n8312), .ZN(n8315) );
  NOR3_X1 U9436 ( .A1(n8316), .A2(n8315), .A3(n9780), .ZN(n8318) );
  OAI22_X1 U9437 ( .A1(n9524), .A2(n9782), .B1(n9569), .B2(n9784), .ZN(n8317)
         );
  NOR2_X1 U9438 ( .A1(n8318), .A2(n8317), .ZN(n9961) );
  NAND2_X1 U9439 ( .A1(n8320), .A2(n8319), .ZN(n8323) );
  NAND2_X1 U9440 ( .A1(n8323), .A2(n8322), .ZN(n8321) );
  OAI21_X1 U9441 ( .B1(n8323), .B2(n8322), .A(n8321), .ZN(n8324) );
  INV_X1 U9442 ( .A(n8324), .ZN(n9962) );
  OAI22_X1 U9443 ( .A1(n10447), .A2(n8325), .B1(n9527), .B2(n10450), .ZN(n8326) );
  AOI21_X1 U9444 ( .B1(n9958), .B2(n9827), .A(n8326), .ZN(n8331) );
  AOI21_X1 U9445 ( .B1(n8327), .B2(n9958), .A(n7137), .ZN(n8328) );
  AND2_X1 U9446 ( .A1(n8329), .A2(n8328), .ZN(n9957) );
  NAND2_X1 U9447 ( .A1(n9957), .A2(n8364), .ZN(n8330) );
  OAI211_X1 U9448 ( .C1(n9962), .C2(n9873), .A(n8331), .B(n8330), .ZN(n8332)
         );
  INV_X1 U9449 ( .A(n8332), .ZN(n8333) );
  OAI21_X1 U9450 ( .B1(n9843), .B2(n9961), .A(n8333), .ZN(P1_U3277) );
  INV_X1 U9451 ( .A(n8571), .ZN(n8334) );
  OAI21_X1 U9452 ( .B1(n8335), .B2(n8334), .A(n8573), .ZN(n8370) );
  OR2_X1 U9453 ( .A1(n8379), .A2(n8372), .ZN(n8574) );
  NAND2_X1 U9454 ( .A1(n8379), .A2(n8372), .ZN(n8575) );
  XNOR2_X1 U9455 ( .A(n8370), .B(n8668), .ZN(n8336) );
  OAI222_X1 U9456 ( .A1(n9341), .A2(n8393), .B1(n9343), .B2(n8337), .C1(n9371), 
        .C2(n8336), .ZN(n10560) );
  INV_X1 U9457 ( .A(n10560), .ZN(n8350) );
  NAND2_X1 U9458 ( .A1(n8338), .A2(n9093), .ZN(n8339) );
  NAND2_X1 U9459 ( .A1(n8341), .A2(n8369), .ZN(n8381) );
  OAI21_X1 U9460 ( .B1(n8341), .B2(n8369), .A(n8381), .ZN(n10562) );
  INV_X1 U9461 ( .A(n8379), .ZN(n10558) );
  OR2_X1 U9462 ( .A1(n8342), .A2(n10558), .ZN(n8343) );
  NAND2_X1 U9463 ( .A1(n8373), .A2(n8343), .ZN(n10559) );
  NAND2_X1 U9464 ( .A1(n9164), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8344) );
  OAI21_X1 U9465 ( .B1(n10471), .B2(n8345), .A(n8344), .ZN(n8346) );
  AOI21_X1 U9466 ( .B1(n9353), .B2(n8379), .A(n8346), .ZN(n8347) );
  OAI21_X1 U9467 ( .B1(n10559), .B2(n10472), .A(n8347), .ZN(n8348) );
  AOI21_X1 U9468 ( .B1(n10562), .B2(n9224), .A(n8348), .ZN(n8349) );
  OAI21_X1 U9469 ( .B1(n9164), .B2(n8350), .A(n8349), .ZN(P2_U3284) );
  INV_X1 U9470 ( .A(n8351), .ZN(n8355) );
  OAI222_X1 U9471 ( .A1(P2_U3152), .A2(n8353), .B1(n7477), .B2(n8355), .C1(
        n8352), .C2(n9503), .ZN(P2_U3332) );
  OAI222_X1 U9472 ( .A1(n8356), .A2(P1_U3084), .B1(n7481), .B2(n8355), .C1(
        n8354), .C2(n8841), .ZN(P1_U3327) );
  INV_X1 U9473 ( .A(n9569), .ZN(n9655) );
  NAND2_X1 U9474 ( .A1(n9952), .A2(n9655), .ZN(n8434) );
  NAND2_X1 U9475 ( .A1(n8439), .A2(n8434), .ZN(n8357) );
  XNOR2_X1 U9476 ( .A(n8357), .B(n8436), .ZN(n9951) );
  XNOR2_X1 U9477 ( .A(n8428), .B(n8436), .ZN(n8360) );
  OAI222_X1 U9478 ( .A1(n9784), .A2(n8784), .B1(n9782), .B2(n9569), .C1(n8360), 
        .C2(n9780), .ZN(n9947) );
  INV_X1 U9479 ( .A(n9949), .ZN(n9574) );
  INV_X1 U9480 ( .A(n8361), .ZN(n8363) );
  NAND2_X1 U9481 ( .A1(n8361), .A2(n9574), .ZN(n8431) );
  INV_X1 U9482 ( .A(n8431), .ZN(n8362) );
  AOI211_X1 U9483 ( .C1(n9949), .C2(n8363), .A(n7137), .B(n8362), .ZN(n9948)
         );
  NAND2_X1 U9484 ( .A1(n9948), .A2(n8364), .ZN(n8366) );
  AOI22_X1 U9485 ( .A1(n9843), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9571), .B2(
        n10008), .ZN(n8365) );
  OAI211_X1 U9486 ( .C1(n9574), .C2(n10442), .A(n8366), .B(n8365), .ZN(n8367)
         );
  AOI21_X1 U9487 ( .B1(n9947), .B2(n10447), .A(n8367), .ZN(n8368) );
  OAI21_X1 U9488 ( .B1(n9951), .B2(n9873), .A(n8368), .ZN(P1_U3275) );
  OR2_X1 U9489 ( .A1(n8396), .A2(n8393), .ZN(n8582) );
  NAND2_X1 U9490 ( .A1(n8396), .A2(n8393), .ZN(n8581) );
  NAND2_X1 U9491 ( .A1(n8582), .A2(n8581), .ZN(n8389) );
  XNOR2_X1 U9492 ( .A(n8390), .B(n8389), .ZN(n8371) );
  OAI222_X1 U9493 ( .A1(n9341), .A2(n8471), .B1(n9343), .B2(n8372), .C1(n8371), 
        .C2(n9371), .ZN(n10570) );
  NAND2_X1 U9494 ( .A1(n8373), .A2(n8396), .ZN(n8374) );
  NAND2_X1 U9495 ( .A1(n8747), .A2(n8374), .ZN(n10569) );
  NAND2_X1 U9496 ( .A1(n9164), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8375) );
  OAI21_X1 U9497 ( .B1(n10471), .B2(n8376), .A(n8375), .ZN(n8377) );
  AOI21_X1 U9498 ( .B1(n8396), .B2(n9353), .A(n8377), .ZN(n8378) );
  OAI21_X1 U9499 ( .B1(n10569), .B2(n10472), .A(n8378), .ZN(n8385) );
  OR2_X1 U9500 ( .A1(n8379), .A2(n9092), .ZN(n8380) );
  NOR2_X1 U9501 ( .A1(n8382), .A2(n8389), .ZN(n10565) );
  INV_X1 U9502 ( .A(n8398), .ZN(n8383) );
  NOR3_X1 U9503 ( .A1(n10565), .A2(n8383), .A3(n10476), .ZN(n8384) );
  AOI211_X1 U9504 ( .C1(n9373), .C2(n10570), .A(n8385), .B(n8384), .ZN(n8386)
         );
  INV_X1 U9505 ( .A(n8386), .ZN(P2_U3283) );
  INV_X1 U9506 ( .A(n8387), .ZN(n8417) );
  OAI222_X1 U9507 ( .A1(P1_U3084), .A2(n4848), .B1(n7481), .B2(n8417), .C1(
        n8388), .C2(n8841), .ZN(P1_U3326) );
  INV_X1 U9508 ( .A(n8389), .ZN(n8669) );
  XNOR2_X1 U9509 ( .A(n10574), .B(n8471), .ZN(n8671) );
  AOI21_X1 U9510 ( .B1(n8391), .B2(n8671), .A(n9371), .ZN(n8395) );
  NAND2_X1 U9511 ( .A1(n8392), .A2(n8584), .ZN(n8474) );
  OAI22_X1 U9512 ( .A1(n8393), .A2(n9343), .B1(n8477), .B2(n9341), .ZN(n8394)
         );
  AOI21_X1 U9513 ( .B1(n8395), .B2(n8474), .A(n8394), .ZN(n10579) );
  NAND2_X1 U9514 ( .A1(n8396), .A2(n9091), .ZN(n8397) );
  OAI21_X1 U9515 ( .B1(n8399), .B2(n8671), .A(n8845), .ZN(n10582) );
  NAND2_X1 U9516 ( .A1(n10582), .A2(n9224), .ZN(n8406) );
  XOR2_X1 U9517 ( .A(n10574), .B(n8747), .Z(n10577) );
  NOR2_X1 U9518 ( .A1(n8400), .A2(n10475), .ZN(n8404) );
  OAI22_X1 U9519 ( .A1(n9373), .A2(n8402), .B1(n8401), .B2(n10471), .ZN(n8403)
         );
  AOI211_X1 U9520 ( .C1(n10577), .C2(n9396), .A(n8404), .B(n8403), .ZN(n8405)
         );
  OAI211_X1 U9521 ( .C1(n9164), .C2(n10579), .A(n8406), .B(n8405), .ZN(
        P2_U3282) );
  OAI21_X1 U9522 ( .B1(n8409), .B2(n8408), .A(n8407), .ZN(n8410) );
  NAND2_X1 U9523 ( .A1(n8410), .A2(n9009), .ZN(n8416) );
  INV_X1 U9524 ( .A(n8411), .ZN(n9383) );
  NAND2_X1 U9525 ( .A1(n9074), .A2(n9383), .ZN(n8412) );
  OAI211_X1 U9526 ( .C1(n9059), .C2(n9344), .A(n8413), .B(n8412), .ZN(n8414)
         );
  AOI21_X1 U9527 ( .B1(n9039), .B2(n9389), .A(n8414), .ZN(n8415) );
  OAI211_X1 U9528 ( .C1(n9385), .C2(n9016), .A(n8416), .B(n8415), .ZN(P2_U3243) );
  OAI222_X1 U9529 ( .A1(n9503), .A2(n8418), .B1(P2_U3152), .B2(n8749), .C1(
        n7477), .C2(n8417), .ZN(P2_U3331) );
  INV_X1 U9530 ( .A(n8419), .ZN(n8468) );
  OAI222_X1 U9531 ( .A1(n9503), .A2(n8420), .B1(P2_U3152), .B2(n6053), .C1(
        n7477), .C2(n8468), .ZN(P2_U3330) );
  INV_X1 U9532 ( .A(n8490), .ZN(n8424) );
  OAI222_X1 U9533 ( .A1(n7481), .A2(n8424), .B1(n8422), .B2(P1_U3084), .C1(
        n8421), .C2(n8841), .ZN(P1_U3324) );
  INV_X1 U9534 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8491) );
  OAI222_X1 U9535 ( .A1(n7477), .A2(n8424), .B1(P2_U3152), .B2(n8423), .C1(
        n8491), .C2(n9503), .ZN(P2_U3329) );
  INV_X1 U9536 ( .A(n8425), .ZN(n8427) );
  XOR2_X1 U9537 ( .A(n8451), .B(n8444), .Z(n8429) );
  INV_X1 U9538 ( .A(n8794), .ZN(n9865) );
  AOI222_X1 U9539 ( .A1(n9869), .A2(n8429), .B1(n9865), .B2(n9866), .C1(n9654), 
        .C2(n9864), .ZN(n9945) );
  INV_X1 U9540 ( .A(n5319), .ZN(n8430) );
  AOI21_X1 U9541 ( .B1(n9942), .B2(n8431), .A(n8430), .ZN(n9943) );
  INV_X1 U9542 ( .A(n9942), .ZN(n9588) );
  INV_X1 U9543 ( .A(n9583), .ZN(n8432) );
  AOI22_X1 U9544 ( .A1(n9843), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8432), .B2(
        n10008), .ZN(n8433) );
  OAI21_X1 U9545 ( .B1(n9588), .B2(n10442), .A(n8433), .ZN(n8446) );
  NAND2_X1 U9546 ( .A1(n9949), .A2(n9654), .ZN(n8435) );
  AND2_X1 U9547 ( .A1(n8434), .A2(n8435), .ZN(n8438) );
  INV_X1 U9548 ( .A(n8435), .ZN(n8437) );
  AOI21_X1 U9549 ( .B1(n8439), .B2(n8438), .A(n4908), .ZN(n8443) );
  INV_X1 U9550 ( .A(n8443), .ZN(n8441) );
  INV_X1 U9551 ( .A(n8453), .ZN(n8442) );
  AOI21_X1 U9552 ( .B1(n8444), .B2(n8443), .A(n8442), .ZN(n9946) );
  NOR2_X1 U9553 ( .A1(n9946), .A2(n9873), .ZN(n8445) );
  AOI211_X1 U9554 ( .C1(n9943), .C2(n10006), .A(n8446), .B(n8445), .ZN(n8447)
         );
  OAI21_X1 U9555 ( .B1(n9843), .B2(n9945), .A(n8447), .ZN(P1_U3274) );
  INV_X1 U9556 ( .A(n8448), .ZN(n8450) );
  XOR2_X1 U9557 ( .A(n8713), .B(n8454), .Z(n8460) );
  INV_X1 U9558 ( .A(n8784), .ZN(n9653) );
  OR2_X1 U9559 ( .A1(n9942), .A2(n9653), .ZN(n8452) );
  AND2_X1 U9560 ( .A1(n8455), .A2(n8454), .ZN(n8456) );
  NOR2_X1 U9561 ( .A1(n8731), .A2(n8456), .ZN(n9940) );
  NAND2_X1 U9562 ( .A1(n9940), .A2(n8457), .ZN(n8459) );
  AOI22_X1 U9563 ( .A1(n9849), .A2(n9866), .B1(n9864), .B2(n9653), .ZN(n8458)
         );
  OAI211_X1 U9564 ( .C1(n9780), .C2(n8460), .A(n8459), .B(n8458), .ZN(n9938)
         );
  INV_X1 U9565 ( .A(n9938), .ZN(n8466) );
  AND2_X1 U9566 ( .A1(n9627), .A2(n5319), .ZN(n8461) );
  OR2_X1 U9567 ( .A1(n8461), .A2(n9856), .ZN(n9937) );
  AOI22_X1 U9568 ( .A1(n9843), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9618), .B2(
        n10008), .ZN(n8463) );
  NAND2_X1 U9569 ( .A1(n9627), .A2(n9827), .ZN(n8462) );
  OAI211_X1 U9570 ( .C1(n9937), .C2(n10443), .A(n8463), .B(n8462), .ZN(n8464)
         );
  AOI21_X1 U9571 ( .B1(n9940), .B2(n10014), .A(n8464), .ZN(n8465) );
  OAI21_X1 U9572 ( .B1(n8466), .B2(n9843), .A(n8465), .ZN(P1_U3273) );
  OAI222_X1 U9573 ( .A1(P1_U3084), .A2(n4847), .B1(n7481), .B2(n8468), .C1(
        n8467), .C2(n8841), .ZN(P1_U3325) );
  INV_X1 U9574 ( .A(n8495), .ZN(n8875) );
  OAI222_X1 U9575 ( .A1(n7481), .A2(n8875), .B1(n8470), .B2(P1_U3084), .C1(
        n8469), .C2(n8841), .ZN(P1_U3323) );
  OR2_X1 U9576 ( .A1(n10574), .A2(n8471), .ZN(n9330) );
  NAND2_X1 U9577 ( .A1(n9474), .A2(n9344), .ZN(n9333) );
  NAND2_X1 U9578 ( .A1(n9467), .A2(n9063), .ZN(n8592) );
  NAND2_X1 U9579 ( .A1(n8593), .A2(n8592), .ZN(n9327) );
  INV_X1 U9580 ( .A(n8478), .ZN(n8472) );
  OR2_X1 U9581 ( .A1(n9477), .A2(n8477), .ZN(n9366) );
  OR2_X1 U9582 ( .A1(n9474), .A2(n9344), .ZN(n8589) );
  AND2_X1 U9583 ( .A1(n9366), .A2(n8589), .ZN(n9332) );
  NAND2_X1 U9584 ( .A1(n8474), .A2(n8473), .ZN(n9310) );
  OR2_X1 U9585 ( .A1(n9462), .A2(n9342), .ZN(n8481) );
  NAND2_X1 U9586 ( .A1(n9462), .A2(n9342), .ZN(n8475) );
  NAND2_X1 U9587 ( .A1(n8481), .A2(n8475), .ZN(n8848) );
  INV_X1 U9588 ( .A(n8476), .ZN(n8479) );
  NAND2_X1 U9589 ( .A1(n9477), .A2(n8477), .ZN(n9331) );
  AND2_X1 U9590 ( .A1(n9331), .A2(n8478), .ZN(n9335) );
  NAND2_X1 U9591 ( .A1(n9310), .A2(n8480), .ZN(n9311) );
  NAND2_X1 U9592 ( .A1(n9311), .A2(n8481), .ZN(n9295) );
  NAND2_X1 U9593 ( .A1(n9459), .A2(n9058), .ZN(n8604) );
  NAND2_X1 U9594 ( .A1(n9295), .A2(n9296), .ZN(n9294) );
  AND2_X1 U9595 ( .A1(n8652), .A2(n9272), .ZN(n8596) );
  NAND2_X1 U9596 ( .A1(n9452), .A2(n9256), .ZN(n8651) );
  NAND2_X1 U9597 ( .A1(n9447), .A2(n9043), .ZN(n8613) );
  NAND2_X1 U9598 ( .A1(n9442), .A2(n9257), .ZN(n8614) );
  NAND2_X1 U9599 ( .A1(n8618), .A2(n8614), .ZN(n8854) );
  NAND2_X1 U9600 ( .A1(n9236), .A2(n8618), .ZN(n9205) );
  NAND2_X1 U9601 ( .A1(n9431), .A2(n9186), .ZN(n8517) );
  AND2_X1 U9602 ( .A1(n9207), .A2(n9206), .ZN(n8484) );
  OAI21_X1 U9603 ( .B1(n9205), .B2(n9221), .A(n8484), .ZN(n8485) );
  NAND2_X1 U9604 ( .A1(n8485), .A2(n8624), .ZN(n9167) );
  NAND2_X1 U9605 ( .A1(n9195), .A2(n9087), .ZN(n8623) );
  INV_X1 U9606 ( .A(n8649), .ZN(n8486) );
  AND2_X1 U9607 ( .A1(n9185), .A2(n8486), .ZN(n8488) );
  INV_X1 U9608 ( .A(n8650), .ZN(n8487) );
  AND2_X1 U9609 ( .A1(n8487), .A2(n9168), .ZN(n8516) );
  NAND2_X1 U9610 ( .A1(n9416), .A2(n9069), .ZN(n8632) );
  INV_X1 U9611 ( .A(n9084), .ZN(n9156) );
  OR2_X1 U9612 ( .A1(n9410), .A2(n9156), .ZN(n8489) );
  NAND2_X1 U9613 ( .A1(n8490), .A2(n5561), .ZN(n8493) );
  OR2_X1 U9614 ( .A1(n8503), .A2(n8491), .ZN(n8492) );
  NAND2_X1 U9615 ( .A1(n9405), .A2(n8866), .ZN(n8639) );
  NOR2_X1 U9616 ( .A1(n8503), .A2(n8873), .ZN(n8494) );
  INV_X1 U9617 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U9618 ( .A1(n5436), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U9619 ( .A1(n8496), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8497) );
  OAI211_X1 U9620 ( .C1(n4846), .C2(n8499), .A(n8498), .B(n8497), .ZN(n9083)
         );
  AND2_X1 U9621 ( .A1(n8755), .A2(n9083), .ZN(n8636) );
  OAI22_X1 U9622 ( .A1(n8500), .A2(n8636), .B1(n8680), .B2(n8752), .ZN(n8502)
         );
  NAND2_X1 U9623 ( .A1(n8500), .A2(n8755), .ZN(n8501) );
  NAND2_X1 U9624 ( .A1(n8502), .A2(n8501), .ZN(n8508) );
  NAND2_X1 U9625 ( .A1(n9997), .A2(n5561), .ZN(n8505) );
  OR2_X1 U9626 ( .A1(n8503), .A2(n6819), .ZN(n8504) );
  INV_X1 U9627 ( .A(n8752), .ZN(n8646) );
  OR2_X1 U9628 ( .A1(n9398), .A2(n8646), .ZN(n8507) );
  INV_X1 U9629 ( .A(n8755), .ZN(n9401) );
  INV_X1 U9630 ( .A(n9083), .ZN(n8506) );
  NAND2_X1 U9631 ( .A1(n9401), .A2(n8506), .ZN(n8641) );
  NOR3_X1 U9632 ( .A1(n8509), .A2(n8510), .A3(n9143), .ZN(n8688) );
  INV_X1 U9633 ( .A(n8510), .ZN(n8512) );
  AOI21_X1 U9634 ( .B1(n8512), .B2(n9143), .A(n8511), .ZN(n8683) );
  NOR2_X1 U9635 ( .A1(n8513), .A2(n8636), .ZN(n8678) );
  INV_X1 U9636 ( .A(n8623), .ZN(n8514) );
  NOR2_X1 U9637 ( .A1(n8649), .A2(n8514), .ZN(n8515) );
  MUX2_X1 U9638 ( .A(n8516), .B(n8515), .S(n8637), .Z(n8631) );
  AND2_X1 U9639 ( .A1(n8517), .A2(n9206), .ZN(n8519) );
  AND2_X1 U9640 ( .A1(n8624), .A2(n8619), .ZN(n8518) );
  MUX2_X1 U9641 ( .A(n8519), .B(n8518), .S(n8637), .Z(n8622) );
  NAND2_X1 U9642 ( .A1(n8653), .A2(n8522), .ZN(n8520) );
  AND2_X1 U9643 ( .A1(n8654), .A2(n8520), .ZN(n8526) );
  NAND3_X1 U9644 ( .A1(n8653), .A2(n8522), .A3(n8521), .ZN(n8523) );
  NAND2_X1 U9645 ( .A1(n8524), .A2(n8523), .ZN(n8525) );
  MUX2_X1 U9646 ( .A(n8526), .B(n8525), .S(n8643), .Z(n8531) );
  MUX2_X1 U9647 ( .A(n8528), .B(n8527), .S(n8637), .Z(n8529) );
  OAI211_X1 U9648 ( .C1(n8531), .C2(n7395), .A(n8530), .B(n8529), .ZN(n8536)
         );
  MUX2_X1 U9649 ( .A(n8533), .B(n8532), .S(n8643), .Z(n8534) );
  NAND3_X1 U9650 ( .A1(n8536), .A2(n8535), .A3(n8534), .ZN(n8541) );
  MUX2_X1 U9651 ( .A(n8538), .B(n8537), .S(n8643), .Z(n8539) );
  NAND3_X1 U9652 ( .A1(n8541), .A2(n8540), .A3(n8539), .ZN(n8545) );
  MUX2_X1 U9653 ( .A(n8543), .B(n8542), .S(n8643), .Z(n8544) );
  INV_X1 U9654 ( .A(n8546), .ZN(n8661) );
  INV_X1 U9655 ( .A(n8548), .ZN(n8551) );
  MUX2_X1 U9656 ( .A(n8549), .B(n9098), .S(n8637), .Z(n8550) );
  MUX2_X1 U9657 ( .A(n8553), .B(n8552), .S(n8643), .Z(n8554) );
  INV_X1 U9658 ( .A(n8559), .ZN(n8556) );
  NAND2_X1 U9659 ( .A1(n8557), .A2(n8566), .ZN(n8570) );
  NAND2_X1 U9660 ( .A1(n8559), .A2(n8558), .ZN(n8562) );
  NAND2_X1 U9661 ( .A1(n8571), .A2(n8560), .ZN(n8561) );
  AOI21_X1 U9662 ( .B1(n8566), .B2(n8562), .A(n8561), .ZN(n8568) );
  AND2_X1 U9663 ( .A1(n8825), .A2(n9096), .ZN(n8565) );
  NAND2_X1 U9664 ( .A1(n8573), .A2(n8563), .ZN(n8564) );
  MUX2_X1 U9665 ( .A(n8568), .B(n8567), .S(n8643), .Z(n8569) );
  NAND3_X1 U9666 ( .A1(n8570), .A2(n8668), .A3(n8569), .ZN(n8580) );
  NAND2_X1 U9667 ( .A1(n8575), .A2(n8571), .ZN(n8572) );
  NAND2_X1 U9668 ( .A1(n8572), .A2(n8574), .ZN(n8578) );
  NAND2_X1 U9669 ( .A1(n8574), .A2(n8573), .ZN(n8576) );
  NAND2_X1 U9670 ( .A1(n8576), .A2(n8575), .ZN(n8577) );
  MUX2_X1 U9671 ( .A(n8578), .B(n8577), .S(n8637), .Z(n8579) );
  INV_X1 U9672 ( .A(n8671), .ZN(n8584) );
  MUX2_X1 U9673 ( .A(n8582), .B(n8581), .S(n8637), .Z(n8583) );
  NAND2_X1 U9674 ( .A1(n9366), .A2(n9331), .ZN(n9386) );
  INV_X1 U9675 ( .A(n9386), .ZN(n9377) );
  NAND2_X1 U9676 ( .A1(n10574), .A2(n8643), .ZN(n8586) );
  OR2_X1 U9677 ( .A1(n10574), .A2(n8643), .ZN(n8585) );
  MUX2_X1 U9678 ( .A(n8586), .B(n8585), .S(n9389), .Z(n8587) );
  MUX2_X1 U9679 ( .A(n9366), .B(n9331), .S(n8637), .Z(n8588) );
  MUX2_X1 U9680 ( .A(n8589), .B(n9333), .S(n8643), .Z(n8590) );
  NAND3_X1 U9681 ( .A1(n8591), .A2(n9339), .A3(n8590), .ZN(n8595) );
  MUX2_X1 U9682 ( .A(n8593), .B(n8592), .S(n8637), .Z(n8594) );
  NAND2_X1 U9683 ( .A1(n8595), .A2(n8594), .ZN(n8598) );
  INV_X1 U9684 ( .A(n9342), .ZN(n9089) );
  MUX2_X1 U9685 ( .A(n9089), .B(n9462), .S(n8637), .Z(n8597) );
  INV_X1 U9686 ( .A(n8597), .ZN(n8600) );
  INV_X1 U9687 ( .A(n8598), .ZN(n8599) );
  NAND3_X1 U9688 ( .A1(n9296), .A2(n8600), .A3(n8599), .ZN(n8601) );
  NAND2_X1 U9689 ( .A1(n8602), .A2(n8601), .ZN(n8607) );
  NAND3_X1 U9690 ( .A1(n8603), .A2(n9462), .A3(n9272), .ZN(n8605) );
  NAND3_X1 U9691 ( .A1(n8605), .A2(n8651), .A3(n8604), .ZN(n8606) );
  AOI22_X1 U9692 ( .A1(n8607), .A2(n8613), .B1(n8643), .B2(n8606), .ZN(n8609)
         );
  NOR2_X1 U9693 ( .A1(n8651), .A2(n8643), .ZN(n8608) );
  OAI211_X1 U9694 ( .C1(n8609), .C2(n8608), .A(n8618), .B(n8610), .ZN(n8617)
         );
  NAND2_X1 U9695 ( .A1(n8610), .A2(n8652), .ZN(n8611) );
  NAND2_X1 U9696 ( .A1(n8611), .A2(n8643), .ZN(n8612) );
  AND2_X1 U9697 ( .A1(n8614), .A2(n8612), .ZN(n8616) );
  AOI21_X1 U9698 ( .B1(n8614), .B2(n8613), .A(n8637), .ZN(n8615) );
  AOI21_X1 U9699 ( .B1(n8619), .B2(n8618), .A(n8637), .ZN(n8621) );
  INV_X1 U9700 ( .A(n9206), .ZN(n8620) );
  INV_X1 U9701 ( .A(n9431), .ZN(n9204) );
  AND2_X1 U9702 ( .A1(n8623), .A2(n8643), .ZN(n8627) );
  OAI211_X1 U9703 ( .C1(n9218), .C2(n8643), .A(n8625), .B(n8624), .ZN(n8626)
         );
  OAI21_X1 U9704 ( .B1(n8628), .B2(n8627), .A(n8626), .ZN(n8630) );
  MUX2_X1 U9705 ( .A(n8649), .B(n8650), .S(n8637), .Z(n8629) );
  MUX2_X1 U9706 ( .A(n8633), .B(n8632), .S(n8643), .Z(n8634) );
  NAND3_X1 U9707 ( .A1(n9410), .A2(n9156), .A3(n8637), .ZN(n8635) );
  INV_X1 U9708 ( .A(n8636), .ZN(n8642) );
  MUX2_X1 U9709 ( .A(n8639), .B(n8638), .S(n8637), .Z(n8640) );
  INV_X1 U9710 ( .A(n9398), .ZN(n8645) );
  MUX2_X1 U9711 ( .A(n8752), .B(n9398), .S(n8643), .Z(n8644) );
  AOI21_X1 U9712 ( .B1(n8646), .B2(n8645), .A(n8644), .ZN(n8647) );
  INV_X1 U9713 ( .A(n8859), .ZN(n9169) );
  NAND2_X1 U9714 ( .A1(n8652), .A2(n8651), .ZN(n9273) );
  INV_X1 U9715 ( .A(n9368), .ZN(n9358) );
  AND2_X1 U9716 ( .A1(n8654), .A2(n8653), .ZN(n10473) );
  NAND4_X1 U9717 ( .A1(n8655), .A2(n10453), .A3(n10473), .A4(n8687), .ZN(n8659) );
  NOR4_X1 U9718 ( .A1(n8659), .A2(n8658), .A3(n8657), .A4(n8656), .ZN(n8662)
         );
  NAND4_X1 U9719 ( .A1(n8662), .A2(n8661), .A3(n7948), .A4(n8660), .ZN(n8666)
         );
  NOR4_X1 U9720 ( .A1(n8666), .A2(n8665), .A3(n8664), .A4(n8663), .ZN(n8667)
         );
  NAND3_X1 U9721 ( .A1(n8669), .A2(n8668), .A3(n8667), .ZN(n8670) );
  NOR4_X1 U9722 ( .A1(n9358), .A2(n8671), .A3(n9386), .A4(n8670), .ZN(n8672)
         );
  NAND4_X1 U9723 ( .A1(n9296), .A2(n9312), .A3(n9339), .A4(n8672), .ZN(n8673)
         );
  NOR4_X1 U9724 ( .A1(n9221), .A2(n9255), .A3(n9273), .A4(n8673), .ZN(n8674)
         );
  NAND4_X1 U9725 ( .A1(n9185), .A2(n9207), .A3(n9237), .A4(n8674), .ZN(n8675)
         );
  NOR4_X1 U9726 ( .A1(n8886), .A2(n9169), .A3(n9154), .A4(n8675), .ZN(n8676)
         );
  NAND4_X1 U9727 ( .A1(n8678), .A2(n8677), .A3(n8676), .A4(n8876), .ZN(n8679)
         );
  XNOR2_X1 U9728 ( .A(n8679), .B(n9180), .ZN(n8681) );
  OAI211_X1 U9729 ( .C1(n8685), .C2(n8687), .A(n8681), .B(n8680), .ZN(n8682)
         );
  NOR4_X1 U9730 ( .A1(n8690), .A2(n9343), .A3(n8689), .A4(n8749), .ZN(n8693)
         );
  OAI21_X1 U9731 ( .B1(n8694), .B2(n8691), .A(P2_B_REG_SCAN_IN), .ZN(n8692) );
  INV_X1 U9732 ( .A(n8695), .ZN(n8696) );
  AOI21_X1 U9733 ( .B1(n8698), .B2(n8697), .A(n8696), .ZN(n10400) );
  OAI22_X1 U9734 ( .A1(n9613), .A2(n10441), .B1(n9623), .B2(n8699), .ZN(n8700)
         );
  AOI21_X1 U9735 ( .B1(n8701), .B2(P1_REG3_REG_0__SCAN_IN), .A(n8700), .ZN(
        n8702) );
  OAI21_X1 U9736 ( .B1(n10400), .B2(n9649), .A(n8702), .ZN(P1_U3230) );
  INV_X1 U9737 ( .A(n9878), .ZN(n9710) );
  INV_X1 U9738 ( .A(n9931), .ZN(n9862) );
  NAND2_X1 U9739 ( .A1(n9710), .A2(n9709), .ZN(n9708) );
  INV_X1 U9740 ( .A(P1_B_REG_SCAN_IN), .ZN(n8705) );
  OR2_X1 U9741 ( .A1(n4848), .A2(n8705), .ZN(n8706) );
  NAND2_X1 U9742 ( .A1(n9866), .A2(n8706), .ZN(n9722) );
  NOR2_X1 U9743 ( .A1(n8707), .A2(n9722), .ZN(n9877) );
  NAND2_X1 U9744 ( .A1(n9877), .A2(n10447), .ZN(n9711) );
  OAI21_X1 U9745 ( .B1(n10447), .B2(n8708), .A(n9711), .ZN(n8709) );
  AOI21_X1 U9746 ( .B1(n9874), .B2(n9827), .A(n8709), .ZN(n8710) );
  OAI21_X1 U9747 ( .B1(n9876), .B2(n10443), .A(n8710), .ZN(P1_U3261) );
  NAND2_X1 U9748 ( .A1(n9804), .A2(n9805), .ZN(n9803) );
  NAND2_X1 U9749 ( .A1(n9803), .A2(n8718), .ZN(n9778) );
  NAND2_X1 U9750 ( .A1(n9778), .A2(n9788), .ZN(n8720) );
  NAND2_X1 U9751 ( .A1(n8720), .A2(n8719), .ZN(n9771) );
  NAND2_X1 U9752 ( .A1(n9771), .A2(n9770), .ZN(n8722) );
  OAI21_X1 U9753 ( .B1(n8726), .B2(n8727), .A(n9719), .ZN(n8728) );
  INV_X1 U9754 ( .A(n9744), .ZN(n9772) );
  INV_X1 U9755 ( .A(n9608), .ZN(n9850) );
  NOR2_X1 U9756 ( .A1(n9931), .A2(n9849), .ZN(n8732) );
  INV_X1 U9757 ( .A(n8813), .ZN(n9867) );
  NAND2_X1 U9758 ( .A1(n8734), .A2(n4916), .ZN(n9789) );
  NAND2_X1 U9759 ( .A1(n8738), .A2(n8737), .ZN(n9716) );
  OAI21_X1 U9760 ( .B1(n8738), .B2(n8737), .A(n9716), .ZN(n9890) );
  OAI22_X1 U9761 ( .A1(n8956), .A2(n10450), .B1(n8739), .B2(n10447), .ZN(n8740) );
  AOI21_X1 U9762 ( .B1(n9885), .B2(n9827), .A(n8740), .ZN(n8744) );
  INV_X1 U9763 ( .A(n9737), .ZN(n8741) );
  NAND2_X1 U9764 ( .A1(n9885), .A2(n8741), .ZN(n8742) );
  NAND2_X1 U9765 ( .A1(n9886), .A2(n10006), .ZN(n8743) );
  OAI211_X1 U9766 ( .C1(n9890), .C2(n9873), .A(n8744), .B(n8743), .ZN(n8745)
         );
  INV_X1 U9767 ( .A(n8745), .ZN(n8746) );
  OAI21_X1 U9768 ( .B1(n9843), .B2(n9888), .A(n8746), .ZN(P1_U3263) );
  INV_X1 U9769 ( .A(n9459), .ZN(n9289) );
  INV_X1 U9770 ( .A(n9452), .ZN(n9271) );
  INV_X1 U9771 ( .A(n9437), .ZN(n9229) );
  OAI21_X1 U9772 ( .B1(n8755), .B2(n8883), .A(n8836), .ZN(n9404) );
  NAND2_X1 U9773 ( .A1(n9393), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8754) );
  INV_X1 U9774 ( .A(n8749), .ZN(n8750) );
  NAND2_X1 U9775 ( .A1(n8750), .A2(P2_B_REG_SCAN_IN), .ZN(n8751) );
  AND2_X1 U9776 ( .A1(n9390), .A2(n8751), .ZN(n8889) );
  NAND2_X1 U9777 ( .A1(n8752), .A2(n8889), .ZN(n9403) );
  NOR2_X1 U9778 ( .A1(n9393), .A2(n9403), .ZN(n8838) );
  INV_X1 U9779 ( .A(n8838), .ZN(n8753) );
  OAI211_X1 U9780 ( .C1(n8755), .C2(n10475), .A(n8754), .B(n8753), .ZN(n8756)
         );
  INV_X1 U9781 ( .A(n8756), .ZN(n8757) );
  OAI21_X1 U9782 ( .B1(n9404), .B2(n10472), .A(n8757), .ZN(P2_U3266) );
  NAND2_X1 U9783 ( .A1(n8762), .A2(n8761), .ZN(n8768) );
  NAND2_X1 U9784 ( .A1(n8768), .A2(n8769), .ZN(n8764) );
  NAND2_X1 U9785 ( .A1(n9958), .A2(n8936), .ZN(n8759) );
  OR2_X1 U9786 ( .A1(n8765), .A2(n8949), .ZN(n8758) );
  NAND2_X1 U9787 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  XNOR2_X1 U9788 ( .A(n8760), .B(n4840), .ZN(n8766) );
  NOR2_X1 U9789 ( .A1(n8762), .A2(n8761), .ZN(n8770) );
  INV_X1 U9790 ( .A(n8770), .ZN(n8763) );
  NAND3_X1 U9791 ( .A1(n8764), .A2(n8766), .A3(n8763), .ZN(n9520) );
  OAI22_X1 U9792 ( .A1(n5064), .A2(n8949), .B1(n8765), .B2(n8236), .ZN(n9522)
         );
  INV_X1 U9793 ( .A(n8766), .ZN(n8767) );
  OAI211_X1 U9794 ( .C1(n8770), .C2(n8769), .A(n8768), .B(n8767), .ZN(n9519)
         );
  INV_X1 U9795 ( .A(n9519), .ZN(n8771) );
  AOI22_X1 U9796 ( .A1(n9952), .A2(n8936), .B1(n8943), .B2(n9655), .ZN(n8772)
         );
  INV_X1 U9797 ( .A(n9952), .ZN(n8773) );
  OAI22_X1 U9798 ( .A1(n8773), .A2(n8949), .B1(n9569), .B2(n8236), .ZN(n9640)
         );
  NAND2_X1 U9799 ( .A1(n9949), .A2(n8936), .ZN(n8775) );
  OR2_X1 U9800 ( .A1(n9582), .A2(n8949), .ZN(n8774) );
  NAND2_X1 U9801 ( .A1(n8775), .A2(n8774), .ZN(n8776) );
  XNOR2_X1 U9802 ( .A(n8776), .B(n4841), .ZN(n8779) );
  NOR2_X1 U9803 ( .A1(n9582), .A2(n8236), .ZN(n8777) );
  AOI21_X1 U9804 ( .B1(n9949), .B2(n8898), .A(n8777), .ZN(n8778) );
  NAND2_X1 U9805 ( .A1(n8779), .A2(n8778), .ZN(n9575) );
  OR2_X1 U9806 ( .A1(n8779), .A2(n8778), .ZN(n8780) );
  AND2_X1 U9807 ( .A1(n9575), .A2(n8780), .ZN(n9564) );
  NAND2_X1 U9808 ( .A1(n9563), .A2(n9575), .ZN(n8791) );
  NAND2_X1 U9809 ( .A1(n9942), .A2(n8936), .ZN(n8782) );
  NAND2_X1 U9810 ( .A1(n9653), .A2(n8943), .ZN(n8781) );
  NAND2_X1 U9811 ( .A1(n8782), .A2(n8781), .ZN(n8783) );
  XNOR2_X1 U9812 ( .A(n8783), .B(n4841), .ZN(n8786) );
  NOR2_X1 U9813 ( .A1(n8784), .A2(n8236), .ZN(n8785) );
  AOI21_X1 U9814 ( .B1(n9942), .B2(n8898), .A(n8785), .ZN(n8787) );
  NAND2_X1 U9815 ( .A1(n8786), .A2(n8787), .ZN(n8792) );
  INV_X1 U9816 ( .A(n8786), .ZN(n8789) );
  INV_X1 U9817 ( .A(n8787), .ZN(n8788) );
  NAND2_X1 U9818 ( .A1(n8789), .A2(n8788), .ZN(n8790) );
  AND2_X1 U9819 ( .A1(n8792), .A2(n8790), .ZN(n9576) );
  NAND2_X1 U9820 ( .A1(n8791), .A2(n9576), .ZN(n9579) );
  NAND2_X1 U9821 ( .A1(n9579), .A2(n8792), .ZN(n8795) );
  AOI22_X1 U9822 ( .A1(n9627), .A2(n8936), .B1(n8898), .B2(n9865), .ZN(n8793)
         );
  XNOR2_X1 U9823 ( .A(n8793), .B(n8947), .ZN(n8796) );
  INV_X1 U9824 ( .A(n9627), .ZN(n9936) );
  OAI22_X1 U9825 ( .A1(n9936), .A2(n8949), .B1(n8794), .B2(n8236), .ZN(n9617)
         );
  NAND2_X1 U9826 ( .A1(n9931), .A2(n8936), .ZN(n8798) );
  NAND2_X1 U9827 ( .A1(n9849), .A2(n8943), .ZN(n8797) );
  NAND2_X1 U9828 ( .A1(n8798), .A2(n8797), .ZN(n8799) );
  XNOR2_X1 U9829 ( .A(n8799), .B(n4841), .ZN(n8802) );
  AND2_X1 U9830 ( .A1(n9849), .A2(n8925), .ZN(n8800) );
  AOI21_X1 U9831 ( .B1(n9931), .B2(n8898), .A(n8800), .ZN(n8801) );
  NOR2_X1 U9832 ( .A1(n8802), .A2(n8801), .ZN(n8811) );
  OAI22_X1 U9833 ( .A1(n9846), .A2(n8950), .B1(n8813), .B2(n7096), .ZN(n8803)
         );
  XNOR2_X1 U9834 ( .A(n8803), .B(n8947), .ZN(n8905) );
  OAI22_X1 U9835 ( .A1(n9846), .A2(n8949), .B1(n8813), .B2(n8236), .ZN(n8904)
         );
  XNOR2_X1 U9836 ( .A(n8905), .B(n8904), .ZN(n8804) );
  XNOR2_X1 U9837 ( .A(n8908), .B(n8804), .ZN(n8809) );
  AOI22_X1 U9838 ( .A1(n9850), .A2(n9642), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8806) );
  NAND2_X1 U9839 ( .A1(n9619), .A2(n9844), .ZN(n8805) );
  OAI211_X1 U9840 ( .C1(n9624), .C2(n9607), .A(n8806), .B(n8805), .ZN(n8807)
         );
  AOI21_X1 U9841 ( .B1(n9926), .B2(n4839), .A(n8807), .ZN(n8808) );
  OAI21_X1 U9842 ( .B1(n8809), .B2(n9649), .A(n8808), .ZN(P1_U3231) );
  NOR2_X1 U9843 ( .A1(n8811), .A2(n4922), .ZN(n8812) );
  XNOR2_X1 U9844 ( .A(n8810), .B(n8812), .ZN(n8818) );
  NAND2_X1 U9845 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9703) );
  OAI21_X1 U9846 ( .B1(n8813), .B2(n9623), .A(n9703), .ZN(n8814) );
  AOI21_X1 U9847 ( .B1(n9641), .B2(n9865), .A(n8814), .ZN(n8815) );
  OAI21_X1 U9848 ( .B1(n9646), .B2(n9859), .A(n8815), .ZN(n8816) );
  AOI21_X1 U9849 ( .B1(n9931), .B2(n4839), .A(n8816), .ZN(n8817) );
  OAI21_X1 U9850 ( .B1(n8818), .B2(n9649), .A(n8817), .ZN(P1_U3217) );
  XNOR2_X1 U9851 ( .A(n8819), .B(n8832), .ZN(n8821) );
  AOI21_X1 U9852 ( .B1(n8821), .B2(n10467), .A(n8820), .ZN(n10524) );
  OAI22_X1 U9853 ( .A1(n9373), .A2(n8823), .B1(n8822), .B2(n10471), .ZN(n8828)
         );
  OAI211_X1 U9854 ( .C1(n8826), .C2(n8825), .A(n10576), .B(n8824), .ZN(n10522)
         );
  NOR2_X1 U9855 ( .A1(n10522), .A2(n9356), .ZN(n8827) );
  AOI211_X1 U9856 ( .C1(n9353), .C2(n10520), .A(n8828), .B(n8827), .ZN(n8835)
         );
  NAND2_X1 U9857 ( .A1(n8831), .A2(n8829), .ZN(n10519) );
  NAND2_X1 U9858 ( .A1(n8831), .A2(n8830), .ZN(n8833) );
  NAND2_X1 U9859 ( .A1(n8833), .A2(n8832), .ZN(n10518) );
  NAND3_X1 U9860 ( .A1(n10519), .A2(n10518), .A3(n9224), .ZN(n8834) );
  OAI211_X1 U9861 ( .C1(n10524), .C2(n9393), .A(n8835), .B(n8834), .ZN(
        P2_U3288) );
  NOR2_X1 U9862 ( .A1(n9373), .A2(n8837), .ZN(n8839) );
  AOI211_X1 U9863 ( .C1(n9398), .C2(n9353), .A(n8839), .B(n8838), .ZN(n8840)
         );
  OAI21_X1 U9864 ( .B1(n9400), .B2(n10472), .A(n8840), .ZN(P2_U3265) );
  OAI222_X1 U9865 ( .A1(n7125), .A2(P1_U3084), .B1(n7481), .B2(n8842), .C1(
        n8841), .C2(n6171), .ZN(P1_U3331) );
  OR2_X1 U9866 ( .A1(n10574), .A2(n9389), .ZN(n8844) );
  NAND2_X1 U9867 ( .A1(n8845), .A2(n8844), .ZN(n9376) );
  OR2_X1 U9868 ( .A1(n9477), .A2(n9090), .ZN(n8846) );
  INV_X1 U9869 ( .A(n9063), .ZN(n9315) );
  OR2_X1 U9870 ( .A1(n9368), .A2(n5320), .ZN(n9301) );
  OR2_X1 U9871 ( .A1(n9301), .A2(n4868), .ZN(n9281) );
  INV_X1 U9872 ( .A(n9344), .ZN(n9391) );
  NAND2_X1 U9873 ( .A1(n9474), .A2(n9391), .ZN(n9324) );
  AND2_X1 U9874 ( .A1(n9327), .A2(n9324), .ZN(n9325) );
  OR2_X1 U9875 ( .A1(n5320), .A2(n9325), .ZN(n9302) );
  AND2_X1 U9876 ( .A1(n8848), .A2(n9302), .ZN(n8849) );
  INV_X1 U9877 ( .A(n9058), .ZN(n9314) );
  NAND2_X1 U9878 ( .A1(n9459), .A2(n9314), .ZN(n8850) );
  NAND2_X1 U9879 ( .A1(n9284), .A2(n8850), .ZN(n9265) );
  NAND2_X1 U9880 ( .A1(n9452), .A2(n9088), .ZN(n8851) );
  OR2_X1 U9881 ( .A1(n9447), .A2(n9275), .ZN(n8852) );
  NAND2_X1 U9882 ( .A1(n9246), .A2(n8852), .ZN(n9233) );
  NOR2_X1 U9883 ( .A1(n9442), .A2(n9219), .ZN(n8853) );
  NAND2_X1 U9884 ( .A1(n9437), .A2(n9209), .ZN(n8855) );
  OR2_X1 U9885 ( .A1(n9431), .A2(n9218), .ZN(n8857) );
  NAND2_X1 U9886 ( .A1(n9198), .A2(n8857), .ZN(n9182) );
  XNOR2_X1 U9887 ( .A(n8877), .B(n5152), .ZN(n9409) );
  INV_X1 U9888 ( .A(n8880), .ZN(n8860) );
  AOI21_X1 U9889 ( .B1(n9410), .B2(n9149), .A(n8860), .ZN(n9411) );
  AOI22_X1 U9890 ( .A1(n8861), .A2(n9382), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9164), .ZN(n8862) );
  OAI21_X1 U9891 ( .B1(n8863), .B2(n10475), .A(n8862), .ZN(n8871) );
  INV_X1 U9892 ( .A(n8864), .ZN(n8865) );
  AOI21_X1 U9893 ( .B1(n8865), .B2(n5152), .A(n9371), .ZN(n8869) );
  OAI22_X1 U9894 ( .A1(n9069), .A2(n9343), .B1(n8866), .B2(n9341), .ZN(n8867)
         );
  AOI21_X1 U9895 ( .B1(n8869), .B2(n8868), .A(n8867), .ZN(n9412) );
  NOR2_X1 U9896 ( .A1(n9412), .A2(n9393), .ZN(n8870) );
  AOI211_X1 U9897 ( .C1(n9396), .C2(n9411), .A(n8871), .B(n8870), .ZN(n8872)
         );
  OAI21_X1 U9898 ( .B1(n9409), .B2(n10476), .A(n8872), .ZN(P2_U3268) );
  XNOR2_X1 U9899 ( .A(n8879), .B(n8878), .ZN(n9408) );
  AOI22_X1 U9900 ( .A1(n8884), .A2(n9382), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9164), .ZN(n8885) );
  OAI21_X1 U9901 ( .B1(n8881), .B2(n10475), .A(n8885), .ZN(n8892) );
  XNOR2_X1 U9902 ( .A(n8887), .B(n8886), .ZN(n8888) );
  INV_X1 U9903 ( .A(n8889), .ZN(n8890) );
  NOR2_X1 U9904 ( .A1(n9407), .A2(n9164), .ZN(n8891) );
  OAI21_X1 U9906 ( .B1(n9408), .B2(n10476), .A(n8893), .ZN(P2_U3267) );
  NOR2_X1 U9907 ( .A1(n8905), .A2(n8904), .ZN(n9542) );
  NAND2_X1 U9908 ( .A1(n9922), .A2(n8936), .ZN(n8895) );
  NAND2_X1 U9909 ( .A1(n9850), .A2(n8943), .ZN(n8894) );
  NAND2_X1 U9910 ( .A1(n8895), .A2(n8894), .ZN(n8896) );
  XNOR2_X1 U9911 ( .A(n8896), .B(n4840), .ZN(n8903) );
  NOR2_X1 U9912 ( .A1(n9608), .A2(n8195), .ZN(n8897) );
  AOI21_X1 U9913 ( .B1(n9922), .B2(n8898), .A(n8897), .ZN(n8902) );
  NAND2_X1 U9914 ( .A1(n8903), .A2(n8902), .ZN(n9548) );
  INV_X1 U9915 ( .A(n9548), .ZN(n8906) );
  OR2_X1 U9916 ( .A1(n9542), .A2(n8906), .ZN(n9598) );
  OAI22_X1 U9917 ( .A1(n9816), .A2(n8949), .B1(n9536), .B2(n8236), .ZN(n8909)
         );
  NAND2_X1 U9918 ( .A1(n9916), .A2(n8936), .ZN(n8900) );
  NAND2_X1 U9919 ( .A1(n9831), .A2(n8898), .ZN(n8899) );
  NAND2_X1 U9920 ( .A1(n8900), .A2(n8899), .ZN(n8901) );
  XNOR2_X1 U9921 ( .A(n8901), .B(n8947), .ZN(n8910) );
  XOR2_X1 U9922 ( .A(n8909), .B(n8910), .Z(n9603) );
  NAND2_X1 U9923 ( .A1(n8905), .A2(n8904), .ZN(n9544) );
  AND2_X1 U9924 ( .A1(n5316), .A2(n9544), .ZN(n9543) );
  OAI21_X1 U9925 ( .B1(n8908), .B2(n9598), .A(n8907), .ZN(n9601) );
  NAND2_X1 U9926 ( .A1(n9601), .A2(n8911), .ZN(n8913) );
  OAI22_X1 U9927 ( .A1(n9802), .A2(n8950), .B1(n9781), .B2(n7096), .ZN(n8912)
         );
  XOR2_X1 U9928 ( .A(n8947), .B(n8912), .Z(n8914) );
  OAI22_X1 U9929 ( .A1(n9802), .A2(n8949), .B1(n9781), .B2(n8195), .ZN(n9534)
         );
  OAI22_X1 U9930 ( .A1(n8917), .A2(n8950), .B1(n8916), .B2(n7096), .ZN(n8915)
         );
  XNOR2_X1 U9931 ( .A(n8915), .B(n8947), .ZN(n8918) );
  OAI22_X1 U9932 ( .A1(n8917), .A2(n8949), .B1(n8916), .B2(n8236), .ZN(n8919)
         );
  XNOR2_X1 U9933 ( .A(n8918), .B(n8919), .ZN(n9590) );
  INV_X1 U9934 ( .A(n8918), .ZN(n8921) );
  INV_X1 U9935 ( .A(n8919), .ZN(n8920) );
  NAND2_X1 U9936 ( .A1(n9901), .A2(n8936), .ZN(n8923) );
  NAND2_X1 U9937 ( .A1(n9759), .A2(n8943), .ZN(n8922) );
  NAND2_X1 U9938 ( .A1(n8923), .A2(n8922), .ZN(n8924) );
  XNOR2_X1 U9939 ( .A(n8924), .B(n8947), .ZN(n9556) );
  NAND2_X1 U9940 ( .A1(n9901), .A2(n8943), .ZN(n8927) );
  NAND2_X1 U9941 ( .A1(n9759), .A2(n8925), .ZN(n8926) );
  NAND2_X1 U9942 ( .A1(n8927), .A2(n8926), .ZN(n9555) );
  NOR2_X1 U9943 ( .A1(n9556), .A2(n9555), .ZN(n8930) );
  INV_X1 U9944 ( .A(n9556), .ZN(n8929) );
  INV_X1 U9945 ( .A(n9555), .ZN(n8928) );
  OAI22_X1 U9946 ( .A1(n9756), .A2(n8949), .B1(n9744), .B2(n8195), .ZN(n8932)
         );
  OAI22_X1 U9947 ( .A1(n9756), .A2(n8950), .B1(n9744), .B2(n8949), .ZN(n8931)
         );
  XNOR2_X1 U9948 ( .A(n8931), .B(n8947), .ZN(n8933) );
  XOR2_X1 U9949 ( .A(n8932), .B(n8933), .Z(n9630) );
  NAND2_X1 U9950 ( .A1(n9631), .A2(n9630), .ZN(n8935) );
  NAND2_X1 U9951 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  NAND2_X1 U9952 ( .A1(n9891), .A2(n8936), .ZN(n8938) );
  NAND2_X1 U9953 ( .A1(n5243), .A2(n8943), .ZN(n8937) );
  NAND2_X1 U9954 ( .A1(n8938), .A2(n8937), .ZN(n8940) );
  XNOR2_X1 U9955 ( .A(n8940), .B(n4840), .ZN(n8945) );
  NOR2_X1 U9956 ( .A1(n8941), .A2(n8195), .ZN(n8942) );
  AOI21_X1 U9957 ( .B1(n9891), .B2(n8943), .A(n8942), .ZN(n8944) );
  NAND2_X1 U9958 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  OAI21_X1 U9959 ( .B1(n8945), .B2(n8944), .A(n8946), .ZN(n9511) );
  OAI22_X1 U9960 ( .A1(n9715), .A2(n8949), .B1(n9745), .B2(n8236), .ZN(n8948)
         );
  XNOR2_X1 U9961 ( .A(n8948), .B(n8947), .ZN(n8952) );
  OAI22_X1 U9962 ( .A1(n9715), .A2(n8950), .B1(n9745), .B2(n8949), .ZN(n8951)
         );
  XNOR2_X1 U9963 ( .A(n8954), .B(n8953), .ZN(n8962) );
  OAI22_X1 U9964 ( .A1(n8956), .A2(n9646), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8955), .ZN(n8957) );
  AOI21_X1 U9965 ( .B1(n9641), .B2(n5243), .A(n8957), .ZN(n8958) );
  OAI21_X1 U9966 ( .B1(n8959), .B2(n9623), .A(n8958), .ZN(n8960) );
  AOI21_X1 U9967 ( .B1(n9885), .B2(n4839), .A(n8960), .ZN(n8961) );
  OAI21_X1 U9968 ( .B1(n8962), .B2(n9649), .A(n8961), .ZN(P1_U3218) );
  XNOR2_X1 U9969 ( .A(n8963), .B(n8964), .ZN(n8969) );
  AOI22_X1 U9970 ( .A1(n9151), .A2(n9074), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8966) );
  NAND2_X1 U9971 ( .A1(n9086), .A2(n9039), .ZN(n8965) );
  OAI211_X1 U9972 ( .C1(n9156), .C2(n9059), .A(n8966), .B(n8965), .ZN(n8967)
         );
  AOI21_X1 U9973 ( .B1(n9416), .B2(n9079), .A(n8967), .ZN(n8968) );
  OAI21_X1 U9974 ( .B1(n8969), .B2(n9081), .A(n8968), .ZN(P2_U3216) );
  OR2_X1 U9975 ( .A1(n8970), .A2(n9049), .ZN(n9047) );
  NAND2_X1 U9976 ( .A1(n9047), .A2(n8971), .ZN(n8973) );
  XNOR2_X1 U9977 ( .A(n8973), .B(n8972), .ZN(n8975) );
  XNOR2_X1 U9978 ( .A(n8975), .B(n8974), .ZN(n8981) );
  NAND2_X1 U9979 ( .A1(n9039), .A2(n9219), .ZN(n8978) );
  INV_X1 U9980 ( .A(n8976), .ZN(n9227) );
  AOI22_X1 U9981 ( .A1(n9074), .A2(n9227), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8977) );
  OAI211_X1 U9982 ( .C1(n9186), .C2(n9059), .A(n8978), .B(n8977), .ZN(n8979)
         );
  AOI21_X1 U9983 ( .B1(n9437), .B2(n9079), .A(n8979), .ZN(n8980) );
  OAI21_X1 U9984 ( .B1(n8981), .B2(n9081), .A(n8980), .ZN(P2_U3218) );
  NAND2_X1 U9985 ( .A1(n8982), .A2(n8983), .ZN(n8984) );
  NAND2_X1 U9986 ( .A1(n8984), .A2(n8985), .ZN(n9036) );
  OAI21_X1 U9987 ( .B1(n8985), .B2(n8984), .A(n9036), .ZN(n8986) );
  NAND2_X1 U9988 ( .A1(n8986), .A2(n9009), .ZN(n8990) );
  INV_X1 U9989 ( .A(n9290), .ZN(n8988) );
  NOR2_X1 U9990 ( .A1(n10188), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9141) );
  AOI22_X1 U9991 ( .A1(n9088), .A2(n9390), .B1(n9089), .B2(n9388), .ZN(n9297)
         );
  NOR2_X1 U9992 ( .A1(n9076), .A2(n9297), .ZN(n8987) );
  AOI211_X1 U9993 ( .C1(n8988), .C2(n9074), .A(n9141), .B(n8987), .ZN(n8989)
         );
  OAI211_X1 U9994 ( .C1(n9289), .C2(n9016), .A(n8990), .B(n8989), .ZN(P2_U3221) );
  XNOR2_X1 U9995 ( .A(n8991), .B(n8992), .ZN(n8998) );
  NAND2_X1 U9996 ( .A1(n9039), .A2(n9088), .ZN(n8995) );
  INV_X1 U9997 ( .A(n8993), .ZN(n9251) );
  AOI22_X1 U9998 ( .A1(n9074), .A2(n9251), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8994) );
  OAI211_X1 U9999 ( .C1(n9257), .C2(n9059), .A(n8995), .B(n8994), .ZN(n8996)
         );
  AOI21_X1 U10000 ( .B1(n9447), .B2(n9079), .A(n8996), .ZN(n8997) );
  OAI21_X1 U10001 ( .B1(n8998), .B2(n9081), .A(n8997), .ZN(P2_U3225) );
  XNOR2_X1 U10002 ( .A(n8999), .B(n9000), .ZN(n9005) );
  AOI22_X1 U10003 ( .A1(n9194), .A2(n9074), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n9002) );
  NAND2_X1 U10004 ( .A1(n9039), .A2(n9218), .ZN(n9001) );
  OAI211_X1 U10005 ( .C1(n9187), .C2(n9059), .A(n9002), .B(n9001), .ZN(n9003)
         );
  AOI21_X1 U10006 ( .B1(n9195), .B2(n9079), .A(n9003), .ZN(n9004) );
  OAI21_X1 U10007 ( .B1(n9005), .B2(n9081), .A(n9004), .ZN(P2_U3227) );
  INV_X1 U10008 ( .A(n9474), .ZN(n9360) );
  OAI21_X1 U10009 ( .B1(n9008), .B2(n9007), .A(n9006), .ZN(n9010) );
  NAND2_X1 U10010 ( .A1(n9010), .A2(n9009), .ZN(n9015) );
  INV_X1 U10011 ( .A(n9361), .ZN(n9013) );
  AOI22_X1 U10012 ( .A1(n9388), .A2(n9090), .B1(n9315), .B2(n9390), .ZN(n9370)
         );
  NOR2_X1 U10013 ( .A1(n9076), .A2(n9370), .ZN(n9011) );
  AOI211_X1 U10014 ( .C1(n9013), .C2(n9074), .A(n9012), .B(n9011), .ZN(n9014)
         );
  OAI211_X1 U10015 ( .C1(n9360), .C2(n9016), .A(n9015), .B(n9014), .ZN(
        P2_U3228) );
  XNOR2_X1 U10016 ( .A(n9018), .B(n9017), .ZN(n9026) );
  NAND2_X1 U10017 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9114) );
  INV_X1 U10018 ( .A(n9114), .ZN(n9021) );
  NOR2_X1 U10019 ( .A1(n9019), .A2(n9351), .ZN(n9020) );
  AOI211_X1 U10020 ( .C1(n9022), .C2(n9089), .A(n9021), .B(n9020), .ZN(n9023)
         );
  OAI21_X1 U10021 ( .B1(n9344), .B2(n9062), .A(n9023), .ZN(n9024) );
  AOI21_X1 U10022 ( .B1(n9467), .B2(n9079), .A(n9024), .ZN(n9025) );
  OAI21_X1 U10023 ( .B1(n9026), .B2(n9081), .A(n9025), .ZN(P2_U3230) );
  XNOR2_X1 U10024 ( .A(n9028), .B(n9027), .ZN(n9034) );
  NAND2_X1 U10025 ( .A1(n9039), .A2(n9209), .ZN(n9031) );
  INV_X1 U10026 ( .A(n9029), .ZN(n9202) );
  AOI22_X1 U10027 ( .A1(n9074), .A2(n9202), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n9030) );
  OAI211_X1 U10028 ( .C1(n9087), .C2(n9059), .A(n9031), .B(n9030), .ZN(n9032)
         );
  AOI21_X1 U10029 ( .B1(n9431), .B2(n9079), .A(n9032), .ZN(n9033) );
  OAI21_X1 U10030 ( .B1(n9034), .B2(n9081), .A(n9033), .ZN(P2_U3231) );
  NAND2_X1 U10031 ( .A1(n9036), .A2(n9035), .ZN(n9038) );
  XNOR2_X1 U10032 ( .A(n9038), .B(n9037), .ZN(n9046) );
  NAND2_X1 U10033 ( .A1(n9039), .A2(n9314), .ZN(n9042) );
  INV_X1 U10034 ( .A(n9040), .ZN(n9269) );
  AOI22_X1 U10035 ( .A1(n9074), .A2(n9269), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n9041) );
  OAI211_X1 U10036 ( .C1(n9043), .C2(n9059), .A(n9042), .B(n9041), .ZN(n9044)
         );
  AOI21_X1 U10037 ( .B1(n9452), .B2(n9079), .A(n9044), .ZN(n9045) );
  OAI21_X1 U10038 ( .B1(n9046), .B2(n9081), .A(n9045), .ZN(P2_U3235) );
  INV_X1 U10039 ( .A(n9047), .ZN(n9048) );
  AOI21_X1 U10040 ( .B1(n8970), .B2(n9049), .A(n9048), .ZN(n9053) );
  AOI22_X1 U10041 ( .A1(n9209), .A2(n9390), .B1(n9388), .B2(n9275), .ZN(n9239)
         );
  AOI22_X1 U10042 ( .A1(n9074), .A2(n9241), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n9050) );
  OAI21_X1 U10043 ( .B1(n9239), .B2(n9076), .A(n9050), .ZN(n9051) );
  AOI21_X1 U10044 ( .B1(n9442), .B2(n9079), .A(n9051), .ZN(n9052) );
  OAI21_X1 U10045 ( .B1(n9053), .B2(n9081), .A(n9052), .ZN(P2_U3237) );
  INV_X1 U10046 ( .A(n8982), .ZN(n9054) );
  AOI21_X1 U10047 ( .B1(n9056), .B2(n9055), .A(n9054), .ZN(n9066) );
  INV_X1 U10048 ( .A(n9057), .ZN(n9306) );
  NOR2_X1 U10049 ( .A1(n10104), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9127) );
  NOR2_X1 U10050 ( .A1(n9059), .A2(n9058), .ZN(n9060) );
  AOI211_X1 U10051 ( .C1(n9306), .C2(n9074), .A(n9127), .B(n9060), .ZN(n9061)
         );
  OAI21_X1 U10052 ( .B1(n9063), .B2(n9062), .A(n9061), .ZN(n9064) );
  AOI21_X1 U10053 ( .B1(n9462), .B2(n9079), .A(n9064), .ZN(n9065) );
  OAI21_X1 U10054 ( .B1(n9066), .B2(n9081), .A(n9065), .ZN(P2_U3240) );
  XNOR2_X1 U10055 ( .A(n9067), .B(n9068), .ZN(n9082) );
  OR2_X1 U10056 ( .A1(n9069), .A2(n9341), .ZN(n9071) );
  OR2_X1 U10057 ( .A1(n9087), .A2(n9343), .ZN(n9070) );
  NAND2_X1 U10058 ( .A1(n9071), .A2(n9070), .ZN(n9171) );
  INV_X1 U10059 ( .A(n9171), .ZN(n9077) );
  INV_X1 U10060 ( .A(n9072), .ZN(n9165) );
  AOI22_X1 U10061 ( .A1(n9165), .A2(n9074), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n9075) );
  OAI21_X1 U10062 ( .B1(n9077), .B2(n9076), .A(n9075), .ZN(n9078) );
  AOI21_X1 U10063 ( .B1(n9422), .B2(n9079), .A(n9078), .ZN(n9080) );
  OAI21_X1 U10064 ( .B1(n9082), .B2(n9081), .A(n9080), .ZN(P2_U3242) );
  MUX2_X1 U10065 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9083), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10066 ( .A(n9084), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9104), .Z(
        P2_U3580) );
  MUX2_X1 U10067 ( .A(n9085), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9104), .Z(
        P2_U3579) );
  MUX2_X1 U10068 ( .A(n9086), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9104), .Z(
        P2_U3578) );
  INV_X1 U10069 ( .A(n9087), .ZN(n9210) );
  MUX2_X1 U10070 ( .A(n9210), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9104), .Z(
        P2_U3577) );
  MUX2_X1 U10071 ( .A(n9209), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9104), .Z(
        P2_U3575) );
  MUX2_X1 U10072 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9088), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10073 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9314), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10074 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9089), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10075 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9315), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10076 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9391), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10077 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9090), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10078 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9389), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10079 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9091), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10080 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9092), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10081 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9093), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10082 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9094), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10083 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n9095), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10084 ( .A(n9096), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9104), .Z(
        P2_U3560) );
  MUX2_X1 U10085 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n9097), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10086 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n9098), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10087 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n9099), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10088 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9100), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10089 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9101), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n9102), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10091 ( .A(n9103), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9104), .Z(
        P2_U3553) );
  MUX2_X1 U10092 ( .A(n9105), .B(P2_DATAO_REG_0__SCAN_IN), .S(n9104), .Z(
        P2_U3552) );
  OAI21_X1 U10093 ( .B1(n9110), .B2(P2_REG1_REG_16__SCAN_IN), .A(n9106), .ZN(
        n9108) );
  XNOR2_X1 U10094 ( .A(n9124), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9107) );
  NOR2_X1 U10095 ( .A1(n9107), .A2(n9108), .ZN(n9123) );
  AOI211_X1 U10096 ( .C1(n9108), .C2(n9107), .A(n9123), .B(n10357), .ZN(n9120)
         );
  AOI21_X1 U10097 ( .B1(n9110), .B2(P2_REG2_REG_16__SCAN_IN), .A(n9109), .ZN(
        n9113) );
  NAND2_X1 U10098 ( .A1(n9124), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9111) );
  OAI21_X1 U10099 ( .B1(n9124), .B2(P2_REG2_REG_17__SCAN_IN), .A(n9111), .ZN(
        n9112) );
  NOR2_X1 U10100 ( .A1(n9113), .A2(n9112), .ZN(n9121) );
  AOI211_X1 U10101 ( .C1(n9113), .C2(n9112), .A(n9121), .B(n10394), .ZN(n9119)
         );
  INV_X1 U10102 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U10103 ( .A1(n10386), .A2(n9124), .ZN(n9115) );
  OAI211_X1 U10104 ( .C1(n9117), .C2(n9116), .A(n9115), .B(n9114), .ZN(n9118)
         );
  OR3_X1 U10105 ( .A1(n9120), .A2(n9119), .A3(n9118), .ZN(P2_U3262) );
  INV_X1 U10106 ( .A(n9122), .ZN(n9136) );
  XNOR2_X1 U10107 ( .A(n9122), .B(n9135), .ZN(n9138) );
  AOI21_X1 U10108 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9124), .A(n9121), .ZN(
        n9137) );
  XNOR2_X1 U10109 ( .A(n9138), .B(n9137), .ZN(n9126) );
  XNOR2_X1 U10110 ( .A(n9122), .B(n9130), .ZN(n9132) );
  AOI21_X1 U10111 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9124), .A(n9123), .ZN(
        n9131) );
  XNOR2_X1 U10112 ( .A(n9132), .B(n9131), .ZN(n9125) );
  AOI22_X1 U10113 ( .A1(n10359), .A2(n9126), .B1(n10391), .B2(n9125), .ZN(
        n9129) );
  AOI21_X1 U10114 ( .B1(n10379), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n9127), .ZN(
        n9128) );
  OAI211_X1 U10115 ( .C1(n9136), .C2(n10356), .A(n9129), .B(n9128), .ZN(
        P2_U3263) );
  AOI22_X1 U10116 ( .A1(n9132), .A2(n9131), .B1(n9136), .B2(n9130), .ZN(n9134)
         );
  XNOR2_X1 U10117 ( .A(n9143), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9133) );
  XNOR2_X1 U10118 ( .A(n9134), .B(n9133), .ZN(n9147) );
  MUX2_X1 U10119 ( .A(n9291), .B(P2_REG2_REG_19__SCAN_IN), .S(n9143), .Z(n9140) );
  AOI22_X1 U10120 ( .A1(n9138), .A2(n9137), .B1(n9136), .B2(n9135), .ZN(n9139)
         );
  XOR2_X1 U10121 ( .A(n9140), .B(n9139), .Z(n9145) );
  AOI21_X1 U10122 ( .B1(n10379), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n9141), .ZN(
        n9142) );
  OAI21_X1 U10123 ( .B1(n10356), .B2(n9143), .A(n9142), .ZN(n9144) );
  AOI21_X1 U10124 ( .B1(n10359), .B2(n9145), .A(n9144), .ZN(n9146) );
  OAI21_X1 U10125 ( .B1(n10357), .B2(n9147), .A(n9146), .ZN(P2_U3264) );
  XOR2_X1 U10126 ( .A(n9154), .B(n9148), .Z(n9420) );
  INV_X1 U10127 ( .A(n4876), .ZN(n9150) );
  AOI21_X1 U10128 ( .B1(n9416), .B2(n9150), .A(n5176), .ZN(n9417) );
  AOI22_X1 U10129 ( .A1(n9151), .A2(n9382), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9164), .ZN(n9152) );
  OAI21_X1 U10130 ( .B1(n9153), .B2(n10475), .A(n9152), .ZN(n9161) );
  AOI21_X1 U10131 ( .B1(n9155), .B2(n9154), .A(n9371), .ZN(n9159) );
  OAI22_X1 U10132 ( .A1(n9156), .A2(n9341), .B1(n9187), .B2(n9343), .ZN(n9157)
         );
  AOI21_X1 U10133 ( .B1(n9159), .B2(n9158), .A(n9157), .ZN(n9419) );
  NOR2_X1 U10134 ( .A1(n9419), .A2(n9393), .ZN(n9160) );
  AOI211_X1 U10135 ( .C1(n9396), .C2(n9417), .A(n9161), .B(n9160), .ZN(n9162)
         );
  OAI21_X1 U10136 ( .B1(n9420), .B2(n10476), .A(n9162), .ZN(P2_U3269) );
  XNOR2_X1 U10137 ( .A(n9163), .B(n9169), .ZN(n9425) );
  AOI211_X1 U10138 ( .C1(n9422), .C2(n9178), .A(n10568), .B(n4876), .ZN(n9421)
         );
  AOI22_X1 U10139 ( .A1(n9165), .A2(n9382), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n9164), .ZN(n9166) );
  OAI21_X1 U10140 ( .B1(n5257), .B2(n10475), .A(n9166), .ZN(n9174) );
  NAND2_X1 U10141 ( .A1(n9167), .A2(n9185), .ZN(n9184) );
  NAND2_X1 U10142 ( .A1(n9184), .A2(n9168), .ZN(n9170) );
  XNOR2_X1 U10143 ( .A(n9170), .B(n9169), .ZN(n9172) );
  NOR2_X1 U10144 ( .A1(n9424), .A2(n9393), .ZN(n9173) );
  AOI211_X1 U10145 ( .C1(n9421), .C2(n9365), .A(n9174), .B(n9173), .ZN(n9175)
         );
  OAI21_X1 U10146 ( .B1(n9425), .B2(n10476), .A(n9175), .ZN(P2_U3270) );
  INV_X1 U10147 ( .A(n9176), .ZN(n9177) );
  AOI21_X1 U10148 ( .B1(n9177), .B2(n9195), .A(n10568), .ZN(n9179) );
  NAND2_X1 U10149 ( .A1(n9179), .A2(n9178), .ZN(n9426) );
  NOR2_X1 U10150 ( .A1(n9426), .A2(n9180), .ZN(n9193) );
  XNOR2_X1 U10151 ( .A(n9182), .B(n9181), .ZN(n9183) );
  INV_X1 U10152 ( .A(n10564), .ZN(n10581) );
  NAND2_X1 U10153 ( .A1(n9183), .A2(n10581), .ZN(n9192) );
  OAI211_X1 U10154 ( .C1(n9185), .C2(n9167), .A(n9184), .B(n10467), .ZN(n9190)
         );
  OAI22_X1 U10155 ( .A1(n9187), .A2(n9341), .B1(n9186), .B2(n9343), .ZN(n9188)
         );
  INV_X1 U10156 ( .A(n9188), .ZN(n9189) );
  AND2_X1 U10157 ( .A1(n9190), .A2(n9189), .ZN(n9191) );
  NAND2_X1 U10158 ( .A1(n9192), .A2(n9191), .ZN(n9428) );
  AOI211_X1 U10159 ( .C1(n9382), .C2(n9194), .A(n9193), .B(n9428), .ZN(n9197)
         );
  AOI22_X1 U10160 ( .A1(n9195), .A2(n9353), .B1(n9393), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9196) );
  OAI21_X1 U10161 ( .B1(n9197), .B2(n9393), .A(n9196), .ZN(P2_U3271) );
  INV_X1 U10162 ( .A(n9198), .ZN(n9199) );
  AOI21_X1 U10163 ( .B1(n9207), .B2(n9200), .A(n9199), .ZN(n9435) );
  XNOR2_X1 U10164 ( .A(n9201), .B(n9204), .ZN(n9432) );
  AOI22_X1 U10165 ( .A1(n9393), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9202), .B2(
        n9382), .ZN(n9203) );
  OAI21_X1 U10166 ( .B1(n9204), .B2(n10475), .A(n9203), .ZN(n9213) );
  OR2_X1 U10167 ( .A1(n9205), .A2(n9221), .ZN(n9215) );
  NAND2_X1 U10168 ( .A1(n9215), .A2(n9206), .ZN(n9208) );
  XNOR2_X1 U10169 ( .A(n9208), .B(n9207), .ZN(n9211) );
  AOI222_X1 U10170 ( .A1(n10467), .A2(n9211), .B1(n9210), .B2(n9390), .C1(
        n9209), .C2(n9388), .ZN(n9434) );
  NOR2_X1 U10171 ( .A1(n9434), .A2(n9393), .ZN(n9212) );
  AOI211_X1 U10172 ( .C1(n9432), .C2(n9396), .A(n9213), .B(n9212), .ZN(n9214)
         );
  OAI21_X1 U10173 ( .B1(n9435), .B2(n10476), .A(n9214), .ZN(P2_U3272) );
  INV_X1 U10174 ( .A(n9205), .ZN(n9217) );
  INV_X1 U10175 ( .A(n9221), .ZN(n9216) );
  OAI21_X1 U10176 ( .B1(n9217), .B2(n9216), .A(n9215), .ZN(n9220) );
  AOI222_X1 U10177 ( .A1(n10467), .A2(n9220), .B1(n9219), .B2(n9388), .C1(
        n9218), .C2(n9390), .ZN(n9440) );
  OR2_X1 U10178 ( .A1(n9222), .A2(n9221), .ZN(n9436) );
  NAND3_X1 U10179 ( .A1(n9436), .A2(n9223), .A3(n9224), .ZN(n9232) );
  INV_X1 U10180 ( .A(n9234), .ZN(n9226) );
  INV_X1 U10181 ( .A(n9201), .ZN(n9225) );
  AOI21_X1 U10182 ( .B1(n9437), .B2(n9226), .A(n9225), .ZN(n9438) );
  AOI22_X1 U10183 ( .A1(n9393), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9227), .B2(
        n9382), .ZN(n9228) );
  OAI21_X1 U10184 ( .B1(n9229), .B2(n10475), .A(n9228), .ZN(n9230) );
  AOI21_X1 U10185 ( .B1(n9438), .B2(n9396), .A(n9230), .ZN(n9231) );
  OAI211_X1 U10186 ( .C1(n9164), .C2(n9440), .A(n9232), .B(n9231), .ZN(
        P2_U3273) );
  XNOR2_X1 U10187 ( .A(n9233), .B(n9237), .ZN(n9446) );
  AOI21_X1 U10188 ( .B1(n9442), .B2(n5317), .A(n9234), .ZN(n9443) );
  INV_X1 U10189 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9235) );
  OAI22_X1 U10190 ( .A1(n5172), .A2(n10475), .B1(n9373), .B2(n9235), .ZN(n9244) );
  OAI211_X1 U10191 ( .C1(n9238), .C2(n9237), .A(n9236), .B(n10467), .ZN(n9240)
         );
  NAND2_X1 U10192 ( .A1(n9241), .A2(n9382), .ZN(n9242) );
  AOI21_X1 U10193 ( .B1(n9445), .B2(n9242), .A(n9393), .ZN(n9243) );
  AOI211_X1 U10194 ( .C1(n9443), .C2(n9396), .A(n9244), .B(n9243), .ZN(n9245)
         );
  OAI21_X1 U10195 ( .B1(n9446), .B2(n10476), .A(n9245), .ZN(P2_U3274) );
  INV_X1 U10196 ( .A(n9246), .ZN(n9247) );
  AOI21_X1 U10197 ( .B1(n9249), .B2(n9248), .A(n9247), .ZN(n9451) );
  INV_X1 U10198 ( .A(n5317), .ZN(n9250) );
  AOI21_X1 U10199 ( .B1(n9447), .B2(n9266), .A(n9250), .ZN(n9448) );
  INV_X1 U10200 ( .A(n9447), .ZN(n9253) );
  AOI22_X1 U10201 ( .A1(n9164), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9251), .B2(
        n9382), .ZN(n9252) );
  OAI21_X1 U10202 ( .B1(n9253), .B2(n10475), .A(n9252), .ZN(n9262) );
  AOI21_X1 U10203 ( .B1(n9254), .B2(n9255), .A(n9371), .ZN(n9260) );
  OAI22_X1 U10204 ( .A1(n9257), .A2(n9341), .B1(n9256), .B2(n9343), .ZN(n9258)
         );
  AOI21_X1 U10205 ( .B1(n9260), .B2(n9259), .A(n9258), .ZN(n9450) );
  NOR2_X1 U10206 ( .A1(n9450), .A2(n9393), .ZN(n9261) );
  AOI211_X1 U10207 ( .C1(n9448), .C2(n9396), .A(n9262), .B(n9261), .ZN(n9263)
         );
  OAI21_X1 U10208 ( .B1(n9451), .B2(n10476), .A(n9263), .ZN(P2_U3275) );
  OAI21_X1 U10209 ( .B1(n9265), .B2(n9273), .A(n9264), .ZN(n9456) );
  INV_X1 U10210 ( .A(n9287), .ZN(n9268) );
  INV_X1 U10211 ( .A(n9266), .ZN(n9267) );
  AOI21_X1 U10212 ( .B1(n9452), .B2(n9268), .A(n9267), .ZN(n9453) );
  AOI22_X1 U10213 ( .A1(n9164), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9269), .B2(
        n9382), .ZN(n9270) );
  OAI21_X1 U10214 ( .B1(n9271), .B2(n10475), .A(n9270), .ZN(n9278) );
  NAND2_X1 U10215 ( .A1(n9294), .A2(n9272), .ZN(n9274) );
  XNOR2_X1 U10216 ( .A(n9274), .B(n9273), .ZN(n9276) );
  AOI222_X1 U10217 ( .A1(n10467), .A2(n9276), .B1(n9275), .B2(n9390), .C1(
        n9314), .C2(n9388), .ZN(n9455) );
  NOR2_X1 U10218 ( .A1(n9455), .A2(n9393), .ZN(n9277) );
  AOI211_X1 U10219 ( .C1(n9453), .C2(n9396), .A(n9278), .B(n9277), .ZN(n9279)
         );
  OAI21_X1 U10220 ( .B1(n10476), .B2(n9456), .A(n9279), .ZN(P2_U3276) );
  OR2_X1 U10221 ( .A1(n9280), .A2(n9281), .ZN(n9283) );
  NAND2_X1 U10222 ( .A1(n9283), .A2(n9282), .ZN(n9286) );
  INV_X1 U10223 ( .A(n9296), .ZN(n9285) );
  OAI21_X1 U10224 ( .B1(n9286), .B2(n9285), .A(n9284), .ZN(n9461) );
  INV_X1 U10225 ( .A(n9305), .ZN(n9288) );
  AOI211_X1 U10226 ( .C1(n9459), .C2(n9288), .A(n10568), .B(n9287), .ZN(n9458)
         );
  NOR2_X1 U10227 ( .A1(n9289), .A2(n10475), .ZN(n9293) );
  OAI22_X1 U10228 ( .A1(n9373), .A2(n9291), .B1(n9290), .B2(n10471), .ZN(n9292) );
  AOI211_X1 U10229 ( .C1(n9458), .C2(n9365), .A(n9293), .B(n9292), .ZN(n9300)
         );
  OAI211_X1 U10230 ( .C1(n9296), .C2(n9295), .A(n9294), .B(n10467), .ZN(n9298)
         );
  NAND2_X1 U10231 ( .A1(n9298), .A2(n9297), .ZN(n9457) );
  NAND2_X1 U10232 ( .A1(n9457), .A2(n9373), .ZN(n9299) );
  OAI211_X1 U10233 ( .C1(n9461), .C2(n10476), .A(n9300), .B(n9299), .ZN(
        P2_U3277) );
  OR2_X1 U10234 ( .A1(n9280), .A2(n9301), .ZN(n9303) );
  AND2_X1 U10235 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  XNOR2_X1 U10236 ( .A(n9304), .B(n9312), .ZN(n9466) );
  AOI21_X1 U10237 ( .B1(n9462), .B2(n9322), .A(n9305), .ZN(n9463) );
  INV_X1 U10238 ( .A(n9462), .ZN(n9308) );
  AOI22_X1 U10239 ( .A1(n9164), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9306), .B2(
        n9382), .ZN(n9307) );
  OAI21_X1 U10240 ( .B1(n9308), .B2(n10475), .A(n9307), .ZN(n9319) );
  AND2_X1 U10241 ( .A1(n9310), .A2(n9309), .ZN(n9313) );
  OAI211_X1 U10242 ( .C1(n9313), .C2(n9312), .A(n9311), .B(n10467), .ZN(n9317)
         );
  AOI22_X1 U10243 ( .A1(n9388), .A2(n9315), .B1(n9314), .B2(n9390), .ZN(n9316)
         );
  NOR2_X1 U10244 ( .A1(n9465), .A2(n9393), .ZN(n9318) );
  AOI211_X1 U10245 ( .C1(n9463), .C2(n9396), .A(n9319), .B(n9318), .ZN(n9320)
         );
  OAI21_X1 U10246 ( .B1(n9466), .B2(n10476), .A(n9320), .ZN(P2_U3278) );
  AOI21_X1 U10247 ( .B1(n5161), .B2(n9467), .A(n10568), .ZN(n9323) );
  NAND2_X1 U10248 ( .A1(n9323), .A2(n9322), .ZN(n9469) );
  AND2_X1 U10249 ( .A1(n9357), .A2(n9324), .ZN(n9328) );
  NAND2_X1 U10250 ( .A1(n9357), .A2(n9325), .ZN(n9326) );
  OAI21_X1 U10251 ( .B1(n9328), .B2(n9327), .A(n9326), .ZN(n9329) );
  NAND2_X1 U10252 ( .A1(n9329), .A2(n10581), .ZN(n9349) );
  NAND2_X1 U10253 ( .A1(n9387), .A2(n9331), .ZN(n9367) );
  NAND2_X1 U10254 ( .A1(n9367), .A2(n9332), .ZN(n9334) );
  AND2_X1 U10255 ( .A1(n9334), .A2(n9333), .ZN(n9340) );
  NAND2_X1 U10256 ( .A1(n9387), .A2(n9335), .ZN(n9337) );
  AND2_X1 U10257 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  OAI211_X1 U10258 ( .C1(n9340), .C2(n9339), .A(n9338), .B(n10467), .ZN(n9347)
         );
  OAI22_X1 U10259 ( .A1(n9344), .A2(n9343), .B1(n9342), .B2(n9341), .ZN(n9345)
         );
  INV_X1 U10260 ( .A(n9345), .ZN(n9346) );
  AND2_X1 U10261 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  NAND2_X1 U10262 ( .A1(n9349), .A2(n9348), .ZN(n9471) );
  NAND2_X1 U10263 ( .A1(n9471), .A2(n9373), .ZN(n9355) );
  NAND2_X1 U10264 ( .A1(n9393), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9350) );
  OAI21_X1 U10265 ( .B1(n10471), .B2(n9351), .A(n9350), .ZN(n9352) );
  AOI21_X1 U10266 ( .B1(n9467), .B2(n9353), .A(n9352), .ZN(n9354) );
  OAI211_X1 U10267 ( .C1(n9469), .C2(n9356), .A(n9355), .B(n9354), .ZN(
        P2_U3279) );
  INV_X1 U10268 ( .A(n9280), .ZN(n9359) );
  OAI21_X1 U10269 ( .B1(n9359), .B2(n9358), .A(n9357), .ZN(n9476) );
  AOI211_X1 U10270 ( .C1(n9474), .C2(n9379), .A(n10568), .B(n9321), .ZN(n9473)
         );
  NOR2_X1 U10271 ( .A1(n9360), .A2(n10475), .ZN(n9364) );
  INV_X1 U10272 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9362) );
  OAI22_X1 U10273 ( .A1(n9373), .A2(n9362), .B1(n9361), .B2(n10471), .ZN(n9363) );
  AOI211_X1 U10274 ( .C1(n9473), .C2(n9365), .A(n9364), .B(n9363), .ZN(n9375)
         );
  NAND2_X1 U10275 ( .A1(n9367), .A2(n9366), .ZN(n9369) );
  XNOR2_X1 U10276 ( .A(n9369), .B(n9368), .ZN(n9372) );
  OAI21_X1 U10277 ( .B1(n9372), .B2(n9371), .A(n9370), .ZN(n9472) );
  NAND2_X1 U10278 ( .A1(n9472), .A2(n9373), .ZN(n9374) );
  OAI211_X1 U10279 ( .C1(n9476), .C2(n10476), .A(n9375), .B(n9374), .ZN(
        P2_U3280) );
  XNOR2_X1 U10280 ( .A(n9376), .B(n9377), .ZN(n9481) );
  INV_X1 U10281 ( .A(n9378), .ZN(n9381) );
  INV_X1 U10282 ( .A(n9379), .ZN(n9380) );
  AOI21_X1 U10283 ( .B1(n9477), .B2(n9381), .A(n9380), .ZN(n9478) );
  AOI22_X1 U10284 ( .A1(n9393), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9383), .B2(
        n9382), .ZN(n9384) );
  OAI21_X1 U10285 ( .B1(n9385), .B2(n10475), .A(n9384), .ZN(n9395) );
  XNOR2_X1 U10286 ( .A(n9387), .B(n9386), .ZN(n9392) );
  AOI222_X1 U10287 ( .A1(n10467), .A2(n9392), .B1(n9391), .B2(n9390), .C1(
        n9389), .C2(n9388), .ZN(n9480) );
  NOR2_X1 U10288 ( .A1(n9480), .A2(n9393), .ZN(n9394) );
  AOI211_X1 U10289 ( .C1(n9478), .C2(n9396), .A(n9395), .B(n9394), .ZN(n9397)
         );
  OAI21_X1 U10290 ( .B1(n9481), .B2(n10476), .A(n9397), .ZN(P2_U3281) );
  NAND2_X1 U10291 ( .A1(n9398), .A2(n10575), .ZN(n9399) );
  MUX2_X1 U10292 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9482), .S(n10584), .Z(
        P2_U3551) );
  NAND2_X1 U10293 ( .A1(n9401), .A2(n10575), .ZN(n9402) );
  OAI211_X1 U10294 ( .C1(n9404), .C2(n10568), .A(n9403), .B(n9402), .ZN(n9483)
         );
  MUX2_X1 U10295 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9483), .S(n10584), .Z(
        P2_U3550) );
  MUX2_X1 U10296 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9484), .S(n10584), .Z(
        P2_U3549) );
  AOI22_X1 U10297 ( .A1(n9411), .A2(n10576), .B1(n10575), .B2(n9410), .ZN(
        n9413) );
  NAND2_X1 U10298 ( .A1(n9415), .A2(n9414), .ZN(n9485) );
  MUX2_X1 U10299 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9485), .S(n10584), .Z(
        P2_U3548) );
  AOI22_X1 U10300 ( .A1(n9417), .A2(n10576), .B1(n10575), .B2(n9416), .ZN(
        n9418) );
  OAI211_X1 U10301 ( .C1(n9420), .C2(n10564), .A(n9419), .B(n9418), .ZN(n9486)
         );
  MUX2_X1 U10302 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9486), .S(n10584), .Z(
        P2_U3547) );
  AOI21_X1 U10303 ( .B1(n10575), .B2(n9422), .A(n9421), .ZN(n9423) );
  OAI211_X1 U10304 ( .C1(n9425), .C2(n10564), .A(n9424), .B(n9423), .ZN(n9487)
         );
  MUX2_X1 U10305 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9487), .S(n10584), .Z(
        P2_U3546) );
  INV_X1 U10306 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9429) );
  OAI21_X1 U10307 ( .B1(n8748), .B2(n10566), .A(n9426), .ZN(n9427) );
  NOR2_X1 U10308 ( .A1(n9428), .A2(n9427), .ZN(n9488) );
  MUX2_X1 U10309 ( .A(n9429), .B(n9488), .S(n10584), .Z(n9430) );
  INV_X1 U10310 ( .A(n9430), .ZN(P2_U3545) );
  AOI22_X1 U10311 ( .A1(n9432), .A2(n10576), .B1(n10575), .B2(n9431), .ZN(
        n9433) );
  OAI211_X1 U10312 ( .C1(n9435), .C2(n10564), .A(n9434), .B(n9433), .ZN(n9491)
         );
  MUX2_X1 U10313 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9491), .S(n10584), .Z(
        P2_U3544) );
  NAND3_X1 U10314 ( .A1(n9436), .A2(n10581), .A3(n9223), .ZN(n9441) );
  AOI22_X1 U10315 ( .A1(n9438), .A2(n10576), .B1(n10575), .B2(n9437), .ZN(
        n9439) );
  NAND3_X1 U10316 ( .A1(n9441), .A2(n9440), .A3(n9439), .ZN(n9492) );
  MUX2_X1 U10317 ( .A(n9492), .B(P2_REG1_REG_23__SCAN_IN), .S(n10583), .Z(
        P2_U3543) );
  AOI22_X1 U10318 ( .A1(n9443), .A2(n10576), .B1(n10575), .B2(n9442), .ZN(
        n9444) );
  OAI211_X1 U10319 ( .C1(n9446), .C2(n10564), .A(n9445), .B(n9444), .ZN(n9493)
         );
  MUX2_X1 U10320 ( .A(n9493), .B(P2_REG1_REG_22__SCAN_IN), .S(n10583), .Z(
        P2_U3542) );
  AOI22_X1 U10321 ( .A1(n9448), .A2(n10576), .B1(n10575), .B2(n9447), .ZN(
        n9449) );
  OAI211_X1 U10322 ( .C1(n9451), .C2(n10564), .A(n9450), .B(n9449), .ZN(n9494)
         );
  MUX2_X1 U10323 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9494), .S(n10584), .Z(
        P2_U3541) );
  AOI22_X1 U10324 ( .A1(n9453), .A2(n10576), .B1(n10575), .B2(n9452), .ZN(
        n9454) );
  OAI211_X1 U10325 ( .C1(n9456), .C2(n10564), .A(n9455), .B(n9454), .ZN(n9495)
         );
  MUX2_X1 U10326 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9495), .S(n10584), .Z(
        P2_U3540) );
  AOI211_X1 U10327 ( .C1(n10575), .C2(n9459), .A(n9458), .B(n9457), .ZN(n9460)
         );
  OAI21_X1 U10328 ( .B1(n9461), .B2(n10564), .A(n9460), .ZN(n9496) );
  MUX2_X1 U10329 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9496), .S(n10584), .Z(
        P2_U3539) );
  AOI22_X1 U10330 ( .A1(n9463), .A2(n10576), .B1(n10575), .B2(n9462), .ZN(
        n9464) );
  OAI211_X1 U10331 ( .C1(n9466), .C2(n10564), .A(n9465), .B(n9464), .ZN(n9497)
         );
  MUX2_X1 U10332 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9497), .S(n10584), .Z(
        P2_U3538) );
  NAND2_X1 U10333 ( .A1(n9467), .A2(n10575), .ZN(n9468) );
  NAND2_X1 U10334 ( .A1(n9469), .A2(n9468), .ZN(n9470) );
  MUX2_X1 U10335 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9498), .S(n10584), .Z(
        P2_U3537) );
  AOI211_X1 U10336 ( .C1(n10575), .C2(n9474), .A(n9473), .B(n9472), .ZN(n9475)
         );
  OAI21_X1 U10337 ( .B1(n9476), .B2(n10564), .A(n9475), .ZN(n9499) );
  MUX2_X1 U10338 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9499), .S(n10584), .Z(
        P2_U3536) );
  AOI22_X1 U10339 ( .A1(n9478), .A2(n10576), .B1(n10575), .B2(n9477), .ZN(
        n9479) );
  OAI211_X1 U10340 ( .C1(n9481), .C2(n10564), .A(n9480), .B(n9479), .ZN(n9500)
         );
  MUX2_X1 U10341 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9500), .S(n10584), .Z(
        P2_U3535) );
  MUX2_X1 U10342 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9482), .S(n10588), .Z(
        P2_U3519) );
  MUX2_X1 U10343 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9483), .S(n10588), .Z(
        P2_U3518) );
  MUX2_X1 U10344 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9484), .S(n10588), .Z(
        P2_U3517) );
  MUX2_X1 U10345 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9485), .S(n10588), .Z(
        P2_U3516) );
  MUX2_X1 U10346 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9486), .S(n10588), .Z(
        P2_U3515) );
  MUX2_X1 U10347 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9487), .S(n10588), .Z(
        P2_U3514) );
  INV_X1 U10348 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9489) );
  MUX2_X1 U10349 ( .A(n9489), .B(n9488), .S(n10588), .Z(n9490) );
  INV_X1 U10350 ( .A(n9490), .ZN(P2_U3513) );
  MUX2_X1 U10351 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9491), .S(n10588), .Z(
        P2_U3512) );
  MUX2_X1 U10352 ( .A(n9492), .B(P2_REG0_REG_23__SCAN_IN), .S(n10585), .Z(
        P2_U3511) );
  MUX2_X1 U10353 ( .A(n9493), .B(P2_REG0_REG_22__SCAN_IN), .S(n10585), .Z(
        P2_U3510) );
  MUX2_X1 U10354 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9494), .S(n10588), .Z(
        P2_U3509) );
  MUX2_X1 U10355 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9495), .S(n10588), .Z(
        P2_U3508) );
  MUX2_X1 U10356 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9496), .S(n10588), .Z(
        P2_U3507) );
  MUX2_X1 U10357 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9497), .S(n10588), .Z(
        P2_U3505) );
  MUX2_X1 U10358 ( .A(n9498), .B(P2_REG0_REG_17__SCAN_IN), .S(n10585), .Z(
        P2_U3502) );
  MUX2_X1 U10359 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9499), .S(n10588), .Z(
        P2_U3499) );
  MUX2_X1 U10360 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9500), .S(n10588), .Z(
        P2_U3496) );
  INV_X1 U10361 ( .A(n9501), .ZN(n9505) );
  NAND3_X1 U10362 ( .A1(n9502), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9504) );
  OAI22_X1 U10363 ( .A1(n9505), .A2(n9504), .B1(n6819), .B2(n9503), .ZN(n9506)
         );
  AOI21_X1 U10364 ( .B1(n9997), .B2(n9507), .A(n9506), .ZN(n9508) );
  INV_X1 U10365 ( .A(n9508), .ZN(P2_U3327) );
  MUX2_X1 U10366 ( .A(n9509), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10367 ( .A1(n9510), .A2(n9511), .ZN(n9512) );
  AOI21_X1 U10368 ( .B1(n9513), .B2(n9512), .A(n9649), .ZN(n9514) );
  INV_X1 U10369 ( .A(n9514), .ZN(n9518) );
  INV_X1 U10370 ( .A(n9745), .ZN(n9652) );
  AOI22_X1 U10371 ( .A1(n9739), .A2(n9619), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9515) );
  OAI21_X1 U10372 ( .B1(n9744), .B2(n9607), .A(n9515), .ZN(n9516) );
  AOI21_X1 U10373 ( .B1(n9652), .B2(n9642), .A(n9516), .ZN(n9517) );
  OAI211_X1 U10374 ( .C1(n9741), .C2(n9613), .A(n9518), .B(n9517), .ZN(
        P1_U3212) );
  NAND2_X1 U10375 ( .A1(n9519), .A2(n9520), .ZN(n9521) );
  XOR2_X1 U10376 ( .A(n9522), .B(n9521), .Z(n9530) );
  OAI21_X1 U10377 ( .B1(n9607), .B2(n9524), .A(n9523), .ZN(n9525) );
  AOI21_X1 U10378 ( .B1(n9642), .B2(n9655), .A(n9525), .ZN(n9526) );
  OAI21_X1 U10379 ( .B1(n9646), .B2(n9527), .A(n9526), .ZN(n9528) );
  AOI21_X1 U10380 ( .B1(n9958), .B2(n4839), .A(n9528), .ZN(n9529) );
  OAI21_X1 U10381 ( .B1(n9530), .B2(n9649), .A(n9529), .ZN(P1_U3213) );
  NAND2_X1 U10382 ( .A1(n9532), .A2(n9531), .ZN(n9533) );
  XOR2_X1 U10383 ( .A(n9534), .B(n9533), .Z(n9541) );
  OAI22_X1 U10384 ( .A1(n9536), .A2(n9607), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9535), .ZN(n9537) );
  AOI21_X1 U10385 ( .B1(n9642), .B2(n9806), .A(n9537), .ZN(n9538) );
  OAI21_X1 U10386 ( .B1(n9646), .B2(n9799), .A(n9538), .ZN(n9539) );
  AOI21_X1 U10387 ( .B1(n9911), .B2(n4839), .A(n9539), .ZN(n9540) );
  OAI21_X1 U10388 ( .B1(n9541), .B2(n9649), .A(n9540), .ZN(P1_U3214) );
  OR2_X1 U10389 ( .A1(n8908), .A2(n9542), .ZN(n9545) );
  NAND2_X1 U10390 ( .A1(n9545), .A2(n9544), .ZN(n9547) );
  NAND2_X1 U10391 ( .A1(n5316), .A2(n9548), .ZN(n9546) );
  AOI22_X1 U10392 ( .A1(n5324), .A2(n9548), .B1(n9547), .B2(n9546), .ZN(n9553)
         );
  AOI22_X1 U10393 ( .A1(n9831), .A2(n9642), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9550) );
  NAND2_X1 U10394 ( .A1(n9867), .A2(n9641), .ZN(n9549) );
  OAI211_X1 U10395 ( .C1(n9646), .C2(n9836), .A(n9550), .B(n9549), .ZN(n9551)
         );
  AOI21_X1 U10396 ( .B1(n9922), .B2(n4839), .A(n9551), .ZN(n9552) );
  OAI21_X1 U10397 ( .B1(n9553), .B2(n9649), .A(n9552), .ZN(P1_U3221) );
  XNOR2_X1 U10398 ( .A(n9556), .B(n9555), .ZN(n9557) );
  XNOR2_X1 U10399 ( .A(n9554), .B(n9557), .ZN(n9562) );
  NAND2_X1 U10400 ( .A1(n9772), .A2(n9642), .ZN(n9559) );
  AOI22_X1 U10401 ( .A1(n9806), .A2(n9641), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9558) );
  OAI211_X1 U10402 ( .C1(n9646), .C2(n9767), .A(n9559), .B(n9558), .ZN(n9560)
         );
  AOI21_X1 U10403 ( .B1(n9901), .B2(n4839), .A(n9560), .ZN(n9561) );
  OAI21_X1 U10404 ( .B1(n9562), .B2(n9649), .A(n9561), .ZN(P1_U3223) );
  INV_X1 U10405 ( .A(n9563), .ZN(n9578) );
  AOI21_X1 U10406 ( .B1(n9565), .B2(n9637), .A(n9564), .ZN(n9566) );
  OAI21_X1 U10407 ( .B1(n9578), .B2(n9566), .A(n9604), .ZN(n9573) );
  AOI21_X1 U10408 ( .B1(n9642), .B2(n9653), .A(n9567), .ZN(n9568) );
  OAI21_X1 U10409 ( .B1(n9569), .B2(n9607), .A(n9568), .ZN(n9570) );
  AOI21_X1 U10410 ( .B1(n9571), .B2(n9619), .A(n9570), .ZN(n9572) );
  OAI211_X1 U10411 ( .C1(n9574), .C2(n9613), .A(n9573), .B(n9572), .ZN(
        P1_U3224) );
  INV_X1 U10412 ( .A(n9575), .ZN(n9577) );
  NOR3_X1 U10413 ( .A1(n9578), .A2(n9577), .A3(n9576), .ZN(n9581) );
  INV_X1 U10414 ( .A(n9579), .ZN(n9580) );
  OAI21_X1 U10415 ( .B1(n9581), .B2(n9580), .A(n9604), .ZN(n9587) );
  NAND2_X1 U10416 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9671) );
  OAI21_X1 U10417 ( .B1(n9607), .B2(n9582), .A(n9671), .ZN(n9585) );
  NOR2_X1 U10418 ( .A1(n9646), .A2(n9583), .ZN(n9584) );
  AOI211_X1 U10419 ( .C1(n9642), .C2(n9865), .A(n9585), .B(n9584), .ZN(n9586)
         );
  OAI211_X1 U10420 ( .C1(n9588), .C2(n9613), .A(n9587), .B(n9586), .ZN(
        P1_U3226) );
  XOR2_X1 U10421 ( .A(n9590), .B(n9589), .Z(n9597) );
  NOR2_X1 U10422 ( .A1(n9591), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9592) );
  AOI21_X1 U10423 ( .B1(n9819), .B2(n9641), .A(n9592), .ZN(n9594) );
  NAND2_X1 U10424 ( .A1(n9785), .A2(n9619), .ZN(n9593) );
  OAI211_X1 U10425 ( .C1(n9783), .C2(n9623), .A(n9594), .B(n9593), .ZN(n9595)
         );
  AOI21_X1 U10426 ( .B1(n9908), .B2(n4839), .A(n9595), .ZN(n9596) );
  OAI21_X1 U10427 ( .B1(n9597), .B2(n9649), .A(n9596), .ZN(P1_U3227) );
  OR2_X1 U10428 ( .A1(n8908), .A2(n9598), .ZN(n9600) );
  AND2_X1 U10429 ( .A1(n9600), .A2(n9599), .ZN(n9602) );
  OAI21_X1 U10430 ( .B1(n9603), .B2(n9602), .A(n9601), .ZN(n9605) );
  NAND2_X1 U10431 ( .A1(n9605), .A2(n9604), .ZN(n9612) );
  NOR2_X1 U10432 ( .A1(n9813), .A2(n9646), .ZN(n9610) );
  OAI22_X1 U10433 ( .A1(n9608), .A2(n9607), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9606), .ZN(n9609) );
  AOI211_X1 U10434 ( .C1(n9642), .C2(n9819), .A(n9610), .B(n9609), .ZN(n9611)
         );
  OAI211_X1 U10435 ( .C1(n9816), .C2(n9613), .A(n9612), .B(n9611), .ZN(
        P1_U3233) );
  NAND2_X1 U10436 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  XOR2_X1 U10437 ( .A(n9617), .B(n9616), .Z(n9629) );
  NAND2_X1 U10438 ( .A1(n9619), .A2(n9618), .ZN(n9622) );
  NOR2_X1 U10439 ( .A1(n9620), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9683) );
  AOI21_X1 U10440 ( .B1(n9641), .B2(n9653), .A(n9683), .ZN(n9621) );
  OAI211_X1 U10441 ( .C1(n9624), .C2(n9623), .A(n9622), .B(n9621), .ZN(n9625)
         );
  AOI21_X1 U10442 ( .B1(n9627), .B2(n4839), .A(n9625), .ZN(n9628) );
  OAI21_X1 U10443 ( .B1(n9629), .B2(n9649), .A(n9628), .ZN(P1_U3236) );
  XNOR2_X1 U10444 ( .A(n9631), .B(n9630), .ZN(n9636) );
  NAND2_X1 U10445 ( .A1(n5243), .A2(n9642), .ZN(n9633) );
  AOI22_X1 U10446 ( .A1(n9759), .A2(n9641), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9632) );
  OAI211_X1 U10447 ( .C1(n9646), .C2(n9753), .A(n9633), .B(n9632), .ZN(n9634)
         );
  AOI21_X1 U10448 ( .B1(n9896), .B2(n4839), .A(n9634), .ZN(n9635) );
  OAI21_X1 U10449 ( .B1(n9636), .B2(n9649), .A(n9635), .ZN(P1_U3238) );
  NAND2_X1 U10450 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  XOR2_X1 U10451 ( .A(n9640), .B(n9639), .Z(n9650) );
  AOI22_X1 U10452 ( .A1(n9641), .A2(n9656), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3084), .ZN(n9644) );
  NAND2_X1 U10453 ( .A1(n9642), .A2(n9654), .ZN(n9643) );
  OAI211_X1 U10454 ( .C1(n9646), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9647)
         );
  AOI21_X1 U10455 ( .B1(n9952), .B2(n4839), .A(n9647), .ZN(n9648) );
  OAI21_X1 U10456 ( .B1(n9650), .B2(n9649), .A(n9648), .ZN(P1_U3239) );
  MUX2_X1 U10457 ( .A(n9651), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9665), .Z(
        P1_U3584) );
  MUX2_X1 U10458 ( .A(n9652), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9665), .Z(
        P1_U3583) );
  MUX2_X1 U10459 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n5243), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9772), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10461 ( .A(n9759), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9665), .Z(
        P1_U3580) );
  MUX2_X1 U10462 ( .A(n9806), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9665), .Z(
        P1_U3579) );
  MUX2_X1 U10463 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9831), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9850), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9867), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10466 ( .A(n9849), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9665), .Z(
        P1_U3574) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9865), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10468 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9653), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9654), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10470 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9655), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9656), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9657), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10473 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9658), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9659), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9660), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10476 ( .A(n9661), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9665), .Z(
        P1_U3561) );
  MUX2_X1 U10477 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9662), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10478 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9663), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n7092), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10480 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9664), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n7129), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10482 ( .A(n7128), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9665), .Z(
        P1_U3555) );
  INV_X1 U10483 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9673) );
  AOI21_X1 U10484 ( .B1(n9675), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9666), .ZN(
        n9669) );
  NAND2_X1 U10485 ( .A1(n9687), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9667) );
  OAI21_X1 U10486 ( .B1(n9687), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9667), .ZN(
        n9668) );
  NOR2_X1 U10487 ( .A1(n9669), .A2(n9668), .ZN(n9686) );
  AOI211_X1 U10488 ( .C1(n9669), .C2(n9668), .A(n9686), .B(n10411), .ZN(n9670)
         );
  AOI21_X1 U10489 ( .B1(n10427), .B2(n9687), .A(n9670), .ZN(n9672) );
  OAI211_X1 U10490 ( .C1(n10420), .C2(n9673), .A(n9672), .B(n9671), .ZN(n9679)
         );
  AOI21_X1 U10491 ( .B1(n9675), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9674), .ZN(
        n9677) );
  XNOR2_X1 U10492 ( .A(n9687), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9676) );
  NOR2_X1 U10493 ( .A1(n9677), .A2(n9676), .ZN(n9680) );
  AOI211_X1 U10494 ( .C1(n9677), .C2(n9676), .A(n9680), .B(n10433), .ZN(n9678)
         );
  OR2_X1 U10495 ( .A1(n9679), .A2(n9678), .ZN(P1_U3258) );
  XOR2_X1 U10496 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9699), .Z(n9682) );
  AOI21_X1 U10497 ( .B1(n9687), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9680), .ZN(
        n9681) );
  NAND2_X1 U10498 ( .A1(n9681), .A2(n9682), .ZN(n9698) );
  OAI21_X1 U10499 ( .B1(n9682), .B2(n9681), .A(n9698), .ZN(n9693) );
  INV_X1 U10500 ( .A(n9699), .ZN(n9685) );
  AOI21_X1 U10501 ( .B1(n10436), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9683), .ZN(
        n9684) );
  OAI21_X1 U10502 ( .B1(n9685), .B2(n10318), .A(n9684), .ZN(n9692) );
  AOI21_X1 U10503 ( .B1(n9687), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9686), .ZN(
        n9690) );
  NAND2_X1 U10504 ( .A1(n9699), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9688) );
  OAI21_X1 U10505 ( .B1(n9699), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9688), .ZN(
        n9689) );
  NOR2_X1 U10506 ( .A1(n9690), .A2(n9689), .ZN(n9695) );
  AOI211_X1 U10507 ( .C1(n9690), .C2(n9689), .A(n9695), .B(n10411), .ZN(n9691)
         );
  AOI211_X1 U10508 ( .C1(n10407), .C2(n9693), .A(n9692), .B(n9691), .ZN(n9694)
         );
  INV_X1 U10509 ( .A(n9694), .ZN(P1_U3259) );
  AOI21_X1 U10510 ( .B1(n9699), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9695), .ZN(
        n9697) );
  MUX2_X1 U10511 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n6197), .S(n9834), .Z(n9696) );
  XNOR2_X1 U10512 ( .A(n9697), .B(n9696), .ZN(n9707) );
  OAI21_X1 U10513 ( .B1(n9699), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9698), .ZN(
        n9701) );
  XNOR2_X1 U10514 ( .A(n9834), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9700) );
  XNOR2_X1 U10515 ( .A(n9701), .B(n9700), .ZN(n9705) );
  NAND2_X1 U10516 ( .A1(n10436), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9702) );
  OAI211_X1 U10517 ( .C1(n10318), .C2(n9834), .A(n9703), .B(n9702), .ZN(n9704)
         );
  AOI21_X1 U10518 ( .B1(n10407), .B2(n9705), .A(n9704), .ZN(n9706) );
  OAI21_X1 U10519 ( .B1(n10411), .B2(n9707), .A(n9706), .ZN(P1_U3260) );
  OAI21_X1 U10520 ( .B1(n9710), .B2(n9709), .A(n9708), .ZN(n9880) );
  OAI21_X1 U10521 ( .B1(n10447), .B2(n9712), .A(n9711), .ZN(n9713) );
  AOI21_X1 U10522 ( .B1(n9878), .B2(n9827), .A(n9713), .ZN(n9714) );
  OAI21_X1 U10523 ( .B1(n9880), .B2(n10443), .A(n9714), .ZN(P1_U3262) );
  NAND2_X1 U10524 ( .A1(n9716), .A2(n4906), .ZN(n9717) );
  XNOR2_X1 U10525 ( .A(n9717), .B(n9720), .ZN(n9881) );
  NAND2_X1 U10526 ( .A1(n9719), .A2(n9718), .ZN(n9721) );
  XNOR2_X1 U10527 ( .A(n9721), .B(n9720), .ZN(n9725) );
  OAI22_X1 U10528 ( .A1(n9745), .A2(n9782), .B1(n9723), .B2(n9722), .ZN(n9724)
         );
  OAI22_X1 U10529 ( .A1(n9727), .A2(n10450), .B1(n9726), .B2(n10447), .ZN(
        n9728) );
  AOI21_X1 U10530 ( .B1(n8704), .B2(n9827), .A(n9728), .ZN(n9732) );
  INV_X1 U10531 ( .A(n8704), .ZN(n9730) );
  NAND2_X1 U10532 ( .A1(n9882), .A2(n10006), .ZN(n9731) );
  OAI211_X1 U10533 ( .C1(n9883), .C2(n9843), .A(n9732), .B(n9731), .ZN(n9733)
         );
  AOI21_X1 U10534 ( .B1(n9881), .B2(n9734), .A(n9733), .ZN(n9735) );
  INV_X1 U10535 ( .A(n9735), .ZN(P1_U3355) );
  XOR2_X1 U10536 ( .A(n9742), .B(n9736), .Z(n9895) );
  INV_X1 U10537 ( .A(n9752), .ZN(n9738) );
  AOI21_X1 U10538 ( .B1(n9891), .B2(n9738), .A(n9737), .ZN(n9892) );
  AOI22_X1 U10539 ( .A1(n9739), .A2(n10008), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n9843), .ZN(n9740) );
  OAI21_X1 U10540 ( .B1(n9741), .B2(n10442), .A(n9740), .ZN(n9749) );
  AOI21_X1 U10541 ( .B1(n9743), .B2(n9742), .A(n9780), .ZN(n9747) );
  OAI22_X1 U10542 ( .A1(n9745), .A2(n9784), .B1(n9744), .B2(n9782), .ZN(n9746)
         );
  AOI21_X1 U10543 ( .B1(n9747), .B2(n5137), .A(n9746), .ZN(n9894) );
  NOR2_X1 U10544 ( .A1(n9894), .A2(n9843), .ZN(n9748) );
  AOI211_X1 U10545 ( .C1(n9892), .C2(n10006), .A(n9749), .B(n9748), .ZN(n9750)
         );
  OAI21_X1 U10546 ( .B1(n9895), .B2(n9873), .A(n9750), .ZN(P1_U3264) );
  XNOR2_X1 U10547 ( .A(n9751), .B(n9757), .ZN(n9900) );
  AOI21_X1 U10548 ( .B1(n9896), .B2(n9766), .A(n9752), .ZN(n9897) );
  INV_X1 U10549 ( .A(n9753), .ZN(n9754) );
  AOI22_X1 U10550 ( .A1(n9754), .A2(n10008), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n9843), .ZN(n9755) );
  OAI21_X1 U10551 ( .B1(n9756), .B2(n10442), .A(n9755), .ZN(n9762) );
  XNOR2_X1 U10552 ( .A(n9758), .B(n9757), .ZN(n9760) );
  AOI222_X1 U10553 ( .A1(n9869), .A2(n9760), .B1(n5243), .B2(n9866), .C1(n9759), .C2(n9864), .ZN(n9899) );
  NOR2_X1 U10554 ( .A1(n9899), .A2(n9843), .ZN(n9761) );
  AOI211_X1 U10555 ( .C1(n9897), .C2(n10006), .A(n9762), .B(n9761), .ZN(n9763)
         );
  OAI21_X1 U10556 ( .B1(n9900), .B2(n9873), .A(n9763), .ZN(P1_U3265) );
  XOR2_X1 U10557 ( .A(n9770), .B(n9764), .Z(n9905) );
  AOI21_X1 U10558 ( .B1(n9901), .B2(n9777), .A(n5063), .ZN(n9902) );
  INV_X1 U10559 ( .A(n9767), .ZN(n9768) );
  AOI22_X1 U10560 ( .A1(n9768), .A2(n10008), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n9843), .ZN(n9769) );
  OAI21_X1 U10561 ( .B1(n8703), .B2(n10442), .A(n9769), .ZN(n9775) );
  XNOR2_X1 U10562 ( .A(n9771), .B(n9770), .ZN(n9773) );
  AOI222_X1 U10563 ( .A1(n9869), .A2(n9773), .B1(n9772), .B2(n9866), .C1(n9806), .C2(n9864), .ZN(n9904) );
  NOR2_X1 U10564 ( .A1(n9904), .A2(n9843), .ZN(n9774) );
  AOI211_X1 U10565 ( .C1(n9902), .C2(n10006), .A(n9775), .B(n9774), .ZN(n9776)
         );
  OAI21_X1 U10566 ( .B1(n9905), .B2(n9873), .A(n9776), .ZN(P1_U3266) );
  AOI211_X1 U10567 ( .C1(n9908), .C2(n9796), .A(n7137), .B(n9765), .ZN(n9907)
         );
  XOR2_X1 U10568 ( .A(n9788), .B(n9778), .Z(n9779) );
  OAI222_X1 U10569 ( .A1(n9784), .A2(n9783), .B1(n9782), .B2(n9781), .C1(n9780), .C2(n9779), .ZN(n9906) );
  AOI21_X1 U10570 ( .B1(n9907), .B2(n9834), .A(n9906), .ZN(n9793) );
  INV_X1 U10571 ( .A(n9785), .ZN(n9787) );
  OAI22_X1 U10572 ( .A1(n9787), .A2(n10450), .B1(n9786), .B2(n10447), .ZN(
        n9791) );
  XOR2_X1 U10573 ( .A(n9789), .B(n9788), .Z(n9910) );
  NOR2_X1 U10574 ( .A1(n9910), .A2(n9873), .ZN(n9790) );
  AOI211_X1 U10575 ( .C1(n9827), .C2(n9908), .A(n9791), .B(n9790), .ZN(n9792)
         );
  OAI21_X1 U10576 ( .B1(n9843), .B2(n9793), .A(n9792), .ZN(P1_U3267) );
  XNOR2_X1 U10577 ( .A(n9794), .B(n9795), .ZN(n9915) );
  INV_X1 U10578 ( .A(n9812), .ZN(n9798) );
  INV_X1 U10579 ( .A(n9796), .ZN(n9797) );
  AOI21_X1 U10580 ( .B1(n9911), .B2(n9798), .A(n9797), .ZN(n9912) );
  INV_X1 U10581 ( .A(n9799), .ZN(n9800) );
  AOI22_X1 U10582 ( .A1(n9800), .A2(n10008), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n9843), .ZN(n9801) );
  OAI21_X1 U10583 ( .B1(n9802), .B2(n10442), .A(n9801), .ZN(n9809) );
  OAI21_X1 U10584 ( .B1(n9805), .B2(n9804), .A(n9803), .ZN(n9807) );
  AOI222_X1 U10585 ( .A1(n9869), .A2(n9807), .B1(n9806), .B2(n9866), .C1(n9831), .C2(n9864), .ZN(n9914) );
  NOR2_X1 U10586 ( .A1(n9914), .A2(n9843), .ZN(n9808) );
  AOI211_X1 U10587 ( .C1(n9912), .C2(n10006), .A(n9809), .B(n9808), .ZN(n9810)
         );
  OAI21_X1 U10588 ( .B1(n9915), .B2(n9873), .A(n9810), .ZN(P1_U3268) );
  XNOR2_X1 U10589 ( .A(n9811), .B(n9817), .ZN(n9920) );
  AOI21_X1 U10590 ( .B1(n9916), .B2(n9833), .A(n9812), .ZN(n9917) );
  INV_X1 U10591 ( .A(n9813), .ZN(n9814) );
  AOI22_X1 U10592 ( .A1(n9814), .A2(n10008), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n9843), .ZN(n9815) );
  OAI21_X1 U10593 ( .B1(n9816), .B2(n10442), .A(n9815), .ZN(n9822) );
  XNOR2_X1 U10594 ( .A(n9818), .B(n9817), .ZN(n9820) );
  AOI222_X1 U10595 ( .A1(n9869), .A2(n9820), .B1(n9819), .B2(n9866), .C1(n9850), .C2(n9864), .ZN(n9919) );
  NOR2_X1 U10596 ( .A1(n9919), .A2(n9843), .ZN(n9821) );
  AOI211_X1 U10597 ( .C1(n9917), .C2(n10006), .A(n9822), .B(n9821), .ZN(n9823)
         );
  OAI21_X1 U10598 ( .B1(n9920), .B2(n9873), .A(n9823), .ZN(P1_U3269) );
  AOI21_X1 U10599 ( .B1(n9830), .B2(n9825), .A(n9824), .ZN(n9826) );
  INV_X1 U10600 ( .A(n9826), .ZN(n9925) );
  AOI22_X1 U10601 ( .A1(n9922), .A2(n9827), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9843), .ZN(n9839) );
  OAI21_X1 U10602 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(n9832) );
  AOI222_X1 U10603 ( .A1(n9869), .A2(n9832), .B1(n9831), .B2(n9866), .C1(n9867), .C2(n9864), .ZN(n9924) );
  AOI211_X1 U10604 ( .C1(n9922), .C2(n9841), .A(n7137), .B(n5061), .ZN(n9921)
         );
  NAND2_X1 U10605 ( .A1(n9921), .A2(n9834), .ZN(n9835) );
  OAI211_X1 U10606 ( .C1(n10450), .C2(n9836), .A(n9924), .B(n9835), .ZN(n9837)
         );
  NAND2_X1 U10607 ( .A1(n9837), .A2(n10447), .ZN(n9838) );
  OAI211_X1 U10608 ( .C1(n9925), .C2(n9873), .A(n9839), .B(n9838), .ZN(
        P1_U3270) );
  XNOR2_X1 U10609 ( .A(n9840), .B(n5119), .ZN(n9930) );
  INV_X1 U10610 ( .A(n9857), .ZN(n9842) );
  AOI21_X1 U10611 ( .B1(n9926), .B2(n9842), .A(n5057), .ZN(n9927) );
  AOI22_X1 U10612 ( .A1(n9844), .A2(n10008), .B1(n9843), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9845) );
  OAI21_X1 U10613 ( .B1(n9846), .B2(n10442), .A(n9845), .ZN(n9853) );
  XNOR2_X1 U10614 ( .A(n9847), .B(n9848), .ZN(n9851) );
  AOI222_X1 U10615 ( .A1(n9869), .A2(n9851), .B1(n9850), .B2(n9866), .C1(n9849), .C2(n9864), .ZN(n9929) );
  NOR2_X1 U10616 ( .A1(n9929), .A2(n9843), .ZN(n9852) );
  AOI211_X1 U10617 ( .C1(n9927), .C2(n10006), .A(n9853), .B(n9852), .ZN(n9854)
         );
  OAI21_X1 U10618 ( .B1(n9873), .B2(n9930), .A(n9854), .ZN(P1_U3271) );
  XNOR2_X1 U10619 ( .A(n9855), .B(n4857), .ZN(n9935) );
  INV_X1 U10620 ( .A(n9856), .ZN(n9858) );
  AOI21_X1 U10621 ( .B1(n9931), .B2(n9858), .A(n9857), .ZN(n9932) );
  INV_X1 U10622 ( .A(n9859), .ZN(n9860) );
  AOI22_X1 U10623 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(n9843), .B1(n9860), .B2(
        n10008), .ZN(n9861) );
  OAI21_X1 U10624 ( .B1(n9862), .B2(n10442), .A(n9861), .ZN(n9871) );
  OAI21_X1 U10625 ( .B1(n4918), .B2(n4857), .A(n9863), .ZN(n9868) );
  AOI222_X1 U10626 ( .A1(n9869), .A2(n9868), .B1(n9867), .B2(n9866), .C1(n9865), .C2(n9864), .ZN(n9934) );
  NOR2_X1 U10627 ( .A1(n9934), .A2(n9843), .ZN(n9870) );
  AOI211_X1 U10628 ( .C1(n9932), .C2(n10006), .A(n9871), .B(n9870), .ZN(n9872)
         );
  OAI21_X1 U10629 ( .B1(n9873), .B2(n9935), .A(n9872), .ZN(P1_U3272) );
  AOI21_X1 U10630 ( .B1(n9874), .B2(n9964), .A(n9877), .ZN(n9875) );
  OAI21_X1 U10631 ( .B1(n9876), .B2(n7137), .A(n9875), .ZN(n9970) );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9970), .S(n4842), .Z(
        P1_U3554) );
  AOI21_X1 U10633 ( .B1(n9878), .B2(n9964), .A(n9877), .ZN(n9879) );
  OAI21_X1 U10634 ( .B1(n9880), .B2(n7137), .A(n9879), .ZN(n9971) );
  MUX2_X1 U10635 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9971), .S(n4842), .Z(
        P1_U3553) );
  NAND2_X1 U10636 ( .A1(n9881), .A2(n10541), .ZN(n9884) );
  MUX2_X1 U10637 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9972), .S(n4842), .Z(
        P1_U3552) );
  AOI22_X1 U10638 ( .A1(n9886), .A2(n9965), .B1(n9964), .B2(n9885), .ZN(n9887)
         );
  MUX2_X1 U10639 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9973), .S(n4842), .Z(
        P1_U3551) );
  AOI22_X1 U10640 ( .A1(n9892), .A2(n9965), .B1(n9964), .B2(n9891), .ZN(n9893)
         );
  OAI211_X1 U10641 ( .C1(n9895), .C2(n10494), .A(n9894), .B(n9893), .ZN(n9974)
         );
  MUX2_X1 U10642 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9974), .S(n4842), .Z(
        P1_U3550) );
  AOI22_X1 U10643 ( .A1(n9897), .A2(n9965), .B1(n9964), .B2(n9896), .ZN(n9898)
         );
  OAI211_X1 U10644 ( .C1(n9900), .C2(n10494), .A(n9899), .B(n9898), .ZN(n9975)
         );
  MUX2_X1 U10645 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9975), .S(n4842), .Z(
        P1_U3549) );
  AOI22_X1 U10646 ( .A1(n9902), .A2(n9965), .B1(n9964), .B2(n9901), .ZN(n9903)
         );
  OAI211_X1 U10647 ( .C1(n9905), .C2(n10494), .A(n9904), .B(n9903), .ZN(n9976)
         );
  MUX2_X1 U10648 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9976), .S(n4842), .Z(
        P1_U3548) );
  AOI211_X1 U10649 ( .C1(n9959), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9909)
         );
  OAI21_X1 U10650 ( .B1(n9910), .B2(n10494), .A(n9909), .ZN(n9977) );
  MUX2_X1 U10651 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9977), .S(n4842), .Z(
        P1_U3547) );
  AOI22_X1 U10652 ( .A1(n9912), .A2(n9965), .B1(n9964), .B2(n9911), .ZN(n9913)
         );
  OAI211_X1 U10653 ( .C1(n9915), .C2(n10494), .A(n9914), .B(n9913), .ZN(n9978)
         );
  MUX2_X1 U10654 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9978), .S(n4842), .Z(
        P1_U3546) );
  AOI22_X1 U10655 ( .A1(n9917), .A2(n9965), .B1(n9964), .B2(n9916), .ZN(n9918)
         );
  OAI211_X1 U10656 ( .C1(n9920), .C2(n10494), .A(n9919), .B(n9918), .ZN(n9979)
         );
  MUX2_X1 U10657 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9979), .S(n4842), .Z(
        P1_U3545) );
  AOI21_X1 U10658 ( .B1(n9959), .B2(n9922), .A(n9921), .ZN(n9923) );
  OAI211_X1 U10659 ( .C1(n9925), .C2(n10494), .A(n9924), .B(n9923), .ZN(n9980)
         );
  MUX2_X1 U10660 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9980), .S(n4842), .Z(
        P1_U3544) );
  AOI22_X1 U10661 ( .A1(n9927), .A2(n9965), .B1(n9964), .B2(n9926), .ZN(n9928)
         );
  OAI211_X1 U10662 ( .C1(n9930), .C2(n10494), .A(n9929), .B(n9928), .ZN(n9981)
         );
  MUX2_X1 U10663 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9981), .S(n4842), .Z(
        P1_U3543) );
  AOI22_X1 U10664 ( .A1(n9932), .A2(n9965), .B1(n9964), .B2(n9931), .ZN(n9933)
         );
  OAI211_X1 U10665 ( .C1(n9935), .C2(n10494), .A(n9934), .B(n9933), .ZN(n9982)
         );
  MUX2_X1 U10666 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9982), .S(n4842), .Z(
        P1_U3542) );
  OAI22_X1 U10667 ( .A1(n9937), .A2(n7137), .B1(n9936), .B2(n10537), .ZN(n9939) );
  AOI211_X1 U10668 ( .C1(n10463), .C2(n9940), .A(n9939), .B(n9938), .ZN(n9941)
         );
  INV_X1 U10669 ( .A(n9941), .ZN(n9983) );
  MUX2_X1 U10670 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9983), .S(n4842), .Z(
        P1_U3541) );
  AOI22_X1 U10671 ( .A1(n9943), .A2(n9965), .B1(n9964), .B2(n9942), .ZN(n9944)
         );
  OAI211_X1 U10672 ( .C1(n9946), .C2(n10494), .A(n9945), .B(n9944), .ZN(n9984)
         );
  MUX2_X1 U10673 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9984), .S(n4842), .Z(
        P1_U3540) );
  AOI211_X1 U10674 ( .C1(n9964), .C2(n9949), .A(n9948), .B(n9947), .ZN(n9950)
         );
  OAI21_X1 U10675 ( .B1(n10494), .B2(n9951), .A(n9950), .ZN(n9985) );
  MUX2_X1 U10676 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9985), .S(n4842), .Z(
        P1_U3539) );
  AOI22_X1 U10677 ( .A1(n9953), .A2(n9965), .B1(n9964), .B2(n9952), .ZN(n9954)
         );
  OAI211_X1 U10678 ( .C1(n9956), .C2(n10494), .A(n9955), .B(n9954), .ZN(n9986)
         );
  MUX2_X1 U10679 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9986), .S(n4842), .Z(
        P1_U3538) );
  AOI21_X1 U10680 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(n9960) );
  OAI211_X1 U10681 ( .C1(n9962), .C2(n10494), .A(n9961), .B(n9960), .ZN(n9987)
         );
  MUX2_X1 U10682 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9987), .S(n4842), .Z(
        P1_U3537) );
  AOI22_X1 U10683 ( .A1(n9966), .A2(n9965), .B1(n9964), .B2(n9963), .ZN(n9967)
         );
  OAI211_X1 U10684 ( .C1(n9969), .C2(n10494), .A(n9968), .B(n9967), .ZN(n9988)
         );
  MUX2_X1 U10685 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9988), .S(n4842), .Z(
        P1_U3536) );
  MUX2_X1 U10686 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9970), .S(n4843), .Z(
        P1_U3522) );
  MUX2_X1 U10687 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9971), .S(n4843), .Z(
        P1_U3521) );
  MUX2_X1 U10688 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9972), .S(n4843), .Z(
        P1_U3520) );
  MUX2_X1 U10689 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9973), .S(n4843), .Z(
        P1_U3519) );
  MUX2_X1 U10690 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9974), .S(n4843), .Z(
        P1_U3518) );
  MUX2_X1 U10691 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9975), .S(n4843), .Z(
        P1_U3517) );
  MUX2_X1 U10692 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9976), .S(n4843), .Z(
        P1_U3516) );
  MUX2_X1 U10693 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9977), .S(n4843), .Z(
        P1_U3515) );
  MUX2_X1 U10694 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9978), .S(n4843), .Z(
        P1_U3514) );
  MUX2_X1 U10695 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9979), .S(n4843), .Z(
        P1_U3513) );
  MUX2_X1 U10696 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9980), .S(n4843), .Z(
        P1_U3512) );
  MUX2_X1 U10697 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9981), .S(n4843), .Z(
        P1_U3511) );
  MUX2_X1 U10698 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9982), .S(n4843), .Z(
        P1_U3510) );
  MUX2_X1 U10699 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9983), .S(n4843), .Z(
        P1_U3508) );
  MUX2_X1 U10700 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9984), .S(n4843), .Z(
        P1_U3505) );
  MUX2_X1 U10701 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9985), .S(n4843), .Z(
        P1_U3502) );
  MUX2_X1 U10702 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9986), .S(n4843), .Z(
        P1_U3499) );
  MUX2_X1 U10703 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9987), .S(n4843), .Z(
        P1_U3496) );
  MUX2_X1 U10704 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9988), .S(n4843), .Z(
        P1_U3493) );
  MUX2_X1 U10705 ( .A(P1_D_REG_0__SCAN_IN), .B(n9990), .S(n9989), .Z(P1_U3440)
         );
  INV_X1 U10706 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9992) );
  NAND3_X1 U10707 ( .A1(n9992), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9994) );
  OAI22_X1 U10708 ( .A1(n9991), .A2(n9994), .B1(n9993), .B2(n8841), .ZN(n9995)
         );
  AOI21_X1 U10709 ( .B1(n9997), .B2(n9996), .A(n9995), .ZN(n9998) );
  INV_X1 U10710 ( .A(n9998), .ZN(P1_U3322) );
  MUX2_X1 U10711 ( .A(n9999), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AND2_X1 U10712 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10000), .ZN(P1_U3321) );
  AND2_X1 U10713 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10000), .ZN(P1_U3320) );
  AND2_X1 U10714 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10000), .ZN(P1_U3319) );
  AND2_X1 U10715 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10000), .ZN(P1_U3318) );
  AND2_X1 U10716 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10000), .ZN(P1_U3317) );
  AND2_X1 U10717 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10000), .ZN(P1_U3316) );
  AND2_X1 U10718 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10000), .ZN(P1_U3315) );
  AND2_X1 U10719 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10000), .ZN(P1_U3314) );
  AND2_X1 U10720 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10000), .ZN(P1_U3313) );
  AND2_X1 U10721 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10000), .ZN(P1_U3312) );
  AND2_X1 U10722 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10000), .ZN(P1_U3311) );
  AND2_X1 U10723 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10000), .ZN(P1_U3310) );
  AND2_X1 U10724 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10000), .ZN(P1_U3309) );
  AND2_X1 U10725 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10000), .ZN(P1_U3308) );
  AND2_X1 U10726 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10000), .ZN(P1_U3307) );
  AND2_X1 U10727 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10000), .ZN(P1_U3306) );
  AND2_X1 U10728 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10000), .ZN(P1_U3305) );
  AND2_X1 U10729 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10000), .ZN(P1_U3304) );
  AND2_X1 U10730 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10000), .ZN(P1_U3303) );
  AND2_X1 U10731 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10000), .ZN(P1_U3302) );
  AND2_X1 U10732 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10000), .ZN(P1_U3301) );
  AND2_X1 U10733 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10000), .ZN(P1_U3300) );
  AND2_X1 U10734 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10000), .ZN(P1_U3299) );
  AND2_X1 U10735 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10000), .ZN(P1_U3298) );
  AND2_X1 U10736 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10000), .ZN(P1_U3297) );
  AND2_X1 U10737 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10000), .ZN(P1_U3296) );
  AND2_X1 U10738 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10000), .ZN(P1_U3295) );
  AND2_X1 U10739 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10000), .ZN(P1_U3294) );
  AND2_X1 U10740 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10000), .ZN(P1_U3293) );
  AND2_X1 U10741 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10000), .ZN(P1_U3292) );
  INV_X1 U10742 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10005) );
  NAND2_X1 U10743 ( .A1(n10002), .A2(n10001), .ZN(n10352) );
  INV_X1 U10744 ( .A(n10003), .ZN(n10004) );
  AOI22_X1 U10745 ( .A1(n10005), .A2(n10352), .B1(n10355), .B2(n10004), .ZN(
        P2_U3438) );
  AND2_X1 U10746 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10352), .ZN(P2_U3326) );
  AND2_X1 U10747 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10352), .ZN(P2_U3325) );
  AND2_X1 U10748 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10352), .ZN(P2_U3324) );
  AND2_X1 U10749 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10352), .ZN(P2_U3323) );
  AND2_X1 U10750 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10352), .ZN(P2_U3322) );
  AND2_X1 U10751 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10352), .ZN(P2_U3321) );
  AND2_X1 U10752 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10352), .ZN(P2_U3320) );
  AND2_X1 U10753 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10352), .ZN(P2_U3319) );
  AND2_X1 U10754 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10352), .ZN(P2_U3318) );
  AND2_X1 U10755 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10352), .ZN(P2_U3317) );
  AND2_X1 U10756 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10352), .ZN(P2_U3316) );
  AND2_X1 U10757 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10352), .ZN(P2_U3315) );
  AND2_X1 U10758 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10352), .ZN(P2_U3314) );
  AND2_X1 U10759 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10352), .ZN(P2_U3313) );
  AND2_X1 U10760 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10352), .ZN(P2_U3312) );
  AND2_X1 U10761 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10352), .ZN(P2_U3311) );
  AND2_X1 U10762 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10352), .ZN(P2_U3310) );
  AND2_X1 U10763 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10352), .ZN(P2_U3309) );
  AND2_X1 U10764 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10352), .ZN(P2_U3308) );
  AND2_X1 U10765 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10352), .ZN(P2_U3307) );
  AND2_X1 U10766 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10352), .ZN(P2_U3306) );
  AND2_X1 U10767 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10352), .ZN(P2_U3305) );
  AND2_X1 U10768 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10352), .ZN(P2_U3304) );
  AND2_X1 U10769 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10352), .ZN(P2_U3303) );
  AND2_X1 U10770 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10352), .ZN(P2_U3302) );
  AND2_X1 U10771 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10352), .ZN(P2_U3301) );
  AND2_X1 U10772 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10352), .ZN(P2_U3300) );
  AND2_X1 U10773 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10352), .ZN(P2_U3299) );
  AND2_X1 U10774 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10352), .ZN(P2_U3298) );
  AND2_X1 U10775 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10352), .ZN(P2_U3297) );
  NAND2_X1 U10776 ( .A1(n10007), .A2(n10006), .ZN(n10011) );
  AOI22_X1 U10777 ( .A1(n9843), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n10009), 
        .B2(n10008), .ZN(n10010) );
  OAI211_X1 U10778 ( .C1(n10012), .C2(n10442), .A(n10011), .B(n10010), .ZN(
        n10013) );
  AOI21_X1 U10779 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(n10016) );
  OAI21_X1 U10780 ( .B1(n10017), .B2(n9843), .A(n10016), .ZN(n10221) );
  OAI22_X1 U10781 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_52), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .ZN(n10018) );
  AOI221_X1 U10782 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .C1(
        keyinput_53), .C2(P2_REG3_REG_9__SCAN_IN), .A(n10018), .ZN(n10098) );
  AOI22_X1 U10783 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_45), .B1(n10117), .B2(keyinput_46), .ZN(n10019) );
  OAI221_X1 U10784 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(
        n10117), .C2(keyinput_46), .A(n10019), .ZN(n10089) );
  INV_X1 U10785 ( .A(keyinput_44), .ZN(n10087) );
  XNOR2_X1 U10786 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n10085)
         );
  INV_X1 U10787 ( .A(keyinput_38), .ZN(n10079) );
  INV_X1 U10788 ( .A(SI_3_), .ZN(n10173) );
  OAI22_X1 U10789 ( .A1(n10169), .A2(keyinput_31), .B1(SI_2_), .B2(keyinput_30), .ZN(n10020) );
  AOI221_X1 U10790 ( .B1(n10169), .B2(keyinput_31), .C1(keyinput_30), .C2(
        SI_2_), .A(n10020), .ZN(n10068) );
  INV_X1 U10791 ( .A(keyinput_28), .ZN(n10066) );
  INV_X1 U10792 ( .A(keyinput_27), .ZN(n10064) );
  INV_X1 U10793 ( .A(keyinput_26), .ZN(n10062) );
  INV_X1 U10794 ( .A(SI_15_), .ZN(n10022) );
  OAI22_X1 U10795 ( .A1(n10022), .A2(keyinput_17), .B1(SI_17_), .B2(
        keyinput_15), .ZN(n10021) );
  AOI221_X1 U10796 ( .B1(n10022), .B2(keyinput_17), .C1(keyinput_15), .C2(
        SI_17_), .A(n10021), .ZN(n10026) );
  OAI22_X1 U10797 ( .A1(n10147), .A2(keyinput_16), .B1(n10024), .B2(
        keyinput_18), .ZN(n10023) );
  AOI221_X1 U10798 ( .B1(n10147), .B2(keyinput_16), .C1(keyinput_18), .C2(
        n10024), .A(n10023), .ZN(n10025) );
  OAI211_X1 U10799 ( .C1(SI_13_), .C2(keyinput_19), .A(n10026), .B(n10025), 
        .ZN(n10027) );
  AOI21_X1 U10800 ( .B1(SI_13_), .B2(keyinput_19), .A(n10027), .ZN(n10055) );
  INV_X1 U10801 ( .A(SI_18_), .ZN(n10143) );
  INV_X1 U10802 ( .A(keyinput_14), .ZN(n10049) );
  INV_X1 U10803 ( .A(keyinput_10), .ZN(n10042) );
  OAI22_X1 U10804 ( .A1(n10029), .A2(keyinput_8), .B1(SI_23_), .B2(keyinput_9), 
        .ZN(n10028) );
  AOI221_X1 U10805 ( .B1(n10029), .B2(keyinput_8), .C1(keyinput_9), .C2(SI_23_), .A(n10028), .ZN(n10039) );
  XNOR2_X1 U10806 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n10037) );
  AOI22_X1 U10807 ( .A1(SI_31_), .A2(keyinput_1), .B1(SI_30_), .B2(keyinput_2), 
        .ZN(n10030) );
  OAI221_X1 U10808 ( .B1(SI_31_), .B2(keyinput_1), .C1(SI_30_), .C2(keyinput_2), .A(n10030), .ZN(n10036) );
  OAI22_X1 U10809 ( .A1(n10032), .A2(keyinput_5), .B1(keyinput_6), .B2(SI_26_), 
        .ZN(n10031) );
  AOI221_X1 U10810 ( .B1(n10032), .B2(keyinput_5), .C1(SI_26_), .C2(keyinput_6), .A(n10031), .ZN(n10035) );
  OAI22_X1 U10811 ( .A1(SI_28_), .A2(keyinput_4), .B1(keyinput_3), .B2(SI_29_), 
        .ZN(n10033) );
  AOI221_X1 U10812 ( .B1(SI_28_), .B2(keyinput_4), .C1(SI_29_), .C2(keyinput_3), .A(n10033), .ZN(n10034) );
  OAI211_X1 U10813 ( .C1(n10037), .C2(n10036), .A(n10035), .B(n10034), .ZN(
        n10038) );
  OAI211_X1 U10814 ( .C1(SI_25_), .C2(keyinput_7), .A(n10039), .B(n10038), 
        .ZN(n10040) );
  AOI21_X1 U10815 ( .B1(SI_25_), .B2(keyinput_7), .A(n10040), .ZN(n10041) );
  AOI221_X1 U10816 ( .B1(SI_22_), .B2(n10042), .C1(n10137), .C2(keyinput_10), 
        .A(n10041), .ZN(n10046) );
  AOI22_X1 U10817 ( .A1(SI_20_), .A2(keyinput_12), .B1(n10044), .B2(
        keyinput_11), .ZN(n10043) );
  OAI221_X1 U10818 ( .B1(SI_20_), .B2(keyinput_12), .C1(n10044), .C2(
        keyinput_11), .A(n10043), .ZN(n10045) );
  AOI211_X1 U10819 ( .C1(SI_19_), .C2(keyinput_13), .A(n10046), .B(n10045), 
        .ZN(n10047) );
  OAI21_X1 U10820 ( .B1(SI_19_), .B2(keyinput_13), .A(n10047), .ZN(n10048) );
  OAI221_X1 U10821 ( .B1(SI_18_), .B2(keyinput_14), .C1(n10143), .C2(n10049), 
        .A(n10048), .ZN(n10054) );
  XOR2_X1 U10822 ( .A(SI_12_), .B(keyinput_20), .Z(n10053) );
  AOI22_X1 U10823 ( .A1(SI_10_), .A2(keyinput_22), .B1(n10051), .B2(
        keyinput_21), .ZN(n10050) );
  OAI221_X1 U10824 ( .B1(SI_10_), .B2(keyinput_22), .C1(n10051), .C2(
        keyinput_21), .A(n10050), .ZN(n10052) );
  AOI211_X1 U10825 ( .C1(n10055), .C2(n10054), .A(n10053), .B(n10052), .ZN(
        n10059) );
  AOI22_X1 U10826 ( .A1(SI_7_), .A2(keyinput_25), .B1(n10057), .B2(keyinput_24), .ZN(n10056) );
  OAI221_X1 U10827 ( .B1(SI_7_), .B2(keyinput_25), .C1(n10057), .C2(
        keyinput_24), .A(n10056), .ZN(n10058) );
  AOI211_X1 U10828 ( .C1(SI_9_), .C2(keyinput_23), .A(n10059), .B(n10058), 
        .ZN(n10060) );
  OAI21_X1 U10829 ( .B1(SI_9_), .B2(keyinput_23), .A(n10060), .ZN(n10061) );
  OAI221_X1 U10830 ( .B1(SI_6_), .B2(n10062), .C1(n10161), .C2(keyinput_26), 
        .A(n10061), .ZN(n10063) );
  OAI221_X1 U10831 ( .B1(SI_5_), .B2(keyinput_27), .C1(n10163), .C2(n10064), 
        .A(n10063), .ZN(n10065) );
  OAI221_X1 U10832 ( .B1(SI_4_), .B2(keyinput_28), .C1(n10166), .C2(n10066), 
        .A(n10065), .ZN(n10067) );
  OAI211_X1 U10833 ( .C1(n10173), .C2(keyinput_29), .A(n10068), .B(n10067), 
        .ZN(n10069) );
  AOI21_X1 U10834 ( .B1(n10173), .B2(keyinput_29), .A(n10069), .ZN(n10077) );
  XOR2_X1 U10835 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .Z(n10071) );
  XNOR2_X1 U10836 ( .A(SI_0_), .B(keyinput_32), .ZN(n10070) );
  NAND2_X1 U10837 ( .A1(n10071), .A2(n10070), .ZN(n10076) );
  OAI22_X1 U10838 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_35), .B1(
        keyinput_37), .B2(P2_REG3_REG_14__SCAN_IN), .ZN(n10072) );
  AOI221_X1 U10839 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_37), .A(n10072), .ZN(n10075) );
  OAI22_X1 U10840 ( .A1(n10176), .A2(keyinput_36), .B1(keyinput_34), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n10073) );
  AOI221_X1 U10841 ( .B1(n10176), .B2(keyinput_36), .C1(P2_STATE_REG_SCAN_IN), 
        .C2(keyinput_34), .A(n10073), .ZN(n10074) );
  OAI211_X1 U10842 ( .C1(n10077), .C2(n10076), .A(n10075), .B(n10074), .ZN(
        n10078) );
  OAI221_X1 U10843 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n10079), .C1(n5894), 
        .C2(keyinput_38), .A(n10078), .ZN(n10084) );
  AOI22_X1 U10844 ( .A1(n10188), .A2(keyinput_41), .B1(keyinput_42), .B2(n5997), .ZN(n10080) );
  OAI221_X1 U10845 ( .B1(n10188), .B2(keyinput_41), .C1(n5997), .C2(
        keyinput_42), .A(n10080), .ZN(n10083) );
  AOI22_X1 U10846 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_43), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .ZN(n10081) );
  OAI221_X1 U10847 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_40), .A(n10081), .ZN(n10082) );
  AOI211_X1 U10848 ( .C1(n10085), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10086) );
  AOI221_X1 U10849 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n10087), .C1(n5438), 
        .C2(keyinput_44), .A(n10086), .ZN(n10088) );
  OAI22_X1 U10850 ( .A1(n10089), .A2(n10088), .B1(keyinput_47), .B2(
        P2_REG3_REG_25__SCAN_IN), .ZN(n10090) );
  AOI21_X1 U10851 ( .B1(keyinput_47), .B2(P2_REG3_REG_25__SCAN_IN), .A(n10090), 
        .ZN(n10096) );
  AOI22_X1 U10852 ( .A1(n5394), .A2(keyinput_49), .B1(keyinput_48), .B2(n10200), .ZN(n10091) );
  OAI221_X1 U10853 ( .B1(n5394), .B2(keyinput_49), .C1(n10200), .C2(
        keyinput_48), .A(n10091), .ZN(n10095) );
  OAI22_X1 U10854 ( .A1(n10093), .A2(keyinput_51), .B1(keyinput_50), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n10092) );
  AOI221_X1 U10855 ( .B1(n10093), .B2(keyinput_51), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_50), .A(n10092), .ZN(n10094) );
  OAI21_X1 U10856 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(n10097) );
  AOI22_X1 U10857 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_54), .B1(n10098), 
        .B2(n10097), .ZN(n10101) );
  AOI22_X1 U10858 ( .A1(n10210), .A2(keyinput_55), .B1(n5667), .B2(keyinput_56), .ZN(n10099) );
  OAI221_X1 U10859 ( .B1(n10210), .B2(keyinput_55), .C1(n5667), .C2(
        keyinput_56), .A(n10099), .ZN(n10100) );
  AOI221_X1 U10860 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n10101), .C1(keyinput_54), .C2(n10101), .A(n10100), .ZN(n10110) );
  AOI22_X1 U10861 ( .A1(n10212), .A2(keyinput_57), .B1(n5612), .B2(keyinput_58), .ZN(n10102) );
  OAI221_X1 U10862 ( .B1(n10212), .B2(keyinput_57), .C1(n5612), .C2(
        keyinput_58), .A(n10102), .ZN(n10109) );
  OAI22_X1 U10863 ( .A1(n10105), .A2(keyinput_61), .B1(n10104), .B2(
        keyinput_60), .ZN(n10103) );
  AOI221_X1 U10864 ( .B1(n10105), .B2(keyinput_61), .C1(keyinput_60), .C2(
        n10104), .A(n10103), .ZN(n10108) );
  OAI22_X1 U10865 ( .A1(n5715), .A2(keyinput_63), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(keyinput_62), .ZN(n10106) );
  AOI221_X1 U10866 ( .B1(n5715), .B2(keyinput_63), .C1(keyinput_62), .C2(
        P2_REG3_REG_26__SCAN_IN), .A(n10106), .ZN(n10107) );
  OAI211_X1 U10867 ( .C1(n10110), .C2(n10109), .A(n10108), .B(n10107), .ZN(
        n10219) );
  XNOR2_X1 U10868 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n10218)
         );
  OAI22_X1 U10869 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_126), .B1(
        keyinput_123), .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n10111) );
  AOI221_X1 U10870 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_126), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_123), .A(n10111), .ZN(n10114) );
  OAI22_X1 U10871 ( .A1(n5715), .A2(keyinput_127), .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .ZN(n10112) );
  AOI221_X1 U10872 ( .B1(n5715), .B2(keyinput_127), .C1(keyinput_124), .C2(
        P2_REG3_REG_18__SCAN_IN), .A(n10112), .ZN(n10113) );
  OAI211_X1 U10873 ( .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_125), .A(n10114), .B(n10113), .ZN(n10115) );
  AOI21_X1 U10874 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .A(n10115), 
        .ZN(n10217) );
  AOI22_X1 U10875 ( .A1(n10117), .A2(keyinput_110), .B1(keyinput_109), .B2(
        n5851), .ZN(n10116) );
  OAI221_X1 U10876 ( .B1(n10117), .B2(keyinput_110), .C1(n5851), .C2(
        keyinput_109), .A(n10116), .ZN(n10196) );
  INV_X1 U10877 ( .A(keyinput_108), .ZN(n10194) );
  INV_X1 U10878 ( .A(keyinput_103), .ZN(n10186) );
  INV_X1 U10879 ( .A(keyinput_102), .ZN(n10183) );
  OAI22_X1 U10880 ( .A1(n5208), .A2(keyinput_97), .B1(keyinput_96), .B2(SI_0_), 
        .ZN(n10118) );
  AOI221_X1 U10881 ( .B1(n5208), .B2(keyinput_97), .C1(SI_0_), .C2(keyinput_96), .A(n10118), .ZN(n10181) );
  INV_X1 U10882 ( .A(keyinput_92), .ZN(n10167) );
  INV_X1 U10883 ( .A(keyinput_91), .ZN(n10164) );
  INV_X1 U10884 ( .A(keyinput_90), .ZN(n10160) );
  INV_X1 U10885 ( .A(SI_7_), .ZN(n10120) );
  OAI22_X1 U10886 ( .A1(n10120), .A2(keyinput_89), .B1(SI_8_), .B2(keyinput_88), .ZN(n10119) );
  AOI221_X1 U10887 ( .B1(n10120), .B2(keyinput_89), .C1(keyinput_88), .C2(
        SI_8_), .A(n10119), .ZN(n10157) );
  INV_X1 U10888 ( .A(keyinput_78), .ZN(n10142) );
  OAI22_X1 U10889 ( .A1(n10122), .A2(keyinput_77), .B1(SI_20_), .B2(
        keyinput_76), .ZN(n10121) );
  AOI221_X1 U10890 ( .B1(n10122), .B2(keyinput_77), .C1(keyinput_76), .C2(
        SI_20_), .A(n10121), .ZN(n10139) );
  INV_X1 U10891 ( .A(keyinput_74), .ZN(n10136) );
  XOR2_X1 U10892 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_64), .Z(n10129) );
  OAI22_X1 U10893 ( .A1(SI_30_), .A2(keyinput_66), .B1(keyinput_65), .B2(
        SI_31_), .ZN(n10123) );
  AOI221_X1 U10894 ( .B1(SI_30_), .B2(keyinput_66), .C1(SI_31_), .C2(
        keyinput_65), .A(n10123), .ZN(n10128) );
  AOI22_X1 U10895 ( .A1(SI_28_), .A2(keyinput_68), .B1(SI_27_), .B2(
        keyinput_69), .ZN(n10124) );
  OAI221_X1 U10896 ( .B1(SI_28_), .B2(keyinput_68), .C1(SI_27_), .C2(
        keyinput_69), .A(n10124), .ZN(n10127) );
  AOI22_X1 U10897 ( .A1(SI_29_), .A2(keyinput_67), .B1(SI_26_), .B2(
        keyinput_70), .ZN(n10125) );
  OAI221_X1 U10898 ( .B1(SI_29_), .B2(keyinput_67), .C1(SI_26_), .C2(
        keyinput_70), .A(n10125), .ZN(n10126) );
  AOI211_X1 U10899 ( .C1(n10129), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10133) );
  AOI22_X1 U10900 ( .A1(SI_25_), .A2(keyinput_71), .B1(n10131), .B2(
        keyinput_73), .ZN(n10130) );
  OAI221_X1 U10901 ( .B1(SI_25_), .B2(keyinput_71), .C1(n10131), .C2(
        keyinput_73), .A(n10130), .ZN(n10132) );
  AOI211_X1 U10902 ( .C1(SI_24_), .C2(keyinput_72), .A(n10133), .B(n10132), 
        .ZN(n10134) );
  OAI21_X1 U10903 ( .B1(SI_24_), .B2(keyinput_72), .A(n10134), .ZN(n10135) );
  OAI221_X1 U10904 ( .B1(SI_22_), .B2(keyinput_74), .C1(n10137), .C2(n10136), 
        .A(n10135), .ZN(n10138) );
  OAI211_X1 U10905 ( .C1(SI_21_), .C2(keyinput_75), .A(n10139), .B(n10138), 
        .ZN(n10140) );
  AOI21_X1 U10906 ( .B1(SI_21_), .B2(keyinput_75), .A(n10140), .ZN(n10141) );
  AOI221_X1 U10907 ( .B1(SI_18_), .B2(keyinput_78), .C1(n10143), .C2(n10142), 
        .A(n10141), .ZN(n10155) );
  AOI22_X1 U10908 ( .A1(SI_14_), .A2(keyinput_82), .B1(n10145), .B2(
        keyinput_79), .ZN(n10144) );
  OAI221_X1 U10909 ( .B1(SI_14_), .B2(keyinput_82), .C1(n10145), .C2(
        keyinput_79), .A(n10144), .ZN(n10149) );
  AOI22_X1 U10910 ( .A1(SI_15_), .A2(keyinput_81), .B1(n10147), .B2(
        keyinput_80), .ZN(n10146) );
  OAI221_X1 U10911 ( .B1(SI_15_), .B2(keyinput_81), .C1(n10147), .C2(
        keyinput_80), .A(n10146), .ZN(n10148) );
  AOI211_X1 U10912 ( .C1(keyinput_83), .C2(SI_13_), .A(n10149), .B(n10148), 
        .ZN(n10150) );
  OAI21_X1 U10913 ( .B1(keyinput_83), .B2(SI_13_), .A(n10150), .ZN(n10154) );
  OAI22_X1 U10914 ( .A1(SI_12_), .A2(keyinput_84), .B1(keyinput_86), .B2(
        SI_10_), .ZN(n10151) );
  AOI221_X1 U10915 ( .B1(SI_12_), .B2(keyinput_84), .C1(SI_10_), .C2(
        keyinput_86), .A(n10151), .ZN(n10153) );
  XNOR2_X1 U10916 ( .A(SI_11_), .B(keyinput_85), .ZN(n10152) );
  OAI211_X1 U10917 ( .C1(n10155), .C2(n10154), .A(n10153), .B(n10152), .ZN(
        n10156) );
  OAI211_X1 U10918 ( .C1(SI_9_), .C2(keyinput_87), .A(n10157), .B(n10156), 
        .ZN(n10158) );
  AOI21_X1 U10919 ( .B1(SI_9_), .B2(keyinput_87), .A(n10158), .ZN(n10159) );
  AOI221_X1 U10920 ( .B1(SI_6_), .B2(keyinput_90), .C1(n10161), .C2(n10160), 
        .A(n10159), .ZN(n10162) );
  AOI221_X1 U10921 ( .B1(SI_5_), .B2(n10164), .C1(n10163), .C2(keyinput_91), 
        .A(n10162), .ZN(n10165) );
  AOI221_X1 U10922 ( .B1(SI_4_), .B2(n10167), .C1(n10166), .C2(keyinput_92), 
        .A(n10165), .ZN(n10171) );
  AOI22_X1 U10923 ( .A1(SI_2_), .A2(keyinput_94), .B1(n10169), .B2(keyinput_95), .ZN(n10168) );
  OAI221_X1 U10924 ( .B1(SI_2_), .B2(keyinput_94), .C1(n10169), .C2(
        keyinput_95), .A(n10168), .ZN(n10170) );
  AOI211_X1 U10925 ( .C1(n10173), .C2(keyinput_93), .A(n10171), .B(n10170), 
        .ZN(n10172) );
  OAI21_X1 U10926 ( .B1(n10173), .B2(keyinput_93), .A(n10172), .ZN(n10180) );
  AOI22_X1 U10927 ( .A1(n10176), .A2(keyinput_100), .B1(n10175), .B2(
        keyinput_101), .ZN(n10174) );
  OAI221_X1 U10928 ( .B1(n10176), .B2(keyinput_100), .C1(n10175), .C2(
        keyinput_101), .A(n10174), .ZN(n10179) );
  AOI22_X1 U10929 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_99), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_98), .ZN(n10177) );
  OAI221_X1 U10930 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_98), .A(n10177), .ZN(n10178) );
  AOI211_X1 U10931 ( .C1(n10181), .C2(n10180), .A(n10179), .B(n10178), .ZN(
        n10182) );
  AOI221_X1 U10932 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n10183), .C1(n5894), 
        .C2(keyinput_102), .A(n10182), .ZN(n10184) );
  AOI221_X1 U10933 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(n10186), .C1(n10185), 
        .C2(keyinput_103), .A(n10184), .ZN(n10192) );
  AOI22_X1 U10934 ( .A1(n5997), .A2(keyinput_106), .B1(n10188), .B2(
        keyinput_105), .ZN(n10187) );
  OAI221_X1 U10935 ( .B1(n5997), .B2(keyinput_106), .C1(n10188), .C2(
        keyinput_105), .A(n10187), .ZN(n10191) );
  AOI22_X1 U10936 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .ZN(n10189) );
  OAI221_X1 U10937 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_104), .A(n10189), .ZN(n10190) );
  NOR3_X1 U10938 ( .A1(n10192), .A2(n10191), .A3(n10190), .ZN(n10193) );
  AOI221_X1 U10939 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n10194), .C1(n5438), 
        .C2(keyinput_108), .A(n10193), .ZN(n10195) );
  OAI22_X1 U10940 ( .A1(keyinput_111), .A2(n10198), .B1(n10196), .B2(n10195), 
        .ZN(n10197) );
  AOI21_X1 U10941 ( .B1(keyinput_111), .B2(n10198), .A(n10197), .ZN(n10204) );
  AOI22_X1 U10942 ( .A1(n10200), .A2(keyinput_112), .B1(n5394), .B2(
        keyinput_113), .ZN(n10199) );
  OAI221_X1 U10943 ( .B1(n10200), .B2(keyinput_112), .C1(n5394), .C2(
        keyinput_113), .A(n10199), .ZN(n10203) );
  OAI22_X1 U10944 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_114), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .ZN(n10201) );
  AOI221_X1 U10945 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_114), .C1(
        keyinput_115), .C2(P2_REG3_REG_24__SCAN_IN), .A(n10201), .ZN(n10202)
         );
  OAI21_X1 U10946 ( .B1(n10204), .B2(n10203), .A(n10202), .ZN(n10208) );
  OAI22_X1 U10947 ( .A1(n7902), .A2(keyinput_117), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_116), .ZN(n10205) );
  AOI221_X1 U10948 ( .B1(n7902), .B2(keyinput_117), .C1(keyinput_116), .C2(
        P2_REG3_REG_4__SCAN_IN), .A(n10205), .ZN(n10207) );
  NOR2_X1 U10949 ( .A1(n5425), .A2(keyinput_118), .ZN(n10206) );
  AOI221_X1 U10950 ( .B1(n10208), .B2(n10207), .C1(keyinput_118), .C2(n5425), 
        .A(n10206), .ZN(n10215) );
  AOI22_X1 U10951 ( .A1(n10210), .A2(keyinput_119), .B1(n5667), .B2(
        keyinput_120), .ZN(n10209) );
  OAI221_X1 U10952 ( .B1(n10210), .B2(keyinput_119), .C1(n5667), .C2(
        keyinput_120), .A(n10209), .ZN(n10214) );
  OAI22_X1 U10953 ( .A1(n10212), .A2(keyinput_121), .B1(keyinput_122), .B2(
        P2_REG3_REG_11__SCAN_IN), .ZN(n10211) );
  AOI221_X1 U10954 ( .B1(n10212), .B2(keyinput_121), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_122), .A(n10211), .ZN(n10213)
         );
  OAI21_X1 U10955 ( .B1(n10215), .B2(n10214), .A(n10213), .ZN(n10216) );
  OAI211_X1 U10956 ( .C1(n10219), .C2(n10218), .A(n10217), .B(n10216), .ZN(
        n10220) );
  XNOR2_X1 U10957 ( .A(n10221), .B(n10220), .ZN(P1_U3280) );
  XOR2_X1 U10958 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U10959 ( .A(n10222), .ZN(n10223) );
  NAND2_X1 U10960 ( .A1(n10224), .A2(n10223), .ZN(n10225) );
  XNOR2_X1 U10961 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10225), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U10962 ( .A(n10227), .B(n10226), .Z(ADD_1071_U54) );
  XOR2_X1 U10963 ( .A(n10229), .B(n10228), .Z(ADD_1071_U53) );
  XNOR2_X1 U10964 ( .A(n10231), .B(n10230), .ZN(ADD_1071_U52) );
  NOR2_X1 U10965 ( .A1(n10233), .A2(n10232), .ZN(n10235) );
  XNOR2_X1 U10966 ( .A(n10235), .B(n10234), .ZN(ADD_1071_U51) );
  XNOR2_X1 U10967 ( .A(n10237), .B(n10236), .ZN(ADD_1071_U50) );
  XNOR2_X1 U10968 ( .A(n10239), .B(n10238), .ZN(ADD_1071_U49) );
  XNOR2_X1 U10969 ( .A(n10241), .B(n10240), .ZN(ADD_1071_U48) );
  XNOR2_X1 U10970 ( .A(n10243), .B(n10242), .ZN(ADD_1071_U47) );
  XOR2_X1 U10971 ( .A(n10245), .B(n10244), .Z(ADD_1071_U63) );
  XOR2_X1 U10972 ( .A(n10247), .B(n10246), .Z(ADD_1071_U62) );
  XNOR2_X1 U10973 ( .A(n10249), .B(n10248), .ZN(ADD_1071_U61) );
  XNOR2_X1 U10974 ( .A(n10251), .B(n10250), .ZN(ADD_1071_U60) );
  XNOR2_X1 U10975 ( .A(n10253), .B(n10252), .ZN(ADD_1071_U59) );
  XNOR2_X1 U10976 ( .A(n10255), .B(n10254), .ZN(ADD_1071_U58) );
  XNOR2_X1 U10977 ( .A(n10257), .B(n10256), .ZN(ADD_1071_U57) );
  XNOR2_X1 U10978 ( .A(n10259), .B(n10258), .ZN(ADD_1071_U56) );
  NOR2_X1 U10979 ( .A1(n10261), .A2(n10260), .ZN(n10262) );
  XOR2_X1 U10980 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10262), .Z(ADD_1071_U55)
         );
  INV_X1 U10981 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10449) );
  INV_X1 U10982 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10440) );
  AOI21_X1 U10983 ( .B1(n10263), .B2(n10440), .A(n4847), .ZN(n10405) );
  OAI21_X1 U10984 ( .B1(n10263), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10405), .ZN(
        n10268) );
  AOI211_X1 U10985 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10405), .A(n10265), .B(
        n10264), .ZN(n10266) );
  AOI21_X1 U10986 ( .B1(n10407), .B2(n7189), .A(n10266), .ZN(n10267) );
  AOI21_X1 U10987 ( .B1(n6371), .B2(n10268), .A(n10267), .ZN(n10269) );
  AOI21_X1 U10988 ( .B1(n10436), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n10269), .ZN(
        n10270) );
  OAI21_X1 U10989 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n10449), .A(n10270), .ZN(
        P1_U3241) );
  AOI22_X1 U10990 ( .A1(n10427), .A2(n10271), .B1(n10436), .B2(
        P1_ADDR_REG_6__SCAN_IN), .ZN(n10282) );
  AOI21_X1 U10991 ( .B1(n10274), .B2(n10273), .A(n10272), .ZN(n10275) );
  NAND2_X1 U10992 ( .A1(n10275), .A2(n10426), .ZN(n10280) );
  OAI211_X1 U10993 ( .C1(n10278), .C2(n10277), .A(n10407), .B(n10276), .ZN(
        n10279) );
  NAND4_X1 U10994 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        P1_U3247) );
  INV_X1 U10995 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10298) );
  AND2_X1 U10996 ( .A1(n10284), .A2(n10283), .ZN(n10285) );
  OR3_X1 U10997 ( .A1(n10411), .A2(n10286), .A3(n10285), .ZN(n10289) );
  INV_X1 U10998 ( .A(n10287), .ZN(n10288) );
  OAI211_X1 U10999 ( .C1(n10318), .C2(n10290), .A(n10289), .B(n10288), .ZN(
        n10291) );
  INV_X1 U11000 ( .A(n10291), .ZN(n10297) );
  AOI21_X1 U11001 ( .B1(n10294), .B2(n10293), .A(n10292), .ZN(n10295) );
  OR2_X1 U11002 ( .A1(n10295), .A2(n10433), .ZN(n10296) );
  OAI211_X1 U11003 ( .C1(n10420), .C2(n10298), .A(n10297), .B(n10296), .ZN(
        P1_U3251) );
  INV_X1 U11004 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10312) );
  OAI21_X1 U11005 ( .B1(n10301), .B2(n10300), .A(n10299), .ZN(n10306) );
  INV_X1 U11006 ( .A(n10302), .ZN(n10303) );
  NOR2_X1 U11007 ( .A1(n10318), .A2(n10303), .ZN(n10304) );
  AOI211_X1 U11008 ( .C1(n10407), .C2(n10306), .A(n10305), .B(n10304), .ZN(
        n10311) );
  OAI211_X1 U11009 ( .C1(n10309), .C2(n10308), .A(n10426), .B(n10307), .ZN(
        n10310) );
  OAI211_X1 U11010 ( .C1(n10420), .C2(n10312), .A(n10311), .B(n10310), .ZN(
        P1_U3253) );
  INV_X1 U11011 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10327) );
  OAI21_X1 U11012 ( .B1(n10315), .B2(n10314), .A(n10313), .ZN(n10321) );
  INV_X1 U11013 ( .A(n10316), .ZN(n10317) );
  NOR2_X1 U11014 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  AOI211_X1 U11015 ( .C1(n10407), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        n10326) );
  OAI211_X1 U11016 ( .C1(n10324), .C2(n10323), .A(n10426), .B(n10322), .ZN(
        n10325) );
  OAI211_X1 U11017 ( .C1(n10420), .C2(n10327), .A(n10326), .B(n10325), .ZN(
        P1_U3254) );
  AOI22_X1 U11018 ( .A1(n10427), .A2(n10328), .B1(n10436), .B2(
        P1_ADDR_REG_5__SCAN_IN), .ZN(n10339) );
  OAI21_X1 U11019 ( .B1(n10331), .B2(n10330), .A(n10329), .ZN(n10332) );
  NAND2_X1 U11020 ( .A1(n10426), .A2(n10332), .ZN(n10337) );
  OAI211_X1 U11021 ( .C1(n10335), .C2(n10334), .A(n10407), .B(n10333), .ZN(
        n10336) );
  NAND4_X1 U11022 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        P1_U3246) );
  AOI22_X1 U11023 ( .A1(n10427), .A2(n10340), .B1(n10436), .B2(
        P1_ADDR_REG_3__SCAN_IN), .ZN(n10351) );
  AOI21_X1 U11024 ( .B1(n10343), .B2(n10342), .A(n10341), .ZN(n10344) );
  NAND2_X1 U11025 ( .A1(n10426), .A2(n10344), .ZN(n10349) );
  OAI211_X1 U11026 ( .C1(n10347), .C2(n10346), .A(n10407), .B(n10345), .ZN(
        n10348) );
  NAND4_X1 U11027 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        P1_U3244) );
  AOI22_X1 U11028 ( .A1(n10355), .A2(n10354), .B1(n10353), .B2(n10352), .ZN(
        P2_U3437) );
  OAI211_X1 U11029 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10357), .A(n10356), .B(
        P2_IR_REG_0__SCAN_IN), .ZN(n10358) );
  AOI21_X1 U11030 ( .B1(n10359), .B2(n5424), .A(n10358), .ZN(n10363) );
  AOI22_X1 U11031 ( .A1(n10359), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n10391), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10362) );
  INV_X1 U11032 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U11033 ( .A1(n10379), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10360) );
  OAI221_X1 U11034 ( .B1(n10363), .B2(n10362), .C1(n10363), .C2(n10361), .A(
        n10360), .ZN(P2_U3245) );
  AOI22_X1 U11035 ( .A1(n10379), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10378) );
  NAND2_X1 U11036 ( .A1(n10365), .A2(n10364), .ZN(n10367) );
  NAND2_X1 U11037 ( .A1(n10367), .A2(n10366), .ZN(n10375) );
  NAND2_X1 U11038 ( .A1(n10386), .A2(n10368), .ZN(n10374) );
  AOI21_X1 U11039 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(n10372) );
  NAND2_X1 U11040 ( .A1(n10391), .A2(n10372), .ZN(n10373) );
  OAI211_X1 U11041 ( .C1(n10375), .C2(n10394), .A(n10374), .B(n10373), .ZN(
        n10376) );
  INV_X1 U11042 ( .A(n10376), .ZN(n10377) );
  NAND2_X1 U11043 ( .A1(n10378), .A2(n10377), .ZN(P2_U3246) );
  AOI22_X1 U11044 ( .A1(n10379), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10398) );
  NAND2_X1 U11045 ( .A1(n10381), .A2(n10380), .ZN(n10384) );
  INV_X1 U11046 ( .A(n10382), .ZN(n10383) );
  NAND2_X1 U11047 ( .A1(n10384), .A2(n10383), .ZN(n10395) );
  NAND2_X1 U11048 ( .A1(n10386), .A2(n10385), .ZN(n10393) );
  AOI21_X1 U11049 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(n10390) );
  NAND2_X1 U11050 ( .A1(n10391), .A2(n10390), .ZN(n10392) );
  OAI211_X1 U11051 ( .C1(n10395), .C2(n10394), .A(n10393), .B(n10392), .ZN(
        n10396) );
  INV_X1 U11052 ( .A(n10396), .ZN(n10397) );
  NAND2_X1 U11053 ( .A1(n10398), .A2(n10397), .ZN(P2_U3247) );
  XNOR2_X1 U11054 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11055 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10421) );
  INV_X1 U11056 ( .A(n10399), .ZN(n10401) );
  MUX2_X1 U11057 ( .A(n10401), .B(n10400), .S(n4848), .Z(n10403) );
  NAND2_X1 U11058 ( .A1(n10403), .A2(n10402), .ZN(n10404) );
  OAI211_X1 U11059 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10405), .A(n10404), .B(
        P1_U4006), .ZN(n10437) );
  OAI211_X1 U11060 ( .C1(n10409), .C2(n10408), .A(n10407), .B(n10406), .ZN(
        n10410) );
  OAI21_X1 U11061 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7495), .A(n10410), .ZN(
        n10416) );
  AOI211_X1 U11062 ( .C1(n10414), .C2(n10413), .A(n10412), .B(n10411), .ZN(
        n10415) );
  AOI211_X1 U11063 ( .C1(n10427), .C2(n10417), .A(n10416), .B(n10415), .ZN(
        n10418) );
  AND2_X1 U11064 ( .A1(n10437), .A2(n10418), .ZN(n10419) );
  OAI21_X1 U11065 ( .B1(n10421), .B2(n10420), .A(n10419), .ZN(P1_U3243) );
  OAI21_X1 U11066 ( .B1(n10424), .B2(n10423), .A(n10422), .ZN(n10425) );
  AOI22_X1 U11067 ( .A1(n10428), .A2(n10427), .B1(n10426), .B2(n10425), .ZN(
        n10439) );
  AOI21_X1 U11068 ( .B1(n10431), .B2(n10430), .A(n10429), .ZN(n10432) );
  NOR2_X1 U11069 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  AOI211_X1 U11070 ( .C1(n10436), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n10435), .B(
        n10434), .ZN(n10438) );
  NAND3_X1 U11071 ( .A1(n10439), .A2(n10438), .A3(n10437), .ZN(P1_U3245) );
  NOR2_X1 U11072 ( .A1(n10447), .A2(n10440), .ZN(n10445) );
  AOI21_X1 U11073 ( .B1(n10443), .B2(n10442), .A(n10441), .ZN(n10444) );
  AOI211_X1 U11074 ( .C1(n10447), .C2(n10446), .A(n10445), .B(n10444), .ZN(
        n10448) );
  OAI21_X1 U11075 ( .B1(n10450), .B2(n10449), .A(n10448), .ZN(P1_U3291) );
  INV_X1 U11076 ( .A(n10451), .ZN(n10455) );
  OAI22_X1 U11077 ( .A1(n10453), .A2(n10564), .B1(n10452), .B2(n10470), .ZN(
        n10454) );
  NOR2_X1 U11078 ( .A1(n10455), .A2(n10454), .ZN(n10457) );
  INV_X1 U11079 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U11080 ( .A1(n10584), .A2(n10457), .B1(n10456), .B2(n10583), .ZN(
        P2_U3520) );
  AOI22_X1 U11081 ( .A1(n10588), .A2(n10457), .B1(n5423), .B2(n10585), .ZN(
        P2_U3451) );
  OAI21_X1 U11082 ( .B1(n10459), .B2(n10537), .A(n10458), .ZN(n10461) );
  AOI211_X1 U11083 ( .C1(n10463), .C2(n10462), .A(n10461), .B(n10460), .ZN(
        n10464) );
  AOI22_X1 U11084 ( .A1(n4842), .A2(n10464), .B1(n6847), .B2(n10542), .ZN(
        P1_U3524) );
  AOI22_X1 U11085 ( .A1(n4843), .A2(n10464), .B1(n6354), .B2(n10543), .ZN(
        P1_U3457) );
  XOR2_X1 U11086 ( .A(n10465), .B(n10473), .Z(n10468) );
  AOI21_X1 U11087 ( .B1(n10468), .B2(n10467), .A(n10466), .ZN(n10483) );
  OAI21_X1 U11088 ( .B1(n10481), .B2(n10470), .A(n10469), .ZN(n10482) );
  OAI22_X1 U11089 ( .A1(n10472), .A2(n10482), .B1(n5438), .B2(n10471), .ZN(
        n10478) );
  XNOR2_X1 U11090 ( .A(n10474), .B(n10473), .ZN(n10480) );
  OAI22_X1 U11091 ( .A1(n10480), .A2(n10476), .B1(n10475), .B2(n10481), .ZN(
        n10477) );
  AOI211_X1 U11092 ( .C1(n9164), .C2(P2_REG2_REG_1__SCAN_IN), .A(n10478), .B(
        n10477), .ZN(n10479) );
  OAI21_X1 U11093 ( .B1(n9164), .B2(n10483), .A(n10479), .ZN(P2_U3295) );
  INV_X1 U11094 ( .A(n10480), .ZN(n10486) );
  OAI22_X1 U11095 ( .A1(n10482), .A2(n10568), .B1(n10481), .B2(n10566), .ZN(
        n10485) );
  INV_X1 U11096 ( .A(n10483), .ZN(n10484) );
  AOI211_X1 U11097 ( .C1(n10581), .C2(n10486), .A(n10485), .B(n10484), .ZN(
        n10487) );
  AOI22_X1 U11098 ( .A1(n10584), .A2(n10487), .B1(n6762), .B2(n10583), .ZN(
        P2_U3521) );
  AOI22_X1 U11099 ( .A1(n10588), .A2(n10487), .B1(n5435), .B2(n10585), .ZN(
        P2_U3454) );
  AOI22_X1 U11100 ( .A1(n10489), .A2(n10576), .B1(n10575), .B2(n10488), .ZN(
        n10490) );
  AND2_X1 U11101 ( .A1(n10491), .A2(n10490), .ZN(n10493) );
  INV_X1 U11102 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U11103 ( .A1(n10584), .A2(n10493), .B1(n10492), .B2(n10583), .ZN(
        P2_U3523) );
  AOI22_X1 U11104 ( .A1(n10588), .A2(n10493), .B1(n5410), .B2(n10585), .ZN(
        P2_U3460) );
  NOR2_X1 U11105 ( .A1(n10495), .A2(n10494), .ZN(n10499) );
  OAI21_X1 U11106 ( .B1(n10497), .B2(n10537), .A(n10496), .ZN(n10498) );
  NOR3_X1 U11107 ( .A1(n10500), .A2(n10499), .A3(n10498), .ZN(n10502) );
  AOI22_X1 U11108 ( .A1(n4842), .A2(n10502), .B1(n6852), .B2(n10542), .ZN(
        P1_U3528) );
  INV_X1 U11109 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U11110 ( .A1(n4843), .A2(n10502), .B1(n10501), .B2(n10543), .ZN(
        P1_U3469) );
  NOR2_X1 U11111 ( .A1(n10503), .A2(n10564), .ZN(n10508) );
  OAI22_X1 U11112 ( .A1(n10505), .A2(n10568), .B1(n10504), .B2(n10566), .ZN(
        n10507) );
  AOI211_X1 U11113 ( .C1(n10508), .C2(n7974), .A(n10507), .B(n10506), .ZN(
        n10510) );
  AOI22_X1 U11114 ( .A1(n10584), .A2(n10510), .B1(n6972), .B2(n10583), .ZN(
        P2_U3526) );
  INV_X1 U11115 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U11116 ( .A1(n10588), .A2(n10510), .B1(n10509), .B2(n10585), .ZN(
        P2_U3469) );
  OAI22_X1 U11117 ( .A1(n10512), .A2(n10568), .B1(n10511), .B2(n10566), .ZN(
        n10514) );
  AOI211_X1 U11118 ( .C1(n10581), .C2(n10515), .A(n10514), .B(n10513), .ZN(
        n10517) );
  AOI22_X1 U11119 ( .A1(n10584), .A2(n10517), .B1(n6976), .B2(n10583), .ZN(
        P2_U3527) );
  INV_X1 U11120 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U11121 ( .A1(n10588), .A2(n10517), .B1(n10516), .B2(n10585), .ZN(
        P2_U3472) );
  NAND3_X1 U11122 ( .A1(n10519), .A2(n10518), .A3(n10581), .ZN(n10523) );
  NAND2_X1 U11123 ( .A1(n10520), .A2(n10575), .ZN(n10521) );
  AND4_X1 U11124 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10526) );
  AOI22_X1 U11125 ( .A1(n10584), .A2(n10526), .B1(n6977), .B2(n10583), .ZN(
        P2_U3528) );
  INV_X1 U11126 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U11127 ( .A1(n10588), .A2(n10526), .B1(n10525), .B2(n10585), .ZN(
        P2_U3475) );
  INV_X1 U11128 ( .A(n10527), .ZN(n10528) );
  OAI22_X1 U11129 ( .A1(n10529), .A2(n10568), .B1(n10528), .B2(n10566), .ZN(
        n10531) );
  AOI211_X1 U11130 ( .C1(n10581), .C2(n10532), .A(n10531), .B(n10530), .ZN(
        n10534) );
  AOI22_X1 U11131 ( .A1(n10584), .A2(n10534), .B1(n10533), .B2(n10583), .ZN(
        P2_U3529) );
  AOI22_X1 U11132 ( .A1(n10588), .A2(n10534), .B1(n5567), .B2(n10585), .ZN(
        P2_U3478) );
  OAI211_X1 U11133 ( .C1(n10538), .C2(n10537), .A(n10536), .B(n10535), .ZN(
        n10539) );
  AOI21_X1 U11134 ( .B1(n10541), .B2(n10540), .A(n10539), .ZN(n10544) );
  AOI22_X1 U11135 ( .A1(n4842), .A2(n10544), .B1(n7208), .B2(n10542), .ZN(
        P1_U3533) );
  AOI22_X1 U11136 ( .A1(n4843), .A2(n10544), .B1(n6282), .B2(n10543), .ZN(
        P1_U3484) );
  NOR2_X1 U11137 ( .A1(n10545), .A2(n10564), .ZN(n10549) );
  OAI22_X1 U11138 ( .A1(n10546), .A2(n10568), .B1(n5171), .B2(n10566), .ZN(
        n10548) );
  AOI211_X1 U11139 ( .C1(n10549), .C2(n8138), .A(n10548), .B(n10547), .ZN(
        n10551) );
  AOI22_X1 U11140 ( .A1(n10584), .A2(n10551), .B1(n7083), .B2(n10583), .ZN(
        P2_U3530) );
  INV_X1 U11141 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U11142 ( .A1(n10588), .A2(n10551), .B1(n10550), .B2(n10585), .ZN(
        P2_U3481) );
  OAI211_X1 U11143 ( .C1(n10554), .C2(n10566), .A(n10553), .B(n10552), .ZN(
        n10555) );
  AOI21_X1 U11144 ( .B1(n10581), .B2(n10556), .A(n10555), .ZN(n10557) );
  AOI22_X1 U11145 ( .A1(n10584), .A2(n10557), .B1(n7195), .B2(n10583), .ZN(
        P2_U3531) );
  AOI22_X1 U11146 ( .A1(n10588), .A2(n10557), .B1(n5615), .B2(n10585), .ZN(
        P2_U3484) );
  OAI22_X1 U11147 ( .A1(n10559), .A2(n10568), .B1(n10558), .B2(n10566), .ZN(
        n10561) );
  AOI211_X1 U11148 ( .C1(n10581), .C2(n10562), .A(n10561), .B(n10560), .ZN(
        n10563) );
  AOI22_X1 U11149 ( .A1(n10584), .A2(n10563), .B1(n7464), .B2(n10583), .ZN(
        P2_U3532) );
  AOI22_X1 U11150 ( .A1(n10588), .A2(n10563), .B1(n5645), .B2(n10585), .ZN(
        P2_U3487) );
  NOR2_X1 U11151 ( .A1(n10565), .A2(n10564), .ZN(n10572) );
  OAI22_X1 U11152 ( .A1(n10569), .A2(n10568), .B1(n10567), .B2(n10566), .ZN(
        n10571) );
  AOI211_X1 U11153 ( .C1(n10572), .C2(n8398), .A(n10571), .B(n10570), .ZN(
        n10573) );
  AOI22_X1 U11154 ( .A1(n10584), .A2(n10573), .B1(n7463), .B2(n10583), .ZN(
        P2_U3533) );
  AOI22_X1 U11155 ( .A1(n10588), .A2(n10573), .B1(n5670), .B2(n10585), .ZN(
        P2_U3490) );
  AOI22_X1 U11156 ( .A1(n10577), .A2(n10576), .B1(n10575), .B2(n10574), .ZN(
        n10578) );
  NAND2_X1 U11157 ( .A1(n10579), .A2(n10578), .ZN(n10580) );
  AOI21_X1 U11158 ( .B1(n10582), .B2(n10581), .A(n10580), .ZN(n10587) );
  AOI22_X1 U11159 ( .A1(n10584), .A2(n10587), .B1(n5689), .B2(n10583), .ZN(
        P2_U3534) );
  INV_X1 U11160 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U11161 ( .A1(n10588), .A2(n10587), .B1(n10586), .B2(n10585), .ZN(
        P2_U3493) );
  XNOR2_X1 U11162 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U4910 ( .A(n6376), .ZN(n6535) );
  CLKBUF_X1 U4919 ( .A(n8939), .Z(n4841) );
  AOI211_X1 U4935 ( .C1(n9406), .C2(n9396), .A(n8892), .B(n8891), .ZN(n8893)
         );
  CLKBUF_X1 U9905 ( .A(n6734), .Z(n4847) );
endmodule

