

module b22_C_SARLock_k_64_2 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6439, n6440, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15226, n15228;

  NAND2_X1 U7188 ( .A1(n7915), .A2(n12658), .ZN(n9645) );
  NAND2_X1 U7189 ( .A1(n7336), .A2(n9326), .ZN(n13222) );
  NOR2_X1 U7190 ( .A1(n9996), .A2(n9995), .ZN(n14849) );
  CLKBUF_X2 U7191 ( .A(n11411), .Z(n12799) );
  INV_X1 U7192 ( .A(n9321), .ZN(n9395) );
  INV_X1 U7193 ( .A(n13290), .ZN(n12116) );
  AOI22_X1 U7194 ( .A1(n9680), .A2(n6450), .B1(n13829), .B2(n14738), .ZN(n9682) );
  CLKBUF_X1 U7195 ( .A(n9679), .Z(n6450) );
  AND2_X2 U7197 ( .A1(n9656), .A2(n9797), .ZN(n9675) );
  AND4_X1 U7199 ( .A1(n8185), .A2(n8184), .A3(n8183), .A4(n8182), .ZN(n11273)
         );
  OR2_X1 U7200 ( .A1(n9044), .A2(n9043), .ZN(n12073) );
  NOR2_X1 U7201 ( .A1(n8169), .A2(n8194), .ZN(n14074) );
  BUF_X1 U7202 ( .A(n14039), .Z(n6651) );
  INV_X1 U7203 ( .A(n8180), .ZN(n8512) );
  NAND2_X1 U7204 ( .A1(n7478), .A2(n13132), .ZN(n13138) );
  XNOR2_X1 U7205 ( .A(n8066), .B(n8067), .ZN(n8072) );
  CLKBUF_X1 U7206 ( .A(n12453), .Z(n6439) );
  NOR2_X1 U7207 ( .A1(n8938), .A2(n8937), .ZN(n12453) );
  INV_X1 U7208 ( .A(n15226), .ZN(n6440) );
  INV_X2 U7209 ( .A(n6440), .ZN(P1_U3086) );
  INV_X1 U7210 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n15226) );
  INV_X2 U7212 ( .A(n15228), .ZN(P1_U4016) );
  AND2_X1 U7213 ( .A1(n12659), .A2(n6510), .ZN(n7089) );
  CLKBUF_X2 U7214 ( .A(n12103), .Z(n12254) );
  INV_X2 U7215 ( .A(n8791), .ZN(n8795) );
  NOR2_X1 U7216 ( .A1(n9797), .A2(n9667), .ZN(n9668) );
  INV_X2 U7217 ( .A(n12688), .ZN(n11411) );
  INV_X1 U7218 ( .A(n12656), .ZN(n6458) );
  NAND2_X1 U7219 ( .A1(n6451), .A2(n12334), .ZN(n9321) );
  INV_X1 U7220 ( .A(n11800), .ZN(n11788) );
  INV_X1 U7221 ( .A(n6646), .ZN(n12486) );
  INV_X1 U7222 ( .A(n13164), .ZN(n9331) );
  AND2_X1 U7223 ( .A1(n6687), .A2(n8979), .ZN(n12235) );
  NOR3_X1 U7224 ( .A1(n14849), .A2(n14848), .A3(n14847), .ZN(n14846) );
  INV_X1 U7225 ( .A(n12073), .ZN(n10736) );
  INV_X1 U7226 ( .A(n13921), .ZN(n13865) );
  NAND2_X1 U7227 ( .A1(n8699), .A2(n8698), .ZN(n8712) );
  NAND2_X1 U7228 ( .A1(n7921), .A2(n7920), .ZN(n12662) );
  XNOR2_X1 U7229 ( .A(n11329), .B(n11330), .ZN(n10897) );
  XNOR2_X1 U7230 ( .A(n7523), .B(n7522), .ZN(n10182) );
  INV_X1 U7231 ( .A(n13925), .ZN(n14407) );
  AND2_X1 U7232 ( .A1(n8313), .A2(n8312), .ZN(n11621) );
  NOR2_X1 U7233 ( .A1(n11866), .A2(n7447), .ZN(n11945) );
  AND2_X1 U7234 ( .A1(n9797), .A2(n9857), .ZN(n10343) );
  XNOR2_X1 U7235 ( .A(n7490), .B(n7489), .ZN(n7491) );
  AND2_X1 U7236 ( .A1(n9267), .A2(n9266), .ZN(n13781) );
  INV_X1 U7237 ( .A(n6481), .ZN(n6448) );
  AND3_X1 U7238 ( .A1(n8052), .A2(n8051), .A3(n8346), .ZN(n6444) );
  AND2_X1 U7239 ( .A1(n13504), .A2(n13407), .ZN(n6445) );
  INV_X1 U7240 ( .A(n7510), .ZN(n6446) );
  OR2_X2 U7242 ( .A1(n10910), .A2(n11330), .ZN(n6688) );
  OAI21_X2 U7243 ( .B1(n12135), .B2(n12134), .A(n12133), .ZN(n12137) );
  AND2_X2 U7244 ( .A1(n6697), .A2(n6696), .ZN(n12135) );
  AND2_X2 U7245 ( .A1(n11023), .A2(n7951), .ZN(n11466) );
  NAND4_X2 U7246 ( .A1(n8098), .A2(n8097), .A3(n8096), .A4(n8095), .ZN(n9679)
         );
  NOR2_X2 U7247 ( .A1(n14449), .A2(n14306), .ZN(n14291) );
  OAI21_X2 U7249 ( .B1(n7917), .B2(n7916), .A(n7918), .ZN(n8902) );
  NOR2_X4 U7250 ( .A1(n13496), .A2(n13763), .ZN(n13482) );
  OAI21_X1 U7251 ( .B1(n11816), .B2(n7064), .A(n7063), .ZN(n11935) );
  NAND2_X1 U7252 ( .A1(n9013), .A2(n6619), .ZN(n13795) );
  INV_X4 U7254 ( .A(n6446), .ZN(n6447) );
  INV_X4 U7255 ( .A(n6448), .ZN(n6449) );
  OAI21_X2 U7256 ( .B1(n13570), .B2(n13361), .A(n13363), .ZN(n13558) );
  NOR2_X2 U7257 ( .A1(n14562), .A2(n14563), .ZN(n14561) );
  NAND2_X4 U7258 ( .A1(n9247), .A2(n9246), .ZN(n14620) );
  OAI21_X2 U7259 ( .B1(n11934), .B2(n7959), .A(n7732), .ZN(n12987) );
  OR2_X2 U7260 ( .A1(n12531), .A2(n10641), .ZN(n8920) );
  NAND2_X2 U7261 ( .A1(n12705), .A2(n7939), .ZN(n12524) );
  AND2_X2 U7262 ( .A1(n12754), .A2(n12753), .ZN(n12784) );
  NOR2_X4 U7263 ( .A1(n13573), .A2(n13715), .ZN(n13561) );
  XNOR2_X2 U7264 ( .A(n14888), .B(n13291), .ZN(n12303) );
  OAI21_X2 U7265 ( .B1(n10764), .B2(n10763), .A(n10765), .ZN(n10767) );
  NAND2_X1 U7266 ( .A1(n10749), .A2(n10748), .ZN(n10764) );
  NOR2_X2 U7267 ( .A1(n14214), .A2(n7112), .ZN(n14215) );
  AOI21_X2 U7268 ( .B1(n8500), .B2(n6840), .A(n6839), .ZN(n8538) );
  NAND2_X2 U7269 ( .A1(n7477), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7474) );
  NAND2_X2 U7270 ( .A1(n7234), .A2(n7237), .ZN(n13448) );
  AND2_X1 U7271 ( .A1(n10523), .A2(n12331), .ZN(n6451) );
  AND2_X1 U7272 ( .A1(n10523), .A2(n12331), .ZN(n13639) );
  NAND2_X2 U7273 ( .A1(n7958), .A2(n7957), .ZN(n11816) );
  OAI21_X2 U7274 ( .B1(n14215), .B2(n12040), .A(n12041), .ZN(n12043) );
  OAI21_X2 U7275 ( .B1(n11070), .B2(n7195), .A(n7191), .ZN(n9719) );
  OAI22_X2 U7276 ( .A1(n10956), .A2(n9701), .B1(n10954), .B2(n10953), .ZN(
        n11070) );
  AND2_X2 U7277 ( .A1(n10896), .A2(n10895), .ZN(n11329) );
  NOR2_X2 U7278 ( .A1(n11414), .A2(n11415), .ZN(n11692) );
  NOR2_X2 U7279 ( .A1(n11311), .A2(n11310), .ZN(n11414) );
  NAND2_X2 U7280 ( .A1(n6961), .A2(n6962), .ZN(n14303) );
  AOI21_X2 U7281 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n10002), .A(n14828), .ZN(
        n9996) );
  XNOR2_X2 U7282 ( .A(n13296), .B(n12076), .ZN(n12297) );
  NOR2_X2 U7283 ( .A1(n9558), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n9557) );
  XNOR2_X2 U7284 ( .A(n12014), .B(n12013), .ZN(n14405) );
  XNOR2_X2 U7285 ( .A(n7122), .B(n8065), .ZN(n14524) );
  NAND2_X4 U7286 ( .A1(n9770), .A2(n8138), .ZN(n14355) );
  XNOR2_X2 U7287 ( .A(n8084), .B(n8083), .ZN(n8138) );
  CLKBUF_X1 U7288 ( .A(n10182), .Z(n6452) );
  CLKBUF_X2 U7289 ( .A(n10182), .Z(n6453) );
  CLKBUF_X2 U7290 ( .A(n10182), .Z(n6454) );
  XNOR2_X1 U7291 ( .A(n7490), .B(n7489), .ZN(n6455) );
  AOI21_X1 U7292 ( .B1(n6975), .B2(n6974), .A(n6606), .ZN(n6973) );
  AOI21_X1 U7293 ( .B1(n6694), .B2(n13635), .A(n13381), .ZN(n13670) );
  NAND2_X1 U7294 ( .A1(n12867), .A2(n7977), .ZN(n12855) );
  AND3_X1 U7295 ( .A1(n6549), .A2(n6786), .A3(n6626), .ZN(n12003) );
  AOI21_X2 U7296 ( .B1(n7449), .B2(n7322), .A(n6559), .ZN(n6826) );
  NAND2_X1 U7297 ( .A1(n8715), .A2(n8714), .ZN(n14404) );
  INV_X2 U7298 ( .A(n13428), .ZN(n13674) );
  NAND2_X4 U7299 ( .A1(n9646), .A2(n12522), .ZN(n12663) );
  XNOR2_X1 U7300 ( .A(n8712), .B(n8711), .ZN(n12250) );
  AOI21_X1 U7301 ( .B1(n13222), .B2(n13151), .A(n13229), .ZN(n9347) );
  INV_X1 U7302 ( .A(n12095), .ZN(n12097) );
  AOI21_X1 U7303 ( .B1(n11318), .B2(n11317), .A(n11316), .ZN(n14957) );
  INV_X2 U7304 ( .A(n15210), .ZN(n13649) );
  INV_X4 U7305 ( .A(n12254), .ZN(n12277) );
  INV_X1 U7306 ( .A(n8352), .ZN(n8487) );
  INV_X1 U7307 ( .A(n13293), .ZN(n12096) );
  INV_X1 U7308 ( .A(n11002), .ZN(n12703) );
  NOR2_X2 U7309 ( .A1(n14986), .A2(n12529), .ZN(n14985) );
  CLKBUF_X2 U7310 ( .A(P2_U3947), .Z(n6457) );
  CLKBUF_X2 U7311 ( .A(n6650), .Z(n6618) );
  INV_X1 U7312 ( .A(n12072), .ZN(n12103) );
  NAND4_X2 U7313 ( .A1(n8123), .A2(n8122), .A3(n8121), .A4(n8120), .ZN(n14740)
         );
  INV_X2 U7315 ( .A(n9027), .ZN(n12239) );
  CLKBUF_X2 U7316 ( .A(n8180), .Z(n8382) );
  AND2_X2 U7317 ( .A1(n8980), .A2(n8979), .ZN(n9026) );
  AND2_X1 U7318 ( .A1(n7480), .A2(n13138), .ZN(n6481) );
  AND2_X2 U7319 ( .A1(n13138), .A2(n12037), .ZN(n12473) );
  OR2_X1 U7320 ( .A1(n10218), .A2(n10827), .ZN(n10216) );
  NAND2_X2 U7321 ( .A1(n14055), .A2(n14524), .ZN(n8113) );
  XNOR2_X1 U7322 ( .A(n9011), .B(n9010), .ZN(n9499) );
  INV_X8 U7323 ( .A(n9014), .ZN(n9842) );
  AND2_X1 U7324 ( .A1(n8063), .A2(n7010), .ZN(n8086) );
  INV_X1 U7325 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7994) );
  NOR2_X1 U7326 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7458) );
  NOR2_X1 U7327 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n7457) );
  INV_X1 U7328 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7311) );
  OAI21_X1 U7329 ( .B1(n14001), .B2(n7161), .A(n7160), .ZN(n7162) );
  AOI21_X1 U7330 ( .B1(n12461), .B2(n12462), .A(n6551), .ZN(n12346) );
  AND2_X1 U7331 ( .A1(n12326), .A2(n12329), .ZN(n12333) );
  NAND2_X1 U7332 ( .A1(n13432), .A2(n6528), .ZN(n13419) );
  OR2_X1 U7333 ( .A1(n12327), .A2(n12334), .ZN(n12326) );
  INV_X1 U7334 ( .A(n7992), .ZN(n6763) );
  XNOR2_X1 U7335 ( .A(n8892), .B(n8890), .ZN(n12443) );
  CLKBUF_X1 U7336 ( .A(n13703), .Z(n6755) );
  NOR2_X1 U7337 ( .A1(n12752), .A2(n13035), .ZN(n12770) );
  XNOR2_X1 U7338 ( .A(n8719), .B(n8718), .ZN(n12232) );
  NOR2_X1 U7339 ( .A1(n13412), .A2(n7236), .ZN(n7235) );
  XNOR2_X1 U7340 ( .A(n6880), .B(n12778), .ZN(n12752) );
  NAND2_X2 U7341 ( .A1(n6632), .A2(n8680), .ZN(n14412) );
  NAND2_X1 U7342 ( .A1(n9434), .A2(n9433), .ZN(n13446) );
  NAND2_X1 U7343 ( .A1(n13981), .A2(n13980), .ZN(n13828) );
  OAI21_X1 U7344 ( .B1(n8712), .B2(n8711), .A(n8713), .ZN(n8719) );
  NAND2_X1 U7345 ( .A1(n13913), .A2(n13823), .ZN(n13981) );
  NAND2_X1 U7346 ( .A1(n9016), .A2(n9015), .ZN(n13681) );
  NAND2_X1 U7347 ( .A1(n9347), .A2(n6802), .ZN(n13232) );
  NAND2_X1 U7348 ( .A1(n12923), .A2(n6533), .ZN(n12910) );
  NAND2_X1 U7349 ( .A1(n12924), .A2(n12925), .ZN(n12923) );
  CLKBUF_X1 U7350 ( .A(n13541), .Z(n6614) );
  NAND2_X1 U7351 ( .A1(n9413), .A2(n9412), .ZN(n13763) );
  NAND2_X1 U7352 ( .A1(n12937), .A2(n7968), .ZN(n12924) );
  OAI21_X1 U7353 ( .B1(n12922), .B2(n7379), .A(n7375), .ZN(n12899) );
  NAND2_X1 U7354 ( .A1(n7881), .A2(n7880), .ZN(n13071) );
  NAND2_X1 U7355 ( .A1(n13205), .A2(n13206), .ZN(n13204) );
  NAND2_X1 U7356 ( .A1(n13192), .A2(n9294), .ZN(n13205) );
  CLKBUF_X1 U7357 ( .A(n12978), .Z(n6766) );
  NAND2_X1 U7358 ( .A1(n7891), .A2(n7879), .ZN(n7890) );
  NAND2_X1 U7359 ( .A1(n13610), .A2(n13391), .ZN(n13605) );
  NAND2_X1 U7360 ( .A1(n13349), .A2(n13348), .ZN(n13629) );
  AND2_X1 U7361 ( .A1(n6793), .A2(n7118), .ZN(n6792) );
  NAND2_X1 U7362 ( .A1(n7057), .A2(n7056), .ZN(n13349) );
  AND2_X1 U7363 ( .A1(n9313), .A2(n9312), .ZN(n13593) );
  NAND2_X1 U7364 ( .A1(n8581), .A2(SI_22_), .ZN(n8600) );
  OR2_X1 U7365 ( .A1(n7823), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U7366 ( .A1(n14016), .A2(n14029), .ZN(n6500) );
  AOI21_X1 U7367 ( .B1(n7194), .B2(n7193), .A(n7192), .ZN(n7191) );
  OR2_X1 U7368 ( .A1(n7821), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7822) );
  INV_X1 U7369 ( .A(n11344), .ZN(n11346) );
  NAND2_X1 U7370 ( .A1(n12377), .A2(n6534), .ZN(n11380) );
  NAND2_X1 U7371 ( .A1(n12379), .A2(n12378), .ZN(n12377) );
  NAND2_X1 U7372 ( .A1(n8400), .A2(n8399), .ZN(n11951) );
  NOR2_X1 U7373 ( .A1(n11477), .A2(n6971), .ZN(n6970) );
  OR2_X1 U7374 ( .A1(n8408), .A2(n8446), .ZN(n8427) );
  NAND2_X1 U7375 ( .A1(n8330), .A2(n8329), .ZN(n14792) );
  NAND2_X1 U7376 ( .A1(n8426), .A2(n8407), .ZN(n8408) );
  OR2_X1 U7377 ( .A1(n10592), .A2(n10593), .ZN(n10679) );
  OAI21_X1 U7378 ( .B1(n7717), .B2(n6894), .A(n6892), .ZN(n7737) );
  NAND2_X1 U7379 ( .A1(n7244), .A2(n7242), .ZN(n8369) );
  NAND2_X1 U7380 ( .A1(n8324), .A2(n8308), .ZN(n10014) );
  NAND2_X1 U7381 ( .A1(n8280), .A2(n8279), .ZN(n11431) );
  NAND2_X1 U7382 ( .A1(n10628), .A2(n10627), .ZN(n10626) );
  AND2_X1 U7383 ( .A1(n9105), .A2(n9104), .ZN(n12109) );
  NAND2_X1 U7384 ( .A1(n10122), .A2(n10121), .ZN(n10120) );
  NAND2_X1 U7385 ( .A1(n9085), .A2(n9084), .ZN(n12102) );
  AND2_X1 U7386 ( .A1(n8198), .A2(n8197), .ZN(n11132) );
  AND2_X1 U7387 ( .A1(n9674), .A2(n9673), .ZN(n10122) );
  AND2_X1 U7388 ( .A1(n9061), .A2(n9060), .ZN(n12087) );
  INV_X1 U7389 ( .A(n10885), .ZN(n12704) );
  INV_X1 U7390 ( .A(n12064), .ZN(n10517) );
  NAND4_X2 U7391 ( .A1(n6498), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(n13294)
         );
  INV_X4 U7392 ( .A(n12228), .ZN(n12276) );
  NAND4_X2 U7393 ( .A1(n9030), .A2(n9028), .A3(n9029), .A4(n9031), .ZN(n12064)
         );
  NAND4_X1 U7394 ( .A1(n9049), .A2(n9048), .A3(n9047), .A4(n9046), .ZN(n13295)
         );
  INV_X1 U7395 ( .A(n6650), .ZN(n12705) );
  NAND4_X2 U7396 ( .A1(n8156), .A2(n8155), .A3(n8154), .A4(n8153), .ZN(n14038)
         );
  NAND2_X2 U7397 ( .A1(n9658), .A2(n9657), .ZN(n13921) );
  NAND3_X1 U7398 ( .A1(n6938), .A2(n6940), .A3(n6707), .ZN(n10281) );
  INV_X1 U7399 ( .A(n7938), .ZN(n12529) );
  BUF_X2 U7400 ( .A(n9321), .Z(n9255) );
  AOI22_X1 U7401 ( .A1(n10274), .A2(n10273), .B1(n6715), .B2(n10272), .ZN(
        n10536) );
  NAND2_X1 U7402 ( .A1(n8163), .A2(n8162), .ZN(n8187) );
  AND3_X1 U7403 ( .A1(n7526), .A2(n7525), .A3(n7524), .ZN(n10606) );
  CLKBUF_X2 U7404 ( .A(n6952), .Z(n6951) );
  NAND2_X1 U7405 ( .A1(n12229), .A2(n10095), .ZN(n13635) );
  NAND2_X2 U7406 ( .A1(n7334), .A2(n12286), .ZN(n13164) );
  AND2_X1 U7407 ( .A1(n12053), .A2(n13788), .ZN(n9045) );
  AND2_X1 U7408 ( .A1(n8138), .A2(n9655), .ZN(n9656) );
  NAND2_X1 U7409 ( .A1(n8821), .A2(n8824), .ZN(n14535) );
  AND2_X2 U7410 ( .A1(n8142), .A2(n8815), .ZN(n14536) );
  CLKBUF_X3 U7411 ( .A(n12473), .Z(n8931) );
  INV_X2 U7412 ( .A(n9038), .ZN(n12249) );
  NAND2_X1 U7413 ( .A1(n10216), .A2(n10179), .ZN(n10177) );
  MUX2_X1 U7414 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8823), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8824) );
  MUX2_X1 U7415 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8140), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8142) );
  INV_X2 U7416 ( .A(n9244), .ZN(n12251) );
  CLKBUF_X3 U7418 ( .A(n7515), .Z(n12487) );
  AND2_X1 U7419 ( .A1(n8221), .A2(n6827), .ZN(n6737) );
  NAND2_X1 U7420 ( .A1(n13783), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8976) );
  AOI22_X1 U7421 ( .A1(n10199), .A2(n12712), .B1(n10211), .B2(n10127), .ZN(
        n10170) );
  CLKBUF_X1 U7422 ( .A(n8072), .Z(n11962) );
  OR2_X1 U7423 ( .A1(n10220), .A2(n10219), .ZN(n10222) );
  XNOR2_X1 U7424 ( .A(n8978), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8979) );
  OR2_X1 U7425 ( .A1(n8189), .A2(n7218), .ZN(n6827) );
  NAND2_X1 U7426 ( .A1(n8817), .A2(n8816), .ZN(n8822) );
  CLKBUF_X1 U7427 ( .A(n12330), .Z(n6756) );
  MUX2_X1 U7428 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8087), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8091) );
  NAND2_X2 U7429 ( .A1(n12687), .A2(n6455), .ZN(n7980) );
  NAND2_X1 U7430 ( .A1(n9008), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9009) );
  CLKBUF_X1 U7431 ( .A(n12687), .Z(n6710) );
  INV_X2 U7432 ( .A(n13134), .ZN(n13140) );
  XNOR2_X1 U7433 ( .A(n7932), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U7434 ( .A1(n14518), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8069) );
  OR2_X1 U7435 ( .A1(n8068), .A2(n8345), .ZN(n8066) );
  NAND2_X1 U7436 ( .A1(n7216), .A2(SI_3_), .ZN(n8186) );
  NAND2_X1 U7437 ( .A1(n8063), .A2(n8060), .ZN(n8479) );
  XNOR2_X1 U7438 ( .A(n7573), .B(n7310), .ZN(n10243) );
  INV_X1 U7439 ( .A(n8429), .ZN(n6983) );
  CLKBUF_X2 U7440 ( .A(n7241), .Z(n9456) );
  XNOR2_X1 U7441 ( .A(n7540), .B(n7551), .ZN(n10185) );
  OR2_X1 U7442 ( .A1(n7554), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U7443 ( .A1(n9020), .A2(n9019), .ZN(n9952) );
  OAI21_X1 U7444 ( .B1(n7537), .B2(n6905), .A(n7566), .ZN(n6904) );
  NOR2_X1 U7445 ( .A1(n8141), .A2(n8061), .ZN(n8062) );
  AND2_X1 U7446 ( .A1(n7568), .A2(n7550), .ZN(n7566) );
  NAND2_X1 U7447 ( .A1(n8124), .A2(n8054), .ZN(n8165) );
  AND3_X1 U7448 ( .A1(n8964), .A2(n8965), .A3(n8963), .ZN(n9002) );
  AND2_X1 U7449 ( .A1(n8050), .A2(n8049), .ZN(n8053) );
  INV_X1 U7450 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8144) );
  NOR2_X2 U7451 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7521) );
  INV_X1 U7452 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9263) );
  INV_X1 U7453 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7468) );
  NOR2_X1 U7454 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8967) );
  NOR2_X1 U7455 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n8968) );
  NOR2_X1 U7456 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8969) );
  NOR2_X1 U7457 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7459) );
  INV_X1 U7458 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8966) );
  INV_X4 U7459 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7460 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7461 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8986) );
  INV_X1 U7462 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9056) );
  INV_X1 U7463 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8193) );
  INV_X2 U7464 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7522) );
  NOR2_X2 U7465 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8124) );
  INV_X1 U7466 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14200) );
  NOR2_X2 U7467 ( .A1(n6761), .A2(n12059), .ZN(n10113) );
  AND4_X1 U7469 ( .A1(n7239), .A2(n9002), .A3(n8998), .A4(n9000), .ZN(n7238)
         );
  NAND2_X1 U7470 ( .A1(n11556), .A2(n12312), .ZN(n7057) );
  OAI22_X1 U7471 ( .A1(n11542), .A2(n11541), .B1(n12150), .B2(n11540), .ZN(
        n11556) );
  OAI21_X2 U7472 ( .B1(n9640), .B2(n12954), .A(n9639), .ZN(n12822) );
  XNOR2_X2 U7473 ( .A(n8696), .B(n8679), .ZN(n13794) );
  NAND2_X1 U7474 ( .A1(n13794), .A2(n8758), .ZN(n6632) );
  XNOR2_X1 U7475 ( .A(n12784), .B(n12785), .ZN(n12756) );
  MUX2_X1 U7476 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13806), .S(n9033), .Z(n12059)
         );
  AOI22_X2 U7477 ( .A1(n12094), .A2(n12093), .B1(n12092), .B2(n12091), .ZN(
        n12101) );
  OAI21_X1 U7478 ( .B1(n7979), .B2(n12659), .A(n12832), .ZN(n7990) );
  OAI21_X2 U7479 ( .B1(n13586), .B2(n13358), .A(n13360), .ZN(n13570) );
  NOR2_X2 U7480 ( .A1(n14536), .A2(n9655), .ZN(n9770) );
  AND2_X2 U7481 ( .A1(n9018), .A2(n8966), .ZN(n9057) );
  NAND2_X2 U7482 ( .A1(n12690), .A2(n12531), .ZN(n12656) );
  CLKBUF_X1 U7483 ( .A(n12103), .Z(n6459) );
  NOR2_X1 U7484 ( .A1(n9656), .A2(n9671), .ZN(n13876) );
  INV_X1 U7485 ( .A(n9862), .ZN(n6460) );
  INV_X1 U7486 ( .A(n9862), .ZN(n6461) );
  INV_X1 U7487 ( .A(n9244), .ZN(n6462) );
  OR2_X2 U7488 ( .A1(n13508), .A2(n13692), .ZN(n13496) );
  AND2_X2 U7489 ( .A1(n12037), .A2(n7479), .ZN(n7510) );
  NAND2_X1 U7490 ( .A1(n7082), .A2(n7081), .ZN(n7080) );
  AND2_X1 U7491 ( .A1(n7307), .A2(n7471), .ZN(n7082) );
  NOR3_X1 U7492 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .A3(
        P3_IR_REG_13__SCAN_IN), .ZN(n7471) );
  OR2_X1 U7493 ( .A1(n9641), .A2(n12837), .ZN(n12676) );
  OR2_X1 U7494 ( .A1(n13674), .A2(n13436), .ZN(n13374) );
  NOR2_X1 U7495 ( .A1(n13386), .A2(n7271), .ZN(n7270) );
  INV_X1 U7496 ( .A(n7273), .ZN(n7271) );
  NAND2_X1 U7497 ( .A1(n8765), .A2(n11977), .ZN(n11976) );
  OR2_X1 U7498 ( .A1(n14412), .A2(n14005), .ZN(n8765) );
  INV_X1 U7499 ( .A(n14320), .ZN(n11990) );
  NAND2_X1 U7500 ( .A1(n12056), .A2(n8071), .ZN(n8180) );
  NAND2_X1 U7501 ( .A1(n11380), .A2(n6521), .ZN(n12358) );
  NAND2_X1 U7502 ( .A1(n6689), .A2(n6509), .ZN(n6936) );
  INV_X1 U7503 ( .A(n6670), .ZN(n11696) );
  AND4_X1 U7504 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n12955)
         );
  NAND2_X1 U7505 ( .A1(n9460), .A2(n9459), .ZN(n9464) );
  INV_X1 U7506 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9459) );
  INV_X1 U7507 ( .A(n9467), .ZN(n9460) );
  AOI21_X1 U7508 ( .B1(n8314), .B2(n8315), .A(n6557), .ZN(n7009) );
  NAND2_X1 U7509 ( .A1(n7021), .A2(n7020), .ZN(n7026) );
  NAND2_X1 U7510 ( .A1(n7027), .A2(n6500), .ZN(n7021) );
  INV_X1 U7511 ( .A(n8444), .ZN(n7027) );
  NAND2_X1 U7512 ( .A1(n7422), .A2(n7421), .ZN(n7420) );
  INV_X1 U7513 ( .A(n12179), .ZN(n7421) );
  INV_X1 U7514 ( .A(n12178), .ZN(n7422) );
  AND2_X1 U7515 ( .A1(n12178), .A2(n12179), .ZN(n7423) );
  NAND2_X1 U7516 ( .A1(n8588), .A2(n8591), .ZN(n6997) );
  AOI21_X1 U7517 ( .B1(n6992), .B2(n6993), .A(n6991), .ZN(n6990) );
  INV_X1 U7518 ( .A(n7232), .ZN(n7231) );
  OAI21_X1 U7519 ( .B1(n8391), .B2(n7233), .A(n8404), .ZN(n7232) );
  AOI21_X1 U7520 ( .B1(n6836), .B2(n6834), .A(n6833), .ZN(n6832) );
  INV_X1 U7521 ( .A(n8367), .ZN(n6834) );
  INV_X1 U7522 ( .A(n7229), .ZN(n6833) );
  AOI21_X1 U7523 ( .B1(n7231), .B2(n7233), .A(n6553), .ZN(n7229) );
  NAND2_X1 U7524 ( .A1(n7126), .A2(n7125), .ZN(n9515) );
  OR2_X1 U7525 ( .A1(n13054), .A2(n12349), .ZN(n9646) );
  OAI21_X1 U7526 ( .B1(n10178), .B2(n6561), .A(n10243), .ZN(n6943) );
  OR2_X1 U7527 ( .A1(n12726), .A2(n14559), .ZN(n6754) );
  NAND2_X1 U7528 ( .A1(n7980), .A2(n9842), .ZN(n7515) );
  AND2_X1 U7529 ( .A1(n7374), .A2(n7489), .ZN(n7373) );
  INV_X1 U7530 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7467) );
  AND2_X1 U7531 ( .A1(n7464), .A2(n7468), .ZN(n7930) );
  INV_X1 U7532 ( .A(n6910), .ZN(n6909) );
  OAI21_X1 U7533 ( .B1(n7752), .B2(n6911), .A(n7784), .ZN(n6910) );
  NAND2_X1 U7534 ( .A1(n7322), .A2(n9428), .ZN(n7320) );
  AND2_X1 U7535 ( .A1(n13264), .A2(n9430), .ZN(n7325) );
  OR2_X1 U7536 ( .A1(n9373), .A2(n13238), .ZN(n9387) );
  AOI21_X1 U7537 ( .B1(n13558), .B2(n13565), .A(n13365), .ZN(n13541) );
  AND2_X1 U7538 ( .A1(n13348), .A2(n11558), .ZN(n12315) );
  NAND2_X1 U7539 ( .A1(n11513), .A2(n14631), .ZN(n11549) );
  INV_X1 U7540 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9010) );
  AND2_X1 U7541 ( .A1(n9189), .A2(n9188), .ZN(n9208) );
  INV_X1 U7542 ( .A(n9767), .ZN(n7190) );
  OR2_X1 U7543 ( .A1(n14740), .A2(n10727), .ZN(n10921) );
  AND2_X1 U7544 ( .A1(n6497), .A2(n11976), .ZN(n7113) );
  INV_X1 U7545 ( .A(n14476), .ZN(n14356) );
  NAND2_X1 U7546 ( .A1(n8696), .A2(n8695), .ZN(n8699) );
  OR2_X1 U7547 ( .A1(n8624), .A2(n8623), .ZN(n8639) );
  NAND2_X1 U7548 ( .A1(n8585), .A2(n8584), .ZN(n8586) );
  NOR2_X1 U7549 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n8057) );
  NOR2_X1 U7550 ( .A1(n6844), .A2(n6841), .ZN(n6840) );
  NOR2_X1 U7551 ( .A1(n6471), .A2(n7257), .ZN(n6839) );
  NOR2_X1 U7552 ( .A1(n7261), .A2(SI_18_), .ZN(n6844) );
  NOR2_X1 U7553 ( .A1(n7296), .A2(n10615), .ZN(n7295) );
  INV_X1 U7554 ( .A(n8845), .ZN(n7296) );
  NAND2_X1 U7555 ( .A1(n13047), .A2(n12817), .ZN(n7358) );
  INV_X1 U7556 ( .A(n7351), .ZN(n7350) );
  OAI21_X1 U7557 ( .B1(n6487), .B2(n7352), .A(n12676), .ZN(n7351) );
  INV_X1 U7558 ( .A(n7353), .ZN(n7352) );
  OR2_X1 U7559 ( .A1(n11331), .A2(n11332), .ZN(n6875) );
  NAND2_X1 U7560 ( .A1(n6875), .A2(n6874), .ZN(n14950) );
  INV_X1 U7561 ( .A(n14947), .ZN(n6874) );
  XNOR2_X1 U7562 ( .A(n11686), .B(n11695), .ZN(n14970) );
  NAND2_X1 U7563 ( .A1(n12717), .A2(n12723), .ZN(n6883) );
  NAND2_X1 U7564 ( .A1(n6882), .A2(n6881), .ZN(n12751) );
  INV_X1 U7565 ( .A(n12721), .ZN(n6881) );
  NAND2_X1 U7566 ( .A1(n12751), .A2(n12750), .ZN(n6880) );
  AOI21_X1 U7567 ( .B1(n9624), .B2(n7087), .A(n6493), .ZN(n7086) );
  INV_X1 U7568 ( .A(n7072), .ZN(n7071) );
  OAI21_X1 U7569 ( .B1(n12618), .B2(n7073), .A(n7966), .ZN(n7072) );
  NAND2_X1 U7570 ( .A1(n7965), .A2(n7076), .ZN(n7073) );
  AND4_X1 U7571 ( .A1(n7666), .A2(n7665), .A3(n7664), .A4(n7663), .ZN(n11390)
         );
  INV_X1 U7572 ( .A(n7946), .ZN(n7062) );
  AND2_X1 U7573 ( .A1(n8009), .A2(n12682), .ZN(n12954) );
  NAND2_X1 U7574 ( .A1(n7980), .A2(n9014), .ZN(n7840) );
  NAND2_X1 U7575 ( .A1(n12676), .A2(n12668), .ZN(n12515) );
  INV_X1 U7576 ( .A(n12663), .ZN(n12833) );
  AND4_X1 U7577 ( .A1(n7929), .A2(n7928), .A3(n7927), .A4(n7926), .ZN(n12857)
         );
  NOR2_X1 U7578 ( .A1(n6548), .A2(n7059), .ZN(n7058) );
  NAND2_X1 U7579 ( .A1(n8936), .A2(n6458), .ZN(n12956) );
  NAND2_X1 U7580 ( .A1(n7818), .A2(n12628), .ZN(n12922) );
  NOR2_X1 U7581 ( .A1(n7817), .A2(n7382), .ZN(n7381) );
  INV_X1 U7582 ( .A(n12616), .ZN(n7382) );
  OR2_X1 U7583 ( .A1(n13032), .A2(n12941), .ZN(n12616) );
  NAND2_X1 U7584 ( .A1(n12965), .A2(n12618), .ZN(n7782) );
  INV_X1 U7585 ( .A(n12487), .ZN(n9629) );
  CLKBUF_X1 U7586 ( .A(n7840), .Z(n6646) );
  NAND2_X1 U7587 ( .A1(n12528), .A2(n10849), .ZN(n15026) );
  NOR2_X1 U7588 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n7306) );
  AND2_X1 U7589 ( .A1(n8003), .A2(n7452), .ZN(n7739) );
  INV_X1 U7590 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7452) );
  NAND2_X1 U7591 ( .A1(n7753), .A2(n7752), .ZN(n7768) );
  INV_X1 U7592 ( .A(n6899), .ZN(n6898) );
  OAI21_X1 U7593 ( .B1(n7651), .B2(n6900), .A(n7670), .ZN(n6899) );
  AND2_X1 U7594 ( .A1(n9320), .A2(n9319), .ZN(n13396) );
  AND2_X1 U7595 ( .A1(n13374), .A2(n12290), .ZN(n13417) );
  NAND2_X1 U7596 ( .A1(n13433), .A2(n13447), .ZN(n13432) );
  INV_X1 U7597 ( .A(n13632), .ZN(n13544) );
  INV_X1 U7598 ( .A(n7049), .ZN(n7048) );
  OAI21_X1 U7599 ( .B1(n13351), .B2(n7050), .A(n13354), .ZN(n7049) );
  NAND2_X1 U7600 ( .A1(n8953), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9299) );
  AND2_X1 U7601 ( .A1(n9861), .A2(n9501), .ZN(n13542) );
  AOI21_X1 U7602 ( .B1(n7270), .B2(n11563), .A(n6518), .ZN(n7269) );
  OAI21_X1 U7603 ( .B1(n11504), .B2(n11503), .A(n11505), .ZN(n11546) );
  XNOR2_X1 U7604 ( .A(n12115), .B(n12116), .ZN(n12305) );
  AND2_X1 U7605 ( .A1(n12329), .A2(n6756), .ZN(n10523) );
  NAND2_X1 U7606 ( .A1(n9033), .A2(n9014), .ZN(n9244) );
  AND2_X1 U7607 ( .A1(n7240), .A2(n9018), .ZN(n7239) );
  AND2_X1 U7608 ( .A1(n8966), .A2(n6809), .ZN(n7240) );
  XNOR2_X1 U7609 ( .A(n8992), .B(P2_IR_REG_21__SCAN_IN), .ZN(n12283) );
  NAND2_X1 U7610 ( .A1(n8991), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8992) );
  INV_X1 U7611 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9006) );
  AND2_X1 U7612 ( .A1(n9769), .A2(n7188), .ZN(n7187) );
  NAND2_X1 U7613 ( .A1(n7189), .A2(n9767), .ZN(n7188) );
  INV_X1 U7614 ( .A(n13959), .ZN(n7189) );
  NAND2_X1 U7615 ( .A1(n9758), .A2(n9757), .ZN(n13957) );
  XNOR2_X1 U7616 ( .A(n9687), .B(n13921), .ZN(n9690) );
  NAND2_X1 U7617 ( .A1(n14002), .A2(n14003), .ZN(n14001) );
  NOR4_X1 U7618 ( .A1(n8786), .A2(n11976), .A3(n12002), .A4(n8785), .ZN(n8788)
         );
  OAI21_X1 U7619 ( .B1(n6981), .B2(n6495), .A(n6980), .ZN(n6977) );
  INV_X1 U7620 ( .A(n14231), .ZN(n6981) );
  NAND2_X1 U7621 ( .A1(n14245), .A2(n12001), .ZN(n14230) );
  NOR2_X1 U7622 ( .A1(n14231), .A2(n6785), .ZN(n6784) );
  INV_X1 U7623 ( .A(n12001), .ZN(n6785) );
  NAND2_X1 U7624 ( .A1(n8603), .A2(n8602), .ZN(n14280) );
  AOI21_X1 U7625 ( .B1(n7103), .B2(n7106), .A(n6542), .ZN(n7100) );
  AOI21_X1 U7626 ( .B1(n6970), .B2(n11152), .A(n6546), .ZN(n6968) );
  INV_X1 U7627 ( .A(n6970), .ZN(n6969) );
  XNOR2_X1 U7628 ( .A(n11488), .B(n11656), .ZN(n11477) );
  NAND2_X1 U7629 ( .A1(n11153), .A2(n11137), .ZN(n11342) );
  AOI21_X1 U7630 ( .B1(n11164), .B2(n6783), .A(n6547), .ZN(n6782) );
  INV_X1 U7631 ( .A(n11135), .ZN(n6783) );
  INV_X1 U7632 ( .A(n8821), .ZN(n7207) );
  AND2_X1 U7633 ( .A1(n6476), .A2(n8065), .ZN(n7206) );
  XNOR2_X1 U7634 ( .A(n8537), .B(n8536), .ZN(n11235) );
  OAI21_X1 U7635 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n9537), .A(n9536), .ZN(
        n9543) );
  AOI21_X1 U7636 ( .B1(n7303), .B2(n7302), .A(n6741), .ZN(n12395) );
  AOI21_X1 U7637 ( .B1(n12425), .B2(n12892), .A(n8893), .ZN(n7302) );
  INV_X1 U7638 ( .A(n7301), .ZN(n6741) );
  INV_X1 U7639 ( .A(n12812), .ZN(n6946) );
  NOR2_X1 U7640 ( .A1(n12844), .A2(n6486), .ZN(n8046) );
  NAND2_X1 U7641 ( .A1(n9478), .A2(n9477), .ZN(n9866) );
  INV_X1 U7642 ( .A(n14225), .ZN(n14418) );
  AND4_X1 U7643 ( .A1(n8693), .A2(n8692), .A3(n8691), .A4(n8690), .ZN(n14401)
         );
  OAI21_X1 U7644 ( .B1(n6463), .B2(n7157), .A(n7154), .ZN(n7159) );
  NAND2_X1 U7645 ( .A1(n12101), .A2(n12100), .ZN(n7425) );
  NAND2_X1 U7646 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  NOR2_X1 U7647 ( .A1(n8314), .A2(n8315), .ZN(n7008) );
  AND2_X1 U7648 ( .A1(n8335), .A2(n6574), .ZN(n6665) );
  MUX2_X1 U7649 ( .A(n12539), .B(n12538), .S(n12656), .Z(n12540) );
  MUX2_X1 U7650 ( .A(n12527), .B(n12526), .S(n6458), .Z(n12543) );
  NAND2_X1 U7651 ( .A1(n6664), .A2(n6663), .ZN(n8376) );
  NAND2_X1 U7652 ( .A1(n8353), .A2(n8355), .ZN(n6663) );
  NAND2_X1 U7653 ( .A1(n8334), .A2(n6665), .ZN(n6664) );
  NAND2_X1 U7654 ( .A1(n6491), .A2(n7006), .ZN(n8334) );
  NAND2_X1 U7655 ( .A1(n7033), .A2(n7032), .ZN(n7030) );
  OAI21_X1 U7656 ( .B1(n7441), .B2(n7440), .A(n7442), .ZN(n12144) );
  NAND2_X1 U7657 ( .A1(n12140), .A2(n7443), .ZN(n7442) );
  INV_X1 U7658 ( .A(n7030), .ZN(n7028) );
  NAND2_X1 U7659 ( .A1(n7031), .A2(n7030), .ZN(n7029) );
  NOR2_X1 U7660 ( .A1(n7033), .A2(n7032), .ZN(n7031) );
  AOI21_X1 U7661 ( .B1(n7023), .B2(n7025), .A(n6556), .ZN(n7022) );
  INV_X1 U7662 ( .A(n12165), .ZN(n7439) );
  OAI21_X1 U7663 ( .B1(n12598), .B2(n12597), .A(n12596), .ZN(n12604) );
  NOR2_X1 U7664 ( .A1(n8550), .A2(n8551), .ZN(n7001) );
  AOI21_X1 U7665 ( .B1(n8550), .B2(n8551), .A(n7003), .ZN(n7002) );
  INV_X1 U7666 ( .A(n8534), .ZN(n7003) );
  NAND2_X1 U7667 ( .A1(n12180), .A2(n7418), .ZN(n7417) );
  INV_X1 U7668 ( .A(n7420), .ZN(n7418) );
  NAND2_X1 U7669 ( .A1(n6489), .A2(n7423), .ZN(n7414) );
  INV_X1 U7670 ( .A(n7423), .ZN(n7419) );
  AOI21_X1 U7671 ( .B1(n6465), .B2(n6997), .A(n6996), .ZN(n6995) );
  NAND2_X1 U7672 ( .A1(n6675), .A2(n6527), .ZN(n12638) );
  INV_X1 U7673 ( .A(n12900), .ZN(n6748) );
  NAND2_X1 U7674 ( .A1(n12189), .A2(n12190), .ZN(n7394) );
  INV_X1 U7675 ( .A(n12189), .ZN(n7392) );
  AND2_X1 U7676 ( .A1(n7408), .A2(n12200), .ZN(n7407) );
  NAND2_X1 U7677 ( .A1(n7411), .A2(n7410), .ZN(n7408) );
  INV_X1 U7678 ( .A(n8683), .ZN(n8686) );
  INV_X1 U7679 ( .A(n13138), .ZN(n7479) );
  AOI21_X1 U7680 ( .B1(n12199), .B2(n7400), .A(n7397), .ZN(n12204) );
  NAND2_X1 U7681 ( .A1(n7399), .A2(n7398), .ZN(n7397) );
  AND2_X1 U7682 ( .A1(n7017), .A2(n8705), .ZN(n7016) );
  NAND2_X1 U7683 ( .A1(n8686), .A2(n8685), .ZN(n7221) );
  AND2_X1 U7684 ( .A1(n7017), .A2(n8706), .ZN(n7013) );
  NAND2_X1 U7685 ( .A1(n7018), .A2(n8717), .ZN(n7017) );
  OR2_X1 U7686 ( .A1(n8620), .A2(n15168), .ZN(n8638) );
  INV_X1 U7687 ( .A(n8451), .ZN(n6831) );
  AOI21_X1 U7688 ( .B1(n6832), .B2(n6829), .A(n6560), .ZN(n6828) );
  NOR2_X1 U7689 ( .A1(n6836), .A2(n8451), .ZN(n6829) );
  NOR2_X1 U7690 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n8049) );
  INV_X1 U7691 ( .A(n7246), .ZN(n7245) );
  OAI21_X1 U7692 ( .B1(n8306), .B2(n7247), .A(n8342), .ZN(n7246) );
  INV_X1 U7693 ( .A(n8323), .ZN(n7247) );
  INV_X1 U7694 ( .A(n6672), .ZN(n9516) );
  OAI21_X1 U7695 ( .B1(n9564), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6555), .ZN(
        n6672) );
  INV_X1 U7696 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9517) );
  INV_X1 U7697 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U7698 ( .A1(n12358), .A2(n8864), .ZN(n8865) );
  OR2_X1 U7699 ( .A1(n12666), .A2(n6458), .ZN(n6677) );
  NAND2_X1 U7700 ( .A1(n12666), .A2(n6679), .ZN(n6678) );
  INV_X1 U7701 ( .A(n12667), .ZN(n6679) );
  NAND2_X1 U7702 ( .A1(n10242), .A2(n10241), .ZN(n10244) );
  NAND2_X1 U7703 ( .A1(n10542), .A2(n10541), .ZN(n10544) );
  NAND2_X1 U7704 ( .A1(n6878), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6877) );
  AND2_X1 U7705 ( .A1(n10544), .A2(n14932), .ZN(n10545) );
  AND2_X1 U7706 ( .A1(n7453), .A2(n7454), .ZN(n7317) );
  INV_X1 U7707 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7454) );
  INV_X1 U7708 ( .A(n7978), .ZN(n7085) );
  INV_X1 U7709 ( .A(n9624), .ZN(n7088) );
  NOR2_X1 U7710 ( .A1(n7795), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7809) );
  NOR2_X1 U7711 ( .A1(n12618), .A2(n7075), .ZN(n7074) );
  INV_X1 U7712 ( .A(n7076), .ZN(n7075) );
  INV_X1 U7713 ( .A(n7365), .ZN(n7364) );
  OAI21_X1 U7714 ( .B1(n12502), .B2(n7366), .A(n12567), .ZN(n7365) );
  INV_X1 U7715 ( .A(n12564), .ZN(n7366) );
  OAI211_X1 U7716 ( .C1(n7980), .C2(n10145), .A(n7509), .B(n7508), .ZN(n8834)
         );
  NAND2_X1 U7717 ( .A1(n7980), .A2(n7065), .ZN(n7508) );
  OR2_X1 U7718 ( .A1(n7515), .A2(n6719), .ZN(n7509) );
  AND2_X1 U7719 ( .A1(n9014), .A2(n7066), .ZN(n7065) );
  OAI21_X1 U7720 ( .B1(n7080), .B2(n7079), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7490) );
  OR2_X1 U7721 ( .A1(n13060), .A2(n8900), .ZN(n12657) );
  NAND2_X1 U7722 ( .A1(n12925), .A2(n12632), .ZN(n7380) );
  OR2_X1 U7723 ( .A1(n13021), .A2(n12902), .ZN(n12635) );
  OR2_X1 U7724 ( .A1(n13098), .A2(n12926), .ZN(n12628) );
  NOR2_X2 U7725 ( .A1(n6740), .A2(n7080), .ZN(n7999) );
  NOR2_X1 U7726 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7450) );
  INV_X1 U7727 ( .A(n7837), .ZN(n6917) );
  NAND2_X1 U7728 ( .A1(n7820), .A2(n7819), .ZN(n7821) );
  AND2_X1 U7729 ( .A1(n8003), .A2(n7461), .ZN(n7464) );
  INV_X1 U7730 ( .A(n7470), .ZN(n7461) );
  INV_X1 U7732 ( .A(n7767), .ZN(n6911) );
  AND2_X1 U7733 ( .A1(n7739), .A2(n7453), .ZN(n7755) );
  NAND2_X1 U7734 ( .A1(n7699), .A2(n7698), .ZN(n7715) );
  AND3_X2 U7735 ( .A1(n7522), .A2(n6709), .A3(n6708), .ZN(n7307) );
  INV_X1 U7736 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n6709) );
  INV_X1 U7737 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n6708) );
  INV_X1 U7738 ( .A(n6485), .ZN(n6813) );
  NOR2_X1 U7739 ( .A1(n11180), .A2(n6815), .ZN(n6812) );
  NAND2_X1 U7740 ( .A1(n12216), .A2(n6469), .ZN(n7388) );
  INV_X1 U7741 ( .A(n12271), .ZN(n12272) );
  NAND2_X1 U7742 ( .A1(n7389), .A2(n12324), .ZN(n7385) );
  XNOR2_X1 U7743 ( .A(n13295), .B(n12073), .ZN(n12296) );
  NAND2_X1 U7744 ( .A1(n7045), .A2(n6484), .ZN(n7044) );
  INV_X1 U7745 ( .A(n6743), .ZN(n7045) );
  AND2_X1 U7746 ( .A1(n9185), .A2(n9184), .ZN(n9189) );
  NOR2_X1 U7747 ( .A1(n9167), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U7748 ( .A1(n9692), .A2(n9691), .ZN(n7182) );
  INV_X1 U7749 ( .A(n9717), .ZN(n7192) );
  INV_X1 U7750 ( .A(n7199), .ZN(n7193) );
  OR2_X1 U7751 ( .A1(n8730), .A2(n10040), .ZN(n8096) );
  AOI21_X1 U7752 ( .B1(n7105), .B2(n7104), .A(n14333), .ZN(n7103) );
  INV_X1 U7753 ( .A(n7108), .ZN(n7104) );
  INV_X1 U7754 ( .A(n11964), .ZN(n6967) );
  INV_X1 U7755 ( .A(n11967), .ZN(n6966) );
  NOR2_X1 U7756 ( .A1(n14663), .A2(n6852), .ZN(n6851) );
  INV_X1 U7757 ( .A(n6853), .ZN(n6852) );
  AND2_X1 U7758 ( .A1(n11788), .A2(n11786), .ZN(n6795) );
  INV_X1 U7759 ( .A(n6959), .ZN(n6958) );
  OAI21_X1 U7760 ( .B1(n11345), .B2(n6960), .A(n11667), .ZN(n6959) );
  INV_X1 U7761 ( .A(n11575), .ZN(n6960) );
  NAND2_X1 U7762 ( .A1(n6845), .A2(n10269), .ZN(n8501) );
  NOR2_X1 U7763 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7012) );
  NAND2_X1 U7764 ( .A1(n6702), .A2(n8458), .ZN(n8497) );
  OAI21_X1 U7765 ( .B1(n8369), .B2(n6835), .A(n6832), .ZN(n8452) );
  OR2_X1 U7766 ( .A1(n8452), .A2(n10011), .ZN(n8426) );
  OAI21_X1 U7767 ( .B1(n8369), .B2(n8368), .A(n8367), .ZN(n8392) );
  XNOR2_X1 U7768 ( .A(n9515), .B(n15098), .ZN(n9564) );
  XNOR2_X1 U7769 ( .A(n9516), .B(n9517), .ZN(n9554) );
  NOR2_X1 U7770 ( .A1(n9527), .A2(n9526), .ZN(n9553) );
  NOR2_X1 U7771 ( .A1(n9578), .A2(n15108), .ZN(n9526) );
  AND2_X1 U7772 ( .A1(n14685), .A2(n7154), .ZN(n7151) );
  INV_X1 U7773 ( .A(n7155), .ZN(n7149) );
  AOI21_X1 U7774 ( .B1(n7151), .B2(n7157), .A(P2_ADDR_REG_14__SCAN_IN), .ZN(
        n7150) );
  INV_X1 U7775 ( .A(n7152), .ZN(n7146) );
  INV_X1 U7776 ( .A(n8870), .ZN(n7285) );
  NAND2_X1 U7777 ( .A1(n11749), .A2(n7284), .ZN(n7283) );
  NAND2_X1 U7778 ( .A1(n11051), .A2(n8857), .ZN(n12379) );
  AOI21_X1 U7779 ( .B1(n8896), .B2(n8895), .A(n8894), .ZN(n7301) );
  NAND2_X1 U7780 ( .A1(n11905), .A2(n12980), .ZN(n7293) );
  INV_X1 U7781 ( .A(n7293), .ZN(n7292) );
  INV_X1 U7782 ( .A(n7291), .ZN(n7290) );
  OAI21_X1 U7783 ( .B1(n7294), .B2(n7292), .A(n12403), .ZN(n7291) );
  NOR2_X1 U7784 ( .A1(n11720), .A2(n11818), .ZN(n7284) );
  NAND2_X1 U7785 ( .A1(n12387), .A2(n8889), .ZN(n8892) );
  NAND3_X1 U7786 ( .A1(n8838), .A2(n10400), .A3(n14990), .ZN(n10399) );
  AND4_X1 U7787 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n12941)
         );
  NAND2_X1 U7788 ( .A1(n6731), .A2(n6944), .ZN(n6938) );
  AND2_X1 U7789 ( .A1(n6613), .A2(n6612), .ZN(n6939) );
  OR2_X1 U7790 ( .A1(n6941), .A2(n10178), .ZN(n6612) );
  NAND2_X1 U7791 ( .A1(n6942), .A2(n6561), .ZN(n6613) );
  NAND2_X1 U7792 ( .A1(n6713), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10287) );
  INV_X1 U7793 ( .A(n6877), .ZN(n6876) );
  OR2_X1 U7794 ( .A1(n14927), .A2(n10545), .ZN(n10546) );
  NAND2_X1 U7795 ( .A1(n10546), .A2(n10547), .ZN(n10910) );
  AND2_X1 U7796 ( .A1(n14950), .A2(n11334), .ZN(n11402) );
  INV_X1 U7797 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11754) );
  NAND2_X1 U7798 ( .A1(n11694), .A2(n11693), .ZN(n6670) );
  NAND2_X1 U7799 ( .A1(n6611), .A2(n6610), .ZN(n11694) );
  INV_X1 U7800 ( .A(n11691), .ZN(n6610) );
  AND2_X1 U7801 ( .A1(n11685), .A2(n11684), .ZN(n11686) );
  AND2_X1 U7802 ( .A1(n6754), .A2(n6753), .ZN(n14565) );
  XNOR2_X1 U7803 ( .A(n6883), .B(n14559), .ZN(n14562) );
  AND2_X1 U7804 ( .A1(n14565), .A2(n14564), .ZN(n14567) );
  OR2_X1 U7805 ( .A1(n14556), .A2(n12739), .ZN(n6934) );
  NAND2_X1 U7806 ( .A1(n6934), .A2(n6933), .ZN(n12754) );
  INV_X1 U7807 ( .A(n12742), .ZN(n6933) );
  NAND2_X1 U7808 ( .A1(n7739), .A2(n7317), .ZN(n7770) );
  AND2_X1 U7809 ( .A1(n7090), .A2(n6510), .ZN(n7979) );
  OR2_X1 U7810 ( .A1(n7866), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U7811 ( .A1(n7827), .A2(n12436), .ZN(n7843) );
  INV_X1 U7812 ( .A(n7828), .ZN(n7827) );
  AND2_X1 U7813 ( .A1(n7071), .A2(n12626), .ZN(n7069) );
  NAND2_X1 U7814 ( .A1(n6766), .A2(n7074), .ZN(n7070) );
  OR2_X1 U7815 ( .A1(n7676), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7693) );
  AND2_X1 U7816 ( .A1(n7659), .A2(n7658), .ZN(n11498) );
  INV_X1 U7817 ( .A(n7093), .ZN(n7092) );
  AOI21_X1 U7818 ( .B1(n7093), .B2(n12567), .A(n6504), .ZN(n7091) );
  NAND2_X1 U7819 ( .A1(n11464), .A2(n7952), .ZN(n11389) );
  NOR2_X1 U7820 ( .A1(n12572), .A2(n7094), .ZN(n7093) );
  INV_X1 U7821 ( .A(n7952), .ZN(n7094) );
  CLKBUF_X1 U7822 ( .A(n11466), .Z(n6711) );
  NAND2_X1 U7823 ( .A1(n6711), .A2(n11465), .ZN(n11464) );
  NAND2_X1 U7824 ( .A1(n10998), .A2(n12560), .ZN(n11029) );
  NAND2_X1 U7825 ( .A1(n11029), .A2(n12502), .ZN(n11031) );
  AND4_X1 U7826 ( .A1(n7613), .A2(n7612), .A3(n7611), .A4(n7610), .ZN(n11391)
         );
  AND4_X1 U7827 ( .A1(n7595), .A2(n7594), .A3(n7593), .A4(n7592), .ZN(n11001)
         );
  AND4_X1 U7828 ( .A1(n7582), .A2(n7581), .A3(n7580), .A4(n7579), .ZN(n11025)
         );
  NOR2_X1 U7829 ( .A1(n7372), .A2(n7369), .ZN(n7368) );
  NAND2_X1 U7830 ( .A1(n12549), .A2(n12550), .ZN(n10627) );
  INV_X1 U7831 ( .A(n10627), .ZN(n12547) );
  NAND2_X1 U7832 ( .A1(n10625), .A2(n12547), .ZN(n10624) );
  INV_X1 U7833 ( .A(n12868), .ZN(n6764) );
  XNOR2_X1 U7834 ( .A(n13008), .B(n12881), .ZN(n12868) );
  AND2_X1 U7835 ( .A1(n12635), .A2(n12636), .ZN(n12915) );
  NAND2_X1 U7836 ( .A1(n7782), .A2(n6526), .ZN(n12950) );
  NAND2_X1 U7837 ( .A1(n12987), .A2(n12988), .ZN(n7342) );
  AND2_X1 U7838 ( .A1(n7344), .A2(n12979), .ZN(n7343) );
  NAND2_X1 U7839 ( .A1(n7345), .A2(n12610), .ZN(n7344) );
  INV_X1 U7840 ( .A(n12988), .ZN(n7345) );
  INV_X1 U7841 ( .A(n12610), .ZN(n7346) );
  AND2_X1 U7842 ( .A1(n12606), .A2(n12610), .ZN(n12988) );
  AND3_X1 U7843 ( .A1(n7607), .A2(n7606), .A3(n7605), .ZN(n15014) );
  NAND2_X1 U7844 ( .A1(n8937), .A2(n6458), .ZN(n12958) );
  OR2_X1 U7845 ( .A1(n12031), .A2(n12030), .ZN(n12034) );
  NAND2_X1 U7846 ( .A1(n7905), .A2(n7904), .ZN(n7917) );
  NAND2_X1 U7847 ( .A1(n7903), .A2(n7902), .ZN(n7905) );
  OAI21_X1 U7848 ( .B1(n7890), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7891), .ZN(
        n7903) );
  OAI21_X1 U7849 ( .B1(n7838), .B2(n6918), .A(n6916), .ZN(n7874) );
  INV_X1 U7850 ( .A(n6919), .ZN(n6918) );
  AOI21_X1 U7851 ( .B1(n6917), .B2(n6919), .A(n6603), .ZN(n6916) );
  NOR2_X1 U7852 ( .A1(n7862), .A2(n6920), .ZN(n6919) );
  NAND2_X1 U7853 ( .A1(n7835), .A2(n7834), .ZN(n7838) );
  NAND2_X1 U7854 ( .A1(n7838), .A2(n7837), .ZN(n7850) );
  NAND2_X1 U7855 ( .A1(n7802), .A2(n7801), .ZN(n7805) );
  NAND2_X1 U7856 ( .A1(n7805), .A2(n7804), .ZN(n7820) );
  AND2_X1 U7857 ( .A1(n7767), .A2(n7751), .ZN(n7752) );
  NAND2_X1 U7858 ( .A1(n7750), .A2(n7749), .ZN(n7753) );
  XNOR2_X1 U7859 ( .A(n7715), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U7860 ( .A1(n7700), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7717) );
  AND2_X1 U7861 ( .A1(n7682), .A2(n7669), .ZN(n7670) );
  INV_X1 U7862 ( .A(n7667), .ZN(n6900) );
  AND2_X1 U7863 ( .A1(n7667), .A2(n7650), .ZN(n7651) );
  NAND2_X1 U7864 ( .A1(n7652), .A2(n7651), .ZN(n7668) );
  NAND2_X1 U7865 ( .A1(n7637), .A2(n7636), .ZN(n7640) );
  NAND2_X1 U7866 ( .A1(n7640), .A2(n7639), .ZN(n7649) );
  OAI21_X1 U7867 ( .B1(n7621), .B2(n7620), .A(n7622), .ZN(n7625) );
  NAND2_X1 U7868 ( .A1(n7625), .A2(n7624), .ZN(n7637) );
  NOR2_X1 U7869 ( .A1(n7615), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7655) );
  NAND2_X1 U7870 ( .A1(n7538), .A2(n7537), .ZN(n7549) );
  INV_X1 U7871 ( .A(n9117), .ZN(n7330) );
  INV_X1 U7872 ( .A(n9097), .ZN(n7333) );
  NAND2_X1 U7873 ( .A1(n13273), .A2(n13271), .ZN(n6799) );
  NAND2_X1 U7874 ( .A1(n6799), .A2(n6798), .ZN(n13192) );
  NOR2_X1 U7875 ( .A1(n9279), .A2(n6797), .ZN(n6798) );
  INV_X1 U7876 ( .A(n13194), .ZN(n6797) );
  NAND2_X1 U7877 ( .A1(n6820), .A2(n6819), .ZN(n9093) );
  AOI21_X1 U7878 ( .B1(n9080), .B2(n10375), .A(n6552), .ZN(n6819) );
  INV_X1 U7879 ( .A(n13294), .ZN(n12088) );
  NAND2_X1 U7880 ( .A1(n13177), .A2(n9367), .ZN(n9382) );
  NAND2_X1 U7881 ( .A1(n8950), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9195) );
  INV_X1 U7882 ( .A(n9172), .ZN(n8950) );
  OR2_X1 U7883 ( .A1(n9299), .A2(n11828), .ZN(n9314) );
  NAND2_X1 U7884 ( .A1(n9410), .A2(n13214), .ZN(n7323) );
  AOI21_X1 U7885 ( .B1(n7326), .B2(n11434), .A(n6817), .ZN(n6816) );
  INV_X1 U7886 ( .A(n9262), .ZN(n6817) );
  NAND2_X1 U7887 ( .A1(n12283), .A2(n10089), .ZN(n12286) );
  INV_X1 U7888 ( .A(n6756), .ZN(n12343) );
  AND2_X1 U7889 ( .A1(n9379), .A2(n9378), .ZN(n13233) );
  NAND2_X1 U7890 ( .A1(n9937), .A2(n9938), .ZN(n9936) );
  NOR2_X1 U7891 ( .A1(n11528), .A2(n11529), .ZN(n11594) );
  NOR2_X1 U7892 ( .A1(n9489), .A2(n13169), .ZN(n13383) );
  AND2_X1 U7893 ( .A1(n9489), .A2(n9436), .ZN(n9502) );
  NAND2_X1 U7894 ( .A1(n13494), .A2(n6519), .ZN(n13477) );
  NAND2_X1 U7895 ( .A1(n6445), .A2(n6631), .ZN(n13494) );
  OAI21_X1 U7896 ( .B1(n13541), .B2(n7054), .A(n7051), .ZN(n13515) );
  NAND2_X1 U7897 ( .A1(n13368), .A2(n7055), .ZN(n7054) );
  INV_X1 U7898 ( .A(n7052), .ZN(n7051) );
  INV_X1 U7899 ( .A(n13366), .ZN(n7055) );
  AND2_X1 U7900 ( .A1(n9385), .A2(n9384), .ZN(n13512) );
  NAND2_X1 U7901 ( .A1(n13703), .A2(n7214), .ZN(n13504) );
  INV_X1 U7902 ( .A(n13405), .ZN(n7215) );
  OAI21_X1 U7903 ( .B1(n13605), .B2(n7265), .A(n7262), .ZN(n13580) );
  AOI21_X1 U7904 ( .B1(n7264), .B2(n7263), .A(n6530), .ZN(n7262) );
  INV_X1 U7905 ( .A(n13394), .ZN(n7263) );
  NOR2_X1 U7906 ( .A1(n13638), .A2(n13775), .ZN(n6699) );
  NOR2_X2 U7907 ( .A1(n13621), .A2(n13730), .ZN(n13600) );
  AND3_X1 U7908 ( .A1(n9288), .A2(n9287), .A3(n9286), .ZN(n13633) );
  XNOR2_X1 U7909 ( .A(n13644), .B(n13350), .ZN(n13645) );
  NAND2_X1 U7910 ( .A1(n13629), .A2(n13645), .ZN(n13628) );
  OR2_X1 U7911 ( .A1(n12157), .A2(n13284), .ZN(n7273) );
  AND2_X1 U7912 ( .A1(n12315), .A2(n11557), .ZN(n7056) );
  AND4_X1 U7913 ( .A1(n9200), .A2(n9199), .A3(n9198), .A4(n9197), .ZN(n12141)
         );
  AOI21_X1 U7914 ( .B1(n7043), .B2(n7042), .A(n6545), .ZN(n7041) );
  INV_X1 U7915 ( .A(n6484), .ZN(n7042) );
  NAND2_X1 U7916 ( .A1(n8948), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9156) );
  INV_X1 U7917 ( .A(n10779), .ZN(n7228) );
  NAND2_X1 U7918 ( .A1(n10761), .A2(n10760), .ZN(n10762) );
  NAND2_X1 U7919 ( .A1(n10762), .A2(n10766), .ZN(n10780) );
  OR2_X1 U7920 ( .A1(n12218), .A2(n10000), .ZN(n9111) );
  INV_X1 U7921 ( .A(n12300), .ZN(n10750) );
  NAND2_X1 U7922 ( .A1(n10421), .A2(n10429), .ZN(n10745) );
  NAND2_X1 U7923 ( .A1(n10116), .A2(n10115), .ZN(n10423) );
  OR2_X1 U7924 ( .A1(n12297), .A2(n10091), .ZN(n10111) );
  INV_X1 U7925 ( .A(n13673), .ZN(n6847) );
  NAND2_X1 U7926 ( .A1(n13674), .A2(n14889), .ZN(n6846) );
  NAND2_X1 U7927 ( .A1(n9400), .A2(n9399), .ZN(n13692) );
  INV_X1 U7928 ( .A(n13552), .ZN(n13710) );
  NAND2_X1 U7929 ( .A1(n9330), .A2(n9329), .ZN(n13715) );
  OR2_X1 U7930 ( .A1(n11538), .A2(n9038), .ZN(n9330) );
  INV_X1 U7931 ( .A(n13604), .ZN(n13730) );
  AND2_X1 U7932 ( .A1(n9192), .A2(n9191), .ZN(n14908) );
  NAND2_X1 U7933 ( .A1(n8977), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U7934 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n13784), .ZN(n6806) );
  NAND2_X1 U7935 ( .A1(n6809), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U7936 ( .A1(n9458), .A2(n9457), .ZN(n9467) );
  INV_X1 U7937 ( .A(n9482), .ZN(n9458) );
  XNOR2_X1 U7938 ( .A(n9226), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11122) );
  INV_X1 U7939 ( .A(n8593), .ZN(n8594) );
  NAND2_X1 U7940 ( .A1(n7187), .A2(n7190), .ZN(n7186) );
  AOI21_X1 U7941 ( .B1(n7212), .B2(n7210), .A(n6505), .ZN(n7209) );
  INV_X1 U7942 ( .A(n7212), .ZN(n7211) );
  INV_X1 U7943 ( .A(n9746), .ZN(n7210) );
  NAND2_X1 U7944 ( .A1(n7180), .A2(n7178), .ZN(n7177) );
  AND2_X1 U7945 ( .A1(n7179), .A2(n7181), .ZN(n7178) );
  NAND2_X1 U7946 ( .A1(n7183), .A2(n7174), .ZN(n10962) );
  NOR2_X1 U7947 ( .A1(n7175), .A2(n7181), .ZN(n7174) );
  INV_X1 U7948 ( .A(n7182), .ZN(n7175) );
  OR2_X1 U7949 ( .A1(n8296), .A2(n8295), .ZN(n8317) );
  NOR2_X1 U7950 ( .A1(n11761), .A2(n7168), .ZN(n7167) );
  INV_X1 U7951 ( .A(n7170), .ZN(n7168) );
  INV_X1 U7952 ( .A(n6953), .ZN(n8548) );
  AOI21_X1 U7953 ( .B1(n7113), .B2(n14217), .A(n6554), .ZN(n6626) );
  AND2_X1 U7954 ( .A1(n8704), .A2(n8703), .ZN(n13925) );
  OR2_X1 U7955 ( .A1(n11979), .A2(n11978), .ZN(n11980) );
  NOR2_X1 U7956 ( .A1(n14219), .A2(n14412), .ZN(n12045) );
  INV_X1 U7957 ( .A(n11976), .ZN(n12041) );
  AOI21_X1 U7958 ( .B1(n12050), .B2(n14254), .A(n12044), .ZN(n6692) );
  NAND2_X1 U7959 ( .A1(n14234), .A2(n14418), .ZN(n14219) );
  NAND2_X1 U7960 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  NAND2_X1 U7961 ( .A1(n11998), .A2(n11997), .ZN(n14245) );
  INV_X1 U7962 ( .A(n14253), .ZN(n11997) );
  AND2_X1 U7963 ( .A1(n11974), .A2(n11995), .ZN(n7121) );
  NOR2_X1 U7964 ( .A1(n14304), .A2(n7117), .ZN(n7116) );
  NAND2_X1 U7965 ( .A1(n14288), .A2(n14287), .ZN(n14286) );
  NOR2_X1 U7966 ( .A1(n6490), .A2(n7109), .ZN(n7108) );
  INV_X1 U7967 ( .A(n11988), .ZN(n7109) );
  INV_X1 U7968 ( .A(n7106), .ZN(n7105) );
  OAI21_X1 U7969 ( .B1(n6490), .B2(n7107), .A(n11989), .ZN(n7106) );
  NAND2_X1 U7970 ( .A1(n7110), .A2(n11988), .ZN(n7107) );
  INV_X1 U7971 ( .A(n11987), .ZN(n7110) );
  NAND2_X1 U7972 ( .A1(n11986), .A2(n11985), .ZN(n14367) );
  NAND2_X1 U7973 ( .A1(n11916), .A2(n6500), .ZN(n11918) );
  OR2_X1 U7974 ( .A1(n11918), .A2(n11930), .ZN(n11965) );
  NAND2_X1 U7975 ( .A1(n11787), .A2(n6795), .ZN(n11801) );
  NAND2_X1 U7976 ( .A1(n11675), .A2(n11674), .ZN(n11787) );
  INV_X1 U7977 ( .A(n14033), .ZN(n11872) );
  INV_X1 U7978 ( .A(n7098), .ZN(n7097) );
  OAI21_X1 U7979 ( .B1(n11355), .B2(n7099), .A(n11666), .ZN(n7098) );
  INV_X1 U7980 ( .A(n11580), .ZN(n7099) );
  NAND2_X1 U7981 ( .A1(n11475), .A2(n11354), .ZN(n11356) );
  NAND2_X1 U7982 ( .A1(n11356), .A2(n11355), .ZN(n11581) );
  NAND2_X1 U7983 ( .A1(n11353), .A2(n11352), .ZN(n11476) );
  NAND2_X1 U7984 ( .A1(n11476), .A2(n11477), .ZN(n11475) );
  INV_X1 U7985 ( .A(n11341), .ZN(n6971) );
  NAND2_X1 U7986 ( .A1(n11342), .A2(n11341), .ZN(n11478) );
  NAND2_X1 U7987 ( .A1(n6782), .A2(n11146), .ZN(n6781) );
  INV_X1 U7988 ( .A(n14483), .ZN(n14400) );
  INV_X1 U7989 ( .A(n8138), .ZN(n10797) );
  INV_X1 U7990 ( .A(n14210), .ZN(n14397) );
  NAND2_X1 U7991 ( .A1(n6864), .A2(n6863), .ZN(n6862) );
  INV_X1 U7992 ( .A(n14403), .ZN(n6863) );
  NAND2_X1 U7993 ( .A1(n8641), .A2(n8640), .ZN(n14425) );
  AND2_X1 U7994 ( .A1(n14537), .A2(n8113), .ZN(n14449) );
  NAND2_X1 U7995 ( .A1(n8525), .A2(n8524), .ZN(n14470) );
  INV_X1 U7996 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8067) );
  INV_X1 U7997 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7208) );
  INV_X1 U7998 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U7999 ( .A1(n8586), .A2(n7277), .ZN(n7274) );
  OR2_X1 U8000 ( .A1(n8538), .A2(n10640), .ZN(n8552) );
  NAND2_X1 U8001 ( .A1(n8539), .A2(n7252), .ZN(n7251) );
  INV_X1 U8002 ( .A(n8552), .ZN(n7250) );
  NAND2_X1 U8003 ( .A1(n8501), .A2(n7261), .ZN(n7260) );
  NAND2_X1 U8004 ( .A1(n6842), .A2(SI_18_), .ZN(n8520) );
  XNOR2_X1 U8005 ( .A(n8405), .B(n8404), .ZN(n10408) );
  NAND2_X1 U8006 ( .A1(n7230), .A2(n8394), .ZN(n8405) );
  NAND2_X1 U8007 ( .A1(n8392), .A2(n8391), .ZN(n7230) );
  XNOR2_X1 U8008 ( .A(n8392), .B(n8391), .ZN(n10358) );
  XNOR2_X1 U8009 ( .A(n8343), .B(n8341), .ZN(n10079) );
  NAND2_X1 U8010 ( .A1(n8324), .A2(n8323), .ZN(n8343) );
  AND2_X1 U8011 ( .A1(n8168), .A2(n8167), .ZN(n8194) );
  NOR2_X1 U8012 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  NOR2_X1 U8013 ( .A1(n9522), .A2(n9521), .ZN(n9576) );
  NAND2_X1 U8014 ( .A1(n9581), .A2(n9580), .ZN(n9582) );
  NAND2_X1 U8015 ( .A1(n9589), .A2(n9588), .ZN(n9590) );
  OR2_X1 U8016 ( .A1(n14680), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7154) );
  AND2_X1 U8017 ( .A1(n14680), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7157) );
  AOI22_X1 U8018 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n10664), .B1(n9543), .B2(
        n9538), .ZN(n9600) );
  OR2_X1 U8019 ( .A1(n14687), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7138) );
  NAND2_X1 U8020 ( .A1(n7136), .A2(n14692), .ZN(n7135) );
  OAI21_X1 U8021 ( .B1(n9610), .B2(n9609), .A(n14552), .ZN(n9618) );
  AND2_X1 U8022 ( .A1(n11380), .A2(n8862), .ZN(n12360) );
  AND4_X1 U8023 ( .A1(n7833), .A2(n7832), .A3(n7831), .A4(n7830), .ZN(n12940)
         );
  INV_X1 U8024 ( .A(n12893), .ZN(n12914) );
  INV_X1 U8025 ( .A(n10582), .ZN(n7297) );
  NAND2_X1 U8026 ( .A1(n8928), .A2(n8927), .ZN(n12464) );
  OR2_X1 U8027 ( .A1(n8897), .A2(n12881), .ZN(n7300) );
  NAND2_X1 U8028 ( .A1(n6888), .A2(n12675), .ZN(n6887) );
  OR2_X1 U8029 ( .A1(n6888), .A2(n8036), .ZN(n6749) );
  AOI21_X1 U8030 ( .B1(n7359), .B2(n7357), .A(n12678), .ZN(n12681) );
  AND2_X1 U8031 ( .A1(n12679), .A2(n7358), .ZN(n7357) );
  INV_X1 U8032 ( .A(n10629), .ZN(n10616) );
  OR2_X1 U8033 ( .A1(n14963), .A2(n14964), .ZN(n6689) );
  XNOR2_X1 U8034 ( .A(n6670), .B(n14965), .ZN(n14963) );
  NAND2_X1 U8035 ( .A1(n6885), .A2(n6884), .ZN(n12717) );
  INV_X1 U8036 ( .A(n11701), .ZN(n6884) );
  INV_X1 U8037 ( .A(n6880), .ZN(n12769) );
  NOR2_X1 U8038 ( .A1(n9642), .A2(n15026), .ZN(n12826) );
  NAND2_X1 U8039 ( .A1(n8906), .A2(n8905), .ZN(n13054) );
  NAND2_X1 U8040 ( .A1(n7826), .A2(n7825), .ZN(n12932) );
  NAND2_X1 U8041 ( .A1(n7794), .A2(n7793), .ZN(n13032) );
  INV_X1 U8042 ( .A(n14580), .ZN(n14998) );
  INV_X1 U8043 ( .A(n13047), .ZN(n13001) );
  NAND2_X1 U8044 ( .A1(n7724), .A2(n7723), .ZN(n12602) );
  AND3_X1 U8045 ( .A1(n7558), .A2(n7557), .A3(n7556), .ZN(n10672) );
  NAND2_X1 U8046 ( .A1(n7349), .A2(n7353), .ZN(n12677) );
  NAND2_X1 U8047 ( .A1(n9645), .A2(n6487), .ZN(n7349) );
  AND2_X1 U8048 ( .A1(n7356), .A2(n7354), .ZN(n12830) );
  INV_X1 U8049 ( .A(n12520), .ZN(n7354) );
  NAND2_X1 U8050 ( .A1(n9645), .A2(n9644), .ZN(n7356) );
  NAND2_X1 U8051 ( .A1(n7852), .A2(n7851), .ZN(n13082) );
  NAND2_X1 U8052 ( .A1(n7774), .A2(n7773), .ZN(n13109) );
  NAND2_X1 U8053 ( .A1(n7760), .A2(n7759), .ZN(n13115) );
  XNOR2_X1 U8054 ( .A(n7465), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12690) );
  XNOR2_X1 U8055 ( .A(n7456), .B(n7455), .ZN(n12808) );
  INV_X1 U8056 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7455) );
  NAND2_X1 U8057 ( .A1(n7318), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7456) );
  AND2_X1 U8058 ( .A1(n6822), .A2(n6470), .ZN(n13163) );
  OR2_X1 U8059 ( .A1(n10637), .A2(n9038), .ZN(n9247) );
  AND2_X1 U8060 ( .A1(n13143), .A2(n9396), .ZN(n13150) );
  XNOR2_X1 U8061 ( .A(n9398), .B(n6767), .ZN(n13143) );
  INV_X1 U8062 ( .A(n9397), .ZN(n6767) );
  INV_X1 U8063 ( .A(n13578), .ZN(n13720) );
  NAND2_X1 U8064 ( .A1(n7319), .A2(n7322), .ZN(n13255) );
  NAND2_X1 U8065 ( .A1(n13215), .A2(n9410), .ZN(n7319) );
  AND2_X1 U8066 ( .A1(n9361), .A2(n9360), .ZN(n13403) );
  INV_X1 U8067 ( .A(n13281), .ZN(n13258) );
  NOR2_X1 U8068 ( .A1(n12333), .A2(n12332), .ZN(n12335) );
  OR2_X1 U8069 ( .A1(n7433), .A2(n12338), .ZN(n7430) );
  INV_X1 U8070 ( .A(n13389), .ZN(n13350) );
  AND2_X1 U8071 ( .A1(n9886), .A2(n9885), .ZN(n14865) );
  OAI21_X1 U8072 ( .B1(n13422), .B2(n6849), .A(n13421), .ZN(n13672) );
  AOI21_X1 U8073 ( .B1(n13438), .B2(n13635), .A(n13437), .ZN(n13679) );
  OAI21_X1 U8074 ( .B1(n11747), .B2(n9038), .A(n9372), .ZN(n13702) );
  NAND2_X1 U8075 ( .A1(n9122), .A2(n9121), .ZN(n12115) );
  OR2_X1 U8076 ( .A1(n9900), .A2(n9038), .ZN(n9122) );
  AND2_X2 U8077 ( .A1(n10103), .A2(n10467), .ZN(n14922) );
  NOR2_X1 U8078 ( .A1(n6522), .A2(n6502), .ZN(n6777) );
  NAND2_X1 U8079 ( .A1(n13446), .A2(n6641), .ZN(n6640) );
  INV_X1 U8080 ( .A(n13330), .ZN(n12334) );
  INV_X1 U8081 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11019) );
  AOI21_X1 U8082 ( .B1(n13888), .B2(n13885), .A(n13918), .ZN(n7160) );
  INV_X1 U8083 ( .A(n13888), .ZN(n7161) );
  INV_X1 U8084 ( .A(n14034), .ZN(n11764) );
  OR2_X1 U8085 ( .A1(n8656), .A2(n9844), .ZN(n6854) );
  AND4_X1 U8086 ( .A1(n8466), .A2(n8465), .A3(n8464), .A4(n8463), .ZN(n14350)
         );
  NAND2_X1 U8087 ( .A1(n13961), .A2(n9767), .ZN(n9768) );
  AND2_X1 U8088 ( .A1(n14697), .A2(n14793), .ZN(n14653) );
  NAND2_X1 U8089 ( .A1(n9792), .A2(n9791), .ZN(n14699) );
  AOI21_X1 U8090 ( .B1(n8803), .B2(n8802), .A(n8801), .ZN(n8812) );
  OR3_X1 U8091 ( .A1(n8810), .A2(n8786), .A3(n8793), .ZN(n8813) );
  INV_X1 U8092 ( .A(n13964), .ZN(n14484) );
  AND4_X1 U8093 ( .A1(n8287), .A2(n8286), .A3(n8285), .A4(n8284), .ZN(n11627)
         );
  AND2_X1 U8094 ( .A1(n10864), .A2(n10863), .ZN(n11204) );
  INV_X1 U8095 ( .A(n14197), .ZN(n6655) );
  OAI21_X1 U8096 ( .B1(n14526), .B2(n8656), .A(n8655), .ZN(n14225) );
  OR2_X1 U8097 ( .A1(n11021), .A2(n8656), .ZN(n8508) );
  NAND2_X1 U8098 ( .A1(n12012), .A2(n12011), .ZN(n12014) );
  XNOR2_X1 U8099 ( .A(n8143), .B(n8144), .ZN(n11239) );
  INV_X1 U8100 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11020) );
  NAND2_X1 U8101 ( .A1(n7158), .A2(n7153), .ZN(n7152) );
  INV_X1 U8102 ( .A(n7154), .ZN(n7153) );
  NAND2_X1 U8103 ( .A1(n7156), .A2(n7158), .ZN(n7155) );
  INV_X1 U8104 ( .A(n7157), .ZN(n7156) );
  OR2_X1 U8105 ( .A1(n14678), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6671) );
  NOR2_X1 U8106 ( .A1(n9603), .A2(n9604), .ZN(n14687) );
  AND2_X1 U8107 ( .A1(n9603), .A2(n9604), .ZN(n14688) );
  INV_X1 U8108 ( .A(n14690), .ZN(n7136) );
  NAND2_X1 U8109 ( .A1(n7138), .A2(n7139), .ZN(n7137) );
  XNOR2_X1 U8110 ( .A(n9618), .B(n9617), .ZN(n14540) );
  NAND2_X1 U8111 ( .A1(n6667), .A2(n6666), .ZN(n8242) );
  NAND2_X1 U8112 ( .A1(n8217), .A2(n8219), .ZN(n6666) );
  NAND2_X1 U8113 ( .A1(n12106), .A2(n12107), .ZN(n7427) );
  OAI21_X1 U8114 ( .B1(n8269), .B2(n8268), .A(n8267), .ZN(n8291) );
  NOR2_X1 U8115 ( .A1(n7008), .A2(n7006), .ZN(n7005) );
  INV_X1 U8116 ( .A(n7008), .ZN(n7004) );
  INV_X1 U8117 ( .A(n12138), .ZN(n7443) );
  INV_X1 U8118 ( .A(n8402), .ZN(n7032) );
  OAI21_X1 U8119 ( .B1(n12543), .B2(n12542), .A(n12541), .ZN(n12548) );
  NAND2_X1 U8120 ( .A1(n12551), .A2(n12552), .ZN(n6744) );
  NAND2_X1 U8121 ( .A1(n8379), .A2(n8378), .ZN(n8380) );
  NAND2_X1 U8122 ( .A1(n8444), .A2(n7019), .ZN(n7024) );
  INV_X1 U8123 ( .A(n7026), .ZN(n7025) );
  NAND2_X1 U8124 ( .A1(n8519), .A2(n6490), .ZN(n6739) );
  OAI21_X1 U8125 ( .B1(n7437), .B2(n7436), .A(n7438), .ZN(n12170) );
  NAND2_X1 U8126 ( .A1(n12167), .A2(n7439), .ZN(n7438) );
  NAND2_X1 U8127 ( .A1(n12608), .A2(n12656), .ZN(n6750) );
  INV_X1 U8128 ( .A(n7001), .ZN(n6998) );
  INV_X1 U8129 ( .A(n8571), .ZN(n6999) );
  INV_X1 U8130 ( .A(n12925), .ZN(n6676) );
  OAI21_X1 U8131 ( .B1(n7416), .B2(n6467), .A(n7414), .ZN(n7413) );
  OAI21_X1 U8132 ( .B1(n8589), .B2(n6465), .A(n6550), .ZN(n8607) );
  INV_X1 U8133 ( .A(n8644), .ZN(n6991) );
  NAND2_X1 U8134 ( .A1(n8631), .A2(n8629), .ZN(n6992) );
  NOR2_X1 U8135 ( .A1(n8629), .A2(n8631), .ZN(n6993) );
  INV_X1 U8136 ( .A(n12198), .ZN(n7412) );
  NOR2_X1 U8137 ( .A1(n6746), .A2(n12512), .ZN(n6745) );
  INV_X1 U8138 ( .A(n12641), .ZN(n6746) );
  NAND2_X1 U8139 ( .A1(n7392), .A2(n7395), .ZN(n7391) );
  NOR2_X1 U8140 ( .A1(n7412), .A2(n12197), .ZN(n7411) );
  AOI21_X1 U8141 ( .B1(n7407), .B2(n7405), .A(n7404), .ZN(n7403) );
  INV_X1 U8142 ( .A(n12201), .ZN(n7404) );
  NOR2_X1 U8143 ( .A1(n7405), .A2(n12200), .ZN(n7409) );
  NAND2_X1 U8144 ( .A1(n6986), .A2(n6987), .ZN(n8683) );
  NAND2_X1 U8145 ( .A1(n8666), .A2(n6988), .ZN(n6987) );
  NAND2_X1 U8146 ( .A1(n7403), .A2(n7406), .ZN(n7399) );
  INV_X1 U8147 ( .A(n7407), .ZN(n7406) );
  NAND2_X1 U8148 ( .A1(n7409), .A2(n7411), .ZN(n7398) );
  INV_X1 U8149 ( .A(n7403), .ZN(n7402) );
  INV_X1 U8150 ( .A(n7409), .ZN(n7401) );
  NAND2_X1 U8151 ( .A1(n8735), .A2(n9655), .ZN(n6984) );
  OR2_X1 U8152 ( .A1(n8735), .A2(n10797), .ZN(n6985) );
  INV_X1 U8153 ( .A(n8394), .ZN(n7233) );
  INV_X1 U8154 ( .A(n9825), .ZN(n7066) );
  NOR2_X1 U8155 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7374) );
  NAND2_X1 U8156 ( .A1(n12058), .A2(n12283), .ZN(n12072) );
  NAND2_X1 U8157 ( .A1(n9657), .A2(n8145), .ZN(n8735) );
  OR2_X1 U8158 ( .A1(n14536), .A2(n11239), .ZN(n8145) );
  NAND2_X1 U8159 ( .A1(n7261), .A2(SI_18_), .ZN(n6843) );
  INV_X1 U8160 ( .A(n8536), .ZN(n7258) );
  NAND2_X1 U8161 ( .A1(n7256), .A2(n8499), .ZN(n6841) );
  NAND2_X1 U8162 ( .A1(n8368), .A2(n8367), .ZN(n6837) );
  OAI21_X1 U8163 ( .B1(n8622), .B2(n9850), .A(n6718), .ZN(n8206) );
  NAND2_X1 U8164 ( .A1(n8622), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6718) );
  INV_X1 U8165 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7493) );
  AOI21_X1 U8166 ( .B1(n9531), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n9530), .ZN(
        n9532) );
  AND2_X1 U8167 ( .A1(n9585), .A2(n9584), .ZN(n9530) );
  OAI21_X1 U8168 ( .B1(n6453), .B2(n10136), .A(n6773), .ZN(n10139) );
  NAND2_X1 U8169 ( .A1(n6452), .A2(n10136), .ZN(n6773) );
  NAND2_X1 U8170 ( .A1(n6877), .A2(n6482), .ZN(n10556) );
  INV_X1 U8171 ( .A(n7089), .ZN(n7087) );
  INV_X1 U8172 ( .A(n12915), .ZN(n7970) );
  NOR2_X1 U8173 ( .A1(n7761), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7776) );
  AND2_X1 U8174 ( .A1(n11814), .A2(n12599), .ZN(n12591) );
  INV_X1 U8175 ( .A(n12550), .ZN(n7372) );
  INV_X1 U8176 ( .A(n12544), .ZN(n7369) );
  NAND2_X1 U8177 ( .A1(n12704), .A2(n10675), .ZN(n12549) );
  NAND2_X1 U8178 ( .A1(n10629), .A2(n10584), .ZN(n12544) );
  NAND2_X1 U8179 ( .A1(n12524), .A2(n12532), .ZN(n10395) );
  INV_X1 U8180 ( .A(n7974), .ZN(n7059) );
  OR2_X1 U8181 ( .A1(n13082), .A2(n12914), .ZN(n12639) );
  NAND2_X1 U8182 ( .A1(n7068), .A2(n7967), .ZN(n7067) );
  INV_X1 U8183 ( .A(n7069), .ZN(n7068) );
  NAND2_X1 U8184 ( .A1(n7078), .A2(n7077), .ZN(n7076) );
  OR2_X1 U8185 ( .A1(n11821), .A2(n8871), .ZN(n12599) );
  NAND2_X1 U8186 ( .A1(n6730), .A2(n8012), .ZN(n8027) );
  NAND2_X1 U8187 ( .A1(n8011), .A2(n11536), .ZN(n6730) );
  INV_X1 U8188 ( .A(n8903), .ZN(n6915) );
  NAND2_X1 U8189 ( .A1(n7874), .A2(n7873), .ZN(n7877) );
  INV_X1 U8190 ( .A(n7849), .ZN(n6920) );
  NAND2_X1 U8191 ( .A1(n7821), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7834) );
  AND2_X1 U8192 ( .A1(n7317), .A2(n7316), .ZN(n7315) );
  INV_X1 U8193 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7316) );
  INV_X1 U8194 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7304) );
  INV_X1 U8195 ( .A(n7548), .ZN(n6905) );
  INV_X1 U8196 ( .A(n13410), .ZN(n7236) );
  OR2_X1 U8197 ( .A1(n9417), .A2(n13257), .ZN(n9435) );
  AOI21_X1 U8198 ( .B1(n6838), .B2(n6517), .A(n7053), .ZN(n7052) );
  INV_X1 U8199 ( .A(n13368), .ZN(n7053) );
  INV_X1 U8200 ( .A(n13535), .ZN(n6838) );
  NAND2_X1 U8201 ( .A1(n13392), .A2(n13394), .ZN(n7266) );
  OR2_X1 U8202 ( .A1(n13720), .A2(n13362), .ZN(n13398) );
  INV_X1 U8203 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15098) );
  AND2_X1 U8204 ( .A1(n12065), .A2(n10089), .ZN(n12058) );
  NAND2_X1 U8205 ( .A1(n9013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9011) );
  AND3_X1 U8206 ( .A1(n8962), .A2(n9056), .A3(n8961), .ZN(n9000) );
  INV_X1 U8207 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8960) );
  NOR2_X1 U8208 ( .A1(n9098), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9102) );
  OR2_X1 U8209 ( .A1(n9071), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U8210 ( .A1(n7197), .A2(n7202), .ZN(n7195) );
  INV_X1 U8211 ( .A(n11425), .ZN(n7202) );
  INV_X1 U8212 ( .A(n11069), .ZN(n7200) );
  OR2_X1 U8213 ( .A1(n9750), .A2(n14011), .ZN(n7212) );
  INV_X1 U8214 ( .A(n11653), .ZN(n7166) );
  NAND2_X1 U8215 ( .A1(n6562), .A2(n7017), .ZN(n7014) );
  NAND2_X1 U8216 ( .A1(n8512), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6954) );
  AOI22_X1 U8217 ( .A1(n14720), .A2(n14719), .B1(P1_REG1_REG_17__SCAN_IN), 
        .B2(n14721), .ZN(n14176) );
  NAND2_X1 U8218 ( .A1(n14231), .A2(n6789), .ZN(n6787) );
  NOR2_X1 U8219 ( .A1(n7111), .A2(n7115), .ZN(n6788) );
  NAND2_X1 U8220 ( .A1(n14425), .A2(n14006), .ZN(n6980) );
  AND2_X1 U8221 ( .A1(n14253), .A2(n11975), .ZN(n6979) );
  INV_X1 U8222 ( .A(n11991), .ZN(n7117) );
  INV_X1 U8223 ( .A(n8562), .ZN(n8563) );
  NOR2_X1 U8224 ( .A1(n14462), .A2(n6867), .ZN(n6866) );
  INV_X1 U8225 ( .A(n6868), .ZN(n6867) );
  NOR2_X1 U8226 ( .A1(n14470), .A2(n14356), .ZN(n6868) );
  OR2_X1 U8227 ( .A1(n6794), .A2(n11674), .ZN(n6793) );
  NOR2_X1 U8228 ( .A1(n7120), .A2(n7119), .ZN(n7118) );
  INV_X1 U8229 ( .A(n11789), .ZN(n7119) );
  INV_X1 U8230 ( .A(n6795), .ZN(n6794) );
  NOR2_X1 U8231 ( .A1(n14643), .A2(n11951), .ZN(n6853) );
  NOR2_X1 U8232 ( .A1(n11768), .A2(n6857), .ZN(n6856) );
  INV_X1 U8233 ( .A(n6858), .ZN(n6857) );
  NOR2_X1 U8234 ( .A1(n14792), .A2(n11488), .ZN(n6858) );
  OR2_X1 U8235 ( .A1(n8317), .A2(n8316), .ZN(n8359) );
  OR2_X1 U8236 ( .A1(n11431), .A2(n8767), .ZN(n11352) );
  AND2_X1 U8237 ( .A1(n11165), .A2(n8769), .ZN(n11272) );
  AND2_X1 U8238 ( .A1(n10926), .A2(n10927), .ZN(n11098) );
  NAND2_X1 U8239 ( .A1(n14404), .A2(n14793), .ZN(n6864) );
  NAND2_X1 U8240 ( .A1(n11740), .A2(n11681), .ZN(n11805) );
  INV_X1 U8241 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8816) );
  AND2_X1 U8242 ( .A1(n7012), .A2(n7011), .ZN(n7010) );
  NOR2_X1 U8243 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8050) );
  NOR2_X1 U8244 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8346) );
  AOI21_X1 U8245 ( .B1(n7245), .B2(n7247), .A(n7243), .ZN(n7242) );
  INV_X1 U8246 ( .A(n8344), .ZN(n7243) );
  NAND2_X1 U8247 ( .A1(n8187), .A2(n8186), .ZN(n8190) );
  NAND2_X1 U8248 ( .A1(n8190), .A2(n8189), .ZN(n8205) );
  OAI21_X1 U8249 ( .B1(n8622), .B2(n9811), .A(n7217), .ZN(n7216) );
  NAND2_X1 U8250 ( .A1(n8622), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7217) );
  INV_X1 U8251 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15097) );
  NOR2_X1 U8252 ( .A1(n9518), .A2(n9519), .ZN(n9520) );
  INV_X1 U8253 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15131) );
  XNOR2_X1 U8254 ( .A(n9520), .B(n15131), .ZN(n9569) );
  OAI22_X1 U8255 ( .A1(n9576), .A2(n9524), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n9523), .ZN(n9525) );
  INV_X1 U8256 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9523) );
  AOI21_X1 U8257 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n9529), .A(n9528), .ZN(
        n9584) );
  NOR2_X1 U8258 ( .A1(n9553), .A2(n9552), .ZN(n9528) );
  OR2_X1 U8259 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n9532), .ZN(n9549) );
  AOI21_X1 U8260 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n9535), .A(n9534), .ZN(
        n9545) );
  NOR2_X1 U8261 ( .A1(n9548), .A2(n9547), .ZN(n9534) );
  AND2_X1 U8262 ( .A1(n8839), .A2(n8837), .ZN(n10400) );
  NAND2_X1 U8263 ( .A1(n6658), .A2(n6539), .ZN(n7303) );
  OR2_X1 U8264 ( .A1(n11905), .A2(n12980), .ZN(n7294) );
  INV_X1 U8265 ( .A(n7303), .ZN(n12423) );
  INV_X1 U8266 ( .A(n11383), .ZN(n7299) );
  INV_X1 U8267 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U8268 ( .A1(n8851), .A2(n6532), .ZN(n11111) );
  NAND2_X1 U8269 ( .A1(n10810), .A2(n10811), .ZN(n8851) );
  NAND2_X1 U8270 ( .A1(n6889), .A2(n6890), .ZN(n6888) );
  NAND2_X1 U8271 ( .A1(n6481), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7511) );
  NAND4_X1 U8272 ( .A1(n7483), .A2(n7481), .A3(n7484), .A4(n7482), .ZN(n14986)
         );
  NAND2_X1 U8273 ( .A1(n7662), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7483) );
  INV_X1 U8274 ( .A(n8919), .ZN(n9654) );
  OR2_X1 U8275 ( .A1(n10203), .A2(n15040), .ZN(n10205) );
  NAND2_X1 U8276 ( .A1(n10186), .A2(n10185), .ZN(n10189) );
  NAND2_X1 U8277 ( .A1(n10285), .A2(n6714), .ZN(n10246) );
  NAND2_X1 U8278 ( .A1(n6716), .A2(n6715), .ZN(n6714) );
  INV_X1 U8279 ( .A(n10244), .ZN(n6716) );
  NAND2_X1 U8280 ( .A1(n10283), .A2(n10284), .ZN(n10554) );
  OAI21_X1 U8281 ( .B1(n10177), .B2(n6561), .A(n6942), .ZN(n10279) );
  NAND2_X1 U8282 ( .A1(n6932), .A2(n6931), .ZN(n6930) );
  INV_X1 U8283 ( .A(n10544), .ZN(n6932) );
  NAND2_X1 U8284 ( .A1(n10557), .A2(n10556), .ZN(n10896) );
  INV_X1 U8285 ( .A(n10556), .ZN(n10558) );
  INV_X1 U8286 ( .A(n12734), .ZN(n6935) );
  INV_X1 U8287 ( .A(n12736), .ZN(n6772) );
  INV_X1 U8288 ( .A(n6754), .ZN(n12727) );
  NAND2_X1 U8289 ( .A1(n7739), .A2(n7315), .ZN(n7791) );
  XNOR2_X1 U8290 ( .A(n12804), .B(n6668), .ZN(n12813) );
  INV_X1 U8291 ( .A(n12805), .ZN(n6668) );
  AND4_X1 U8292 ( .A1(n12477), .A2(n9637), .A3(n9636), .A4(n9635), .ZN(n12493)
         );
  OR2_X1 U8293 ( .A1(n7909), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7924) );
  OR2_X1 U8294 ( .A1(n7895), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U8295 ( .A1(n7854), .A2(n7853), .ZN(n7866) );
  INV_X1 U8296 ( .A(n7855), .ZN(n7854) );
  NAND2_X1 U8297 ( .A1(n7810), .A2(n7809), .ZN(n7828) );
  NAND2_X1 U8298 ( .A1(n7743), .A2(n11908), .ZN(n7761) );
  AND2_X1 U8299 ( .A1(n7709), .A2(n11754), .ZN(n7726) );
  INV_X1 U8300 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7725) );
  AND2_X1 U8301 ( .A1(n7726), .A2(n7725), .ZN(n7743) );
  INV_X1 U8302 ( .A(n12591), .ZN(n12506) );
  NOR2_X1 U8303 ( .A1(n7693), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7709) );
  INV_X1 U8304 ( .A(n7956), .ZN(n14583) );
  OR2_X1 U8305 ( .A1(n7660), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U8306 ( .A1(n7630), .A2(n7629), .ZN(n7660) );
  AOI21_X1 U8307 ( .B1(n7364), .B2(n7366), .A(n7362), .ZN(n7361) );
  INV_X1 U8308 ( .A(n12570), .ZN(n7362) );
  INV_X1 U8309 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10551) );
  NOR2_X1 U8310 ( .A1(n7590), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7608) );
  AND2_X1 U8311 ( .A1(n7608), .A2(n10551), .ZN(n7630) );
  OR2_X1 U8312 ( .A1(n7577), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7590) );
  AND2_X1 U8313 ( .A1(n12560), .A2(n12558), .ZN(n12498) );
  NAND2_X1 U8314 ( .A1(n10495), .A2(n12544), .ZN(n10625) );
  INV_X1 U8315 ( .A(n7943), .ZN(n12534) );
  NAND2_X1 U8316 ( .A1(n14986), .A2(n7938), .ZN(n14990) );
  CLKBUF_X1 U8317 ( .A(n10395), .Z(n6779) );
  INV_X1 U8318 ( .A(n8834), .ZN(n7939) );
  NAND2_X1 U8319 ( .A1(n6558), .A2(n7360), .ZN(n7353) );
  INV_X1 U8320 ( .A(n12522), .ZN(n7355) );
  AND2_X1 U8321 ( .A1(n12657), .A2(n12658), .ZN(n12854) );
  OAI21_X1 U8322 ( .B1(n12878), .B2(n12644), .A(n12645), .ZN(n12864) );
  NAND2_X1 U8323 ( .A1(n7060), .A2(n7974), .ZN(n12880) );
  INV_X1 U8324 ( .A(n12644), .ZN(n12879) );
  AOI21_X1 U8325 ( .B1(n7378), .B2(n7377), .A(n7376), .ZN(n7375) );
  INV_X1 U8326 ( .A(n12632), .ZN(n7377) );
  INV_X1 U8327 ( .A(n12635), .ZN(n7376) );
  OAI21_X1 U8328 ( .B1(n6766), .B2(n7965), .A(n7076), .ZN(n12967) );
  AOI21_X1 U8329 ( .B1(n7343), .B2(n7346), .A(n7340), .ZN(n7339) );
  INV_X1 U8330 ( .A(n12618), .ZN(n12966) );
  NOR2_X1 U8331 ( .A1(n14602), .A2(n8871), .ZN(n7064) );
  OR2_X1 U8332 ( .A1(n11821), .A2(n14577), .ZN(n7063) );
  INV_X1 U8333 ( .A(n12954), .ZN(n14991) );
  INV_X1 U8334 ( .A(n12958), .ZN(n14988) );
  INV_X1 U8335 ( .A(n15026), .ZN(n15015) );
  INV_X1 U8336 ( .A(n8027), .ZN(n9907) );
  OAI22_X2 U8337 ( .A1(n8027), .A2(P3_D_REG_0__SCAN_IN), .B1(n8013), .B2(n8012), .ZN(n10347) );
  INV_X1 U8338 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7473) );
  NAND2_X1 U8339 ( .A1(n6912), .A2(n6913), .ZN(n12031) );
  AOI21_X1 U8340 ( .B1(n6914), .B2(n6479), .A(n6605), .ZN(n6913) );
  NAND2_X1 U8341 ( .A1(n7488), .A2(n7487), .ZN(n12687) );
  NAND2_X1 U8342 ( .A1(n6645), .A2(n6643), .ZN(n7487) );
  NAND2_X1 U8343 ( .A1(n6644), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6643) );
  OAI21_X1 U8344 ( .B1(n7486), .B2(n7485), .A(P3_IR_REG_28__SCAN_IN), .ZN(
        n6645) );
  NAND2_X1 U8345 ( .A1(n7999), .A2(n7472), .ZN(n7996) );
  NAND4_X1 U8346 ( .A1(n7467), .A2(n7994), .A3(n7468), .A4(n7466), .ZN(n7469)
         );
  INV_X1 U8347 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7466) );
  XNOR2_X1 U8348 ( .A(n7994), .B(n7995), .ZN(n10130) );
  OAI21_X1 U8349 ( .B1(n7993), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U8350 ( .A1(n7930), .A2(n7467), .ZN(n7993) );
  NAND2_X1 U8351 ( .A1(n7931), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7932) );
  AND2_X1 U8352 ( .A1(n7849), .A2(n7836), .ZN(n7837) );
  XNOR2_X1 U8353 ( .A(n7463), .B(P3_IR_REG_20__SCAN_IN), .ZN(n8035) );
  AND2_X1 U8354 ( .A1(n7315), .A2(n7314), .ZN(n7313) );
  INV_X1 U8355 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7314) );
  AND2_X1 U8356 ( .A1(n7819), .A2(n7803), .ZN(n7804) );
  AOI21_X1 U8357 ( .B1(n6909), .B2(n6911), .A(n6908), .ZN(n6907) );
  INV_X1 U8358 ( .A(n7786), .ZN(n6908) );
  NOR2_X1 U8359 ( .A1(n7758), .A2(n7757), .ZN(n12740) );
  INV_X1 U8360 ( .A(n6893), .ZN(n6892) );
  INV_X1 U8361 ( .A(n7719), .ZN(n6894) );
  AND2_X1 U8362 ( .A1(n7749), .A2(n7735), .ZN(n7736) );
  NAND2_X1 U8363 ( .A1(n6897), .A2(n6895), .ZN(n7686) );
  AOI21_X1 U8364 ( .B1(n6898), .B2(n6900), .A(n6896), .ZN(n6895) );
  NAND2_X1 U8365 ( .A1(n7652), .A2(n6898), .ZN(n6897) );
  INV_X1 U8366 ( .A(n7682), .ZN(n6896) );
  AND2_X1 U8367 ( .A1(n7698), .A2(n7684), .ZN(n7685) );
  NAND2_X1 U8368 ( .A1(n7686), .A2(n7685), .ZN(n7699) );
  AND2_X1 U8369 ( .A1(n7648), .A2(n7638), .ZN(n7639) );
  AND2_X1 U8370 ( .A1(n7636), .A2(n7623), .ZN(n7624) );
  OR2_X1 U8371 ( .A1(n7614), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U8372 ( .A1(n7599), .A2(n7598), .ZN(n7621) );
  AND2_X1 U8373 ( .A1(n7622), .A2(n7601), .ZN(n7619) );
  NOR2_X1 U8374 ( .A1(n7583), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7603) );
  INV_X1 U8375 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U8376 ( .A1(n7552), .A2(n7551), .ZN(n7554) );
  AND2_X1 U8377 ( .A1(n7521), .A2(n7522), .ZN(n7552) );
  INV_X1 U8378 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U8379 ( .A1(n6826), .A2(n7321), .ZN(n6821) );
  AND2_X1 U8380 ( .A1(n9261), .A2(n9240), .ZN(n7326) );
  OR2_X1 U8381 ( .A1(n11435), .A2(n11434), .ZN(n7327) );
  NAND2_X1 U8382 ( .A1(n13204), .A2(n7337), .ZN(n7336) );
  NOR2_X1 U8383 ( .A1(n13245), .A2(n7338), .ZN(n7337) );
  INV_X1 U8384 ( .A(n9309), .ZN(n7338) );
  NAND2_X1 U8385 ( .A1(n12343), .A2(n12334), .ZN(n7334) );
  NAND2_X1 U8386 ( .A1(n8956), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9373) );
  OAI21_X1 U8387 ( .B1(n10981), .B2(n6814), .A(n6810), .ZN(n11299) );
  NAND2_X1 U8388 ( .A1(n9183), .A2(n6811), .ZN(n6814) );
  AOI22_X1 U8389 ( .A1(n6813), .A2(n6812), .B1(n6811), .B2(n6599), .ZN(n6810)
         );
  NOR2_X1 U8390 ( .A1(n13150), .A2(n7449), .ZN(n13215) );
  NAND2_X1 U8391 ( .A1(n11299), .A2(n11300), .ZN(n11298) );
  XNOR2_X1 U8392 ( .A(n13164), .B(n6761), .ZN(n10435) );
  NAND2_X1 U8393 ( .A1(n10373), .A2(n7332), .ZN(n10819) );
  AND2_X1 U8394 ( .A1(n12343), .A2(n12283), .ZN(n9861) );
  AND2_X1 U8395 ( .A1(n7385), .A2(n7387), .ZN(n6757) );
  AND2_X1 U8396 ( .A1(n12264), .A2(n7388), .ZN(n7387) );
  NAND2_X1 U8397 ( .A1(n12273), .A2(n12274), .ZN(n7386) );
  NAND2_X1 U8398 ( .A1(n12272), .A2(n12324), .ZN(n12275) );
  NAND2_X1 U8399 ( .A1(n12235), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U8400 ( .A1(n9936), .A2(n6523), .ZN(n9887) );
  NAND2_X1 U8401 ( .A1(n13301), .A2(n6529), .ZN(n14830) );
  NOR2_X1 U8402 ( .A1(n13312), .A2(n6704), .ZN(n13314) );
  NOR2_X1 U8403 ( .A1(n13318), .A2(n6705), .ZN(n6704) );
  INV_X1 U8404 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U8405 ( .A1(n14862), .A2(n14861), .ZN(n14860) );
  INV_X1 U8406 ( .A(n9310), .ZN(n9005) );
  AND2_X1 U8407 ( .A1(n9497), .A2(n9496), .ZN(n13436) );
  NAND2_X1 U8408 ( .A1(n13515), .A2(n13516), .ZN(n13514) );
  NAND2_X1 U8409 ( .A1(n13507), .A2(n13512), .ZN(n13508) );
  INV_X1 U8410 ( .A(n13645), .ZN(n7267) );
  AND3_X1 U8411 ( .A1(n9303), .A2(n9302), .A3(n9301), .ZN(n13393) );
  NAND2_X1 U8412 ( .A1(n8952), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9284) );
  OR2_X1 U8413 ( .A1(n9230), .A2(n9229), .ZN(n9249) );
  OR2_X1 U8414 ( .A1(n9249), .A2(n9248), .ZN(n9271) );
  NAND2_X1 U8415 ( .A1(n7057), .A2(n11557), .ZN(n11559) );
  AND4_X1 U8416 ( .A1(n9219), .A2(n9218), .A3(n9217), .A4(n9216), .ZN(n12150)
         );
  OR2_X1 U8417 ( .A1(n9195), .A2(n9194), .ZN(n9214) );
  NAND2_X1 U8418 ( .A1(n8951), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9230) );
  INV_X1 U8419 ( .A(n9214), .ZN(n8951) );
  NOR2_X1 U8420 ( .A1(n7039), .A2(n12311), .ZN(n7038) );
  INV_X1 U8421 ( .A(n7041), .ZN(n7039) );
  OR2_X1 U8422 ( .A1(n9156), .A2(n8949), .ZN(n9172) );
  CLKBUF_X1 U8423 ( .A(n11290), .Z(n6743) );
  INV_X1 U8424 ( .A(n12307), .ZN(n6629) );
  XNOR2_X1 U8425 ( .A(n10995), .B(n13289), .ZN(n12307) );
  INV_X1 U8426 ( .A(n12305), .ZN(n6774) );
  AND4_X1 U8427 ( .A1(n9146), .A2(n9145), .A3(n9144), .A4(n9143), .ZN(n12123)
         );
  INV_X1 U8428 ( .A(n13542), .ZN(n13630) );
  NOR2_X2 U8429 ( .A1(n10754), .A2(n12102), .ZN(n10773) );
  NAND2_X1 U8430 ( .A1(n10450), .A2(n10420), .ZN(n10421) );
  XNOR2_X1 U8431 ( .A(n12343), .B(n12286), .ZN(n7335) );
  NAND2_X1 U8432 ( .A1(n10517), .A2(n12063), .ZN(n12062) );
  NAND2_X1 U8433 ( .A1(n12248), .A2(n12247), .ZN(n13336) );
  INV_X1 U8434 ( .A(n13593), .ZN(n13725) );
  NAND2_X1 U8435 ( .A1(n13628), .A2(n13351), .ZN(n13614) );
  NAND2_X1 U8436 ( .A1(n7044), .A2(n7043), .ZN(n11367) );
  NAND2_X1 U8437 ( .A1(n6462), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6801) );
  CLKBUF_X1 U8438 ( .A(n12058), .Z(n14901) );
  CLKBUF_X1 U8439 ( .A(n9499), .Z(n9500) );
  OR2_X1 U8440 ( .A1(n9456), .A2(n9455), .ZN(n9482) );
  XNOR2_X1 U8441 ( .A(n8997), .B(n8996), .ZN(n12330) );
  INV_X1 U8442 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8996) );
  NAND2_X1 U8443 ( .A1(n8995), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8997) );
  AND2_X1 U8444 ( .A1(n9190), .A2(n9205), .ZN(n10597) );
  OR2_X1 U8445 ( .A1(n9119), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9137) );
  OR2_X1 U8446 ( .A1(n9137), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9167) );
  NOR2_X1 U8447 ( .A1(n9059), .A2(n9058), .ZN(n9883) );
  AND2_X2 U8448 ( .A1(n6622), .A2(n6621), .ZN(n9018) );
  INV_X1 U8449 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6622) );
  INV_X1 U8450 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6621) );
  NOR2_X1 U8451 ( .A1(n8527), .A2(n8526), .ZN(n8545) );
  OR2_X1 U8452 ( .A1(n8510), .A2(n8509), .ZN(n8527) );
  AOI21_X1 U8453 ( .B1(n13813), .B2(n13812), .A(n13918), .ZN(n13888) );
  INV_X1 U8454 ( .A(n7195), .ZN(n7194) );
  NAND2_X1 U8455 ( .A1(n11070), .A2(n7199), .ZN(n7196) );
  NOR2_X1 U8456 ( .A1(n13938), .A2(n7205), .ZN(n7204) );
  INV_X1 U8457 ( .A(n13827), .ZN(n7205) );
  AND2_X1 U8458 ( .A1(n13875), .A2(n13873), .ZN(n13947) );
  AND2_X1 U8459 ( .A1(n8467), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8469) );
  AND2_X1 U8460 ( .A1(n13946), .A2(n13861), .ZN(n13969) );
  NAND2_X1 U8461 ( .A1(n7172), .A2(n7171), .ZN(n7170) );
  INV_X1 U8462 ( .A(n9722), .ZN(n7172) );
  XNOR2_X1 U8463 ( .A(n9678), .B(n13921), .ZN(n9681) );
  OAI21_X1 U8464 ( .B1(n9766), .B2(n7190), .A(n7187), .ZN(n13909) );
  NAND2_X1 U8465 ( .A1(n8609), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U8466 ( .A1(n13949), .A2(n13875), .ZN(n14002) );
  OR2_X1 U8467 ( .A1(n8419), .A2(n8418), .ZN(n8435) );
  NOR2_X1 U8468 ( .A1(n8435), .A2(n14013), .ZN(n8467) );
  AND4_X1 U8469 ( .A1(n8441), .A2(n8440), .A3(n8439), .A4(n8438), .ZN(n11920)
         );
  NAND4_X1 U8470 ( .A1(n8077), .A2(n8076), .A3(n8075), .A4(n8074), .ZN(n14039)
         );
  OR2_X1 U8471 ( .A1(n8689), .A2(n11194), .ZN(n8075) );
  INV_X1 U8472 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14058) );
  INV_X1 U8473 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15108) );
  OR2_X1 U8474 ( .A1(n8277), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8278) );
  NOR2_X1 U8475 ( .A1(n14404), .A2(n12018), .ZN(n14208) );
  NOR2_X1 U8476 ( .A1(n6483), .A2(n14425), .ZN(n14234) );
  AND2_X1 U8477 ( .A1(n14264), .A2(n11975), .ZN(n14252) );
  AND2_X1 U8478 ( .A1(n14264), .A2(n6979), .ZN(n14259) );
  XNOR2_X1 U8479 ( .A(n14251), .B(n14276), .ZN(n14253) );
  NAND3_X1 U8480 ( .A1(n14352), .A2(n6865), .A3(n6866), .ZN(n14306) );
  AOI21_X1 U8481 ( .B1(n6464), .B2(n14335), .A(n6540), .ZN(n6962) );
  NAND2_X1 U8482 ( .A1(n14352), .A2(n6866), .ZN(n14321) );
  NAND2_X1 U8483 ( .A1(n14352), .A2(n14476), .ZN(n14353) );
  AOI21_X1 U8484 ( .B1(n6501), .B2(n11930), .A(n6966), .ZN(n6965) );
  AND2_X1 U8485 ( .A1(n11740), .A2(n6570), .ZN(n14372) );
  NAND2_X1 U8486 ( .A1(n11740), .A2(n6851), .ZN(n11919) );
  NAND2_X1 U8487 ( .A1(n7096), .A2(n7095), .ZN(n11734) );
  AOI21_X1 U8488 ( .B1(n7097), .B2(n7099), .A(n6543), .ZN(n7095) );
  NAND2_X1 U8489 ( .A1(n11356), .A2(n7097), .ZN(n7096) );
  AOI21_X1 U8490 ( .B1(n6958), .B2(n6960), .A(n6544), .ZN(n6956) );
  NAND2_X1 U8491 ( .A1(n11484), .A2(n6856), .ZN(n11741) );
  NAND2_X1 U8492 ( .A1(n11576), .A2(n11575), .ZN(n11668) );
  NAND2_X1 U8493 ( .A1(n11346), .A2(n11345), .ZN(n11576) );
  OR2_X1 U8494 ( .A1(n10014), .A2(n8656), .ZN(n8313) );
  NOR2_X1 U8495 ( .A1(n11254), .A2(n11431), .ZN(n11484) );
  NAND2_X1 U8496 ( .A1(n11484), .A2(n11621), .ZN(n11485) );
  NOR2_X1 U8497 ( .A1(n11447), .A2(n10727), .ZN(n10926) );
  AND3_X1 U8498 ( .A1(n12018), .A2(n14370), .A3(n12006), .ZN(n14406) );
  NAND2_X1 U8499 ( .A1(n7114), .A2(n6497), .ZN(n12039) );
  AND2_X1 U8500 ( .A1(n7113), .A2(n7114), .ZN(n12038) );
  NAND2_X1 U8501 ( .A1(n6791), .A2(n7112), .ZN(n7114) );
  INV_X1 U8502 ( .A(n14355), .ZN(n14370) );
  AND2_X1 U8503 ( .A1(n9770), .A2(n9771), .ZN(n14793) );
  AND2_X1 U8504 ( .A1(n7207), .A2(n6512), .ZN(n8068) );
  XNOR2_X1 U8505 ( .A(n8825), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U8506 ( .A1(n6492), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8825) );
  AND2_X1 U8507 ( .A1(n8639), .A2(n8625), .ZN(n13802) );
  NAND2_X1 U8508 ( .A1(n8063), .A2(n7012), .ZN(n8505) );
  OR2_X1 U8509 ( .A1(n8370), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8371) );
  INV_X1 U8510 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8054) );
  OAI21_X1 U8511 ( .B1(n8130), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6776), .ZN(
        n8104) );
  NAND2_X1 U8512 ( .A1(n8130), .A2(n8102), .ZN(n6776) );
  NAND2_X1 U8513 ( .A1(n9514), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n7128) );
  NAND2_X1 U8514 ( .A1(n7131), .A2(n9577), .ZN(n9579) );
  NAND2_X1 U8515 ( .A1(n14548), .A2(n14547), .ZN(n7131) );
  INV_X1 U8516 ( .A(n6673), .ZN(n9586) );
  OAI21_X1 U8517 ( .B1(n14549), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6511), .ZN(
        n6673) );
  NAND2_X1 U8518 ( .A1(n7141), .A2(n9592), .ZN(n9594) );
  NAND2_X1 U8519 ( .A1(n14551), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7141) );
  AOI21_X1 U8520 ( .B1(n7150), .B2(n7147), .A(n7146), .ZN(n7145) );
  NOR2_X1 U8521 ( .A1(n7150), .A2(n7149), .ZN(n7148) );
  INV_X1 U8522 ( .A(n7151), .ZN(n7147) );
  OAI21_X1 U8523 ( .B1(n7279), .B2(n7278), .A(n7282), .ZN(n11881) );
  AND2_X1 U8524 ( .A1(n7283), .A2(n11750), .ZN(n7282) );
  OR2_X1 U8525 ( .A1(n8901), .A2(n12696), .ZN(n6674) );
  NAND2_X1 U8526 ( .A1(n7842), .A2(n7841), .ZN(n13021) );
  NAND2_X1 U8527 ( .A1(n8869), .A2(n11633), .ZN(n11722) );
  NAND2_X1 U8528 ( .A1(n7289), .A2(n7293), .ZN(n12405) );
  NAND2_X1 U8529 ( .A1(n6712), .A2(n7294), .ZN(n7289) );
  NAND2_X1 U8530 ( .A1(n7288), .A2(n7286), .ZN(n12415) );
  AOI21_X1 U8531 ( .B1(n7290), .B2(n7292), .A(n7287), .ZN(n7286) );
  INV_X1 U8532 ( .A(n12404), .ZN(n7287) );
  NAND2_X1 U8533 ( .A1(n12377), .A2(n8859), .ZN(n11382) );
  NAND2_X1 U8534 ( .A1(n7281), .A2(n7280), .ZN(n11751) );
  INV_X1 U8535 ( .A(n7284), .ZN(n7280) );
  OR2_X1 U8536 ( .A1(n11722), .A2(n8870), .ZN(n7281) );
  NAND2_X1 U8537 ( .A1(n8913), .A2(n8912), .ZN(n12449) );
  NAND2_X1 U8538 ( .A1(n8851), .A2(n8850), .ZN(n11113) );
  OR2_X1 U8539 ( .A1(n8938), .A2(n8936), .ZN(n12455) );
  CLKBUF_X1 U8540 ( .A(n11907), .Z(n6712) );
  INV_X1 U8541 ( .A(n12693), .ZN(n6682) );
  AND4_X1 U8542 ( .A1(n7988), .A2(n7987), .A3(n7986), .A4(n7985), .ZN(n12349)
         );
  NAND4_X1 U8543 ( .A1(n7900), .A2(n7899), .A3(n7898), .A4(n7897), .ZN(n12881)
         );
  NAND4_X1 U8544 ( .A1(n7889), .A2(n7888), .A3(n7887), .A4(n7886), .ZN(n12892)
         );
  INV_X1 U8545 ( .A(n12903), .ZN(n12697) );
  INV_X1 U8546 ( .A(n12941), .ZN(n12969) );
  INV_X1 U8547 ( .A(n12955), .ZN(n12981) );
  NAND4_X1 U8548 ( .A1(n7681), .A2(n7680), .A3(n7679), .A4(n7678), .ZN(n14576)
         );
  INV_X1 U8549 ( .A(n11391), .ZN(n12700) );
  INV_X1 U8550 ( .A(n11001), .ZN(n12701) );
  INV_X1 U8551 ( .A(n11025), .ZN(n12702) );
  CLKBUF_X1 U8552 ( .A(n14986), .Z(n6657) );
  OR2_X2 U8553 ( .A1(n13127), .A2(n9654), .ZN(n12706) );
  AND2_X1 U8554 ( .A1(n6939), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U8555 ( .A1(n6937), .A2(n6940), .ZN(n10238) );
  AND2_X1 U8556 ( .A1(n6938), .A2(n6939), .ZN(n6937) );
  NAND2_X1 U8557 ( .A1(n6878), .A2(n6482), .ZN(n14931) );
  INV_X1 U8558 ( .A(n10546), .ZN(n10550) );
  INV_X1 U8559 ( .A(n6875), .ZN(n14948) );
  NAND2_X1 U8560 ( .A1(n6873), .A2(n6872), .ZN(n11685) );
  INV_X1 U8561 ( .A(n11407), .ZN(n6872) );
  INV_X1 U8562 ( .A(n6936), .ZN(n12735) );
  NAND2_X1 U8563 ( .A1(n6648), .A2(n6506), .ZN(n6882) );
  INV_X1 U8564 ( .A(n6883), .ZN(n12718) );
  INV_X1 U8565 ( .A(n6934), .ZN(n12743) );
  NOR2_X1 U8566 ( .A1(n12706), .A2(n10128), .ZN(n14936) );
  NAND2_X1 U8567 ( .A1(n7894), .A2(n7893), .ZN(n13008) );
  NAND2_X1 U8568 ( .A1(n12923), .A2(n7969), .ZN(n12912) );
  NAND2_X1 U8569 ( .A1(n7070), .A2(n7071), .ZN(n12951) );
  NAND2_X1 U8570 ( .A1(n11464), .A2(n7093), .ZN(n11393) );
  AND2_X1 U8571 ( .A1(n7644), .A2(n7643), .ZN(n12574) );
  NAND2_X1 U8572 ( .A1(n11031), .A2(n12564), .ZN(n11463) );
  NAND2_X1 U8573 ( .A1(n10626), .A2(n7946), .ZN(n10883) );
  NAND2_X1 U8574 ( .A1(n10624), .A2(n12550), .ZN(n10887) );
  NAND2_X1 U8575 ( .A1(n10354), .A2(n12675), .ZN(n14580) );
  AND3_X1 U8576 ( .A1(n7576), .A2(n7575), .A3(n7574), .ZN(n11011) );
  NAND2_X1 U8577 ( .A1(n12480), .A2(n12479), .ZN(n13047) );
  NAND2_X1 U8578 ( .A1(n7908), .A2(n7907), .ZN(n13060) );
  NAND2_X1 U8579 ( .A1(n7865), .A2(n7864), .ZN(n13077) );
  OAI21_X1 U8580 ( .B1(n12922), .B2(n12925), .A(n12632), .ZN(n12916) );
  NAND2_X1 U8581 ( .A1(n7808), .A2(n7807), .ZN(n13098) );
  NAND2_X1 U8582 ( .A1(n12950), .A2(n12616), .ZN(n12936) );
  OAI21_X1 U8583 ( .B1(n12987), .B2(n7346), .A(n7343), .ZN(n12975) );
  NAND2_X1 U8584 ( .A1(n7342), .A2(n12610), .ZN(n12976) );
  NAND2_X1 U8585 ( .A1(n7742), .A2(n7741), .ZN(n13122) );
  INV_X1 U8586 ( .A(n11011), .ZN(n11014) );
  NAND2_X1 U8587 ( .A1(n10130), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13127) );
  INV_X1 U8588 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13129) );
  OAI21_X1 U8589 ( .B1(n8902), .B2(n6479), .A(n8903), .ZN(n9627) );
  NAND2_X1 U8590 ( .A1(n7850), .A2(n7849), .ZN(n7863) );
  INV_X1 U8591 ( .A(n12531), .ZN(n10849) );
  INV_X1 U8592 ( .A(SI_20_), .ZN(n10640) );
  INV_X1 U8593 ( .A(n8035), .ZN(n10641) );
  INV_X1 U8594 ( .A(SI_17_), .ZN(n10233) );
  NAND2_X1 U8595 ( .A1(n7768), .A2(n7767), .ZN(n7785) );
  INV_X1 U8596 ( .A(SI_16_), .ZN(n10077) );
  INV_X1 U8597 ( .A(SI_15_), .ZN(n10015) );
  NAND2_X1 U8598 ( .A1(n7720), .A2(n7719), .ZN(n7734) );
  NAND2_X1 U8599 ( .A1(n7717), .A2(n7716), .ZN(n7720) );
  INV_X1 U8600 ( .A(SI_12_), .ZN(n9854) );
  INV_X1 U8601 ( .A(SI_11_), .ZN(n9847) );
  OAI21_X1 U8602 ( .B1(n7652), .B2(n6900), .A(n6898), .ZN(n7683) );
  NAND2_X1 U8603 ( .A1(n7668), .A2(n7667), .ZN(n7671) );
  XNOR2_X1 U8604 ( .A(n7657), .B(n7656), .ZN(n14944) );
  NAND2_X1 U8605 ( .A1(n7549), .A2(n7548), .ZN(n7567) );
  INV_X1 U8606 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10142) );
  AOI21_X1 U8607 ( .B1(n7332), .B2(n7331), .A(n7330), .ZN(n7329) );
  INV_X1 U8608 ( .A(n7332), .ZN(n7328) );
  NAND2_X1 U8609 ( .A1(n7327), .A2(n9240), .ZN(n11612) );
  INV_X1 U8610 ( .A(n13512), .ZN(n13698) );
  NAND2_X1 U8611 ( .A1(n10981), .A2(n6485), .ZN(n11079) );
  NAND2_X1 U8612 ( .A1(n10981), .A2(n9166), .ZN(n11078) );
  NOR2_X1 U8613 ( .A1(n13163), .A2(n13162), .ZN(n13168) );
  NAND2_X1 U8614 ( .A1(n13232), .A2(n6531), .ZN(n13177) );
  NAND2_X1 U8615 ( .A1(n13232), .A2(n9350), .ZN(n13176) );
  AND2_X1 U8616 ( .A1(n9212), .A2(n9211), .ZN(n14631) );
  AND2_X1 U8617 ( .A1(n9283), .A2(n9282), .ZN(n13390) );
  AND2_X1 U8618 ( .A1(n6799), .A2(n6800), .ZN(n13193) );
  INV_X1 U8619 ( .A(n9279), .ZN(n6800) );
  NAND2_X1 U8620 ( .A1(n9093), .A2(n10363), .ZN(n10373) );
  NOR2_X1 U8621 ( .A1(n13215), .A2(n13214), .ZN(n13213) );
  NAND2_X1 U8622 ( .A1(n13215), .A2(n13214), .ZN(n6771) );
  OR2_X1 U8623 ( .A1(n10376), .A2(n10375), .ZN(n10382) );
  AND2_X1 U8624 ( .A1(n9346), .A2(n9345), .ZN(n13247) );
  INV_X1 U8625 ( .A(n13702), .ZN(n13526) );
  XNOR2_X1 U8626 ( .A(n9382), .B(n9380), .ZN(n13235) );
  NAND2_X1 U8627 ( .A1(n11079), .A2(n9183), .ZN(n11182) );
  NAND2_X1 U8628 ( .A1(n13204), .A2(n9309), .ZN(n13246) );
  NAND2_X1 U8629 ( .A1(n10373), .A2(n9097), .ZN(n10821) );
  NAND2_X1 U8630 ( .A1(n6824), .A2(n6826), .ZN(n13254) );
  NAND2_X1 U8631 ( .A1(n13150), .A2(n7322), .ZN(n6824) );
  NAND2_X1 U8632 ( .A1(n9506), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13276) );
  NAND2_X1 U8633 ( .A1(n9488), .A2(n13651), .ZN(n13281) );
  AND2_X1 U8634 ( .A1(n12287), .A2(n12339), .ZN(n7432) );
  NAND2_X1 U8635 ( .A1(n9441), .A2(n9440), .ZN(n13456) );
  INV_X1 U8636 ( .A(n13396), .ZN(n13359) );
  INV_X1 U8637 ( .A(n12150), .ZN(n13285) );
  INV_X1 U8638 ( .A(n12123), .ZN(n13289) );
  INV_X1 U8639 ( .A(n12108), .ZN(n13291) );
  OR2_X1 U8640 ( .A1(n12220), .A2(n9062), .ZN(n9063) );
  NAND2_X1 U8641 ( .A1(n12235), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9049) );
  CLKBUF_X2 U8642 ( .A(n13296), .Z(n6734) );
  NAND2_X1 U8643 ( .A1(n13303), .A2(n13302), .ZN(n13301) );
  NAND2_X1 U8644 ( .A1(n10679), .A2(n6703), .ZN(n10681) );
  OR2_X1 U8645 ( .A1(n10680), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6703) );
  NOR2_X1 U8646 ( .A1(n11594), .A2(n6706), .ZN(n11599) );
  AND2_X1 U8647 ( .A1(n11595), .A2(n11596), .ZN(n6706) );
  AND2_X1 U8648 ( .A1(n12253), .A2(n12252), .ZN(n13428) );
  NAND2_X1 U8649 ( .A1(n13477), .A2(n13410), .ZN(n13451) );
  AND2_X1 U8650 ( .A1(n13494), .A2(n13409), .ZN(n13479) );
  NAND2_X1 U8651 ( .A1(n6755), .A2(n13405), .ZN(n13506) );
  AOI21_X1 U8652 ( .B1(n6614), .B2(n13367), .A(n13366), .ZN(n13522) );
  AND2_X1 U8653 ( .A1(n9352), .A2(n9351), .ZN(n13552) );
  AND2_X1 U8654 ( .A1(n9328), .A2(n9327), .ZN(n13578) );
  AND2_X1 U8655 ( .A1(n9298), .A2(n9297), .ZN(n13604) );
  NAND2_X1 U8656 ( .A1(n7268), .A2(n7269), .ZN(n13646) );
  INV_X1 U8657 ( .A(n13781), .ZN(n13644) );
  NAND2_X1 U8658 ( .A1(n7272), .A2(n7273), .ZN(n13387) );
  OR2_X1 U8659 ( .A1(n11564), .A2(n11563), .ZN(n7272) );
  INV_X1 U8660 ( .A(n14631), .ZN(n11540) );
  NAND2_X1 U8661 ( .A1(n15210), .A2(n12334), .ZN(n13641) );
  OAI21_X1 U8662 ( .B1(n10762), .B2(n7228), .A(n7226), .ZN(n10983) );
  NAND2_X1 U8663 ( .A1(n10780), .A2(n10779), .ZN(n10781) );
  OR2_X1 U8664 ( .A1(n9898), .A2(n9038), .ZN(n9105) );
  NAND2_X1 U8665 ( .A1(n10745), .A2(n10744), .ZN(n10746) );
  NAND2_X1 U8666 ( .A1(n9487), .A2(n14881), .ZN(n13651) );
  AND2_X1 U8667 ( .A1(n14922), .A2(n13666), .ZN(n6925) );
  INV_X1 U8668 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U8669 ( .A1(n9228), .A2(n9227), .ZN(n12157) );
  AND2_X1 U8670 ( .A1(n14915), .A2(n13666), .ZN(n6926) );
  AOI21_X2 U8671 ( .B1(n12217), .B2(n12249), .A(n6604), .ZN(n13755) );
  OR2_X1 U8672 ( .A1(n13675), .A2(n13734), .ZN(n6627) );
  INV_X1 U8673 ( .A(n13672), .ZN(n6848) );
  INV_X1 U8674 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6634) );
  INV_X1 U8675 ( .A(n13390), .ZN(n13775) );
  NAND2_X2 U8676 ( .A1(n9171), .A2(n9170), .ZN(n13655) );
  AND2_X2 U8677 ( .A1(n10467), .A2(n10466), .ZN(n14915) );
  AND2_X1 U8678 ( .A1(n9504), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14881) );
  INV_X1 U8679 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8974) );
  INV_X1 U8680 ( .A(n8979), .ZN(n13788) );
  NAND2_X1 U8681 ( .A1(n6805), .A2(n6538), .ZN(n6619) );
  NAND2_X1 U8682 ( .A1(n9465), .A2(n9464), .ZN(n13799) );
  NAND2_X1 U8683 ( .A1(n9371), .A2(n9370), .ZN(n11747) );
  NAND2_X1 U8684 ( .A1(n8600), .A2(n7276), .ZN(n9371) );
  INV_X1 U8685 ( .A(n12283), .ZN(n12329) );
  INV_X1 U8686 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10836) );
  INV_X1 U8687 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n15113) );
  INV_X1 U8688 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10920) );
  INV_X1 U8689 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10638) );
  XNOR2_X1 U8690 ( .A(n9243), .B(n9242), .ZN(n11524) );
  INV_X1 U8691 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n15054) );
  INV_X1 U8692 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10109) );
  INV_X1 U8693 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10082) );
  INV_X1 U8694 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9897) );
  INV_X1 U8695 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9860) );
  INV_X1 U8696 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9895) );
  INV_X1 U8697 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9843) );
  AOI21_X1 U8698 ( .B1(n11070), .B2(n11069), .A(n7201), .ZN(n11188) );
  INV_X1 U8699 ( .A(n14640), .ZN(n6608) );
  NAND2_X1 U8700 ( .A1(n6593), .A2(n11651), .ZN(n11652) );
  NAND2_X1 U8701 ( .A1(n7184), .A2(n7185), .ZN(n13913) );
  AND2_X1 U8702 ( .A1(n7186), .A2(n13820), .ZN(n7185) );
  NAND2_X1 U8703 ( .A1(n7196), .A2(n7197), .ZN(n11426) );
  INV_X1 U8704 ( .A(n9758), .ZN(n14650) );
  INV_X1 U8705 ( .A(n14036), .ZN(n11274) );
  NAND2_X1 U8706 ( .A1(n10962), .A2(n7173), .ZN(n10956) );
  NAND2_X1 U8707 ( .A1(n7177), .A2(n6536), .ZN(n7173) );
  INV_X1 U8708 ( .A(n10965), .ZN(n7176) );
  NAND2_X1 U8709 ( .A1(n7177), .A2(n6488), .ZN(n10964) );
  INV_X1 U8710 ( .A(n11448), .ZN(n10718) );
  NAND2_X1 U8711 ( .A1(n11652), .A2(n7170), .ZN(n11760) );
  INV_X1 U8712 ( .A(n14699), .ZN(n14655) );
  XNOR2_X1 U8713 ( .A(n7213), .B(n9750), .ZN(n14012) );
  NAND2_X1 U8714 ( .A1(n14639), .A2(n9746), .ZN(n7213) );
  AND2_X1 U8715 ( .A1(n10795), .A2(n9802), .ZN(n14704) );
  AND2_X1 U8716 ( .A1(n9772), .A2(n10031), .ZN(n14483) );
  AND4_X1 U8717 ( .A1(n8301), .A2(n8300), .A3(n8299), .A4(n8298), .ZN(n11656)
         );
  INV_X1 U8718 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10164) );
  INV_X1 U8719 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10166) );
  INV_X1 U8720 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10162) );
  NAND2_X1 U8721 ( .A1(n6952), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8185) );
  OR2_X1 U8722 ( .A1(n8689), .A2(n10796), .ZN(n8121) );
  OAI21_X1 U8723 ( .B1(n14079), .B2(n14075), .A(n10025), .ZN(n14090) );
  NOR2_X1 U8724 ( .A1(n10320), .A2(n10321), .ZN(n10479) );
  NAND2_X1 U8725 ( .A1(n8760), .A2(n8759), .ZN(n14392) );
  NAND2_X1 U8726 ( .A1(n8726), .A2(n8725), .ZN(n14210) );
  XNOR2_X1 U8727 ( .A(n12017), .B(n12016), .ZN(n14398) );
  NAND2_X1 U8728 ( .A1(n11982), .A2(n11981), .ZN(n11983) );
  AOI21_X1 U8729 ( .B1(n12042), .B2(n12043), .A(n14795), .ZN(n6693) );
  INV_X1 U8730 ( .A(n6791), .ZN(n14213) );
  INV_X1 U8731 ( .A(n6790), .ZN(n14229) );
  NAND2_X1 U8732 ( .A1(n14286), .A2(n11995), .ZN(n14269) );
  NAND2_X1 U8733 ( .A1(n14317), .A2(n11991), .ZN(n14305) );
  NAND2_X1 U8734 ( .A1(n7101), .A2(n7100), .ZN(n14319) );
  NAND2_X1 U8735 ( .A1(n6963), .A2(n6464), .ZN(n14315) );
  AND2_X1 U8736 ( .A1(n6963), .A2(n6496), .ZN(n14316) );
  OR2_X1 U8737 ( .A1(n14334), .A2(n14335), .ZN(n6963) );
  NAND2_X1 U8738 ( .A1(n7102), .A2(n7105), .ZN(n14336) );
  NAND2_X1 U8739 ( .A1(n14367), .A2(n7108), .ZN(n7102) );
  OAI21_X1 U8740 ( .B1(n14367), .B2(n7110), .A(n11988), .ZN(n14347) );
  NAND2_X1 U8741 ( .A1(n8461), .A2(n8460), .ZN(n14385) );
  NAND2_X1 U8742 ( .A1(n11965), .A2(n11964), .ZN(n14369) );
  NAND2_X1 U8743 ( .A1(n11801), .A2(n11789), .ZN(n11926) );
  AND2_X1 U8744 ( .A1(n11787), .A2(n11786), .ZN(n11802) );
  NAND2_X1 U8745 ( .A1(n11581), .A2(n11580), .ZN(n11582) );
  OAI21_X1 U8746 ( .B1(n11356), .B2(n7099), .A(n7097), .ZN(n11672) );
  NAND2_X1 U8747 ( .A1(n11342), .A2(n6970), .ZN(n11480) );
  OAI21_X1 U8748 ( .B1(n11262), .B2(n11146), .A(n6782), .ZN(n11241) );
  NAND2_X1 U8749 ( .A1(n11161), .A2(n11164), .ZN(n11163) );
  NAND2_X1 U8750 ( .A1(n11262), .A2(n11135), .ZN(n11161) );
  INV_X1 U8751 ( .A(n14384), .ZN(n14364) );
  INV_X1 U8752 ( .A(n14357), .ZN(n14387) );
  AND2_X1 U8753 ( .A1(n14377), .A2(n11239), .ZN(n14357) );
  NAND2_X1 U8754 ( .A1(n14262), .A2(n10805), .ZN(n14337) );
  NAND2_X1 U8755 ( .A1(n9796), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9905) );
  AND2_X1 U8756 ( .A1(n6512), .A2(n8067), .ZN(n6972) );
  NAND2_X1 U8757 ( .A1(n6870), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8080) );
  AND2_X1 U8758 ( .A1(n8062), .A2(n7206), .ZN(n6869) );
  NAND2_X1 U8759 ( .A1(n8600), .A2(n7274), .ZN(n8619) );
  OR2_X1 U8760 ( .A1(n7250), .A2(n7251), .ZN(n8553) );
  INV_X1 U8761 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8083) );
  NAND2_X1 U8762 ( .A1(n8082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8084) );
  INV_X1 U8763 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n15074) );
  NAND2_X1 U8764 ( .A1(n7259), .A2(n8520), .ZN(n8521) );
  INV_X1 U8765 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10652) );
  INV_X1 U8766 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10918) );
  INV_X1 U8767 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n15067) );
  XNOR2_X1 U8768 ( .A(n8414), .B(n8413), .ZN(n11207) );
  INV_X1 U8769 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10107) );
  INV_X1 U8770 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10080) );
  INV_X1 U8771 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10013) );
  INV_X1 U8772 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9987) );
  OR2_X1 U8773 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  INV_X1 U8774 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9899) );
  INV_X1 U8775 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9852) );
  AND2_X1 U8776 ( .A1(n7123), .A2(n6566), .ZN(n15214) );
  OR2_X1 U8777 ( .A1(n15221), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n7123) );
  XNOR2_X1 U8778 ( .A(n9574), .B(n7132), .ZN(n14548) );
  INV_X1 U8779 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7132) );
  XNOR2_X1 U8780 ( .A(n9579), .B(n7130), .ZN(n15219) );
  XNOR2_X1 U8781 ( .A(n9582), .B(n9583), .ZN(n14549) );
  XNOR2_X1 U8782 ( .A(n9586), .B(n7129), .ZN(n14550) );
  INV_X1 U8783 ( .A(n9587), .ZN(n7129) );
  XNOR2_X1 U8784 ( .A(n9590), .B(n7142), .ZN(n14551) );
  INV_X1 U8785 ( .A(n9591), .ZN(n7142) );
  XNOR2_X1 U8786 ( .A(n9594), .B(n7140), .ZN(n14677) );
  INV_X1 U8787 ( .A(n9593), .ZN(n7140) );
  OAI21_X1 U8788 ( .B1(n7133), .B2(n7134), .A(n6466), .ZN(n14553) );
  NAND2_X1 U8789 ( .A1(n7139), .A2(n7135), .ZN(n7134) );
  INV_X1 U8790 ( .A(n7138), .ZN(n7133) );
  NAND2_X1 U8791 ( .A1(n10579), .A2(n8845), .ZN(n10614) );
  OR2_X1 U8792 ( .A1(n12692), .A2(n12691), .ZN(n6680) );
  INV_X1 U8793 ( .A(n6689), .ZN(n14962) );
  NOR2_X1 U8794 ( .A1(n12797), .A2(n12796), .ZN(n6717) );
  NAND2_X1 U8795 ( .A1(n6669), .A2(n6478), .ZN(n12843) );
  OR2_X1 U8796 ( .A1(n12829), .A2(n13043), .ZN(n9647) );
  NOR2_X1 U8797 ( .A1(n6588), .A2(n6725), .ZN(n6724) );
  NOR2_X1 U8798 ( .A1(n15051), .A2(n8047), .ZN(n6725) );
  OR2_X1 U8799 ( .A1(n12829), .A2(n13125), .ZN(n9651) );
  NOR2_X1 U8800 ( .A1(n6589), .A2(n6722), .ZN(n6721) );
  NOR2_X1 U8801 ( .A1(n15039), .A2(n8032), .ZN(n6722) );
  NAND2_X1 U8802 ( .A1(n9486), .A2(n9485), .ZN(n9513) );
  OAI21_X1 U8803 ( .B1(n13759), .B2(n13258), .A(n9510), .ZN(n9511) );
  OAI21_X1 U8804 ( .B1(n13213), .B2(n6770), .A(n6768), .ZN(P2_U3201) );
  INV_X1 U8805 ( .A(n6769), .ZN(n6768) );
  NAND2_X1 U8806 ( .A1(n6771), .A2(n9485), .ZN(n6770) );
  OAI21_X1 U8807 ( .B1(n13500), .B2(n13258), .A(n13221), .ZN(n6769) );
  AND2_X1 U8808 ( .A1(n12344), .A2(n7430), .ZN(n7429) );
  AOI21_X1 U8809 ( .B1(n13327), .B2(n14865), .A(n6752), .ZN(n13331) );
  OAI211_X1 U8810 ( .C1(n13670), .C2(n13649), .A(n7254), .B(n7253), .ZN(
        P2_U3236) );
  NAND2_X1 U8811 ( .A1(n7255), .A2(n13656), .ZN(n7254) );
  AOI21_X1 U8812 ( .B1(n6522), .B2(n13658), .A(n13415), .ZN(n7253) );
  OR2_X1 U8813 ( .A1(n14922), .A2(n7035), .ZN(n7034) );
  NAND2_X1 U8814 ( .A1(n13756), .A2(n14922), .ZN(n7036) );
  INV_X1 U8815 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7035) );
  NAND2_X1 U8816 ( .A1(n6639), .A2(n6636), .ZN(P2_U3526) );
  AOI21_X1 U8817 ( .B1(n13446), .B2(n13742), .A(n6637), .ZN(n6636) );
  NOR2_X1 U8818 ( .A1(n14922), .A2(n6638), .ZN(n6637) );
  OR2_X1 U8819 ( .A1(n14915), .A2(n6728), .ZN(n6727) );
  INV_X1 U8820 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U8821 ( .A1(n6635), .A2(n6537), .ZN(P2_U3494) );
  NAND2_X1 U8822 ( .A1(n13758), .A2(n14915), .ZN(n6635) );
  OR2_X1 U8823 ( .A1(n14915), .A2(n6634), .ZN(n6633) );
  XNOR2_X1 U8824 ( .A(n7162), .B(n13928), .ZN(n13935) );
  OR4_X1 U8825 ( .A1(n9806), .A2(n9805), .A3(n9804), .A4(n9803), .ZN(P1_U3238)
         );
  AOI21_X1 U8826 ( .B1(n6655), .B2(n11239), .A(n6654), .ZN(n6653) );
  OR2_X1 U8827 ( .A1(n14196), .A2(n11239), .ZN(n6656) );
  OAI21_X1 U8828 ( .B1(n14199), .B2(n14200), .A(n14198), .ZN(n6654) );
  NAND2_X1 U8829 ( .A1(n14811), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6859) );
  OAI21_X1 U8830 ( .B1(n6974), .B2(n6861), .A(n14813), .ZN(n6860) );
  NOR2_X1 U8831 ( .A1(n14405), .A2(n14795), .ZN(n6861) );
  INV_X1 U8832 ( .A(n14405), .ZN(n6660) );
  NOR2_X1 U8833 ( .A1(n6463), .A2(n14680), .ZN(n14679) );
  OAI21_X1 U8834 ( .B1(n6463), .B2(n7155), .A(n7152), .ZN(n14683) );
  INV_X1 U8835 ( .A(n7137), .ZN(n14691) );
  XNOR2_X1 U8836 ( .A(n7144), .B(n7143), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8837 ( .A(n9623), .B(n6607), .ZN(n7143) );
  OAI21_X1 U8838 ( .B1(n14540), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6515), .ZN(
        n7144) );
  INV_X1 U8839 ( .A(n14333), .ZN(n14335) );
  BUF_X1 U8840 ( .A(n12072), .Z(n12228) );
  INV_X1 U8841 ( .A(n9675), .ZN(n9684) );
  AND2_X1 U8842 ( .A1(n13183), .A2(n7323), .ZN(n7322) );
  AND2_X2 U8843 ( .A1(n6671), .A2(n6516), .ZN(n6463) );
  AND2_X1 U8844 ( .A1(n14320), .A2(n6496), .ZN(n6464) );
  NOR2_X1 U8845 ( .A1(n8591), .A2(n8588), .ZN(n6465) );
  NAND2_X1 U8846 ( .A1(n14690), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n6466) );
  INV_X1 U8847 ( .A(n13681), .ZN(n13411) );
  AND2_X1 U8848 ( .A1(n12180), .A2(n7419), .ZN(n6467) );
  AND2_X1 U8849 ( .A1(n13645), .A2(n13352), .ZN(n6468) );
  AND2_X1 U8850 ( .A1(n12208), .A2(n7390), .ZN(n6469) );
  AND2_X1 U8851 ( .A1(n6821), .A2(n6524), .ZN(n6470) );
  INV_X1 U8852 ( .A(n11180), .ZN(n6811) );
  AND2_X1 U8853 ( .A1(n7258), .A2(n6843), .ZN(n6471) );
  INV_X1 U8854 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U8855 ( .A1(n15097), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6472) );
  AND2_X1 U8856 ( .A1(n13781), .A2(n13389), .ZN(n6473) );
  AND2_X1 U8857 ( .A1(n6803), .A2(n9326), .ZN(n6474) );
  AND2_X1 U8858 ( .A1(n6821), .A2(n7324), .ZN(n6475) );
  AND2_X1 U8859 ( .A1(n8064), .A2(n7208), .ZN(n6476) );
  NAND2_X1 U8860 ( .A1(n12207), .A2(n12209), .ZN(n6477) );
  INV_X1 U8861 ( .A(n12991), .ZN(n7077) );
  OR2_X1 U8862 ( .A1(n15002), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8863 ( .A1(n7335), .A2(n12334), .ZN(n10088) );
  NOR2_X1 U8864 ( .A1(n14522), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6479) );
  OR2_X1 U8865 ( .A1(n14915), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6480) );
  INV_X1 U8866 ( .A(n9045), .ZN(n12220) );
  INV_X1 U8867 ( .A(n9680), .ZN(n13920) );
  INV_X1 U8868 ( .A(n14932), .ZN(n6931) );
  INV_X1 U8869 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7485) );
  NAND2_X1 U8870 ( .A1(n13957), .A2(n13958), .ZN(n9766) );
  NAND2_X1 U8871 ( .A1(n12234), .A2(n12233), .ZN(n13335) );
  NAND2_X1 U8872 ( .A1(n10555), .A2(n14932), .ZN(n6482) );
  NAND2_X1 U8873 ( .A1(n8520), .A2(n7260), .ZN(n8537) );
  INV_X1 U8874 ( .A(n7491), .ZN(n12688) );
  NAND2_X1 U8875 ( .A1(n7649), .A2(n7648), .ZN(n7652) );
  INV_X1 U8876 ( .A(n8179), .ZN(n6952) );
  INV_X1 U8877 ( .A(n13414), .ZN(n13375) );
  OR2_X1 U8878 ( .A1(n14271), .A2(n14251), .ZN(n6483) );
  OR2_X1 U8879 ( .A1(n12130), .A2(n12131), .ZN(n6484) );
  AND2_X1 U8880 ( .A1(n9178), .A2(n9166), .ZN(n6485) );
  INV_X1 U8881 ( .A(n11146), .ZN(n11164) );
  AND2_X1 U8882 ( .A1(n8770), .A2(n11148), .ZN(n11146) );
  AND2_X1 U8883 ( .A1(n6763), .A2(n15023), .ZN(n6486) );
  AND2_X1 U8884 ( .A1(n7360), .A2(n9644), .ZN(n6487) );
  INV_X1 U8885 ( .A(n9695), .ZN(n7181) );
  OR2_X1 U8886 ( .A1(n7182), .A2(n9695), .ZN(n6488) );
  AND2_X1 U8887 ( .A1(n12181), .A2(n7420), .ZN(n6489) );
  AND2_X1 U8888 ( .A1(n14356), .A2(n14484), .ZN(n6490) );
  NAND2_X1 U8889 ( .A1(n14265), .A2(n14270), .ZN(n14264) );
  NAND2_X1 U8890 ( .A1(n7007), .A2(n7004), .ZN(n6491) );
  OR2_X1 U8891 ( .A1(n8821), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n6492) );
  NOR2_X1 U8892 ( .A1(n9625), .A2(n12349), .ZN(n6493) );
  OR2_X1 U8893 ( .A1(n12132), .A2(n13288), .ZN(n6494) );
  XNOR2_X1 U8894 ( .A(n14225), .B(n14025), .ZN(n14217) );
  INV_X1 U8895 ( .A(n14217), .ZN(n7112) );
  AND2_X1 U8896 ( .A1(n12000), .A2(n14276), .ZN(n6495) );
  NAND2_X1 U8897 ( .A1(n14470), .A2(n14475), .ZN(n6496) );
  OR2_X1 U8898 ( .A1(n14418), .A2(n13952), .ZN(n6497) );
  INV_X1 U8899 ( .A(n14663), .ZN(n14016) );
  XNOR2_X1 U8900 ( .A(n7998), .B(n7997), .ZN(n11592) );
  NAND2_X1 U8901 ( .A1(n12235), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6498) );
  NOR2_X1 U8902 ( .A1(n14259), .A2(n6495), .ZN(n6499) );
  NOR2_X1 U8903 ( .A1(n11968), .A2(n6967), .ZN(n6501) );
  NAND2_X1 U8904 ( .A1(n8482), .A2(n8481), .ZN(n14654) );
  AND2_X1 U8905 ( .A1(n13335), .A2(n14889), .ZN(n6502) );
  OR2_X1 U8906 ( .A1(n10909), .A2(n11330), .ZN(n6503) );
  AND2_X1 U8907 ( .A1(n12699), .A2(n12574), .ZN(n6504) );
  AND2_X1 U8908 ( .A1(n9750), .A2(n14011), .ZN(n6505) );
  NAND2_X1 U8909 ( .A1(n8627), .A2(n8626), .ZN(n14251) );
  OR2_X1 U8910 ( .A1(n12737), .A2(n12718), .ZN(n6506) );
  XNOR2_X1 U8911 ( .A(n8724), .B(n8723), .ZN(n12217) );
  AND2_X1 U8912 ( .A1(n10909), .A2(n11330), .ZN(n6507) );
  OR2_X1 U8913 ( .A1(n14402), .A2(n6862), .ZN(n6508) );
  OR2_X1 U8914 ( .A1(n8479), .A2(n8141), .ZN(n8815) );
  INV_X1 U8915 ( .A(n12512), .ZN(n12891) );
  OR2_X1 U8916 ( .A1(n11695), .A2(n11696), .ZN(n6509) );
  NAND2_X1 U8917 ( .A1(n13060), .A2(n12871), .ZN(n6510) );
  INV_X1 U8918 ( .A(n8667), .ZN(n6988) );
  NAND2_X1 U8919 ( .A1(n13828), .A2(n13827), .ZN(n13936) );
  OR2_X1 U8920 ( .A1(n9583), .A2(n9582), .ZN(n6511) );
  AND2_X1 U8921 ( .A1(n7206), .A2(n8079), .ZN(n6512) );
  AND2_X1 U8922 ( .A1(n6832), .A2(n6831), .ZN(n6513) );
  INV_X1 U8923 ( .A(n8333), .ZN(n7006) );
  AND3_X1 U8924 ( .A1(n12548), .A2(n12547), .A3(n12546), .ZN(n6514) );
  OR2_X1 U8925 ( .A1(n9618), .A2(n9617), .ZN(n6515) );
  NAND2_X1 U8926 ( .A1(n8557), .A2(n8556), .ZN(n8585) );
  NAND2_X1 U8927 ( .A1(n8351), .A2(n8350), .ZN(n11768) );
  OR2_X1 U8928 ( .A1(n9598), .A2(n9597), .ZN(n6516) );
  OR2_X1 U8929 ( .A1(n13367), .A2(n13366), .ZN(n6517) );
  AND2_X1 U8930 ( .A1(n14620), .A2(n13388), .ZN(n6518) );
  AND2_X1 U8931 ( .A1(n13478), .A2(n13409), .ZN(n6519) );
  AND2_X1 U8932 ( .A1(n7074), .A2(n7967), .ZN(n6520) );
  AND2_X1 U8933 ( .A1(n8544), .A2(n8543), .ZN(n14322) );
  AND2_X1 U8934 ( .A1(n8862), .A2(n12359), .ZN(n6521) );
  NOR2_X1 U8935 ( .A1(n13382), .A2(n6927), .ZN(n6522) );
  OR2_X1 U8936 ( .A1(n9948), .A2(n9884), .ZN(n6523) );
  INV_X1 U8937 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8345) );
  NOR2_X1 U8938 ( .A1(n9444), .A2(n6825), .ZN(n6524) );
  AND2_X1 U8939 ( .A1(n8091), .A2(n8139), .ZN(n9655) );
  NAND2_X1 U8940 ( .A1(n7412), .A2(n12197), .ZN(n7410) );
  INV_X1 U8941 ( .A(n7410), .ZN(n7405) );
  INV_X1 U8942 ( .A(n8606), .ZN(n6996) );
  OR2_X1 U8943 ( .A1(n8113), .A2(n14057), .ZN(n6525) );
  INV_X1 U8944 ( .A(n6944), .ZN(n6941) );
  AND2_X1 U8945 ( .A1(n12952), .A2(n12615), .ZN(n6526) );
  NAND2_X1 U8946 ( .A1(n8081), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8143) );
  AND2_X1 U8947 ( .A1(n12915), .A2(n12634), .ZN(n6527) );
  AND2_X1 U8948 ( .A1(n13417), .A2(n13418), .ZN(n6528) );
  OR2_X1 U8949 ( .A1(n13298), .A2(n10772), .ZN(n6529) );
  AND2_X1 U8950 ( .A1(n13593), .A2(n13396), .ZN(n6530) );
  AND2_X1 U8951 ( .A1(n9362), .A2(n9350), .ZN(n6531) );
  AND2_X1 U8952 ( .A1(n8852), .A2(n8850), .ZN(n6532) );
  AND2_X1 U8953 ( .A1(n7970), .A2(n7969), .ZN(n6533) );
  AND2_X1 U8954 ( .A1(n7299), .A2(n8859), .ZN(n6534) );
  NAND2_X1 U8955 ( .A1(n12186), .A2(n12185), .ZN(n6535) );
  AND2_X1 U8956 ( .A1(n6488), .A2(n7176), .ZN(n6536) );
  AND2_X1 U8957 ( .A1(n6640), .A2(n6633), .ZN(n6537) );
  AND2_X1 U8958 ( .A1(n6806), .A2(n6808), .ZN(n6538) );
  INV_X1 U8959 ( .A(n13352), .ZN(n7050) );
  INV_X1 U8960 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8079) );
  OR2_X1 U8961 ( .A1(n8892), .A2(n8891), .ZN(n6539) );
  AND2_X1 U8962 ( .A1(n14322), .A2(n14027), .ZN(n6540) );
  AND3_X1 U8963 ( .A1(n9101), .A2(n8960), .A3(n9135), .ZN(n8998) );
  INV_X1 U8964 ( .A(n7322), .ZN(n7321) );
  AND2_X1 U8965 ( .A1(n7070), .A2(n7069), .ZN(n6541) );
  NOR2_X1 U8966 ( .A1(n14470), .A2(n14361), .ZN(n6542) );
  NOR2_X1 U8967 ( .A1(n11768), .A2(n14033), .ZN(n6543) );
  NOR2_X1 U8968 ( .A1(n11768), .A2(n11872), .ZN(n6544) );
  NOR2_X1 U8969 ( .A1(n13655), .A2(n11366), .ZN(n6545) );
  NOR2_X1 U8970 ( .A1(n11621), .A2(n11343), .ZN(n6546) );
  INV_X1 U8971 ( .A(n6836), .ZN(n6835) );
  AND2_X1 U8972 ( .A1(n7231), .A2(n6837), .ZN(n6836) );
  MUX2_X1 U8973 ( .A(n14022), .B(n14404), .S(n8795), .Z(n8716) );
  INV_X1 U8974 ( .A(n8716), .ZN(n7018) );
  AND2_X1 U8975 ( .A1(n11175), .A2(n11274), .ZN(n6547) );
  INV_X1 U8976 ( .A(n7257), .ZN(n7256) );
  NOR2_X1 U8977 ( .A1(n8535), .A2(SI_19_), .ZN(n7257) );
  AND2_X1 U8978 ( .A1(n13071), .A2(n12892), .ZN(n6548) );
  OR2_X1 U8979 ( .A1(n7111), .A2(n6787), .ZN(n6549) );
  INV_X1 U8980 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7472) );
  AND2_X1 U8981 ( .A1(n12309), .A2(n6494), .ZN(n7043) );
  AND2_X1 U8982 ( .A1(n6997), .A2(n6996), .ZN(n6550) );
  INV_X1 U8983 ( .A(n7115), .ZN(n6789) );
  AND2_X1 U8984 ( .A1(n14425), .A2(n14255), .ZN(n7115) );
  AND2_X1 U8985 ( .A1(n8899), .A2(n8900), .ZN(n6551) );
  AND2_X1 U8986 ( .A1(n10364), .A2(n9082), .ZN(n6552) );
  AND2_X1 U8987 ( .A1(n8406), .A2(n9964), .ZN(n6553) );
  AND2_X1 U8988 ( .A1(n13895), .A2(n14005), .ZN(n6554) );
  INV_X1 U8989 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9850) );
  OR2_X1 U8990 ( .A1(n9515), .A2(n15098), .ZN(n6555) );
  NOR2_X1 U8991 ( .A1(n8766), .A2(n8795), .ZN(n6556) );
  INV_X1 U8992 ( .A(n7379), .ZN(n7378) );
  NAND2_X1 U8993 ( .A1(n12636), .A2(n7380), .ZN(n7379) );
  AND2_X1 U8994 ( .A1(n8293), .A2(n11352), .ZN(n6557) );
  INV_X1 U8995 ( .A(n7265), .ZN(n7264) );
  NAND2_X1 U8996 ( .A1(n13395), .A2(n7266), .ZN(n7265) );
  OR2_X1 U8997 ( .A1(n7355), .A2(n12520), .ZN(n6558) );
  OAI21_X1 U8998 ( .B1(n13329), .B2(n13328), .A(n14820), .ZN(n6752) );
  INV_X1 U8999 ( .A(n9183), .ZN(n6815) );
  NAND2_X1 U9000 ( .A1(n7325), .A2(n7320), .ZN(n6559) );
  INV_X1 U9001 ( .A(n7416), .ZN(n7415) );
  NAND2_X1 U9002 ( .A1(n7417), .A2(n12182), .ZN(n7416) );
  NAND2_X1 U9003 ( .A1(n8450), .A2(n8449), .ZN(n6560) );
  AND2_X1 U9004 ( .A1(n10240), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6561) );
  NOR2_X1 U9005 ( .A1(n7018), .A2(n8717), .ZN(n6562) );
  AND2_X1 U9006 ( .A1(n12216), .A2(n6477), .ZN(n6563) );
  INV_X1 U9007 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6809) );
  INV_X1 U9008 ( .A(n14685), .ZN(n7158) );
  AND2_X1 U9009 ( .A1(n7127), .A2(n6472), .ZN(n6564) );
  OR2_X1 U9010 ( .A1(n9709), .A2(n9710), .ZN(n6565) );
  OR2_X1 U9011 ( .A1(n9566), .A2(n9565), .ZN(n6566) );
  AND2_X1 U9012 ( .A1(n7100), .A2(n11990), .ZN(n6567) );
  AND2_X1 U9013 ( .A1(n6781), .A2(n11240), .ZN(n6568) );
  AND2_X1 U9014 ( .A1(n10744), .A2(n10420), .ZN(n6569) );
  AND2_X1 U9015 ( .A1(n6851), .A2(n11924), .ZN(n6570) );
  AND2_X1 U9016 ( .A1(n11749), .A2(n7285), .ZN(n6571) );
  NOR2_X1 U9017 ( .A1(n7001), .A2(n6999), .ZN(n6572) );
  AND2_X1 U9018 ( .A1(n7267), .A2(n7269), .ZN(n6573) );
  AND2_X1 U9019 ( .A1(n12616), .A2(n12622), .ZN(n12952) );
  INV_X1 U9020 ( .A(n8204), .ZN(n7218) );
  NAND2_X1 U9021 ( .A1(n6850), .A2(SI_4_), .ZN(n8204) );
  OR2_X1 U9022 ( .A1(n8355), .A2(n8353), .ZN(n6574) );
  AND2_X1 U9023 ( .A1(n10910), .A2(n10909), .ZN(n6575) );
  OR2_X1 U9024 ( .A1(n11867), .A2(n11868), .ZN(n7169) );
  OR2_X1 U9025 ( .A1(n8219), .A2(n8217), .ZN(n6576) );
  AND2_X1 U9026 ( .A1(n7383), .A2(n7386), .ZN(n6577) );
  OR2_X1 U9027 ( .A1(n8666), .A2(n6988), .ZN(n6578) );
  AND2_X1 U9028 ( .A1(n7137), .A2(n7136), .ZN(n6579) );
  NAND2_X1 U9029 ( .A1(n14058), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6580) );
  AND2_X1 U9030 ( .A1(n6979), .A2(n6980), .ZN(n6581) );
  NAND2_X1 U9031 ( .A1(n12139), .A2(n12138), .ZN(n6582) );
  NAND2_X1 U9032 ( .A1(n12166), .A2(n12165), .ZN(n6583) );
  AND2_X1 U9033 ( .A1(n6847), .A2(n6846), .ZN(n6584) );
  INV_X1 U9034 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n6644) );
  OR2_X1 U9035 ( .A1(n7415), .A2(n6489), .ZN(n6585) );
  INV_X1 U9036 ( .A(n7324), .ZN(n6825) );
  OR2_X1 U9037 ( .A1(n9431), .A2(n9432), .ZN(n7324) );
  INV_X1 U9038 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7011) );
  INV_X1 U9039 ( .A(n7203), .ZN(n7201) );
  NAND2_X1 U9040 ( .A1(n9705), .A2(n9706), .ZN(n7203) );
  INV_X1 U9041 ( .A(n10243), .ZN(n6715) );
  INV_X1 U9042 ( .A(SI_18_), .ZN(n10269) );
  NAND2_X1 U9043 ( .A1(n6609), .A2(n6608), .ZN(n14639) );
  INV_X1 U9044 ( .A(n13493), .ZN(n6631) );
  AND2_X1 U9045 ( .A1(n14352), .A2(n6868), .ZN(n6586) );
  NAND2_X1 U9046 ( .A1(n11740), .A2(n6853), .ZN(n6587) );
  INV_X1 U9047 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8100) );
  AND2_X1 U9048 ( .A1(n12662), .A2(n8048), .ZN(n6588) );
  INV_X1 U9049 ( .A(n12611), .ZN(n7340) );
  AND2_X1 U9050 ( .A1(n12662), .A2(n13121), .ZN(n6589) );
  AND2_X1 U9051 ( .A1(n11652), .A2(n7167), .ZN(n6590) );
  NAND2_X1 U9052 ( .A1(n8985), .A2(n8984), .ZN(n13472) );
  INV_X1 U9053 ( .A(n12190), .ZN(n7395) );
  AND2_X1 U9054 ( .A1(n7040), .A2(n7041), .ZN(n6591) );
  AND2_X1 U9055 ( .A1(n7782), .A2(n12615), .ZN(n6592) );
  AND2_X1 U9056 ( .A1(n11650), .A2(n11653), .ZN(n6593) );
  AND2_X1 U9057 ( .A1(n7044), .A2(n6494), .ZN(n6594) );
  NAND2_X1 U9058 ( .A1(n9766), .A2(n13959), .ZN(n13961) );
  OR2_X1 U9059 ( .A1(n8617), .A2(n11106), .ZN(n6595) );
  AND2_X1 U9060 ( .A1(n7708), .A2(n7707), .ZN(n14602) );
  INV_X1 U9061 ( .A(n14602), .ZN(n11821) );
  OR2_X1 U9062 ( .A1(n8618), .A2(SI_23_), .ZN(n6596) );
  AND2_X1 U9063 ( .A1(n7450), .A2(n7304), .ZN(n6597) );
  INV_X1 U9064 ( .A(n13627), .ZN(n13656) );
  INV_X1 U9065 ( .A(n12311), .ZN(n7046) );
  NAND2_X1 U9066 ( .A1(n10382), .A2(n9080), .ZN(n10362) );
  NOR2_X1 U9067 ( .A1(n10822), .A2(n7333), .ZN(n7332) );
  AND2_X1 U9068 ( .A1(n11484), .A2(n6858), .ZN(n6598) );
  NAND2_X1 U9069 ( .A1(n8560), .A2(n8559), .ZN(n14455) );
  INV_X1 U9070 ( .A(n14455), .ZN(n6865) );
  AND2_X1 U9071 ( .A1(n9202), .A2(n9201), .ZN(n6599) );
  INV_X1 U9072 ( .A(n6701), .ZN(n11287) );
  AND2_X1 U9073 ( .A1(n7196), .A2(n7194), .ZN(n6600) );
  AND2_X1 U9074 ( .A1(n7327), .A2(n7326), .ZN(n6601) );
  AND2_X1 U9075 ( .A1(n6876), .A2(n6482), .ZN(n6602) );
  AND2_X1 U9076 ( .A1(n11748), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6603) );
  AND3_X1 U9077 ( .A1(n8969), .A2(n8968), .A3(n8967), .ZN(n9479) );
  INV_X1 U9078 ( .A(n13780), .ZN(n6641) );
  OR2_X1 U9079 ( .A1(n10717), .A2(n10345), .ZN(n14811) );
  INV_X1 U9080 ( .A(n10363), .ZN(n7331) );
  INV_X2 U9081 ( .A(n14800), .ZN(n14802) );
  OR2_X1 U9082 ( .A1(n10717), .A2(n10793), .ZN(n14800) );
  NAND2_X1 U9083 ( .A1(n8373), .A2(n8372), .ZN(n11889) );
  INV_X1 U9084 ( .A(n11889), .ZN(n6855) );
  INV_X1 U9085 ( .A(n13749), .ZN(n13742) );
  AND2_X1 U9086 ( .A1(n10338), .A2(n10337), .ZN(n14795) );
  INV_X1 U9087 ( .A(n14795), .ZN(n14489) );
  AND2_X1 U9088 ( .A1(n12251), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6604) );
  INV_X1 U9089 ( .A(n12737), .ZN(n14559) );
  AND4_X2 U9090 ( .A1(n8045), .A2(n8044), .A3(n10353), .A4(n8043), .ZN(n15051)
         );
  INV_X1 U9091 ( .A(n12785), .ZN(n12778) );
  INV_X2 U9092 ( .A(n15037), .ZN(n15039) );
  INV_X1 U9093 ( .A(n13655), .ZN(n6700) );
  NAND2_X1 U9094 ( .A1(n10457), .A2(n12087), .ZN(n10458) );
  INV_X1 U9095 ( .A(n10458), .ZN(n6921) );
  AND2_X1 U9096 ( .A1(n9628), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6605) );
  AND2_X1 U9097 ( .A1(n14800), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6606) );
  NOR2_X1 U9098 ( .A1(n9626), .A2(n6915), .ZN(n6914) );
  INV_X1 U9099 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6955) );
  INV_X1 U9100 ( .A(n11239), .ZN(n14195) );
  NOR2_X1 U9101 ( .A1(n11836), .A2(P2_U3088), .ZN(n12339) );
  XOR2_X1 U9102 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n6607) );
  INV_X1 U9103 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7124) );
  INV_X1 U9104 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7130) );
  NAND2_X1 U9105 ( .A1(n13052), .A2(n15002), .ZN(n6669) );
  AND2_X2 U9106 ( .A1(n10355), .A2(n14580), .ZN(n15004) );
  INV_X1 U9107 ( .A(n9671), .ZN(n9797) );
  OAI21_X2 U9108 ( .B1(n14639), .B2(n7211), .A(n7209), .ZN(n9758) );
  INV_X1 U9109 ( .A(n14641), .ZN(n6609) );
  NOR2_X1 U9110 ( .A1(n7088), .A2(n7085), .ZN(n7084) );
  AND4_X2 U9111 ( .A1(n7502), .A2(n7504), .A3(n7505), .A4(n7503), .ZN(n6650)
         );
  INV_X1 U9112 ( .A(n11692), .ZN(n6611) );
  NOR2_X1 U9113 ( .A1(n14929), .A2(n14928), .ZN(n14927) );
  NOR2_X1 U9114 ( .A1(n11307), .A2(n11308), .ZN(n14943) );
  NOR2_X1 U9115 ( .A1(n10911), .A2(n11397), .ZN(n11307) );
  NOR2_X1 U9116 ( .A1(n14943), .A2(n14942), .ZN(n14941) );
  XNOR2_X1 U9117 ( .A(n11412), .B(n11413), .ZN(n11310) );
  AOI21_X2 U9118 ( .B1(n6976), .B2(n14795), .A(n14800), .ZN(n6975) );
  NAND2_X1 U9119 ( .A1(n12003), .A2(n12002), .ZN(n12015) );
  NAND2_X1 U9120 ( .A1(n11290), .A2(n7043), .ZN(n7040) );
  NAND2_X1 U9121 ( .A1(n6775), .A2(n6774), .ZN(n10987) );
  NAND3_X1 U9122 ( .A1(n7014), .A2(n7015), .A3(n6615), .ZN(n8739) );
  NAND3_X1 U9123 ( .A1(n7013), .A2(n7222), .A3(n7221), .ZN(n6615) );
  OAI21_X1 U9124 ( .B1(n12547), .B2(n7372), .A(n12552), .ZN(n7371) );
  INV_X1 U9125 ( .A(n10402), .ZN(n14989) );
  AND2_X1 U9126 ( .A1(n7514), .A2(n7512), .ZN(n6616) );
  NAND2_X1 U9127 ( .A1(n7363), .A2(n7361), .ZN(n11399) );
  NAND2_X1 U9128 ( .A1(n14594), .A2(n12592), .ZN(n14584) );
  AND3_X2 U9129 ( .A1(n6616), .A2(n7513), .A3(n7511), .ZN(n10402) );
  NAND2_X1 U9130 ( .A1(n7341), .A2(n7339), .ZN(n12965) );
  NAND2_X1 U9131 ( .A1(n10886), .A2(n12553), .ZN(n10999) );
  NAND2_X1 U9132 ( .A1(n6617), .A2(n12582), .ZN(n14596) );
  NAND2_X1 U9133 ( .A1(n11497), .A2(n12580), .ZN(n6617) );
  NAND2_X1 U9134 ( .A1(n14584), .A2(n14583), .ZN(n14582) );
  NAND2_X1 U9135 ( .A1(n7370), .A2(n7367), .ZN(n10886) );
  OAI21_X1 U9136 ( .B1(n11815), .B2(n12594), .A(n12599), .ZN(n11934) );
  NAND2_X1 U9137 ( .A1(n11494), .A2(n12577), .ZN(n11493) );
  NAND2_X1 U9138 ( .A1(n10497), .A2(n7945), .ZN(n10628) );
  NAND2_X1 U9139 ( .A1(n7949), .A2(n7948), .ZN(n11004) );
  NAND2_X1 U9140 ( .A1(n11004), .A2(n7950), .ZN(n11024) );
  NAND2_X1 U9141 ( .A1(n11937), .A2(n7961), .ZN(n12989) );
  NAND2_X1 U9142 ( .A1(n6652), .A2(n7067), .ZN(n12939) );
  NAND2_X1 U9143 ( .A1(n7298), .A2(n7297), .ZN(n10579) );
  NAND2_X1 U9144 ( .A1(n11111), .A2(n8855), .ZN(n11053) );
  NAND2_X1 U9145 ( .A1(n11632), .A2(n12362), .ZN(n8869) );
  NAND2_X1 U9146 ( .A1(n12433), .A2(n8887), .ZN(n12389) );
  INV_X1 U9147 ( .A(n12037), .ZN(n7480) );
  OAI21_X1 U9148 ( .B1(n14401), .B2(n13925), .A(n12015), .ZN(n12017) );
  INV_X1 U9149 ( .A(n7113), .ZN(n7111) );
  OAI21_X1 U9150 ( .B1(n12101), .B2(n12100), .A(n12098), .ZN(n12099) );
  NAND2_X1 U9151 ( .A1(n7393), .A2(n7391), .ZN(n12194) );
  AOI21_X1 U9152 ( .B1(n6620), .B2(n6585), .A(n7413), .ZN(n12186) );
  AOI21_X1 U9153 ( .B1(n12114), .B2(n12113), .A(n12112), .ZN(n12120) );
  NAND2_X1 U9154 ( .A1(n12298), .A2(n10451), .ZN(n10450) );
  NAND4_X1 U9155 ( .A1(n9025), .A2(n9023), .A3(n9022), .A4(n9024), .ZN(n13296)
         );
  AOI21_X1 U9156 ( .B1(n7268), .B2(n6573), .A(n6473), .ZN(n13611) );
  AOI21_X1 U9157 ( .B1(n13554), .B2(n13540), .A(n13404), .ZN(n13534) );
  OAI22_X1 U9158 ( .A1(n13416), .A2(n13417), .B1(n13428), .B2(n13436), .ZN(
        n6690) );
  AOI22_X1 U9159 ( .A1(n12156), .A2(n12155), .B1(n12154), .B2(n12151), .ZN(
        n12162) );
  INV_X1 U9160 ( .A(n9295), .ZN(n6623) );
  NAND2_X1 U9161 ( .A1(n6623), .A2(n8988), .ZN(n9310) );
  OAI21_X1 U9162 ( .B1(n12194), .B2(n12192), .A(n12191), .ZN(n12196) );
  INV_X1 U9163 ( .A(n12171), .ZN(n6625) );
  OR2_X1 U9164 ( .A1(n12176), .A2(n12177), .ZN(n6620) );
  AOI21_X1 U9165 ( .B1(n12170), .B2(n12169), .A(n12168), .ZN(n12171) );
  OAI22_X1 U9166 ( .A1(n12105), .A2(n12228), .B1(n12104), .B2(n12276), .ZN(
        n12106) );
  NAND2_X1 U9167 ( .A1(n8205), .A2(n8204), .ZN(n8222) );
  INV_X1 U9168 ( .A(n12172), .ZN(n6624) );
  NAND2_X1 U9169 ( .A1(n7402), .A2(n7401), .ZN(n7400) );
  NAND2_X1 U9170 ( .A1(n6625), .A2(n6624), .ZN(n12175) );
  INV_X1 U9171 ( .A(n13671), .ZN(n7255) );
  NAND2_X1 U9172 ( .A1(n11564), .A2(n7270), .ZN(n7268) );
  NAND2_X1 U9173 ( .A1(n6630), .A2(n6629), .ZN(n11037) );
  NAND2_X1 U9174 ( .A1(n8105), .A2(n8106), .ZN(n8129) );
  INV_X1 U9175 ( .A(n7227), .ZN(n7226) );
  AOI22_X1 U9176 ( .A1(n13413), .A2(n13448), .B1(n13446), .B2(n13456), .ZN(
        n13416) );
  AND2_X1 U9177 ( .A1(n12060), .A2(n12061), .ZN(n6628) );
  AOI22_X1 U9178 ( .A1(n12080), .A2(n12079), .B1(n12083), .B2(n12084), .ZN(
        n12082) );
  NAND2_X1 U9179 ( .A1(n8638), .A2(n8621), .ZN(n8624) );
  NAND2_X1 U9180 ( .A1(n8552), .A2(n7251), .ZN(n8557) );
  OAI22_X1 U9181 ( .A1(n8650), .A2(n8649), .B1(SI_25_), .B2(n8648), .ZN(n8653)
         );
  NAND3_X1 U9182 ( .A1(n6627), .A2(n6848), .A3(n6584), .ZN(n13757) );
  NAND2_X1 U9183 ( .A1(n8159), .A2(n8158), .ZN(n8163) );
  NAND2_X1 U9184 ( .A1(n11286), .A2(n11285), .ZN(n11363) );
  INV_X1 U9185 ( .A(n10984), .ZN(n6630) );
  NAND2_X1 U9186 ( .A1(n8129), .A2(n8128), .ZN(n8135) );
  NAND2_X1 U9187 ( .A1(n6736), .A2(n8223), .ZN(n8227) );
  OAI21_X1 U9188 ( .B1(n11546), .B2(n11545), .A(n11547), .ZN(n11564) );
  NAND2_X1 U9189 ( .A1(n13534), .A2(n13535), .ZN(n13703) );
  NAND2_X1 U9190 ( .A1(n6628), .A2(n12062), .ZN(n12071) );
  NAND3_X1 U9191 ( .A1(n7225), .A2(n10982), .A3(n7224), .ZN(n10984) );
  NAND2_X1 U9192 ( .A1(n13402), .A2(n13401), .ZN(n13554) );
  NAND2_X1 U9193 ( .A1(n12127), .A2(n12126), .ZN(n6696) );
  NAND2_X1 U9194 ( .A1(n8456), .A2(n8455), .ZN(n8476) );
  AOI21_X1 U9195 ( .B1(n11207), .B2(n11904), .A(n11204), .ZN(n11839) );
  NOR2_X1 U9196 ( .A1(n10656), .A2(n10655), .ZN(n10850) );
  NAND2_X1 U9197 ( .A1(n6656), .A2(n6653), .ZN(P1_U3262) );
  XNOR2_X1 U9198 ( .A(n14181), .B(n14180), .ZN(n14189) );
  AOI21_X1 U9199 ( .B1(n14119), .B2(n10028), .A(n10027), .ZN(n10305) );
  NOR2_X1 U9200 ( .A1(n11841), .A2(n11840), .ZN(n14165) );
  NAND2_X1 U9201 ( .A1(n14106), .A2(n14107), .ZN(n14105) );
  AOI21_X1 U9202 ( .B1(n10308), .B2(n10309), .A(n14152), .ZN(n10312) );
  OAI211_X2 U9203 ( .C1(n9038), .C2(n9903), .A(n9021), .B(n6801), .ZN(n12076)
         );
  AND2_X2 U9204 ( .A1(n11370), .A2(n14908), .ZN(n11513) );
  AND2_X2 U9205 ( .A1(n6701), .A2(n6700), .ZN(n11370) );
  NAND2_X1 U9206 ( .A1(n10425), .A2(n10424), .ZN(n10453) );
  NAND2_X1 U9207 ( .A1(n13452), .A2(n13372), .ZN(n13433) );
  NAND2_X1 U9208 ( .A1(n13758), .A2(n14922), .ZN(n6639) );
  NAND2_X1 U9209 ( .A1(n10987), .A2(n10986), .ZN(n11038) );
  NAND2_X1 U9210 ( .A1(n10428), .A2(n10427), .ZN(n10747) );
  NAND2_X1 U9211 ( .A1(n7047), .A2(n7048), .ZN(n13597) );
  NAND2_X1 U9212 ( .A1(n13471), .A2(n13371), .ZN(n13453) );
  NAND2_X1 U9213 ( .A1(n13514), .A2(n13369), .ZN(n13490) );
  NAND2_X1 U9214 ( .A1(n10783), .A2(n10782), .ZN(n10784) );
  NAND2_X1 U9215 ( .A1(n12435), .A2(n12434), .ZN(n12433) );
  NAND2_X1 U9216 ( .A1(n12372), .A2(n12371), .ZN(n12370) );
  NAND2_X1 U9217 ( .A1(n12415), .A2(n12414), .ZN(n12413) );
  NAND2_X1 U9218 ( .A1(n8865), .A2(n8866), .ZN(n11632) );
  NAND2_X1 U9219 ( .A1(n6642), .A2(n8842), .ZN(n10581) );
  NAND2_X1 U9220 ( .A1(n10604), .A2(n10605), .ZN(n6642) );
  NAND2_X1 U9221 ( .A1(n12450), .A2(n8882), .ZN(n12372) );
  NAND2_X1 U9222 ( .A1(n6733), .A2(n12303), .ZN(n10783) );
  AOI21_X1 U9224 ( .B1(n12175), .B2(n12174), .A(n12173), .ZN(n12176) );
  NAND2_X1 U9225 ( .A1(n12135), .A2(n12134), .ZN(n12136) );
  NAND2_X1 U9226 ( .A1(n7494), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7498) );
  INV_X1 U9227 ( .A(n6882), .ZN(n12722) );
  INV_X1 U9228 ( .A(n14561), .ZN(n6648) );
  NOR2_X1 U9229 ( .A1(n10897), .A2(n15047), .ZN(n11331) );
  NAND2_X1 U9230 ( .A1(n6879), .A2(n6931), .ZN(n6878) );
  INV_X1 U9231 ( .A(n7260), .ZN(n7259) );
  INV_X1 U9232 ( .A(n10246), .ZN(n6713) );
  NAND2_X1 U9233 ( .A1(n8520), .A2(n8501), .ZN(n8503) );
  INV_X1 U9234 ( .A(n6845), .ZN(n6842) );
  NAND2_X1 U9235 ( .A1(n7101), .A2(n6567), .ZN(n14317) );
  INV_X1 U9236 ( .A(n6692), .ZN(n6691) );
  XNOR2_X1 U9237 ( .A(n6717), .B(n12800), .ZN(n12815) );
  NAND2_X1 U9238 ( .A1(n6649), .A2(n7519), .ZN(n7533) );
  NAND2_X1 U9239 ( .A1(n7517), .A2(n7518), .ZN(n6649) );
  NAND2_X1 U9240 ( .A1(n7877), .A2(n7876), .ZN(n7878) );
  NAND2_X1 U9241 ( .A1(n12034), .A2(n12033), .ZN(n12483) );
  INV_X1 U9242 ( .A(n12492), .ZN(n13046) );
  NAND2_X1 U9243 ( .A1(n7789), .A2(n7788), .ZN(n7802) );
  NAND2_X1 U9244 ( .A1(n7737), .A2(n7736), .ZN(n7750) );
  NAND2_X1 U9245 ( .A1(n7834), .A2(n7822), .ZN(n7823) );
  NAND2_X1 U9246 ( .A1(n12685), .A2(n12686), .ZN(n6891) );
  NAND2_X1 U9247 ( .A1(n12443), .A2(n12914), .ZN(n6658) );
  AND2_X1 U9248 ( .A1(n8174), .A2(n8772), .ZN(n10723) );
  NAND2_X2 U9249 ( .A1(n11970), .A2(n11969), .ZN(n14334) );
  NAND2_X1 U9250 ( .A1(n10930), .A2(n10929), .ZN(n10932) );
  NAND2_X1 U9251 ( .A1(n12043), .A2(n11977), .ZN(n11979) );
  NAND2_X1 U9252 ( .A1(n11145), .A2(n11144), .ZN(n11271) );
  AOI21_X1 U9253 ( .B1(n14303), .B2(n14304), .A(n11971), .ZN(n14285) );
  NAND2_X1 U9254 ( .A1(n11167), .A2(n11148), .ZN(n11246) );
  NAND2_X2 U9255 ( .A1(n11493), .A2(n7953), .ZN(n14589) );
  OAI21_X2 U9256 ( .B1(n11466), .B2(n7092), .A(n7091), .ZN(n11494) );
  AOI21_X2 U9257 ( .B1(n10509), .B2(n7943), .A(n7446), .ZN(n10498) );
  NAND2_X1 U9258 ( .A1(n10881), .A2(n7947), .ZN(n11000) );
  OAI22_X2 U9259 ( .A1(n12901), .A2(n7973), .B1(n12914), .B2(n7972), .ZN(
        n12890) );
  NAND2_X1 U9260 ( .A1(n7991), .A2(n6762), .ZN(n12844) );
  NAND2_X1 U9261 ( .A1(n7964), .A2(n7963), .ZN(n12978) );
  NAND2_X1 U9262 ( .A1(n12855), .A2(n7978), .ZN(n7090) );
  NAND2_X1 U9263 ( .A1(n12890), .A2(n12512), .ZN(n7060) );
  NAND2_X1 U9264 ( .A1(n12978), .A2(n6520), .ZN(n6652) );
  NAND2_X1 U9265 ( .A1(n12910), .A2(n7971), .ZN(n12901) );
  NAND2_X1 U9266 ( .A1(n12495), .A2(n10496), .ZN(n10495) );
  NAND2_X1 U9267 ( .A1(n10506), .A2(n12537), .ZN(n10496) );
  NAND2_X1 U9268 ( .A1(n10725), .A2(n10724), .ZN(n10930) );
  NOR2_X1 U9269 ( .A1(n14039), .A2(n11448), .ZN(n8173) );
  NAND2_X1 U9270 ( .A1(n6957), .A2(n6956), .ZN(n11736) );
  NOR2_X2 U9271 ( .A1(n8196), .A2(n8195), .ZN(n14093) );
  NAND2_X1 U9272 ( .A1(n6978), .A2(n6977), .ZN(n14214) );
  NAND2_X1 U9273 ( .A1(n6860), .A2(n6859), .ZN(P1_U3557) );
  INV_X1 U9274 ( .A(n7371), .ZN(n7370) );
  NAND2_X1 U9275 ( .A1(n6973), .A2(n6659), .ZN(P1_U3525) );
  NAND2_X1 U9276 ( .A1(n6975), .A2(n6660), .ZN(n6659) );
  OR2_X1 U9277 ( .A1(n8570), .A2(n8571), .ZN(n8572) );
  NAND2_X1 U9278 ( .A1(n8303), .A2(n8302), .ZN(n8307) );
  INV_X1 U9279 ( .A(n8401), .ZN(n7033) );
  OR2_X1 U9280 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND2_X1 U9281 ( .A1(n8495), .A2(n8494), .ZN(n8519) );
  NAND2_X1 U9282 ( .A1(n7022), .A2(n6661), .ZN(n6735) );
  NAND2_X1 U9283 ( .A1(n7023), .A2(n8403), .ZN(n6661) );
  NAND2_X1 U9284 ( .A1(n6662), .A2(n7002), .ZN(n7000) );
  NAND3_X1 U9285 ( .A1(n8531), .A2(n6739), .A3(n14333), .ZN(n6662) );
  NAND2_X1 U9286 ( .A1(n8186), .A2(n6760), .ZN(n8161) );
  NAND3_X1 U9287 ( .A1(n7220), .A2(n7016), .A3(n7219), .ZN(n7015) );
  NAND2_X1 U9288 ( .A1(n8148), .A2(n8149), .ZN(n8150) );
  NAND3_X1 U9289 ( .A1(n8203), .A2(n8202), .A3(n6576), .ZN(n6667) );
  NAND2_X1 U9290 ( .A1(n6444), .A2(n8053), .ZN(n8429) );
  NAND2_X1 U9291 ( .A1(n10903), .A2(n10904), .ZN(n11318) );
  NOR2_X2 U9292 ( .A1(n11409), .A2(n11410), .ZN(n11707) );
  NAND2_X1 U9293 ( .A1(n12726), .A2(n14559), .ZN(n6753) );
  NAND2_X1 U9294 ( .A1(n6947), .A2(n6946), .ZN(n6945) );
  AOI21_X1 U9295 ( .B1(n12778), .B2(n12777), .A(n12776), .ZN(n12803) );
  OAI21_X1 U9296 ( .B1(n12762), .B2(n12761), .A(n12760), .ZN(n12764) );
  NAND2_X1 U9297 ( .A1(n10626), .A2(n7061), .ZN(n10881) );
  NAND2_X1 U9298 ( .A1(n6765), .A2(n6764), .ZN(n12867) );
  NAND2_X1 U9299 ( .A1(n7976), .A2(n7975), .ZN(n12869) );
  NAND2_X1 U9300 ( .A1(n13756), .A2(n14915), .ZN(n6729) );
  NOR2_X2 U9301 ( .A1(n14557), .A2(n14558), .ZN(n14556) );
  XNOR2_X2 U9302 ( .A(n12738), .B(n12737), .ZN(n14557) );
  NOR2_X1 U9303 ( .A1(n14553), .A2(n14554), .ZN(n9610) );
  XNOR2_X1 U9304 ( .A(n6949), .B(n12811), .ZN(n6948) );
  INV_X1 U9305 ( .A(n10177), .ZN(n6731) );
  AOI21_X1 U9306 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n14944), .A(n14941), .ZN(
        n11412) );
  NOR2_X1 U9307 ( .A1(n12786), .A2(n12787), .ZN(n12790) );
  NAND2_X1 U9308 ( .A1(n11365), .A2(n11364), .ZN(n11504) );
  NAND2_X1 U9309 ( .A1(n7226), .A2(n7228), .ZN(n7224) );
  NAND3_X1 U9310 ( .A1(n13670), .A2(n7037), .A3(n6777), .ZN(n13756) );
  OAI21_X1 U9311 ( .B1(n10766), .B2(n7228), .A(n12305), .ZN(n7227) );
  NAND2_X1 U9312 ( .A1(n12370), .A2(n8885), .ZN(n12435) );
  OAI21_X1 U9313 ( .B1(n12346), .B2(n12345), .A(n6674), .ZN(n8909) );
  NAND2_X1 U9314 ( .A1(n12537), .A2(n12536), .ZN(n7943) );
  NAND2_X1 U9315 ( .A1(n12452), .A2(n12451), .ZN(n12450) );
  NAND2_X1 U9316 ( .A1(n10616), .A2(n10828), .ZN(n12545) );
  NAND2_X1 U9317 ( .A1(n10612), .A2(n8847), .ZN(n10810) );
  NAND2_X1 U9318 ( .A1(n10579), .A2(n7295), .ZN(n10612) );
  INV_X1 U9319 ( .A(n12869), .ZN(n6765) );
  NAND3_X1 U9320 ( .A1(n12631), .A2(n12630), .A3(n6676), .ZN(n6675) );
  NAND3_X1 U9321 ( .A1(n6678), .A2(n6677), .A3(n12676), .ZN(n12673) );
  NAND3_X1 U9322 ( .A1(n6749), .A2(n6887), .A3(n6891), .ZN(n6886) );
  AOI21_X1 U9323 ( .B1(n12579), .B2(n12578), .A(n12577), .ZN(n12585) );
  AOI21_X1 U9324 ( .B1(n6751), .B2(n6750), .A(n7340), .ZN(n12614) );
  OAI21_X1 U9325 ( .B1(n6514), .B2(n6744), .A(n12555), .ZN(n12559) );
  OR3_X1 U9326 ( .A1(n12563), .A2(n12562), .A3(n12561), .ZN(n12568) );
  NAND2_X2 U9327 ( .A1(n7090), .A2(n7089), .ZN(n12832) );
  NAND2_X1 U9328 ( .A1(n6681), .A2(n6680), .ZN(P3_U3296) );
  OAI21_X1 U9329 ( .B1(n6886), .B2(n12684), .A(n6682), .ZN(n6681) );
  NAND2_X1 U9330 ( .A1(n13004), .A2(n6683), .ZN(P3_U3487) );
  INV_X1 U9331 ( .A(n6684), .ZN(n6683) );
  OAI21_X1 U9332 ( .B1(n13057), .B2(n13043), .A(n13003), .ZN(n6684) );
  NAND2_X1 U9333 ( .A1(n13056), .A2(n6685), .ZN(P3_U3455) );
  INV_X1 U9334 ( .A(n6686), .ZN(n6685) );
  OAI21_X1 U9335 ( .B1(n13057), .B2(n13125), .A(n13055), .ZN(n6686) );
  NAND2_X1 U9336 ( .A1(n6747), .A2(n6745), .ZN(n12642) );
  NAND2_X1 U9337 ( .A1(n12609), .A2(n12988), .ZN(n6751) );
  OAI21_X1 U9338 ( .B1(n12665), .B2(n12664), .A(n12833), .ZN(n12666) );
  INV_X1 U9339 ( .A(n8980), .ZN(n6687) );
  XNOR2_X2 U9340 ( .A(n8976), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U9341 ( .A1(n11881), .A2(n11880), .ZN(n11879) );
  XNOR2_X1 U9342 ( .A(n13376), .B(n13375), .ZN(n6694) );
  NAND2_X1 U9343 ( .A1(n13357), .A2(n13356), .ZN(n13586) );
  INV_X1 U9344 ( .A(n6943), .ZN(n6942) );
  NOR2_X1 U9345 ( .A1(n12755), .A2(n12756), .ZN(n12786) );
  NAND2_X1 U9346 ( .A1(n7040), .A2(n7038), .ZN(n11507) );
  NAND2_X1 U9347 ( .A1(n6950), .A2(n12809), .ZN(n6949) );
  NOR2_X1 U9348 ( .A1(n12790), .A2(n12789), .ZN(n12810) );
  NAND2_X2 U9349 ( .A1(n7555), .A2(n7583), .ZN(n10240) );
  NAND2_X1 U9350 ( .A1(n7255), .A2(n14623), .ZN(n7037) );
  XNOR2_X1 U9351 ( .A(n6690), .B(n13375), .ZN(n13671) );
  NAND2_X1 U9352 ( .A1(n6720), .A2(n6719), .ZN(n6738) );
  NOR2_X2 U9353 ( .A1(n6693), .A2(n6691), .ZN(n14414) );
  NAND2_X1 U9354 ( .A1(n8833), .A2(n10396), .ZN(n8838) );
  NAND2_X1 U9355 ( .A1(n12524), .A2(n14985), .ZN(n8833) );
  INV_X1 U9356 ( .A(n10581), .ZN(n7298) );
  NAND2_X1 U9357 ( .A1(n11040), .A2(n11039), .ZN(n11290) );
  NAND2_X1 U9358 ( .A1(n12297), .A2(n10094), .ZN(n10116) );
  NAND2_X1 U9359 ( .A1(n13223), .A2(n13152), .ZN(n6802) );
  NAND2_X1 U9360 ( .A1(n6695), .A2(n13255), .ZN(n13191) );
  NAND2_X1 U9361 ( .A1(n13186), .A2(n13185), .ZN(n6695) );
  NAND2_X1 U9362 ( .A1(n6738), .A2(n8128), .ZN(n8108) );
  NAND2_X1 U9363 ( .A1(n12129), .A2(n12128), .ZN(n6697) );
  NAND2_X1 U9364 ( .A1(n12149), .A2(n12148), .ZN(n12152) );
  NAND2_X1 U9365 ( .A1(n12282), .A2(n12281), .ZN(n12337) );
  NAND2_X1 U9366 ( .A1(n6698), .A2(n7394), .ZN(n7393) );
  NAND2_X1 U9367 ( .A1(n7396), .A2(n6535), .ZN(n6698) );
  NAND2_X1 U9368 ( .A1(n7384), .A2(n6577), .ZN(n12282) );
  NAND2_X1 U9369 ( .A1(n13443), .A2(n13428), .ZN(n13426) );
  INV_X1 U9370 ( .A(n6699), .ZN(n13621) );
  NAND2_X1 U9371 ( .A1(n7036), .A2(n7034), .ZN(P2_U3528) );
  NOR2_X2 U9372 ( .A1(n11044), .A2(n12130), .ZN(n6701) );
  NAND2_X2 U9373 ( .A1(n13591), .A2(n13578), .ZN(n13573) );
  INV_X1 U9374 ( .A(n6928), .ZN(n6927) );
  NAND3_X1 U9375 ( .A1(n12836), .A2(n12835), .A3(n14991), .ZN(n12840) );
  AOI21_X1 U9376 ( .B1(n6948), .B2(n12710), .A(n6945), .ZN(n12814) );
  NAND2_X1 U9377 ( .A1(n8476), .A2(n8475), .ZN(n6702) );
  NAND2_X1 U9378 ( .A1(n8275), .A2(n8274), .ZN(n8303) );
  NOR2_X1 U9379 ( .A1(n10256), .A2(n10257), .ZN(n10589) );
  NOR2_X1 U9380 ( .A1(n11527), .A2(n11526), .ZN(n11593) );
  NOR2_X1 U9381 ( .A1(n6561), .A2(n10243), .ZN(n6944) );
  AOI21_X1 U9382 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n11122), .A(n11119), .ZN(
        n11525) );
  NAND2_X1 U9383 ( .A1(n14596), .A2(n14595), .ZN(n14594) );
  NAND2_X1 U9384 ( .A1(n12853), .A2(n12657), .ZN(n7915) );
  NAND2_X1 U9385 ( .A1(n6763), .A2(n15029), .ZN(n6762) );
  NAND2_X1 U9386 ( .A1(n11879), .A2(n8875), .ZN(n11907) );
  INV_X1 U9387 ( .A(n12857), .ZN(n12696) );
  INV_X1 U9388 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7310) );
  NAND2_X1 U9389 ( .A1(n12832), .A2(n9624), .ZN(n12835) );
  NAND2_X1 U9390 ( .A1(n7347), .A2(n7501), .ZN(n7938) );
  OAI22_X1 U9391 ( .A1(n7840), .A2(n9818), .B1(n7980), .B2(n10142), .ZN(n7348)
         );
  NOR2_X1 U9392 ( .A1(n14969), .A2(n11687), .ZN(n11690) );
  NOR2_X1 U9393 ( .A1(n11403), .A2(n11404), .ZN(n11408) );
  NAND2_X1 U9394 ( .A1(n6732), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7523) );
  OAI21_X1 U9395 ( .B1(n6454), .B2(n15042), .A(n6871), .ZN(n10147) );
  AOI22_X1 U9396 ( .A1(n8744), .A2(n8743), .B1(n8742), .B2(n8741), .ZN(n8810)
         );
  NAND3_X1 U9397 ( .A1(n6500), .A2(n7029), .A3(n11800), .ZN(n7020) );
  INV_X1 U9398 ( .A(SI_1_), .ZN(n6719) );
  INV_X1 U9399 ( .A(n8101), .ZN(n6720) );
  OAI21_X1 U9400 ( .B1(n8519), .B2(n11989), .A(n8518), .ZN(n8531) );
  NAND2_X1 U9401 ( .A1(n7872), .A2(n12648), .ZN(n12878) );
  NAND2_X1 U9402 ( .A1(n6723), .A2(n6721), .ZN(P3_U3454) );
  OR2_X1 U9403 ( .A1(n8046), .A2(n15037), .ZN(n6723) );
  NAND2_X1 U9404 ( .A1(n6726), .A2(n6724), .ZN(P3_U3486) );
  OR2_X1 U9405 ( .A1(n8046), .A2(n15049), .ZN(n6726) );
  NAND2_X1 U9406 ( .A1(n12864), .A2(n12868), .ZN(n12866) );
  NAND2_X1 U9407 ( .A1(n6729), .A2(n6727), .ZN(P2_U3496) );
  AND2_X2 U9408 ( .A1(n7480), .A2(n7479), .ZN(n7662) );
  NAND2_X1 U9409 ( .A1(n13490), .A2(n13493), .ZN(n13489) );
  OAI21_X2 U9410 ( .B1(n10347), .B2(n8920), .A(n8831), .ZN(n8835) );
  INV_X1 U9411 ( .A(n7521), .ZN(n6732) );
  NAND2_X1 U9412 ( .A1(n10543), .A2(n6930), .ZN(n14929) );
  INV_X1 U9413 ( .A(n12810), .ZN(n6950) );
  AND2_X4 U9414 ( .A1(n8980), .A2(n13788), .ZN(n9027) );
  INV_X1 U9415 ( .A(n10767), .ZN(n6733) );
  NAND2_X1 U9416 ( .A1(n8307), .A2(n8306), .ZN(n8324) );
  AOI21_X2 U9417 ( .B1(n12041), .B2(n12039), .A(n12038), .ZN(n14415) );
  NAND2_X1 U9418 ( .A1(n7426), .A2(n7427), .ZN(n12111) );
  NAND2_X1 U9419 ( .A1(n6758), .A2(n6757), .ZN(n7384) );
  NAND2_X1 U9420 ( .A1(n8135), .A2(n8134), .ZN(n8159) );
  NAND2_X1 U9421 ( .A1(n8261), .A2(n8260), .ZN(n8271) );
  NAND2_X1 U9422 ( .A1(n6735), .A2(n8486), .ZN(n8495) );
  NAND2_X1 U9423 ( .A1(n6742), .A2(n6737), .ZN(n6736) );
  INV_X1 U9424 ( .A(n8108), .ZN(n8105) );
  NAND2_X1 U9425 ( .A1(n8682), .A2(n8681), .ZN(n7222) );
  NAND2_X1 U9426 ( .A1(n13640), .A2(n13781), .ZN(n13638) );
  NOR2_X2 U9427 ( .A1(n13462), .A2(n13446), .ZN(n13443) );
  AND2_X2 U9428 ( .A1(n13552), .A2(n13561), .ZN(n13547) );
  AND2_X2 U9429 ( .A1(n13600), .A2(n13593), .ZN(n13591) );
  AND2_X2 U9430 ( .A1(n10113), .A2(n10736), .ZN(n10457) );
  NOR2_X2 U9431 ( .A1(n10787), .A2(n12115), .ZN(n7445) );
  OR2_X1 U9432 ( .A1(n11187), .A2(n7203), .ZN(n7198) );
  NOR2_X2 U9433 ( .A1(n14535), .A2(n8827), .ZN(n9671) );
  NAND2_X1 U9434 ( .A1(n8002), .A2(n7308), .ZN(n6740) );
  NAND2_X1 U9435 ( .A1(n14582), .A2(n12593), .ZN(n11815) );
  NAND2_X1 U9436 ( .A1(n7238), .A2(n7434), .ZN(n9013) );
  NOR2_X2 U9437 ( .A1(n9455), .A2(n8972), .ZN(n7434) );
  NAND2_X1 U9438 ( .A1(n10453), .A2(n10426), .ZN(n10428) );
  NAND2_X1 U9439 ( .A1(n8187), .A2(n6759), .ZN(n6742) );
  NAND2_X1 U9440 ( .A1(n11507), .A2(n11506), .ZN(n11542) );
  INV_X1 U9441 ( .A(n6976), .ZN(n6974) );
  NAND2_X1 U9442 ( .A1(n8986), .A2(n9263), .ZN(n8999) );
  NAND2_X1 U9443 ( .A1(n6830), .A2(n6828), .ZN(n8456) );
  XNOR2_X2 U9444 ( .A(n7474), .B(n13129), .ZN(n12037) );
  NAND2_X1 U9445 ( .A1(n12679), .A2(n12673), .ZN(n6889) );
  NAND3_X1 U9446 ( .A1(n12638), .A2(n12637), .A3(n6748), .ZN(n6747) );
  NAND2_X1 U9447 ( .A1(n12813), .A2(n14936), .ZN(n6947) );
  NAND2_X1 U9448 ( .A1(n12413), .A2(n8880), .ZN(n12452) );
  NAND3_X1 U9449 ( .A1(n12206), .A2(n12205), .A3(n6563), .ZN(n6758) );
  AND2_X1 U9450 ( .A1(n8204), .A2(n8186), .ZN(n6759) );
  OR2_X1 U9451 ( .A1(n7216), .A2(SI_3_), .ZN(n6760) );
  BUF_X2 U9452 ( .A(n12076), .Z(n6761) );
  NAND2_X1 U9453 ( .A1(n6818), .A2(n6816), .ZN(n9278) );
  INV_X1 U9454 ( .A(n11613), .ZN(n9261) );
  OAI21_X1 U9455 ( .B1(n8130), .B2(n8100), .A(n8099), .ZN(n8101) );
  AOI21_X2 U9456 ( .B1(n6936), .B2(n6935), .A(n6772), .ZN(n12738) );
  INV_X1 U9457 ( .A(n10784), .ZN(n6775) );
  NOR2_X1 U9458 ( .A1(n12770), .A2(n12771), .ZN(n12773) );
  NOR2_X1 U9459 ( .A1(n14970), .A2(n14971), .ZN(n14969) );
  INV_X1 U9460 ( .A(n11690), .ZN(n6885) );
  INV_X1 U9461 ( .A(n11408), .ZN(n6873) );
  XNOR2_X2 U9462 ( .A(n7507), .B(n7506), .ZN(n10145) );
  NAND2_X1 U9463 ( .A1(n6778), .A2(n14200), .ZN(n7497) );
  NAND3_X1 U9464 ( .A1(n7495), .A2(n7496), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n6778) );
  AND2_X2 U9465 ( .A1(n7521), .A2(n7451), .ZN(n7308) );
  NAND2_X1 U9466 ( .A1(n10773), .A2(n12109), .ZN(n10787) );
  NAND2_X1 U9467 ( .A1(n13887), .A2(n13888), .ZN(n13919) );
  AOI21_X1 U9468 ( .B1(n7990), .B2(n14991), .A(n7989), .ZN(n7991) );
  NAND2_X1 U9469 ( .A1(n12473), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U9470 ( .A1(n11262), .A2(n6782), .ZN(n6780) );
  NAND2_X1 U9471 ( .A1(n6568), .A2(n6780), .ZN(n11243) );
  AOI21_X2 U9472 ( .B1(n14398), .B2(n14799), .A(n6508), .ZN(n6976) );
  NAND2_X1 U9473 ( .A1(n14317), .A2(n7116), .ZN(n11993) );
  NAND2_X1 U9474 ( .A1(n14245), .A2(n6784), .ZN(n6790) );
  NAND2_X1 U9475 ( .A1(n6788), .A2(n14230), .ZN(n6786) );
  OAI21_X1 U9476 ( .B1(n11675), .B2(n6794), .A(n6792), .ZN(n11929) );
  NAND2_X1 U9477 ( .A1(n6796), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7122) );
  NAND4_X1 U9478 ( .A1(n8062), .A2(n6983), .A3(n6982), .A4(n6476), .ZN(n6796)
         );
  NAND3_X1 U9479 ( .A1(n6983), .A2(n8062), .A3(n6982), .ZN(n8821) );
  AND2_X2 U9480 ( .A1(n6983), .A2(n6982), .ZN(n8063) );
  INV_X1 U9481 ( .A(n8063), .ZN(n8477) );
  NAND2_X1 U9482 ( .A1(n7336), .A2(n6474), .ZN(n13223) );
  INV_X1 U9483 ( .A(n13151), .ZN(n6803) );
  INV_X1 U9484 ( .A(n9456), .ZN(n7435) );
  NAND3_X1 U9485 ( .A1(n6807), .A2(n6804), .A3(P2_IR_REG_27__SCAN_IN), .ZN(
        n6805) );
  INV_X1 U9486 ( .A(n9456), .ZN(n6807) );
  NAND2_X1 U9487 ( .A1(n7435), .A2(n6804), .ZN(n9012) );
  NAND2_X1 U9488 ( .A1(n11435), .A2(n7326), .ZN(n6818) );
  NAND2_X1 U9489 ( .A1(n10376), .A2(n9080), .ZN(n6820) );
  INV_X1 U9490 ( .A(n13150), .ZN(n6823) );
  NAND2_X1 U9491 ( .A1(n6822), .A2(n6475), .ZN(n9445) );
  NAND2_X1 U9492 ( .A1(n6823), .A2(n6826), .ZN(n6822) );
  NAND2_X1 U9493 ( .A1(n8369), .A2(n6513), .ZN(n6830) );
  NAND2_X1 U9494 ( .A1(n8500), .A2(n8499), .ZN(n6845) );
  AOI21_X1 U9495 ( .B1(n13432), .B2(n13418), .A(n13417), .ZN(n6849) );
  INV_X4 U9496 ( .A(n7499), .ZN(n8622) );
  OAI21_X1 U9497 ( .B1(n6850), .B2(SI_4_), .A(n8204), .ZN(n8188) );
  MUX2_X1 U9498 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7499), .Z(n6850) );
  OAI211_X2 U9499 ( .C1(n8157), .C2(n9807), .A(n6525), .B(n6854), .ZN(n10727)
         );
  AND3_X1 U9500 ( .A1(n8116), .A2(n8115), .A3(n8114), .ZN(n11449) );
  NAND4_X1 U9501 ( .A1(n8116), .A2(n8115), .A3(n8114), .A4(n11448), .ZN(n11447) );
  NAND3_X1 U9502 ( .A1(n11484), .A2(n6856), .A3(n6855), .ZN(n11677) );
  NAND2_X1 U9503 ( .A1(n8063), .A2(n6869), .ZN(n6870) );
  NAND2_X1 U9504 ( .A1(n10146), .A2(n10147), .ZN(n10184) );
  NAND2_X1 U9505 ( .A1(n6454), .A2(n15042), .ZN(n6871) );
  NAND2_X1 U9506 ( .A1(n10184), .A2(n10183), .ZN(n10186) );
  INV_X1 U9507 ( .A(n10555), .ZN(n6879) );
  NAND2_X1 U9508 ( .A1(n12671), .A2(n12672), .ZN(n6890) );
  NAND2_X1 U9509 ( .A1(n12491), .A2(n12490), .ZN(n12671) );
  OAI21_X1 U9510 ( .B1(n7716), .B2(n6894), .A(n7733), .ZN(n6893) );
  NAND3_X1 U9511 ( .A1(n6902), .A2(n6901), .A3(n7568), .ZN(n7571) );
  NAND2_X1 U9512 ( .A1(n6903), .A2(n6905), .ZN(n6901) );
  NAND2_X1 U9513 ( .A1(n6903), .A2(n7538), .ZN(n6902) );
  INV_X1 U9514 ( .A(n6904), .ZN(n6903) );
  NAND2_X1 U9515 ( .A1(n7753), .A2(n6909), .ZN(n6906) );
  NAND2_X1 U9516 ( .A1(n6906), .A2(n6907), .ZN(n7789) );
  NAND2_X1 U9517 ( .A1(n8902), .A2(n6914), .ZN(n6912) );
  NAND2_X1 U9518 ( .A1(n6921), .A2(n12097), .ZN(n10754) );
  NAND2_X1 U9519 ( .A1(n6922), .A2(n6480), .ZN(n13750) );
  NAND2_X1 U9520 ( .A1(n13664), .A2(n6926), .ZN(n6922) );
  NAND2_X1 U9521 ( .A1(n6923), .A2(n6924), .ZN(n13665) );
  NAND2_X1 U9522 ( .A1(n13664), .A2(n6925), .ZN(n6923) );
  OR2_X1 U9523 ( .A1(n14922), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6924) );
  NOR2_X2 U9524 ( .A1(n11566), .A2(n14620), .ZN(n13640) );
  OR2_X2 U9525 ( .A1(n11549), .A2(n12157), .ZN(n11566) );
  AND2_X2 U9526 ( .A1(n13547), .A2(n13526), .ZN(n13507) );
  AOI21_X1 U9527 ( .B1(n13426), .B2(n13335), .A(n13620), .ZN(n6928) );
  NAND2_X2 U9528 ( .A1(n13795), .A2(n9499), .ZN(n9033) );
  NAND2_X1 U9529 ( .A1(n10910), .A2(n6507), .ZN(n6929) );
  NAND2_X1 U9530 ( .A1(n10177), .A2(n6942), .ZN(n6940) );
  NAND2_X1 U9531 ( .A1(n10177), .A2(n10178), .ZN(n10237) );
  NAND2_X1 U9532 ( .A1(n6951), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U9533 ( .A1(n6952), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U9534 ( .A1(n6951), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8255) );
  NAND2_X1 U9535 ( .A1(n6951), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U9536 ( .A1(n6951), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U9537 ( .A1(n6951), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U9538 ( .A1(n6951), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U9539 ( .A1(n6951), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U9540 ( .A1(n6951), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U9541 ( .A1(n6951), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U9542 ( .A1(n6951), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U9543 ( .A1(n6951), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U9544 ( .A1(n6951), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U9545 ( .A1(n6951), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U9546 ( .A1(n6951), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U9547 ( .A1(n6951), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8665) );
  NAND2_X1 U9548 ( .A1(n6951), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U9549 ( .A1(n6951), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8693) );
  OAI21_X1 U9550 ( .B1(n8179), .B2(n6955), .A(n6954), .ZN(n6953) );
  NAND2_X1 U9551 ( .A1(n11346), .A2(n6958), .ZN(n6957) );
  NAND2_X1 U9552 ( .A1(n14334), .A2(n6464), .ZN(n6961) );
  NAND2_X1 U9553 ( .A1(n11918), .A2(n6501), .ZN(n6964) );
  NAND2_X1 U9554 ( .A1(n6964), .A2(n6965), .ZN(n14349) );
  OAI21_X1 U9555 ( .B1(n11153), .B2(n6969), .A(n6968), .ZN(n11344) );
  NAND2_X1 U9556 ( .A1(n7207), .A2(n6972), .ZN(n14518) );
  NAND2_X1 U9557 ( .A1(n14264), .A2(n6581), .ZN(n6978) );
  NAND2_X1 U9558 ( .A1(n8376), .A2(n8377), .ZN(n8375) );
  NOR2_X2 U9559 ( .A1(n8165), .A2(n8056), .ZN(n6982) );
  NAND2_X1 U9560 ( .A1(n8242), .A2(n8243), .ZN(n8241) );
  NAND2_X2 U9561 ( .A1(n6985), .A2(n6984), .ZN(n8352) );
  NAND3_X1 U9562 ( .A1(n8646), .A2(n8647), .A3(n6578), .ZN(n6986) );
  NAND2_X1 U9563 ( .A1(n8630), .A2(n6992), .ZN(n6989) );
  OAI21_X1 U9564 ( .B1(n8630), .B2(n6993), .A(n6992), .ZN(n8645) );
  NAND2_X1 U9565 ( .A1(n6989), .A2(n6990), .ZN(n8643) );
  NAND2_X1 U9566 ( .A1(n8589), .A2(n6997), .ZN(n6994) );
  NAND2_X1 U9567 ( .A1(n6994), .A2(n6995), .ZN(n8605) );
  AND2_X1 U9568 ( .A1(n7000), .A2(n6998), .ZN(n8570) );
  NAND2_X1 U9569 ( .A1(n7000), .A2(n6572), .ZN(n8569) );
  NAND2_X1 U9570 ( .A1(n8294), .A2(n7009), .ZN(n7007) );
  NAND2_X1 U9571 ( .A1(n7007), .A2(n7005), .ZN(n8332) );
  NAND3_X1 U9572 ( .A1(n7029), .A2(n11800), .A3(n7028), .ZN(n7019) );
  AOI21_X1 U9573 ( .B1(n7026), .B2(n7024), .A(n8445), .ZN(n7023) );
  NAND2_X1 U9574 ( .A1(n13629), .A2(n6468), .ZN(n7047) );
  NAND2_X1 U9575 ( .A1(n7060), .A2(n7058), .ZN(n7976) );
  NOR2_X1 U9576 ( .A1(n12552), .A2(n7062), .ZN(n7061) );
  INV_X1 U9577 ( .A(n11935), .ZN(n7960) );
  INV_X1 U9578 ( .A(n13115), .ZN(n7078) );
  NAND3_X1 U9579 ( .A1(n8002), .A2(n7374), .A3(n7308), .ZN(n7079) );
  NAND3_X1 U9580 ( .A1(n7308), .A2(n7081), .A3(n7307), .ZN(n7688) );
  AND2_X2 U9581 ( .A1(n7309), .A2(n7450), .ZN(n7081) );
  NAND2_X1 U9582 ( .A1(n7083), .A2(n7086), .ZN(n9632) );
  NAND2_X1 U9583 ( .A1(n12855), .A2(n7084), .ZN(n7083) );
  OAI21_X1 U9584 ( .B1(n14589), .B2(n14576), .A(n11639), .ZN(n7955) );
  NAND2_X1 U9585 ( .A1(n12939), .A2(n12938), .ZN(n12937) );
  NAND2_X1 U9586 ( .A1(n7960), .A2(n7959), .ZN(n11937) );
  NAND2_X1 U9587 ( .A1(n10498), .A2(n7944), .ZN(n10497) );
  NAND2_X1 U9588 ( .A1(n7941), .A2(n7940), .ZN(n10509) );
  NAND2_X1 U9589 ( .A1(n14367), .A2(n7103), .ZN(n7101) );
  INV_X1 U9590 ( .A(n11927), .ZN(n7120) );
  NAND2_X1 U9591 ( .A1(n14286), .A2(n7121), .ZN(n14267) );
  NAND2_X1 U9592 ( .A1(n15215), .A2(n15214), .ZN(n9567) );
  XNOR2_X1 U9593 ( .A(n9566), .B(n9565), .ZN(n15221) );
  XNOR2_X1 U9594 ( .A(n9555), .B(n7124), .ZN(n15215) );
  XNOR2_X1 U9595 ( .A(n9554), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U9596 ( .A1(n9557), .A2(n7128), .ZN(n7127) );
  NAND2_X1 U9597 ( .A1(n9562), .A2(n6580), .ZN(n7125) );
  NAND3_X1 U9598 ( .A1(n7127), .A2(n6580), .A3(n6472), .ZN(n7126) );
  INV_X1 U9599 ( .A(n14688), .ZN(n7139) );
  OAI21_X1 U9600 ( .B1(n6463), .B2(n7148), .A(n7145), .ZN(n9603) );
  INV_X1 U9601 ( .A(n7159), .ZN(n14684) );
  NAND2_X1 U9602 ( .A1(n14001), .A2(n13886), .ZN(n13887) );
  NAND3_X1 U9603 ( .A1(n11622), .A2(n11650), .A3(n7165), .ZN(n7163) );
  NAND2_X1 U9604 ( .A1(n7163), .A2(n7164), .ZN(n11866) );
  OR2_X1 U9605 ( .A1(n7169), .A2(n7167), .ZN(n7164) );
  NOR2_X1 U9606 ( .A1(n7169), .A2(n7166), .ZN(n7165) );
  INV_X1 U9607 ( .A(n9723), .ZN(n7171) );
  NAND2_X1 U9608 ( .A1(n7180), .A2(n7179), .ZN(n7183) );
  INV_X1 U9609 ( .A(n7183), .ZN(n14698) );
  INV_X1 U9610 ( .A(n14701), .ZN(n7179) );
  INV_X1 U9611 ( .A(n14700), .ZN(n7180) );
  NAND2_X1 U9612 ( .A1(n9766), .A2(n7187), .ZN(n7184) );
  AND2_X1 U9613 ( .A1(n7198), .A2(n6565), .ZN(n7197) );
  NOR2_X1 U9614 ( .A1(n11187), .A2(n7200), .ZN(n7199) );
  NAND2_X1 U9615 ( .A1(n13828), .A2(n7204), .ZN(n13937) );
  NAND2_X1 U9616 ( .A1(n13937), .A2(n13990), .ZN(n13842) );
  NOR2_X1 U9617 ( .A1(n13516), .A2(n7215), .ZN(n7214) );
  NAND3_X1 U9618 ( .A1(n8686), .A2(n7223), .A3(n8685), .ZN(n7219) );
  NAND3_X1 U9619 ( .A1(n8682), .A2(n7223), .A3(n8681), .ZN(n7220) );
  INV_X1 U9620 ( .A(n8706), .ZN(n7223) );
  NAND2_X1 U9621 ( .A1(n10762), .A2(n7226), .ZN(n7225) );
  NAND2_X1 U9622 ( .A1(n13477), .A2(n7235), .ZN(n7234) );
  NAND2_X1 U9623 ( .A1(n13681), .A2(n13472), .ZN(n7237) );
  NAND4_X1 U9624 ( .A1(n9057), .A2(n9002), .A3(n9000), .A4(n8998), .ZN(n7241)
         );
  NAND2_X1 U9625 ( .A1(n8307), .A2(n7245), .ZN(n7244) );
  NAND2_X1 U9626 ( .A1(n12301), .A2(n10744), .ZN(n7248) );
  NAND2_X1 U9627 ( .A1(n10450), .A2(n6569), .ZN(n7249) );
  NAND3_X1 U9628 ( .A1(n7249), .A2(n7248), .A3(n10750), .ZN(n10761) );
  NAND2_X1 U9629 ( .A1(n8552), .A2(n8539), .ZN(n8541) );
  INV_X1 U9630 ( .A(n8540), .ZN(n7252) );
  INV_X1 U9631 ( .A(n8502), .ZN(n7261) );
  OAI21_X1 U9632 ( .B1(n13605), .B2(n13392), .A(n13394), .ZN(n13584) );
  NAND2_X1 U9633 ( .A1(n7275), .A2(n6596), .ZN(n8620) );
  NAND3_X1 U9634 ( .A1(n8600), .A2(n7274), .A3(n6595), .ZN(n7275) );
  INV_X1 U9635 ( .A(n7274), .ZN(n7276) );
  NAND2_X1 U9636 ( .A1(n8600), .A2(n8586), .ZN(n9369) );
  INV_X1 U9637 ( .A(n9368), .ZN(n7277) );
  NAND2_X1 U9638 ( .A1(n11633), .A2(n6571), .ZN(n7279) );
  INV_X1 U9639 ( .A(n8869), .ZN(n7278) );
  NAND2_X1 U9640 ( .A1(n11907), .A2(n7290), .ZN(n7288) );
  OAI21_X2 U9641 ( .B1(n12395), .B2(n12396), .A(n7300), .ZN(n12461) );
  AND2_X1 U9642 ( .A1(n7450), .A2(n7306), .ZN(n7305) );
  NAND4_X1 U9643 ( .A1(n7307), .A2(n7308), .A3(n7309), .A4(n6597), .ZN(n7703)
         );
  AND4_X2 U9644 ( .A1(n7307), .A2(n7308), .A3(n7309), .A4(n7305), .ZN(n8003)
         );
  AND3_X2 U9645 ( .A1(n7312), .A2(n7311), .A3(n7310), .ZN(n7309) );
  INV_X1 U9646 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7312) );
  NAND2_X1 U9647 ( .A1(n7739), .A2(n7313), .ZN(n7318) );
  AND2_X1 U9648 ( .A1(n12330), .A2(n13330), .ZN(n12065) );
  OAI21_X1 U9649 ( .B1(n9093), .B2(n7328), .A(n7329), .ZN(n9134) );
  OR2_X2 U9650 ( .A1(n7241), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U9651 ( .A1(n12987), .A2(n7343), .ZN(n7341) );
  INV_X1 U9652 ( .A(n7348), .ZN(n7347) );
  OAI21_X1 U9653 ( .B1(n9645), .B2(n7352), .A(n7350), .ZN(n7359) );
  INV_X1 U9654 ( .A(n12521), .ZN(n7360) );
  NAND2_X1 U9655 ( .A1(n11029), .A2(n7364), .ZN(n7363) );
  NAND2_X1 U9656 ( .A1(n10495), .A2(n7368), .ZN(n7367) );
  AND2_X2 U9657 ( .A1(n7999), .A2(n7373), .ZN(n7486) );
  NAND2_X1 U9658 ( .A1(n12950), .A2(n7381), .ZN(n7818) );
  NAND2_X1 U9659 ( .A1(n12275), .A2(n7385), .ZN(n7383) );
  OAI22_X1 U9660 ( .A1(n12273), .A2(n12274), .B1(n12265), .B2(n12266), .ZN(
        n7389) );
  INV_X1 U9661 ( .A(n12207), .ZN(n7390) );
  NAND2_X1 U9662 ( .A1(n12188), .A2(n12187), .ZN(n7396) );
  NAND3_X1 U9663 ( .A1(n12099), .A2(n7425), .A3(n7424), .ZN(n7426) );
  OR2_X1 U9664 ( .A1(n12106), .A2(n12107), .ZN(n7424) );
  NOR2_X1 U9665 ( .A1(n12111), .A2(n12110), .ZN(n12112) );
  NAND2_X1 U9666 ( .A1(n12288), .A2(n7432), .ZN(n7431) );
  NAND3_X1 U9667 ( .A1(n7431), .A2(n7429), .A3(n7428), .ZN(P2_U3328) );
  NAND3_X1 U9668 ( .A1(n12336), .A2(n12337), .A3(n12339), .ZN(n7428) );
  INV_X1 U9669 ( .A(n12339), .ZN(n7433) );
  NAND2_X1 U9670 ( .A1(n12163), .A2(n6583), .ZN(n7436) );
  INV_X1 U9671 ( .A(n12164), .ZN(n7437) );
  NAND2_X1 U9672 ( .A1(n12136), .A2(n6582), .ZN(n7440) );
  INV_X1 U9673 ( .A(n12137), .ZN(n7441) );
  NOR2_X2 U9674 ( .A1(n13335), .A2(n13426), .ZN(n13382) );
  NAND2_X1 U9675 ( .A1(n12012), .A2(n11980), .ZN(n11984) );
  NAND2_X1 U9676 ( .A1(n8772), .A2(n8771), .ZN(n10719) );
  INV_X1 U9677 ( .A(n8689), .ZN(n8708) );
  OR2_X1 U9678 ( .A1(n8689), .A2(n11455), .ZN(n8097) );
  OR2_X1 U9679 ( .A1(n9679), .A2(n11449), .ZN(n8772) );
  NAND2_X1 U9680 ( .A1(n8086), .A2(n8085), .ZN(n8088) );
  INV_X1 U9681 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7496) );
  INV_X1 U9682 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7492) );
  INV_X1 U9683 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9135) );
  CLKBUF_X1 U9684 ( .A(n11622), .Z(n11651) );
  INV_X1 U9685 ( .A(n8088), .ZN(n8090) );
  OR2_X1 U9686 ( .A1(n14535), .A2(P1_B_REG_SCAN_IN), .ZN(n9774) );
  NAND2_X1 U9687 ( .A1(n8639), .A2(n8638), .ZN(n8650) );
  AND2_X1 U9688 ( .A1(n9671), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9672) );
  AND2_X1 U9689 ( .A1(n10523), .A2(n12285), .ZN(n14889) );
  BUF_X1 U9690 ( .A(n7477), .Z(n13132) );
  NAND3_X1 U9691 ( .A1(n7493), .A2(n7492), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7494) );
  INV_X1 U9692 ( .A(n14251), .ZN(n12000) );
  INV_X1 U9693 ( .A(n9656), .ZN(n9658) );
  INV_X1 U9694 ( .A(n9655), .ZN(n11573) );
  AOI21_X1 U9695 ( .B1(n13868), .B2(n10718), .A(n9672), .ZN(n9673) );
  NAND2_X1 U9696 ( .A1(n7475), .A2(n7473), .ZN(n7477) );
  INV_X1 U9697 ( .A(n12808), .ZN(n12680) );
  OR2_X1 U9698 ( .A1(n12808), .A2(n8035), .ZN(n14996) );
  NAND2_X1 U9699 ( .A1(n8810), .A2(n8809), .ZN(n8811) );
  XNOR2_X1 U9700 ( .A(n9278), .B(n9276), .ZN(n13273) );
  OR2_X1 U9701 ( .A1(n10847), .A2(n6646), .ZN(n7842) );
  OR2_X1 U9702 ( .A1(n10639), .A2(n6646), .ZN(n7826) );
  OR2_X1 U9703 ( .A1(n10270), .A2(n6646), .ZN(n7794) );
  OAI21_X1 U9704 ( .B1(n13163), .B2(n9513), .A(n9512), .ZN(P2_U3186) );
  NOR2_X1 U9705 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9569), .ZN(n9521) );
  AND2_X1 U9706 ( .A1(n9001), .A2(n9000), .ZN(n9003) );
  INV_X1 U9707 ( .A(n7999), .ZN(n8006) );
  NAND2_X1 U9708 ( .A1(n8585), .A2(n8582), .ZN(n8581) );
  INV_X2 U9709 ( .A(n8622), .ZN(n9014) );
  AND2_X1 U9710 ( .A1(n9462), .A2(n9012), .ZN(n9478) );
  NAND2_X1 U9711 ( .A1(n9445), .A2(n9444), .ZN(n9486) );
  INV_X2 U9712 ( .A(n9026), .ZN(n9492) );
  NAND2_X1 U9713 ( .A1(n8719), .A2(n8718), .ZN(n8757) );
  INV_X1 U9714 ( .A(n13336), .ZN(n13751) );
  NAND2_X1 U9715 ( .A1(n8757), .A2(n8746), .ZN(n8724) );
  AOI22_X1 U9716 ( .A1(n10412), .A2(n10411), .B1(n9683), .B2(n9682), .ZN(
        n10488) );
  INV_X1 U9717 ( .A(n12495), .ZN(n7944) );
  AND2_X1 U9718 ( .A1(n7693), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7444) );
  INV_X1 U9719 ( .A(n13097), .ZN(n13121) );
  AND2_X1 U9720 ( .A1(n10402), .A2(n7942), .ZN(n7446) );
  AND2_X1 U9721 ( .A1(n9734), .A2(n9733), .ZN(n7447) );
  AND2_X1 U9722 ( .A1(n9014), .A2(P1_U3086), .ZN(n11861) );
  INV_X1 U9723 ( .A(n12315), .ZN(n11565) );
  INV_X1 U9724 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9004) );
  OR2_X1 U9725 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10143), .ZN(n7448) );
  INV_X1 U9726 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8249) );
  AND2_X1 U9727 ( .A1(n9842), .A2(P1_U3086), .ZN(n10409) );
  AND3_X1 U9728 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(n8794) );
  INV_X1 U9729 ( .A(n11137), .ZN(n11152) );
  NAND2_X2 U9730 ( .A1(n12022), .A2(n14374), .ZN(n14377) );
  NAND2_X2 U9731 ( .A1(n10522), .A2(n13651), .ZN(n15210) );
  INV_X1 U9732 ( .A(n13272), .ZN(n9485) );
  INV_X1 U9733 ( .A(n14651), .ZN(n9757) );
  INV_X1 U9734 ( .A(n11914), .ZN(n11930) );
  AND2_X1 U9735 ( .A1(n9398), .A2(n9397), .ZN(n7449) );
  AND2_X1 U9736 ( .A1(n12067), .A2(n12066), .ZN(n12068) );
  AOI22_X1 U9737 ( .A1(n6734), .A2(n6459), .B1(n12076), .B2(n12228), .ZN(
        n12079) );
  AOI22_X1 U9738 ( .A1(n13295), .A2(n12103), .B1(n12073), .B2(n12228), .ZN(
        n12083) );
  OR2_X1 U9739 ( .A1(n12084), .A2(n12083), .ZN(n12085) );
  OAI22_X1 U9740 ( .A1(n12088), .A2(n12228), .B1(n12087), .B2(n12254), .ZN(
        n12090) );
  OAI22_X1 U9741 ( .A1(n14897), .A2(n12277), .B1(n12123), .B2(n12276), .ZN(
        n12125) );
  AOI22_X1 U9742 ( .A1(n13655), .A2(n12277), .B1(n12276), .B2(n13287), .ZN(
        n12138) );
  NAND2_X1 U9743 ( .A1(n12162), .A2(n12161), .ZN(n12163) );
  AOI22_X1 U9744 ( .A1(n14620), .A2(n12277), .B1(n12254), .B2(n13388), .ZN(
        n12165) );
  OAI22_X1 U9745 ( .A1(n13578), .A2(n12276), .B1(n13247), .B2(n12277), .ZN(
        n12184) );
  MUX2_X1 U9746 ( .A(n14255), .B(n14425), .S(n8795), .Z(n8644) );
  OAI22_X1 U9747 ( .A1(n13526), .A2(n12276), .B1(n13233), .B2(n12277), .ZN(
        n12197) );
  INV_X1 U9748 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8055) );
  INV_X1 U9749 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8962) );
  INV_X1 U9750 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7453) );
  INV_X1 U9751 ( .A(n9387), .ZN(n8957) );
  OR4_X1 U9752 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9451) );
  XNOR2_X1 U9753 ( .A(n14210), .B(n14021), .ZN(n8787) );
  INV_X1 U9754 ( .A(n8446), .ZN(n8448) );
  INV_X1 U9755 ( .A(n12507), .ZN(n7959) );
  INV_X1 U9756 ( .A(n9354), .ZN(n8956) );
  INV_X1 U9757 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U9758 ( .A1(n8957), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9401) );
  INV_X1 U9759 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9248) );
  INV_X1 U9760 ( .A(n9314), .ZN(n8954) );
  INV_X1 U9761 ( .A(n9271), .ZN(n8952) );
  XNOR2_X1 U9762 ( .A(n14392), .B(n8794), .ZN(n8786) );
  INV_X1 U9763 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8316) );
  INV_X1 U9764 ( .A(n14276), .ZN(n11999) );
  INV_X1 U9765 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U9766 ( .A1(n11271), .A2(n11272), .ZN(n11270) );
  INV_X1 U9767 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8064) );
  INV_X1 U9768 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U9769 ( .A1(n8130), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8099) );
  INV_X1 U9770 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7559) );
  INV_X1 U9771 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7489) );
  INV_X1 U9772 ( .A(n7884), .ZN(n7883) );
  OR2_X1 U9773 ( .A1(n7843), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7855) );
  INV_X1 U9774 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12416) );
  INV_X1 U9775 ( .A(n12498), .ZN(n7948) );
  NOR2_X1 U9776 ( .A1(n8027), .A2(n8026), .ZN(n8040) );
  INV_X1 U9777 ( .A(n7930), .ZN(n7931) );
  AND2_X1 U9778 ( .A1(n7585), .A2(n7569), .ZN(n7570) );
  OR2_X1 U9779 ( .A1(n9435), .A2(n9507), .ZN(n9489) );
  OR2_X1 U9780 ( .A1(n9401), .A2(n13218), .ZN(n9415) );
  OR2_X1 U9781 ( .A1(n9341), .A2(n8955), .ZN(n9354) );
  INV_X1 U9782 ( .A(n12235), .ZN(n12218) );
  NAND2_X1 U9783 ( .A1(n8954), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9341) );
  AND2_X1 U9784 ( .A1(n10523), .A2(n12295), .ZN(n15201) );
  INV_X1 U9785 ( .A(n6456), .ZN(n13924) );
  OR2_X1 U9786 ( .A1(n8687), .A2(n13929), .ZN(n12021) );
  INV_X1 U9787 ( .A(n8575), .ZN(n8576) );
  NOR2_X1 U9788 ( .A1(n8359), .A2(n8358), .ZN(n8383) );
  NAND2_X1 U9789 ( .A1(n12000), .A2(n11999), .ZN(n12001) );
  INV_X2 U9790 ( .A(n8656), .ZN(n8758) );
  INV_X1 U9791 ( .A(n10719), .ZN(n11446) );
  INV_X1 U9792 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8065) );
  INV_X1 U9793 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8167) );
  INV_X1 U9794 ( .A(n8165), .ZN(n8168) );
  AOI22_X1 U9795 ( .A1(n9600), .A2(n9539), .B1(P1_ADDR_REG_14__SCAN_IN), .B2(
        n11714), .ZN(n9601) );
  INV_X1 U9796 ( .A(n8832), .ZN(n12422) );
  OR2_X1 U9797 ( .A1(n13127), .A2(n8919), .ZN(n10131) );
  INV_X1 U9798 ( .A(n12871), .ZN(n8900) );
  INV_X1 U9799 ( .A(n12980), .ZN(n12409) );
  AND2_X1 U9800 ( .A1(n8008), .A2(n8013), .ZN(n8919) );
  INV_X1 U9801 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n11908) );
  INV_X1 U9802 ( .A(n9638), .ZN(n9639) );
  NAND2_X1 U9803 ( .A1(n7883), .A2(n7882), .ZN(n7895) );
  NAND2_X1 U9804 ( .A1(n12416), .A2(n7776), .ZN(n7795) );
  INV_X1 U9805 ( .A(n14996), .ZN(n12675) );
  OR2_X1 U9806 ( .A1(n12817), .A2(n12816), .ZN(n13044) );
  AND2_X1 U9807 ( .A1(n12620), .A2(n12615), .ZN(n12618) );
  AND2_X1 U9808 ( .A1(n12592), .A2(n12583), .ZN(n14595) );
  INV_X1 U9809 ( .A(n12690), .ZN(n12528) );
  AND2_X1 U9810 ( .A1(n7801), .A2(n7787), .ZN(n7788) );
  AND2_X1 U9811 ( .A1(n7733), .A2(n7718), .ZN(n7719) );
  OR2_X1 U9812 ( .A1(n13423), .A2(n9492), .ZN(n9497) );
  INV_X1 U9813 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U9814 ( .A1(n13379), .A2(n13542), .B1(n13378), .B2(n13377), .ZN(
        n13380) );
  NAND2_X1 U9815 ( .A1(n15210), .A2(n15201), .ZN(n13603) );
  INV_X1 U9816 ( .A(n13639), .ZN(n13620) );
  INV_X1 U9817 ( .A(n14901), .ZN(n14903) );
  NAND2_X1 U9818 ( .A1(n9500), .A2(n9861), .ZN(n13632) );
  INV_X1 U9819 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9457) );
  AND2_X1 U9820 ( .A1(n13968), .A2(n13851), .ZN(n13898) );
  INV_X1 U9821 ( .A(n14024), .ZN(n14005) );
  INV_X1 U9822 ( .A(n9684), .ZN(n13868) );
  INV_X1 U9823 ( .A(n8072), .ZN(n8071) );
  INV_X1 U9824 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14123) );
  INV_X1 U9825 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14138) );
  OR2_X1 U9826 ( .A1(n10662), .A2(n10661), .ZN(n10853) );
  INV_X1 U9827 ( .A(n11974), .ZN(n14270) );
  INV_X1 U9828 ( .A(n14739), .ZN(n14474) );
  INV_X1 U9829 ( .A(n11355), .ZN(n11345) );
  INV_X1 U9830 ( .A(n11621), .ZN(n11488) );
  OR2_X1 U9831 ( .A1(n11265), .A2(n14765), .ZN(n11253) );
  NAND2_X1 U9832 ( .A1(n11445), .A2(n10720), .ZN(n10722) );
  NAND2_X2 U9833 ( .A1(n9770), .A2(n9794), .ZN(n14374) );
  AND2_X1 U9834 ( .A1(n8138), .A2(n14195), .ZN(n11196) );
  INV_X1 U9835 ( .A(n14322), .ZN(n14462) );
  INV_X1 U9836 ( .A(n11768), .ZN(n14669) );
  NAND2_X1 U9837 ( .A1(n14536), .A2(n9655), .ZN(n10334) );
  XNOR2_X1 U9838 ( .A(n8535), .B(SI_19_), .ZN(n8536) );
  INV_X1 U9839 ( .A(n8163), .ZN(n8160) );
  INV_X1 U9840 ( .A(n8135), .ZN(n8132) );
  OAI21_X1 U9841 ( .B1(n9625), .B2(n12459), .A(n8942), .ZN(n8943) );
  INV_X1 U9842 ( .A(n12455), .ZN(n12463) );
  NOR2_X1 U9843 ( .A1(n10131), .A2(n15026), .ZN(n10354) );
  AND4_X1 U9844 ( .A1(n12477), .A2(n12476), .A3(n12475), .A4(n12474), .ZN(
        n12817) );
  AND4_X1 U9845 ( .A1(n7871), .A2(n7870), .A3(n7869), .A4(n7868), .ZN(n12903)
         );
  AND4_X1 U9846 ( .A1(n7848), .A2(n7847), .A3(n7846), .A4(n7845), .ZN(n12902)
         );
  AND4_X1 U9847 ( .A1(n7697), .A2(n7696), .A3(n7695), .A4(n7694), .ZN(n11818)
         );
  INV_X1 U9848 ( .A(n14966), .ZN(n14954) );
  INV_X1 U9849 ( .A(n12956), .ZN(n14987) );
  INV_X1 U9850 ( .A(n12997), .ZN(n14599) );
  INV_X1 U9851 ( .A(n13027), .ZN(n8048) );
  AND2_X1 U9852 ( .A1(n8042), .A2(n8041), .ZN(n10353) );
  AND2_X1 U9853 ( .A1(n12971), .A2(n12970), .ZN(n13107) );
  OR2_X1 U9854 ( .A1(n15029), .A2(n15023), .ZN(n15032) );
  NOR2_X1 U9855 ( .A1(n14996), .A2(n12690), .ZN(n15023) );
  INV_X1 U9856 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7997) );
  OR2_X1 U9857 ( .A1(n13199), .A2(n13630), .ZN(n13277) );
  INV_X1 U9858 ( .A(n13276), .ZN(n13240) );
  INV_X1 U9859 ( .A(n12109), .ZN(n14888) );
  AND2_X1 U9860 ( .A1(n9394), .A2(n9393), .ZN(n13406) );
  AND3_X1 U9861 ( .A1(n9275), .A2(n9274), .A3(n9273), .ZN(n13389) );
  AND2_X1 U9862 ( .A1(n9886), .A2(n9873), .ZN(n14868) );
  INV_X1 U9863 ( .A(n13380), .ZN(n13381) );
  INV_X1 U9864 ( .A(n13347), .ZN(n13454) );
  AND2_X1 U9865 ( .A1(n13369), .A2(n12294), .ZN(n13516) );
  INV_X1 U9866 ( .A(n12306), .ZN(n11283) );
  INV_X1 U9867 ( .A(n13641), .ZN(n13658) );
  AND2_X1 U9868 ( .A1(n10088), .A2(n14903), .ZN(n13734) );
  INV_X1 U9869 ( .A(n13734), .ZN(n14623) );
  AND2_X1 U9870 ( .A1(n9478), .A2(n9470), .ZN(n14873) );
  INV_X1 U9871 ( .A(n11863), .ZN(n8819) );
  AND3_X1 U9872 ( .A1(n8549), .A2(n8548), .A3(n8547), .ZN(n13939) );
  AND3_X1 U9873 ( .A1(n8517), .A2(n8516), .A3(n8515), .ZN(n13964) );
  INV_X1 U9874 ( .A(n14190), .ZN(n14724) );
  INV_X1 U9875 ( .A(n12016), .ZN(n12013) );
  INV_X1 U9876 ( .A(n11278), .ZN(n14254) );
  AND2_X1 U9877 ( .A1(n14377), .A2(n10798), .ZN(n14384) );
  INV_X1 U9878 ( .A(n14793), .ZN(n14775) );
  INV_X1 U9879 ( .A(n14799), .ZN(n14753) );
  NAND2_X1 U9880 ( .A1(n11278), .A2(n14430), .ZN(n14799) );
  NAND3_X1 U9881 ( .A1(n9774), .A2(n9773), .A3(n9789), .ZN(n10714) );
  INV_X1 U9882 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n9558) );
  AND2_X1 U9883 ( .A1(n10134), .A2(n10133), .ZN(n14923) );
  INV_X1 U9884 ( .A(n12662), .ZN(n12848) );
  NAND2_X1 U9885 ( .A1(n8915), .A2(n10354), .ZN(n12459) );
  AND4_X1 U9886 ( .A1(n12477), .A2(n8934), .A3(n8933), .A4(n8932), .ZN(n12837)
         );
  INV_X1 U9887 ( .A(n12902), .ZN(n12927) );
  INV_X1 U9888 ( .A(n11390), .ZN(n14590) );
  INV_X1 U9889 ( .A(n14936), .ZN(n14975) );
  OR2_X1 U9890 ( .A1(n10141), .A2(n10135), .ZN(n14983) );
  OR2_X1 U9891 ( .A1(n10141), .A2(n12688), .ZN(n14977) );
  OR2_X1 U9892 ( .A1(n15004), .A2(n10623), .ZN(n12997) );
  INV_X1 U9893 ( .A(n15004), .ZN(n15002) );
  NAND2_X1 U9894 ( .A1(n15051), .A2(n15032), .ZN(n13043) );
  INV_X1 U9895 ( .A(n15051), .ZN(n15049) );
  NAND2_X1 U9896 ( .A1(n15051), .A2(n15015), .ZN(n13027) );
  OR2_X1 U9897 ( .A1(n15037), .A2(n14603), .ZN(n13125) );
  AND3_X1 U9898 ( .A1(n15036), .A2(n15035), .A3(n15034), .ZN(n15050) );
  AND2_X2 U9899 ( .A1(n8031), .A2(n8030), .ZN(n15037) );
  OR2_X1 U9900 ( .A1(n15037), .A2(n15026), .ZN(n13097) );
  INV_X1 U9901 ( .A(SI_24_), .ZN(n15168) );
  INV_X1 U9902 ( .A(SI_13_), .ZN(n9964) );
  NAND2_X1 U9903 ( .A1(n7618), .A2(n7617), .ZN(n10908) );
  INV_X1 U9904 ( .A(n13261), .ZN(n13278) );
  NAND2_X1 U9905 ( .A1(n9498), .A2(n9484), .ZN(n13272) );
  INV_X1 U9906 ( .A(n13436), .ZN(n13379) );
  INV_X1 U9907 ( .A(n13403), .ZN(n13524) );
  INV_X1 U9908 ( .A(n14865), .ZN(n11825) );
  OR2_X1 U9909 ( .A1(n9886), .A2(P2_U3088), .ZN(n14857) );
  NAND2_X1 U9910 ( .A1(n15210), .A2(n10695), .ZN(n13627) );
  INV_X1 U9911 ( .A(n14922), .ZN(n14920) );
  INV_X1 U9912 ( .A(n13446), .ZN(n13759) );
  NOR2_X1 U9913 ( .A1(n14878), .A2(n14873), .ZN(n14874) );
  INV_X1 U9914 ( .A(n14874), .ZN(n14875) );
  INV_X1 U9915 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n15180) );
  INV_X1 U9916 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10448) );
  NAND2_X1 U9917 ( .A1(n9799), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14707) );
  INV_X1 U9918 ( .A(n14449), .ZN(n14300) );
  INV_X1 U9919 ( .A(n14653), .ZN(n14015) );
  INV_X1 U9920 ( .A(n8794), .ZN(n14204) );
  INV_X1 U9921 ( .A(n13939), .ZN(n14027) );
  INV_X1 U9922 ( .A(n11920), .ZN(n14029) );
  INV_X1 U9923 ( .A(n14194), .ZN(n14729) );
  INV_X1 U9924 ( .A(n14733), .ZN(n14199) );
  INV_X1 U9925 ( .A(n14337), .ZN(n14391) );
  INV_X2 U9926 ( .A(n14811), .ZN(n14813) );
  AND2_X1 U9927 ( .A1(n14780), .A2(n14779), .ZN(n14809) );
  AND2_X1 U9928 ( .A1(n14771), .A2(n14770), .ZN(n14808) );
  INV_X1 U9929 ( .A(n9905), .ZN(n9857) );
  INV_X1 U9930 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10835) );
  INV_X1 U9931 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10359) );
  XNOR2_X1 U9932 ( .A(n9622), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n9623) );
  INV_X1 U9933 ( .A(n12706), .ZN(P3_U3897) );
  NOR2_X1 U9934 ( .A1(n9866), .A2(n9653), .ZN(P2_U3947) );
  INV_X1 U9935 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8032) );
  NOR2_X1 U9936 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7451) );
  NAND3_X1 U9937 ( .A1(n7459), .A2(n7458), .A3(n7457), .ZN(n7470) );
  INV_X1 U9938 ( .A(n7464), .ZN(n7462) );
  NAND2_X1 U9939 ( .A1(n7462), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U9940 ( .A1(n7993), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7465) );
  NOR2_X2 U9941 ( .A1(n7470), .A2(n7469), .ZN(n8002) );
  AND2_X2 U9942 ( .A1(n7486), .A2(n6644), .ZN(n7475) );
  INV_X1 U9943 ( .A(n7475), .ZN(n7488) );
  NAND2_X1 U9944 ( .A1(n7488), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7476) );
  NAND2_X1 U9945 ( .A1(n7510), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U9946 ( .A1(n12473), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7482) );
  NAND2_X1 U9947 ( .A1(n6481), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7481) );
  INV_X1 U9948 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7495) );
  NAND2_X2 U9949 ( .A1(n7498), .A2(n7497), .ZN(n8130) );
  INV_X2 U9950 ( .A(n8130), .ZN(n7499) );
  INV_X1 U9951 ( .A(SI_0_), .ZN(n9817) );
  OR2_X1 U9952 ( .A1(n7515), .A2(n9817), .ZN(n7501) );
  INV_X1 U9953 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U9954 ( .A1(n8102), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7516) );
  INV_X1 U9955 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U9956 ( .A1(n8103), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7500) );
  AND2_X1 U9957 ( .A1(n7516), .A2(n7500), .ZN(n9818) );
  NAND2_X1 U9958 ( .A1(n7510), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7505) );
  NAND2_X1 U9959 ( .A1(n7662), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U9960 ( .A1(n6481), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7502) );
  INV_X1 U9961 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U9962 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7506) );
  XNOR2_X1 U9963 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7518) );
  XNOR2_X1 U9964 ( .A(n7516), .B(n7518), .ZN(n9825) );
  NAND2_X1 U9965 ( .A1(n6650), .A2(n8834), .ZN(n12532) );
  NAND2_X1 U9966 ( .A1(n8833), .A2(n12532), .ZN(n10507) );
  NAND2_X1 U9967 ( .A1(n7510), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7514) );
  NAND2_X1 U9968 ( .A1(n7662), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7513) );
  NAND2_X1 U9969 ( .A1(n12473), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7512) );
  OR2_X1 U9970 ( .A1(n12487), .A2(SI_2_), .ZN(n7526) );
  INV_X1 U9971 ( .A(n7516), .ZN(n7517) );
  INV_X1 U9972 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U9973 ( .A1(n9902), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U9974 ( .A1(n9843), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7534) );
  INV_X1 U9975 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U9976 ( .A1(n9807), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7520) );
  AND2_X1 U9977 ( .A1(n7534), .A2(n7520), .ZN(n7532) );
  XNOR2_X1 U9978 ( .A(n7533), .B(n7532), .ZN(n9826) );
  OR2_X1 U9979 ( .A1(n7840), .A2(n9826), .ZN(n7525) );
  INV_X2 U9980 ( .A(n7980), .ZN(n10129) );
  NAND2_X1 U9981 ( .A1(n10129), .A2(n6453), .ZN(n7524) );
  NAND2_X1 U9982 ( .A1(n10402), .A2(n10606), .ZN(n12537) );
  INV_X1 U9983 ( .A(n10606), .ZN(n7942) );
  NAND2_X1 U9984 ( .A1(n14989), .A2(n7942), .ZN(n12536) );
  NAND2_X1 U9985 ( .A1(n10507), .A2(n12534), .ZN(n10506) );
  NAND2_X1 U9986 ( .A1(n7510), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7531) );
  INV_X1 U9987 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U9988 ( .A1(n7662), .A2(n7527), .ZN(n7530) );
  NAND2_X1 U9989 ( .A1(n12473), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U9990 ( .A1(n6481), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7528) );
  AND4_X2 U9991 ( .A1(n7531), .A2(n7530), .A3(n7529), .A4(n7528), .ZN(n10629)
         );
  OR2_X1 U9992 ( .A1(n12487), .A2(SI_3_), .ZN(n7543) );
  NAND2_X1 U9993 ( .A1(n7533), .A2(n7532), .ZN(n7535) );
  NAND2_X1 U9994 ( .A1(n7535), .A2(n7534), .ZN(n7538) );
  NAND2_X1 U9995 ( .A1(n9895), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7548) );
  INV_X1 U9996 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U9997 ( .A1(n9811), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7536) );
  AND2_X1 U9998 ( .A1(n7548), .A2(n7536), .ZN(n7537) );
  OR2_X1 U9999 ( .A1(n7538), .A2(n7537), .ZN(n7539) );
  NAND2_X1 U10000 ( .A1(n7549), .A2(n7539), .ZN(n9829) );
  OR2_X1 U10001 ( .A1(n7840), .A2(n9829), .ZN(n7542) );
  OR2_X1 U10002 ( .A1(n7552), .A2(n7485), .ZN(n7540) );
  NAND2_X1 U10003 ( .A1(n10129), .A2(n10185), .ZN(n7541) );
  AND3_X2 U10004 ( .A1(n7543), .A2(n7542), .A3(n7541), .ZN(n10584) );
  INV_X1 U10005 ( .A(n10584), .ZN(n10828) );
  AND2_X1 U10006 ( .A1(n12544), .A2(n12545), .ZN(n12495) );
  NAND2_X1 U10007 ( .A1(n6449), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7547) );
  NAND2_X1 U10008 ( .A1(n6447), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7546) );
  XNOR2_X1 U10009 ( .A(P3_REG3_REG_4__SCAN_IN), .B(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n10633) );
  NAND2_X1 U10010 ( .A1(n8930), .A2(n10633), .ZN(n7545) );
  NAND2_X1 U10011 ( .A1(n8931), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7544) );
  AND4_X2 U10012 ( .A1(n7547), .A2(n7546), .A3(n7545), .A4(n7544), .ZN(n10885)
         );
  OR2_X1 U10013 ( .A1(n12487), .A2(SI_4_), .ZN(n7558) );
  NAND2_X1 U10014 ( .A1(n10162), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7568) );
  INV_X1 U10015 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U10016 ( .A1(n9840), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7550) );
  XNOR2_X1 U10017 ( .A(n7567), .B(n7566), .ZN(n9819) );
  OR2_X1 U10018 ( .A1(n7840), .A2(n9819), .ZN(n7557) );
  NAND2_X1 U10019 ( .A1(n7554), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7553) );
  MUX2_X1 U10020 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7553), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7555) );
  NAND2_X1 U10021 ( .A1(n10129), .A2(n10240), .ZN(n7556) );
  NAND2_X1 U10022 ( .A1(n10885), .A2(n10672), .ZN(n12550) );
  INV_X1 U10023 ( .A(n10672), .ZN(n10675) );
  NAND2_X1 U10024 ( .A1(n6449), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7565) );
  NAND2_X1 U10025 ( .A1(n6447), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7564) );
  NOR2_X1 U10026 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7560) );
  NAND2_X1 U10027 ( .A1(n7560), .A2(n7559), .ZN(n7577) );
  OR2_X1 U10028 ( .A1(n7560), .A2(n7559), .ZN(n7561) );
  NAND2_X1 U10029 ( .A1(n7577), .A2(n7561), .ZN(n10888) );
  NAND2_X1 U10030 ( .A1(n8930), .A2(n10888), .ZN(n7563) );
  NAND2_X1 U10031 ( .A1(n8931), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7562) );
  AND4_X2 U10032 ( .A1(n7565), .A2(n7564), .A3(n7563), .A4(n7562), .ZN(n11002)
         );
  OR2_X1 U10033 ( .A1(n12487), .A2(SI_5_), .ZN(n7576) );
  NAND2_X1 U10034 ( .A1(n9860), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U10035 ( .A1(n9850), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7569) );
  NAND2_X1 U10036 ( .A1(n7571), .A2(n7570), .ZN(n7586) );
  OR2_X1 U10037 ( .A1(n7571), .A2(n7570), .ZN(n7572) );
  NAND2_X1 U10038 ( .A1(n7586), .A2(n7572), .ZN(n9808) );
  OR2_X1 U10039 ( .A1(n7840), .A2(n9808), .ZN(n7575) );
  NAND2_X1 U10040 ( .A1(n7583), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U10041 ( .A1(n10129), .A2(n10243), .ZN(n7574) );
  NAND2_X1 U10042 ( .A1(n11002), .A2(n11011), .ZN(n12553) );
  NAND2_X1 U10043 ( .A1(n12703), .A2(n11014), .ZN(n12556) );
  AND2_X2 U10044 ( .A1(n12553), .A2(n12556), .ZN(n12552) );
  NAND2_X1 U10045 ( .A1(n6449), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7582) );
  NAND2_X1 U10046 ( .A1(n6447), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U10047 ( .A1(n7577), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7578) );
  NAND2_X1 U10048 ( .A1(n7590), .A2(n7578), .ZN(n11117) );
  NAND2_X1 U10049 ( .A1(n8930), .A2(n11117), .ZN(n7580) );
  NAND2_X1 U10050 ( .A1(n8931), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7579) );
  OR2_X1 U10051 ( .A1(n7603), .A2(n7485), .ZN(n7584) );
  XNOR2_X1 U10052 ( .A(n7584), .B(n7602), .ZN(n10552) );
  NAND2_X1 U10053 ( .A1(n7586), .A2(n7585), .ZN(n7597) );
  XNOR2_X1 U10054 ( .A(n9897), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7587) );
  XNOR2_X1 U10055 ( .A(n7597), .B(n7587), .ZN(n9816) );
  OR2_X1 U10056 ( .A1(n6646), .A2(n9816), .ZN(n7589) );
  INV_X1 U10057 ( .A(SI_6_), .ZN(n9815) );
  OR2_X1 U10058 ( .A1(n12487), .A2(n9815), .ZN(n7588) );
  OAI211_X1 U10059 ( .C1(n7980), .C2(n10552), .A(n7589), .B(n7588), .ZN(n11066) );
  NAND2_X1 U10060 ( .A1(n11025), .A2(n11066), .ZN(n12560) );
  INV_X1 U10061 ( .A(n11066), .ZN(n11110) );
  NAND2_X1 U10062 ( .A1(n12702), .A2(n11110), .ZN(n12558) );
  NAND2_X1 U10063 ( .A1(n10999), .A2(n12498), .ZN(n10998) );
  NAND2_X1 U10064 ( .A1(n6449), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U10065 ( .A1(n6447), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7594) );
  AND2_X1 U10066 ( .A1(n7590), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7591) );
  OR2_X1 U10067 ( .A1(n7591), .A2(n7608), .ZN(n11057) );
  NAND2_X1 U10068 ( .A1(n8930), .A2(n11057), .ZN(n7593) );
  NAND2_X1 U10069 ( .A1(n8931), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7592) );
  NAND2_X1 U10070 ( .A1(n9852), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7596) );
  NAND2_X1 U10071 ( .A1(n7597), .A2(n7596), .ZN(n7599) );
  NAND2_X1 U10072 ( .A1(n9897), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7598) );
  NAND2_X1 U10073 ( .A1(n9899), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7622) );
  INV_X1 U10074 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7600) );
  NAND2_X1 U10075 ( .A1(n7600), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7601) );
  XNOR2_X1 U10076 ( .A(n7621), .B(n7619), .ZN(n9822) );
  OR2_X1 U10077 ( .A1(n6646), .A2(n9822), .ZN(n7607) );
  OR2_X1 U10078 ( .A1(n12487), .A2(SI_7_), .ZN(n7606) );
  NAND2_X1 U10079 ( .A1(n7603), .A2(n7602), .ZN(n7614) );
  NAND2_X1 U10080 ( .A1(n7614), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7604) );
  XNOR2_X1 U10081 ( .A(n7604), .B(n7311), .ZN(n14932) );
  NAND2_X1 U10082 ( .A1(n10129), .A2(n14932), .ZN(n7605) );
  NAND2_X1 U10083 ( .A1(n11001), .A2(n15014), .ZN(n12564) );
  INV_X1 U10084 ( .A(n15014), .ZN(n11055) );
  NAND2_X1 U10085 ( .A1(n12701), .A2(n11055), .ZN(n12565) );
  NAND2_X1 U10086 ( .A1(n12564), .A2(n12565), .ZN(n12561) );
  INV_X1 U10087 ( .A(n12561), .ZN(n12502) );
  NAND2_X1 U10088 ( .A1(n6449), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U10089 ( .A1(n6447), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7612) );
  NOR2_X1 U10090 ( .A1(n7608), .A2(n10551), .ZN(n7609) );
  OR2_X1 U10091 ( .A1(n7630), .A2(n7609), .ZN(n12382) );
  NAND2_X1 U10092 ( .A1(n8930), .A2(n12382), .ZN(n7611) );
  NAND2_X1 U10093 ( .A1(n8931), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7610) );
  INV_X1 U10094 ( .A(n7655), .ZN(n7618) );
  NAND2_X1 U10095 ( .A1(n7615), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7616) );
  MUX2_X1 U10096 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7616), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n7617) );
  INV_X1 U10097 ( .A(n7619), .ZN(n7620) );
  NAND2_X1 U10098 ( .A1(n9987), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7636) );
  NAND2_X1 U10099 ( .A1(n10166), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7623) );
  OR2_X1 U10100 ( .A1(n7625), .A2(n7624), .ZN(n7626) );
  NAND2_X1 U10101 ( .A1(n7637), .A2(n7626), .ZN(n9814) );
  OR2_X1 U10102 ( .A1(n6646), .A2(n9814), .ZN(n7628) );
  INV_X1 U10103 ( .A(SI_8_), .ZN(n9813) );
  OR2_X1 U10104 ( .A1(n12487), .A2(n9813), .ZN(n7627) );
  OAI211_X1 U10105 ( .C1(n7980), .C2(n10908), .A(n7628), .B(n7627), .ZN(n12381) );
  NAND2_X1 U10106 ( .A1(n11391), .A2(n12381), .ZN(n12570) );
  INV_X1 U10107 ( .A(n12381), .ZN(n11471) );
  NAND2_X1 U10108 ( .A1(n12700), .A2(n11471), .ZN(n12569) );
  NAND2_X1 U10109 ( .A1(n12570), .A2(n12569), .ZN(n11465) );
  INV_X1 U10110 ( .A(n11465), .ZN(n12567) );
  NAND2_X1 U10111 ( .A1(n6449), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U10112 ( .A1(n6447), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7634) );
  OR2_X1 U10113 ( .A1(n7630), .A2(n7629), .ZN(n7631) );
  NAND2_X1 U10114 ( .A1(n7660), .A2(n7631), .ZN(n11395) );
  NAND2_X1 U10115 ( .A1(n8930), .A2(n11395), .ZN(n7633) );
  NAND2_X1 U10116 ( .A1(n8931), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7632) );
  NAND4_X1 U10117 ( .A1(n7635), .A2(n7634), .A3(n7633), .A4(n7632), .ZN(n12699) );
  NAND2_X1 U10118 ( .A1(n10013), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7648) );
  NAND2_X1 U10119 ( .A1(n10164), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7638) );
  OR2_X1 U10120 ( .A1(n7640), .A2(n7639), .ZN(n7641) );
  NAND2_X1 U10121 ( .A1(n7649), .A2(n7641), .ZN(n9833) );
  NAND2_X1 U10122 ( .A1(n9833), .A2(n12486), .ZN(n7644) );
  INV_X1 U10123 ( .A(SI_9_), .ZN(n9832) );
  OR2_X1 U10124 ( .A1(n7655), .A2(n7485), .ZN(n7642) );
  XNOR2_X1 U10125 ( .A(n7642), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11330) );
  INV_X1 U10126 ( .A(n11330), .ZN(n10898) );
  AOI22_X1 U10127 ( .A1(n9629), .A2(n9832), .B1(n10898), .B2(n10129), .ZN(
        n7643) );
  INV_X1 U10128 ( .A(n12574), .ZN(n15027) );
  NAND2_X1 U10129 ( .A1(n12699), .A2(n15027), .ZN(n7645) );
  NAND2_X1 U10130 ( .A1(n11399), .A2(n7645), .ZN(n7647) );
  INV_X1 U10131 ( .A(n12699), .ZN(n8860) );
  NAND2_X1 U10132 ( .A1(n8860), .A2(n12574), .ZN(n7646) );
  NAND2_X1 U10133 ( .A1(n7647), .A2(n7646), .ZN(n11497) );
  NAND2_X1 U10134 ( .A1(n10080), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U10135 ( .A1(n10082), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7650) );
  OR2_X1 U10136 ( .A1(n7652), .A2(n7651), .ZN(n7653) );
  NAND2_X1 U10137 ( .A1(n7668), .A2(n7653), .ZN(n9835) );
  NAND2_X1 U10138 ( .A1(n9835), .A2(n12486), .ZN(n7659) );
  INV_X1 U10139 ( .A(SI_10_), .ZN(n9834) );
  INV_X1 U10140 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7654) );
  NAND2_X1 U10141 ( .A1(n7655), .A2(n7654), .ZN(n7673) );
  NAND2_X1 U10142 ( .A1(n7673), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7657) );
  INV_X1 U10143 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7656) );
  AOI22_X1 U10144 ( .A1(n9629), .A2(n9834), .B1(n10129), .B2(n14944), .ZN(
        n7658) );
  INV_X1 U10145 ( .A(n11498), .ZN(n12365) );
  NAND2_X1 U10146 ( .A1(n6449), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7666) );
  NAND2_X1 U10147 ( .A1(n7510), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7665) );
  NAND2_X1 U10148 ( .A1(n7660), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U10149 ( .A1(n7676), .A2(n7661), .ZN(n12364) );
  NAND2_X1 U10150 ( .A1(n8930), .A2(n12364), .ZN(n7664) );
  NAND2_X1 U10151 ( .A1(n8931), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7663) );
  NAND2_X1 U10152 ( .A1(n12365), .A2(n14590), .ZN(n12580) );
  NAND2_X1 U10153 ( .A1(n11498), .A2(n11390), .ZN(n12582) );
  NAND2_X1 U10154 ( .A1(n10107), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7682) );
  NAND2_X1 U10155 ( .A1(n10109), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7669) );
  OR2_X1 U10156 ( .A1(n7671), .A2(n7670), .ZN(n7672) );
  NAND2_X1 U10157 ( .A1(n7683), .A2(n7672), .ZN(n9848) );
  OAI21_X1 U10158 ( .B1(n7673), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7674) );
  XNOR2_X1 U10159 ( .A(n7674), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11413) );
  OAI22_X1 U10160 ( .A1(n11413), .A2(n7980), .B1(n12487), .B2(SI_11_), .ZN(
        n7675) );
  AOI21_X1 U10161 ( .B1(n9848), .B2(n12486), .A(n7675), .ZN(n11639) );
  INV_X1 U10162 ( .A(n11639), .ZN(n14597) );
  NAND2_X1 U10163 ( .A1(n6447), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U10164 ( .A1(n7676), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U10165 ( .A1(n7693), .A2(n7677), .ZN(n14593) );
  NAND2_X1 U10166 ( .A1(n8930), .A2(n14593), .ZN(n7680) );
  NAND2_X1 U10167 ( .A1(n8931), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U10168 ( .A1(n6449), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7678) );
  OR2_X1 U10169 ( .A1(n14597), .A2(n14576), .ZN(n12592) );
  NAND2_X1 U10170 ( .A1(n14597), .A2(n14576), .ZN(n12583) );
  NAND2_X1 U10171 ( .A1(n10359), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7698) );
  NAND2_X1 U10172 ( .A1(n15054), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7684) );
  OR2_X1 U10173 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  NAND2_X1 U10174 ( .A1(n7699), .A2(n7687), .ZN(n9855) );
  OR2_X1 U10175 ( .A1(n9855), .A2(n6646), .ZN(n7692) );
  NAND2_X1 U10176 ( .A1(n7688), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7689) );
  MUX2_X1 U10177 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7689), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7690) );
  AND2_X1 U10178 ( .A1(n7690), .A2(n7703), .ZN(n11416) );
  AOI22_X1 U10179 ( .A1(n9629), .A2(SI_12_), .B1(n10129), .B2(n11416), .ZN(
        n7691) );
  NAND2_X1 U10180 ( .A1(n7692), .A2(n7691), .ZN(n14585) );
  NAND2_X1 U10181 ( .A1(n6447), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7697) );
  NOR2_X1 U10182 ( .A1(n7709), .A2(n7444), .ZN(n14579) );
  INV_X1 U10183 ( .A(n14579), .ZN(n11724) );
  NAND2_X1 U10184 ( .A1(n8930), .A2(n11724), .ZN(n7696) );
  NAND2_X1 U10185 ( .A1(n8931), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U10186 ( .A1(n6449), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7694) );
  OR2_X1 U10187 ( .A1(n14585), .A2(n11818), .ZN(n12589) );
  NAND2_X1 U10188 ( .A1(n14585), .A2(n11818), .ZN(n12593) );
  NAND2_X1 U10189 ( .A1(n12589), .A2(n12593), .ZN(n7956) );
  INV_X1 U10190 ( .A(n7700), .ZN(n7701) );
  NAND2_X1 U10191 ( .A1(n7701), .A2(n10448), .ZN(n7702) );
  NAND2_X1 U10192 ( .A1(n7717), .A2(n7702), .ZN(n9965) );
  OR2_X1 U10193 ( .A1(n9965), .A2(n6646), .ZN(n7708) );
  NAND2_X1 U10194 ( .A1(n7703), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7704) );
  MUX2_X1 U10195 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7704), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n7705) );
  INV_X1 U10196 ( .A(n7705), .ZN(n7706) );
  NOR2_X1 U10197 ( .A1(n7706), .A2(n8003), .ZN(n11695) );
  AOI22_X1 U10198 ( .A1(n9629), .A2(SI_13_), .B1(n10129), .B2(n11695), .ZN(
        n7707) );
  NAND2_X1 U10199 ( .A1(n6447), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U10200 ( .A1(n6449), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7713) );
  NOR2_X1 U10201 ( .A1(n7709), .A2(n11754), .ZN(n7710) );
  OR2_X1 U10202 ( .A1(n7726), .A2(n7710), .ZN(n11753) );
  NAND2_X1 U10203 ( .A1(n8930), .A2(n11753), .ZN(n7712) );
  NAND2_X1 U10204 ( .A1(n8931), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7711) );
  NAND4_X1 U10205 ( .A1(n7714), .A2(n7713), .A3(n7712), .A4(n7711), .ZN(n14577) );
  INV_X1 U10206 ( .A(n14577), .ZN(n8871) );
  AND2_X1 U10207 ( .A1(n11821), .A2(n8871), .ZN(n12594) );
  NAND2_X1 U10208 ( .A1(n7715), .A2(n8395), .ZN(n7716) );
  NAND2_X1 U10209 ( .A1(n15067), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U10210 ( .A1(n10638), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7718) );
  OR2_X1 U10211 ( .A1(n7720), .A2(n7719), .ZN(n7721) );
  NAND2_X1 U10212 ( .A1(n7734), .A2(n7721), .ZN(n10012) );
  OR2_X1 U10213 ( .A1(n10012), .A2(n6646), .ZN(n7724) );
  OR2_X1 U10214 ( .A1(n8003), .A2(n7485), .ZN(n7722) );
  XNOR2_X1 U10215 ( .A(n7722), .B(P3_IR_REG_14__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U10216 ( .A1(n9629), .A2(SI_14_), .B1(n10129), .B2(n11698), .ZN(
        n7723) );
  NAND2_X1 U10217 ( .A1(n6449), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U10218 ( .A1(n6447), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7730) );
  NOR2_X1 U10219 ( .A1(n7726), .A2(n7725), .ZN(n7727) );
  OR2_X1 U10220 ( .A1(n7743), .A2(n7727), .ZN(n11958) );
  NAND2_X1 U10221 ( .A1(n8930), .A2(n11958), .ZN(n7729) );
  NAND2_X1 U10222 ( .A1(n8931), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7728) );
  NAND4_X1 U10223 ( .A1(n7731), .A2(n7730), .A3(n7729), .A4(n7728), .ZN(n12990) );
  XNOR2_X1 U10224 ( .A(n12602), .B(n12990), .ZN(n12507) );
  INV_X1 U10225 ( .A(n12990), .ZN(n12603) );
  NAND2_X1 U10226 ( .A1(n12602), .A2(n12603), .ZN(n7732) );
  NAND2_X1 U10227 ( .A1(n10918), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U10228 ( .A1(n10920), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7735) );
  OR2_X1 U10229 ( .A1(n7737), .A2(n7736), .ZN(n7738) );
  NAND2_X1 U10230 ( .A1(n7750), .A2(n7738), .ZN(n10016) );
  OR2_X1 U10231 ( .A1(n10016), .A2(n6646), .ZN(n7742) );
  OR2_X1 U10232 ( .A1(n7739), .A2(n7485), .ZN(n7740) );
  XNOR2_X1 U10233 ( .A(n7740), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U10234 ( .A1(n9629), .A2(SI_15_), .B1(n10129), .B2(n12737), .ZN(
        n7741) );
  NAND2_X1 U10235 ( .A1(n6449), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U10236 ( .A1(n6447), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7747) );
  OR2_X1 U10237 ( .A1(n7743), .A2(n11908), .ZN(n7744) );
  NAND2_X1 U10238 ( .A1(n7761), .A2(n7744), .ZN(n12993) );
  NAND2_X1 U10239 ( .A1(n8930), .A2(n12993), .ZN(n7746) );
  NAND2_X1 U10240 ( .A1(n12473), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7745) );
  NAND4_X1 U10241 ( .A1(n7748), .A2(n7747), .A3(n7746), .A4(n7745), .ZN(n12980) );
  OR2_X1 U10242 ( .A1(n13122), .A2(n12409), .ZN(n12606) );
  NAND2_X1 U10243 ( .A1(n13122), .A2(n12409), .ZN(n12610) );
  NAND2_X1 U10244 ( .A1(n10652), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U10245 ( .A1(n15113), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7751) );
  OR2_X1 U10246 ( .A1(n7753), .A2(n7752), .ZN(n7754) );
  NAND2_X1 U10247 ( .A1(n7768), .A2(n7754), .ZN(n10078) );
  OR2_X1 U10248 ( .A1(n10078), .A2(n6646), .ZN(n7760) );
  NOR2_X1 U10249 ( .A1(n7755), .A2(n7485), .ZN(n7756) );
  MUX2_X1 U10250 ( .A(n7485), .B(n7756), .S(P3_IR_REG_16__SCAN_IN), .Z(n7758)
         );
  INV_X1 U10251 ( .A(n7770), .ZN(n7757) );
  AOI22_X1 U10252 ( .A1(n9629), .A2(SI_16_), .B1(n10129), .B2(n12740), .ZN(
        n7759) );
  NAND2_X1 U10253 ( .A1(n6447), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U10254 ( .A1(n7761), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7762) );
  INV_X1 U10255 ( .A(n7776), .ZN(n7775) );
  NAND2_X1 U10256 ( .A1(n7762), .A2(n7775), .ZN(n12984) );
  NAND2_X1 U10257 ( .A1(n12984), .A2(n8930), .ZN(n7765) );
  NAND2_X1 U10258 ( .A1(n6449), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U10259 ( .A1(n8931), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7763) );
  NAND4_X1 U10260 ( .A1(n7766), .A2(n7765), .A3(n7764), .A4(n7763), .ZN(n12991) );
  XNOR2_X1 U10261 ( .A(n13115), .B(n12991), .ZN(n12979) );
  NAND2_X1 U10262 ( .A1(n13115), .A2(n7077), .ZN(n12611) );
  NAND2_X1 U10263 ( .A1(n10835), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U10264 ( .A1(n10836), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U10265 ( .A1(n7786), .A2(n7769), .ZN(n7783) );
  XNOR2_X1 U10266 ( .A(n7785), .B(n7783), .ZN(n10231) );
  NAND2_X1 U10267 ( .A1(n10231), .A2(n12486), .ZN(n7774) );
  NAND2_X1 U10268 ( .A1(n7770), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7771) );
  MUX2_X1 U10269 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7771), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n7772) );
  AND2_X1 U10270 ( .A1(n7772), .A2(n7791), .ZN(n12785) );
  AOI22_X1 U10271 ( .A1(n9629), .A2(SI_17_), .B1(n10129), .B2(n12785), .ZN(
        n7773) );
  NAND2_X1 U10272 ( .A1(n6447), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7781) );
  NAND2_X1 U10273 ( .A1(n6449), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U10274 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(n7775), .ZN(n7777) );
  NAND2_X1 U10275 ( .A1(n7777), .A2(n7795), .ZN(n12972) );
  NAND2_X1 U10276 ( .A1(n8930), .A2(n12972), .ZN(n7779) );
  NAND2_X1 U10277 ( .A1(n8931), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7778) );
  OR2_X1 U10278 ( .A1(n13109), .A2(n12955), .ZN(n12620) );
  NAND2_X1 U10279 ( .A1(n13109), .A2(n12955), .ZN(n12615) );
  INV_X1 U10280 ( .A(n7783), .ZN(n7784) );
  NAND2_X1 U10281 ( .A1(n11020), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7801) );
  NAND2_X1 U10282 ( .A1(n11019), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7787) );
  OR2_X1 U10283 ( .A1(n7789), .A2(n7788), .ZN(n7790) );
  NAND2_X1 U10284 ( .A1(n7802), .A2(n7790), .ZN(n10270) );
  NAND2_X1 U10285 ( .A1(n7791), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7792) );
  XNOR2_X1 U10286 ( .A(n7792), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U10287 ( .A1(n9629), .A2(SI_18_), .B1(n12802), .B2(n10129), .ZN(
        n7793) );
  NAND2_X1 U10288 ( .A1(n6447), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10289 ( .A1(n12473), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U10290 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(n7795), .ZN(n7796) );
  INV_X1 U10291 ( .A(n7809), .ZN(n7811) );
  NAND2_X1 U10292 ( .A1(n7796), .A2(n7811), .ZN(n12959) );
  NAND2_X1 U10293 ( .A1(n8930), .A2(n12959), .ZN(n7798) );
  NAND2_X1 U10294 ( .A1(n6449), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U10295 ( .A1(n13032), .A2(n12941), .ZN(n12622) );
  INV_X1 U10296 ( .A(n12952), .ZN(n12626) );
  INV_X1 U10297 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U10298 ( .A1(n11237), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7819) );
  INV_X1 U10299 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11236) );
  NAND2_X1 U10300 ( .A1(n11236), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7803) );
  OR2_X1 U10301 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  NAND2_X1 U10302 ( .A1(n7820), .A2(n7806), .ZN(n10416) );
  NAND2_X1 U10303 ( .A1(n10416), .A2(n12486), .ZN(n7808) );
  INV_X1 U10304 ( .A(SI_19_), .ZN(n10417) );
  AOI22_X1 U10305 ( .A1(n12808), .A2(n10129), .B1(n9629), .B2(n10417), .ZN(
        n7807) );
  NAND2_X1 U10306 ( .A1(n6449), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U10307 ( .A1(n6447), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n7815) );
  INV_X1 U10308 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7810) );
  NAND2_X1 U10309 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n7811), .ZN(n7812) );
  NAND2_X1 U10310 ( .A1(n7828), .A2(n7812), .ZN(n12946) );
  NAND2_X1 U10311 ( .A1(n8930), .A2(n12946), .ZN(n7814) );
  NAND2_X1 U10312 ( .A1(n8931), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n7813) );
  NAND4_X1 U10313 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n12926) );
  NAND2_X1 U10314 ( .A1(n13098), .A2(n12926), .ZN(n12629) );
  INV_X1 U10315 ( .A(n12629), .ZN(n7817) );
  NAND2_X1 U10316 ( .A1(n7823), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10317 ( .A1(n7835), .A2(n7824), .ZN(n10639) );
  OR2_X1 U10318 ( .A1(n12487), .A2(n10640), .ZN(n7825) );
  NAND2_X1 U10319 ( .A1(n6449), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U10320 ( .A1(n6447), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n7832) );
  INV_X1 U10321 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12436) );
  NAND2_X1 U10322 ( .A1(n7828), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U10323 ( .A1(n7843), .A2(n7829), .ZN(n12931) );
  NAND2_X1 U10324 ( .A1(n8930), .A2(n12931), .ZN(n7831) );
  NAND2_X1 U10325 ( .A1(n8931), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n7830) );
  XNOR2_X1 U10326 ( .A(n12932), .B(n12940), .ZN(n12925) );
  OR2_X1 U10327 ( .A1(n12932), .A2(n12940), .ZN(n12632) );
  INV_X1 U10328 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U10329 ( .A1(n11572), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U10330 ( .A1(n15180), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7836) );
  OR2_X1 U10331 ( .A1(n7838), .A2(n7837), .ZN(n7839) );
  NAND2_X1 U10332 ( .A1(n7850), .A2(n7839), .ZN(n10847) );
  INV_X1 U10333 ( .A(SI_21_), .ZN(n10848) );
  OR2_X1 U10334 ( .A1(n12487), .A2(n10848), .ZN(n7841) );
  NAND2_X1 U10335 ( .A1(n6449), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U10336 ( .A1(n6447), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n7847) );
  NAND2_X1 U10337 ( .A1(n7843), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10338 ( .A1(n7855), .A2(n7844), .ZN(n12917) );
  NAND2_X1 U10339 ( .A1(n8930), .A2(n12917), .ZN(n7846) );
  NAND2_X1 U10340 ( .A1(n8931), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10341 ( .A1(n13021), .A2(n12902), .ZN(n12636) );
  INV_X1 U10342 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11748) );
  XNOR2_X1 U10343 ( .A(n11748), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n7862) );
  XNOR2_X1 U10344 ( .A(n7863), .B(n7862), .ZN(n10950) );
  NAND2_X1 U10345 ( .A1(n10950), .A2(n12486), .ZN(n7852) );
  NAND2_X1 U10346 ( .A1(n9629), .A2(SI_22_), .ZN(n7851) );
  NAND2_X1 U10347 ( .A1(n6449), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U10348 ( .A1(n6447), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n7859) );
  INV_X1 U10349 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n7853) );
  NAND2_X1 U10350 ( .A1(n7855), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10351 ( .A1(n7866), .A2(n7856), .ZN(n12907) );
  NAND2_X1 U10352 ( .A1(n8930), .A2(n12907), .ZN(n7858) );
  NAND2_X1 U10353 ( .A1(n8931), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7857) );
  NAND4_X1 U10354 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n7857), .ZN(n12893) );
  NAND2_X1 U10355 ( .A1(n13082), .A2(n12914), .ZN(n12640) );
  NAND2_X1 U10356 ( .A1(n12899), .A2(n12640), .ZN(n7861) );
  NAND2_X1 U10357 ( .A1(n7861), .A2(n12639), .ZN(n12889) );
  XNOR2_X1 U10358 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n7873) );
  XNOR2_X1 U10359 ( .A(n7874), .B(n7873), .ZN(n11104) );
  NAND2_X1 U10360 ( .A1(n11104), .A2(n12486), .ZN(n7865) );
  INV_X1 U10361 ( .A(SI_23_), .ZN(n11106) );
  OR2_X1 U10362 ( .A1(n12487), .A2(n11106), .ZN(n7864) );
  NAND2_X1 U10363 ( .A1(n6449), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10364 ( .A1(n6447), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U10365 ( .A1(n7866), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U10366 ( .A1(n7884), .A2(n7867), .ZN(n12896) );
  NAND2_X1 U10367 ( .A1(n8930), .A2(n12896), .ZN(n7869) );
  NAND2_X1 U10368 ( .A1(n8931), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n7868) );
  XNOR2_X1 U10369 ( .A(n13077), .B(n12903), .ZN(n12512) );
  NAND2_X1 U10370 ( .A1(n12889), .A2(n12891), .ZN(n7872) );
  OR2_X1 U10371 ( .A1(n13077), .A2(n12903), .ZN(n12648) );
  INV_X1 U10372 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10373 ( .A1(n7875), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7876) );
  INV_X1 U10374 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13804) );
  OR2_X2 U10375 ( .A1(n7878), .A2(n13804), .ZN(n7891) );
  NAND2_X1 U10376 ( .A1(n7878), .A2(n13804), .ZN(n7879) );
  INV_X1 U10377 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14532) );
  XNOR2_X1 U10378 ( .A(n7890), .B(n14532), .ZN(n11359) );
  NAND2_X1 U10379 ( .A1(n11359), .A2(n12486), .ZN(n7881) );
  OR2_X1 U10380 ( .A1(n12487), .A2(n15168), .ZN(n7880) );
  NAND2_X1 U10381 ( .A1(n6481), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U10382 ( .A1(n6447), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n7888) );
  INV_X1 U10383 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U10384 ( .A1(n7884), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U10385 ( .A1(n7895), .A2(n7885), .ZN(n12886) );
  NAND2_X1 U10386 ( .A1(n8930), .A2(n12886), .ZN(n7887) );
  NAND2_X1 U10387 ( .A1(n8931), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n7886) );
  INV_X1 U10388 ( .A(n12892), .ZN(n12399) );
  OR2_X1 U10389 ( .A1(n13071), .A2(n12399), .ZN(n12647) );
  NAND2_X1 U10390 ( .A1(n13071), .A2(n12399), .ZN(n12645) );
  NAND2_X1 U10391 ( .A1(n12647), .A2(n12645), .ZN(n12644) );
  INV_X1 U10392 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13801) );
  XNOR2_X1 U10393 ( .A(n13801), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n7892) );
  XNOR2_X1 U10394 ( .A(n7903), .B(n7892), .ZN(n11534) );
  NAND2_X1 U10395 ( .A1(n11534), .A2(n12486), .ZN(n7894) );
  NAND2_X1 U10396 ( .A1(n9629), .A2(SI_25_), .ZN(n7893) );
  NAND2_X1 U10397 ( .A1(n6449), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10398 ( .A1(n6447), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n7899) );
  NAND2_X1 U10399 ( .A1(n7895), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U10400 ( .A1(n7909), .A2(n7896), .ZN(n12875) );
  NAND2_X1 U10401 ( .A1(n8930), .A2(n12875), .ZN(n7898) );
  NAND2_X1 U10402 ( .A1(n8931), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n7897) );
  INV_X1 U10403 ( .A(n12881), .ZN(n12651) );
  NAND2_X1 U10404 ( .A1(n13008), .A2(n12651), .ZN(n7901) );
  NAND2_X1 U10405 ( .A1(n12866), .A2(n7901), .ZN(n12853) );
  NAND2_X1 U10406 ( .A1(n13801), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7902) );
  INV_X1 U10407 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14529) );
  NAND2_X1 U10408 ( .A1(n14529), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7904) );
  INV_X1 U10409 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13797) );
  XNOR2_X1 U10410 ( .A(n13797), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n7906) );
  XNOR2_X1 U10411 ( .A(n7917), .B(n7906), .ZN(n11589) );
  NAND2_X1 U10412 ( .A1(n11589), .A2(n12486), .ZN(n7908) );
  INV_X1 U10413 ( .A(SI_26_), .ZN(n11591) );
  OR2_X1 U10414 ( .A1(n12487), .A2(n11591), .ZN(n7907) );
  NAND2_X1 U10415 ( .A1(n6447), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U10416 ( .A1(n6449), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10417 ( .A1(n7909), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7910) );
  NAND2_X1 U10418 ( .A1(n7924), .A2(n7910), .ZN(n12861) );
  NAND2_X1 U10419 ( .A1(n8930), .A2(n12861), .ZN(n7912) );
  NAND2_X1 U10420 ( .A1(n8931), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n7911) );
  NAND4_X1 U10421 ( .A1(n7914), .A2(n7913), .A3(n7912), .A4(n7911), .ZN(n12871) );
  NAND2_X1 U10422 ( .A1(n13060), .A2(n8900), .ZN(n12658) );
  INV_X1 U10423 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14525) );
  AND2_X1 U10424 ( .A1(n14525), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10425 ( .A1(n13797), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7918) );
  XNOR2_X1 U10426 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n7919) );
  XNOR2_X1 U10427 ( .A(n8902), .B(n7919), .ZN(n11663) );
  NAND2_X1 U10428 ( .A1(n11663), .A2(n12486), .ZN(n7921) );
  INV_X1 U10429 ( .A(SI_27_), .ZN(n11664) );
  OR2_X1 U10430 ( .A1(n12487), .A2(n11664), .ZN(n7920) );
  NAND2_X1 U10431 ( .A1(n6449), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U10432 ( .A1(n6447), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n7928) );
  INV_X1 U10433 ( .A(n7924), .ZN(n7923) );
  INV_X1 U10434 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n7922) );
  NAND2_X1 U10435 ( .A1(n7923), .A2(n7922), .ZN(n7983) );
  NAND2_X1 U10436 ( .A1(n7924), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U10437 ( .A1(n7983), .A2(n7925), .ZN(n12845) );
  NAND2_X1 U10438 ( .A1(n8930), .A2(n12845), .ZN(n7927) );
  NAND2_X1 U10439 ( .A1(n8931), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7926) );
  XNOR2_X2 U10440 ( .A(n12662), .B(n12857), .ZN(n12659) );
  XNOR2_X1 U10441 ( .A(n9645), .B(n12659), .ZN(n7992) );
  NAND2_X1 U10442 ( .A1(n12808), .A2(n10641), .ZN(n8036) );
  INV_X1 U10443 ( .A(n8036), .ZN(n12674) );
  NAND2_X1 U10444 ( .A1(n12808), .A2(n10849), .ZN(n7935) );
  OR2_X1 U10445 ( .A1(n12531), .A2(n8035), .ZN(n7933) );
  XNOR2_X1 U10446 ( .A(n12690), .B(n7933), .ZN(n7934) );
  NAND2_X1 U10447 ( .A1(n7935), .A2(n7934), .ZN(n8916) );
  NAND3_X1 U10448 ( .A1(n12674), .A2(n8916), .A3(n15026), .ZN(n7937) );
  AND2_X1 U10449 ( .A1(n12690), .A2(n8035), .ZN(n7936) );
  NAND2_X1 U10450 ( .A1(n12808), .A2(n7936), .ZN(n8033) );
  NAND2_X1 U10451 ( .A1(n7937), .A2(n8033), .ZN(n15029) );
  INV_X1 U10452 ( .A(n15029), .ZN(n14995) );
  NAND2_X1 U10453 ( .A1(n10395), .A2(n14990), .ZN(n7941) );
  NAND2_X1 U10454 ( .A1(n6618), .A2(n7939), .ZN(n7940) );
  NAND2_X1 U10455 ( .A1(n10616), .A2(n10584), .ZN(n7945) );
  NAND2_X1 U10456 ( .A1(n12704), .A2(n10672), .ZN(n7946) );
  NAND2_X1 U10457 ( .A1(n11002), .A2(n11014), .ZN(n7947) );
  INV_X1 U10458 ( .A(n11000), .ZN(n7949) );
  NAND2_X1 U10459 ( .A1(n12702), .A2(n11066), .ZN(n7950) );
  NAND2_X1 U10460 ( .A1(n11024), .A2(n12561), .ZN(n11023) );
  NAND2_X1 U10461 ( .A1(n12701), .A2(n15014), .ZN(n7951) );
  NAND2_X1 U10462 ( .A1(n11391), .A2(n11471), .ZN(n7952) );
  XNOR2_X1 U10463 ( .A(n12699), .B(n12574), .ZN(n12572) );
  NAND2_X1 U10464 ( .A1(n12582), .A2(n12580), .ZN(n12577) );
  NAND2_X1 U10465 ( .A1(n11498), .A2(n14590), .ZN(n7953) );
  NAND2_X1 U10466 ( .A1(n14589), .A2(n14576), .ZN(n7954) );
  NAND2_X1 U10467 ( .A1(n7955), .A2(n7954), .ZN(n14575) );
  NAND2_X1 U10468 ( .A1(n14575), .A2(n7956), .ZN(n7958) );
  INV_X1 U10469 ( .A(n11818), .ZN(n14591) );
  NAND2_X1 U10470 ( .A1(n14585), .A2(n14591), .ZN(n7957) );
  NAND2_X1 U10471 ( .A1(n12602), .A2(n12990), .ZN(n7961) );
  OR2_X1 U10472 ( .A1(n13122), .A2(n12980), .ZN(n7962) );
  NAND2_X1 U10473 ( .A1(n12989), .A2(n7962), .ZN(n7964) );
  NAND2_X1 U10474 ( .A1(n13122), .A2(n12980), .ZN(n7963) );
  AND2_X1 U10475 ( .A1(n13115), .A2(n12991), .ZN(n7965) );
  NAND2_X1 U10476 ( .A1(n13109), .A2(n12981), .ZN(n7966) );
  OR2_X1 U10477 ( .A1(n13032), .A2(n12969), .ZN(n7967) );
  NAND2_X1 U10478 ( .A1(n12628), .A2(n12629), .ZN(n12938) );
  INV_X1 U10479 ( .A(n12926), .ZN(n12957) );
  OR2_X1 U10480 ( .A1(n13098), .A2(n12957), .ZN(n7968) );
  INV_X1 U10481 ( .A(n12940), .ZN(n12698) );
  NAND2_X1 U10482 ( .A1(n12932), .A2(n12698), .ZN(n7969) );
  OR2_X1 U10483 ( .A1(n13021), .A2(n12927), .ZN(n7971) );
  NOR2_X1 U10484 ( .A1(n13082), .A2(n12893), .ZN(n7973) );
  INV_X1 U10485 ( .A(n13082), .ZN(n7972) );
  NAND2_X1 U10486 ( .A1(n13077), .A2(n12697), .ZN(n7974) );
  OR2_X1 U10487 ( .A1(n13071), .A2(n12892), .ZN(n7975) );
  NAND2_X1 U10488 ( .A1(n13008), .A2(n12881), .ZN(n7977) );
  OR2_X1 U10489 ( .A1(n12871), .A2(n13060), .ZN(n7978) );
  NAND2_X1 U10490 ( .A1(n12680), .A2(n12690), .ZN(n8009) );
  NAND2_X1 U10491 ( .A1(n12531), .A2(n8035), .ZN(n12682) );
  INV_X1 U10492 ( .A(n6710), .ZN(n10128) );
  NAND2_X1 U10493 ( .A1(n10128), .A2(n12688), .ZN(n10135) );
  NAND2_X1 U10494 ( .A1(n10135), .A2(n7980), .ZN(n8937) );
  INV_X1 U10495 ( .A(n8937), .ZN(n8936) );
  NAND2_X1 U10496 ( .A1(n6449), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U10497 ( .A1(n6447), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7987) );
  INV_X1 U10498 ( .A(n7983), .ZN(n7982) );
  INV_X1 U10499 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n7981) );
  NAND2_X1 U10500 ( .A1(n7982), .A2(n7981), .ZN(n8929) );
  NAND2_X1 U10501 ( .A1(n7983), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U10502 ( .A1(n8929), .A2(n7984), .ZN(n12841) );
  NAND2_X1 U10503 ( .A1(n8930), .A2(n12841), .ZN(n7986) );
  NAND2_X1 U10504 ( .A1(n8931), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7985) );
  OAI22_X1 U10505 ( .A1(n8900), .A2(n12956), .B1(n12349), .B2(n12958), .ZN(
        n7989) );
  NOR2_X1 U10506 ( .A1(n8036), .A2(n12656), .ZN(n10156) );
  NAND2_X1 U10507 ( .A1(n7996), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U10508 ( .A1(n8006), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8000) );
  MUX2_X1 U10509 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8000), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8001) );
  NAND2_X1 U10510 ( .A1(n8001), .A2(n7996), .ZN(n11536) );
  NOR2_X1 U10511 ( .A1(n11592), .A2(n11536), .ZN(n8008) );
  NAND2_X1 U10512 ( .A1(n8003), .A2(n8002), .ZN(n8004) );
  NAND2_X1 U10513 ( .A1(n8004), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8005) );
  MUX2_X1 U10514 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8005), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8007) );
  NAND2_X1 U10515 ( .A1(n8007), .A2(n8006), .ZN(n11361) );
  INV_X1 U10516 ( .A(n11361), .ZN(n8013) );
  INV_X1 U10517 ( .A(n10131), .ZN(n8910) );
  NAND2_X1 U10518 ( .A1(n10156), .A2(n8910), .ZN(n12689) );
  NOR2_X1 U10519 ( .A1(n10131), .A2(n8920), .ZN(n8010) );
  INV_X1 U10520 ( .A(n8009), .ZN(n8921) );
  NAND2_X1 U10521 ( .A1(n8010), .A2(n8921), .ZN(n8911) );
  NAND2_X1 U10522 ( .A1(n12689), .A2(n8911), .ZN(n8028) );
  XNOR2_X1 U10523 ( .A(n11361), .B(P3_B_REG_SCAN_IN), .ZN(n8011) );
  INV_X1 U10524 ( .A(n11592), .ZN(n8012) );
  INV_X1 U10525 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n15111) );
  NAND2_X1 U10526 ( .A1(n9907), .A2(n15111), .ZN(n8015) );
  NAND2_X1 U10527 ( .A1(n11592), .A2(n11536), .ZN(n8014) );
  NAND2_X1 U10528 ( .A1(n8015), .A2(n8014), .ZN(n10348) );
  OR2_X1 U10529 ( .A1(n10347), .A2(n10348), .ZN(n8043) );
  NOR2_X1 U10530 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .ZN(
        n8019) );
  NOR4_X1 U10531 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8018) );
  NOR4_X1 U10532 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n8017) );
  NOR4_X1 U10533 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n8016) );
  NAND4_X1 U10534 ( .A1(n8019), .A2(n8018), .A3(n8017), .A4(n8016), .ZN(n8025)
         );
  NOR4_X1 U10535 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8023) );
  NOR4_X1 U10536 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8022) );
  NOR4_X1 U10537 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8021) );
  NOR4_X1 U10538 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8020) );
  NAND4_X1 U10539 ( .A1(n8023), .A2(n8022), .A3(n8021), .A4(n8020), .ZN(n8024)
         );
  NOR2_X1 U10540 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  NOR2_X1 U10541 ( .A1(n8043), .A2(n8040), .ZN(n8918) );
  NAND2_X1 U10542 ( .A1(n8028), .A2(n8918), .ZN(n8031) );
  NAND2_X1 U10543 ( .A1(n10347), .A2(n10348), .ZN(n8041) );
  OR2_X1 U10544 ( .A1(n8041), .A2(n8040), .ZN(n8935) );
  NAND2_X1 U10545 ( .A1(n8910), .A2(n8916), .ZN(n8029) );
  OR2_X1 U10546 ( .A1(n8935), .A2(n8029), .ZN(n8030) );
  INV_X1 U10547 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10548 ( .A1(n8033), .A2(n12656), .ZN(n10350) );
  OR2_X1 U10549 ( .A1(n10350), .A2(n10348), .ZN(n8034) );
  NAND2_X1 U10550 ( .A1(n8036), .A2(n6458), .ZN(n10351) );
  AND2_X1 U10551 ( .A1(n8034), .A2(n10351), .ZN(n8045) );
  OAI22_X1 U10552 ( .A1(n12680), .A2(n12528), .B1(n8035), .B2(n15026), .ZN(
        n8037) );
  NAND2_X1 U10553 ( .A1(n8037), .A2(n8036), .ZN(n8038) );
  NAND2_X1 U10554 ( .A1(n8038), .A2(n12656), .ZN(n8039) );
  NAND2_X1 U10555 ( .A1(n8039), .A2(n10348), .ZN(n8044) );
  NOR2_X1 U10556 ( .A1(n10131), .A2(n8040), .ZN(n8042) );
  NOR2_X1 U10557 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n8052) );
  NOR2_X1 U10558 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8051) );
  NAND3_X1 U10559 ( .A1(n8167), .A2(n8193), .A3(n8055), .ZN(n8056) );
  NOR2_X1 U10560 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n8058) );
  NAND4_X1 U10561 ( .A1(n8058), .A2(n8057), .A3(n7011), .A4(n8144), .ZN(n8141)
         );
  NAND3_X1 U10562 ( .A1(n8060), .A2(n8059), .A3(n8816), .ZN(n8061) );
  XNOR2_X2 U10563 ( .A(n8069), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8070) );
  AND2_X2 U10564 ( .A1(n8072), .A2(n8070), .ZN(n8093) );
  NAND2_X1 U10565 ( .A1(n8093), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8077) );
  INV_X1 U10566 ( .A(n8070), .ZN(n12056) );
  INV_X1 U10567 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9667) );
  OR2_X1 U10568 ( .A1(n8180), .A2(n9667), .ZN(n8076) );
  NAND2_X4 U10569 ( .A1(n8070), .A2(n8071), .ZN(n8689) );
  INV_X1 U10570 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11194) );
  NAND2_X2 U10571 ( .A1(n11962), .A2(n12056), .ZN(n8179) );
  INV_X1 U10572 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8073) );
  OR2_X1 U10573 ( .A1(n8179), .A2(n8073), .ZN(n8074) );
  INV_X1 U10574 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14711) );
  NOR2_X1 U10575 ( .A1(n9842), .A2(n9817), .ZN(n8078) );
  XNOR2_X1 U10576 ( .A(n8078), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14538) );
  XNOR2_X2 U10577 ( .A(n8080), .B(n8079), .ZN(n14055) );
  MUX2_X1 U10578 ( .A(n14711), .B(n14538), .S(n8113), .Z(n11448) );
  NAND2_X1 U10579 ( .A1(n6651), .A2(n11448), .ZN(n8092) );
  INV_X1 U10580 ( .A(n8086), .ZN(n8081) );
  NAND2_X1 U10581 ( .A1(n8143), .A2(n8144), .ZN(n8082) );
  NOR2_X1 U10582 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n8085) );
  NAND2_X1 U10583 ( .A1(n8088), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8087) );
  INV_X1 U10584 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10585 ( .A1(n8090), .A2(n8089), .ZN(n8139) );
  NAND2_X1 U10586 ( .A1(n8092), .A2(n9656), .ZN(n8118) );
  NAND2_X1 U10587 ( .A1(n8512), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8098) );
  INV_X1 U10588 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11455) );
  INV_X4 U10589 ( .A(n8093), .ZN(n8730) );
  INV_X1 U10590 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10040) );
  INV_X1 U10591 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8094) );
  OR2_X1 U10592 ( .A1(n8179), .A2(n8094), .ZN(n8095) );
  NAND2_X2 U10593 ( .A1(n8113), .A2(n9842), .ZN(n8157) );
  OR2_X1 U10594 ( .A1(n8157), .A2(n8100), .ZN(n8116) );
  NAND2_X2 U10595 ( .A1(n8113), .A2(n9014), .ZN(n8656) );
  NAND2_X1 U10596 ( .A1(n8101), .A2(SI_1_), .ZN(n8128) );
  NOR2_X1 U10597 ( .A1(n8104), .A2(n9817), .ZN(n8106) );
  INV_X1 U10598 ( .A(n8106), .ZN(n8107) );
  NAND2_X1 U10599 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  NAND2_X1 U10600 ( .A1(n8129), .A2(n8109), .ZN(n9903) );
  OR2_X1 U10601 ( .A1(n8656), .A2(n9903), .ZN(n8115) );
  NAND2_X1 U10602 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8110) );
  MUX2_X1 U10603 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8110), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8112) );
  INV_X1 U10604 ( .A(n8124), .ZN(n8111) );
  NAND2_X1 U10605 ( .A1(n8112), .A2(n8111), .ZN(n10042) );
  OR2_X1 U10606 ( .A1(n8113), .A2(n10042), .ZN(n8114) );
  INV_X1 U10607 ( .A(n8173), .ZN(n8117) );
  NAND3_X1 U10608 ( .A1(n8118), .A2(n8772), .A3(n8117), .ZN(n8146) );
  NAND2_X1 U10609 ( .A1(n8512), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8123) );
  INV_X1 U10610 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10039) );
  OR2_X1 U10611 ( .A1(n8730), .A2(n10039), .ZN(n8122) );
  INV_X1 U10612 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10796) );
  INV_X1 U10613 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8119) );
  OR2_X1 U10614 ( .A1(n8179), .A2(n8119), .ZN(n8120) );
  NOR2_X1 U10615 ( .A1(n8124), .A2(n8345), .ZN(n8125) );
  MUX2_X1 U10616 ( .A(n8345), .B(n8125), .S(P1_IR_REG_2__SCAN_IN), .Z(n8126)
         );
  INV_X1 U10617 ( .A(n8126), .ZN(n8127) );
  NAND2_X1 U10618 ( .A1(n8127), .A2(n8165), .ZN(n14057) );
  MUX2_X1 U10619 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8130), .Z(n8131) );
  NAND2_X1 U10620 ( .A1(n8131), .A2(SI_2_), .ZN(n8158) );
  OAI21_X1 U10621 ( .B1(n8131), .B2(SI_2_), .A(n8158), .ZN(n8133) );
  NAND2_X1 U10622 ( .A1(n8132), .A2(n8133), .ZN(n8136) );
  INV_X1 U10623 ( .A(n8133), .ZN(n8134) );
  NAND2_X1 U10624 ( .A1(n8136), .A2(n8159), .ZN(n9844) );
  NAND2_X1 U10625 ( .A1(n14740), .A2(n10727), .ZN(n8137) );
  NAND2_X2 U10626 ( .A1(n10921), .A2(n8137), .ZN(n10724) );
  NAND2_X1 U10627 ( .A1(n9679), .A2(n11449), .ZN(n8771) );
  NAND2_X1 U10628 ( .A1(n8139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U10629 ( .A1(n14536), .A2(n11239), .ZN(n9657) );
  NAND4_X1 U10630 ( .A1(n8146), .A2(n10724), .A3(n8771), .A4(n8352), .ZN(n8151) );
  INV_X1 U10631 ( .A(n10727), .ZN(n10799) );
  OR2_X1 U10632 ( .A1(n14740), .A2(n10799), .ZN(n10929) );
  NAND2_X1 U10633 ( .A1(n10929), .A2(n8352), .ZN(n8149) );
  NAND2_X1 U10634 ( .A1(n14740), .A2(n10799), .ZN(n8147) );
  NAND2_X1 U10635 ( .A1(n8147), .A2(n8487), .ZN(n8148) );
  NAND2_X1 U10636 ( .A1(n8151), .A2(n8150), .ZN(n8172) );
  NAND2_X1 U10637 ( .A1(n8512), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8156) );
  OR2_X1 U10638 ( .A1(n8689), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8155) );
  INV_X1 U10639 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10038) );
  OR2_X1 U10640 ( .A1(n8730), .A2(n10038), .ZN(n8154) );
  INV_X1 U10641 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8152) );
  OR2_X1 U10642 ( .A1(n8179), .A2(n8152), .ZN(n8153) );
  NAND2_X1 U10643 ( .A1(n8160), .A2(n8161), .ZN(n8164) );
  INV_X1 U10644 ( .A(n8161), .ZN(n8162) );
  NAND2_X1 U10645 ( .A1(n8164), .A2(n8187), .ZN(n9896) );
  OR2_X1 U10646 ( .A1(n9896), .A2(n8656), .ZN(n8171) );
  INV_X2 U10647 ( .A(n8113), .ZN(n8522) );
  NOR2_X1 U10648 ( .A1(n8168), .A2(n8345), .ZN(n8166) );
  MUX2_X1 U10649 ( .A(n8345), .B(n8166), .S(P1_IR_REG_3__SCAN_IN), .Z(n8169)
         );
  NAND2_X1 U10650 ( .A1(n8522), .A2(n14074), .ZN(n8170) );
  OAI211_X1 U10651 ( .C1(n8157), .C2(n9811), .A(n8171), .B(n8170), .ZN(n14694)
         );
  XNOR2_X1 U10652 ( .A(n14038), .B(n14694), .ZN(n10931) );
  NAND2_X1 U10653 ( .A1(n8172), .A2(n10931), .ZN(n8178) );
  NAND2_X1 U10654 ( .A1(n8173), .A2(n8771), .ZN(n8174) );
  NAND4_X1 U10655 ( .A1(n10723), .A2(n8487), .A3(n10931), .A4(n10724), .ZN(
        n8177) );
  INV_X1 U10656 ( .A(n14694), .ZN(n10927) );
  NAND3_X1 U10657 ( .A1(n8487), .A2(n10927), .A3(n14038), .ZN(n8176) );
  NOR2_X1 U10658 ( .A1(n14038), .A2(n10927), .ZN(n11090) );
  NAND2_X1 U10659 ( .A1(n11090), .A2(n8791), .ZN(n8175) );
  NAND4_X1 U10660 ( .A1(n8178), .A2(n8177), .A3(n8176), .A4(n8175), .ZN(n8201)
         );
  INV_X1 U10661 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n8181) );
  OR2_X1 U10662 ( .A1(n8382), .A2(n8181), .ZN(n8184) );
  XNOR2_X1 U10663 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11100) );
  OR2_X1 U10664 ( .A1(n8689), .A2(n11100), .ZN(n8183) );
  INV_X1 U10665 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11097) );
  OR2_X1 U10666 ( .A1(n8730), .A2(n11097), .ZN(n8182) );
  INV_X1 U10667 ( .A(n8188), .ZN(n8189) );
  OR2_X1 U10668 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  AND2_X1 U10669 ( .A1(n8205), .A2(n8191), .ZN(n9839) );
  NAND2_X1 U10670 ( .A1(n9839), .A2(n8758), .ZN(n8198) );
  INV_X2 U10671 ( .A(n8157), .ZN(n8523) );
  NOR2_X1 U10672 ( .A1(n8194), .A2(n8345), .ZN(n8192) );
  MUX2_X1 U10673 ( .A(n8345), .B(n8192), .S(P1_IR_REG_4__SCAN_IN), .Z(n8196)
         );
  NAND2_X1 U10674 ( .A1(n8194), .A2(n8193), .ZN(n8430) );
  INV_X1 U10675 ( .A(n8430), .ZN(n8195) );
  AOI22_X1 U10676 ( .A1(n8523), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8522), .B2(
        n14093), .ZN(n8197) );
  MUX2_X1 U10677 ( .A(n11273), .B(n11132), .S(n8487), .Z(n8200) );
  INV_X1 U10678 ( .A(n11132), .ZN(n11143) );
  INV_X1 U10679 ( .A(n11273), .ZN(n9693) );
  MUX2_X1 U10680 ( .A(n11143), .B(n9693), .S(n8487), .Z(n8199) );
  OAI21_X1 U10681 ( .B1(n8201), .B2(n8200), .A(n8199), .ZN(n8203) );
  NAND2_X1 U10682 ( .A1(n8201), .A2(n8200), .ZN(n8202) );
  NAND2_X1 U10683 ( .A1(n8206), .A2(SI_5_), .ZN(n8223) );
  OAI21_X1 U10684 ( .B1(n8206), .B2(SI_5_), .A(n8223), .ZN(n8220) );
  XNOR2_X1 U10685 ( .A(n8222), .B(n8220), .ZN(n9849) );
  NAND2_X1 U10686 ( .A1(n9849), .A2(n8758), .ZN(n8209) );
  NAND2_X1 U10687 ( .A1(n8430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8207) );
  XNOR2_X1 U10688 ( .A(n8207), .B(P1_IR_REG_5__SCAN_IN), .ZN(n14109) );
  AOI22_X1 U10689 ( .A1(n8523), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8522), .B2(
        n14109), .ZN(n8208) );
  NAND2_X1 U10690 ( .A1(n8209), .A2(n8208), .ZN(n11268) );
  AOI21_X1 U10691 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8210) );
  AND3_X1 U10692 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8235) );
  NOR2_X1 U10693 ( .A1(n8210), .A2(n8235), .ZN(n11267) );
  NAND2_X1 U10694 ( .A1(n8708), .A2(n11267), .ZN(n8216) );
  INV_X1 U10695 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8211) );
  OR2_X1 U10696 ( .A1(n8382), .A2(n8211), .ZN(n8215) );
  INV_X1 U10697 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n8212) );
  OR2_X1 U10698 ( .A1(n8179), .A2(n8212), .ZN(n8214) );
  INV_X1 U10699 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10047) );
  OR2_X1 U10700 ( .A1(n8730), .A2(n10047), .ZN(n8213) );
  NAND4_X1 U10701 ( .A1(n8216), .A2(n8215), .A3(n8214), .A4(n8213), .ZN(n14037) );
  MUX2_X1 U10702 ( .A(n11268), .B(n14037), .S(n8487), .Z(n8218) );
  MUX2_X1 U10703 ( .A(n14037), .B(n11268), .S(n8487), .Z(n8217) );
  INV_X1 U10704 ( .A(n8218), .ZN(n8219) );
  INV_X1 U10705 ( .A(n8220), .ZN(n8221) );
  MUX2_X1 U10706 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8622), .Z(n8224) );
  NAND2_X1 U10707 ( .A1(n8224), .A2(SI_6_), .ZN(n8256) );
  OAI21_X1 U10708 ( .B1(n8224), .B2(SI_6_), .A(n8256), .ZN(n8225) );
  INV_X1 U10709 ( .A(n8225), .ZN(n8226) );
  NAND2_X1 U10710 ( .A1(n8227), .A2(n8226), .ZN(n8257) );
  OR2_X1 U10711 ( .A1(n8227), .A2(n8226), .ZN(n8228) );
  NAND2_X1 U10712 ( .A1(n8257), .A2(n8228), .ZN(n9898) );
  OR2_X1 U10713 ( .A1(n9898), .A2(n8656), .ZN(n8234) );
  NOR2_X1 U10714 ( .A1(n8430), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n8231) );
  OR2_X1 U10715 ( .A1(n8231), .A2(n8345), .ZN(n8229) );
  MUX2_X1 U10716 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8229), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n8232) );
  INV_X1 U10717 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8230) );
  NAND2_X1 U10718 ( .A1(n8231), .A2(n8230), .ZN(n8277) );
  AND2_X1 U10719 ( .A1(n8232), .A2(n8277), .ZN(n14125) );
  AOI22_X1 U10720 ( .A1(n8523), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8522), .B2(
        n14125), .ZN(n8233) );
  NAND2_X1 U10721 ( .A1(n8234), .A2(n8233), .ZN(n14765) );
  INV_X1 U10722 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14118) );
  OR2_X1 U10723 ( .A1(n8382), .A2(n14118), .ZN(n8238) );
  NAND2_X1 U10724 ( .A1(n8235), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8250) );
  OAI21_X1 U10725 ( .B1(n8235), .B2(P1_REG3_REG_6__SCAN_IN), .A(n8250), .ZN(
        n11174) );
  OR2_X1 U10726 ( .A1(n8689), .A2(n11174), .ZN(n8237) );
  INV_X1 U10727 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11172) );
  OR2_X1 U10728 ( .A1(n8730), .A2(n11172), .ZN(n8236) );
  NAND4_X1 U10729 ( .A1(n8239), .A2(n8238), .A3(n8237), .A4(n8236), .ZN(n14036) );
  MUX2_X1 U10730 ( .A(n14765), .B(n14036), .S(n8352), .Z(n8243) );
  MUX2_X1 U10731 ( .A(n14765), .B(n14036), .S(n8795), .Z(n8240) );
  NAND2_X1 U10732 ( .A1(n8241), .A2(n8240), .ZN(n8247) );
  INV_X1 U10733 ( .A(n8242), .ZN(n8245) );
  INV_X1 U10734 ( .A(n8243), .ZN(n8244) );
  NAND2_X1 U10735 ( .A1(n8247), .A2(n8246), .ZN(n8269) );
  INV_X1 U10736 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8248) );
  OR2_X1 U10737 ( .A1(n8382), .A2(n8248), .ZN(n8254) );
  AND2_X1 U10738 ( .A1(n8250), .A2(n8249), .ZN(n8251) );
  NOR2_X1 U10739 ( .A1(n8250), .A2(n8249), .ZN(n8282) );
  OR2_X1 U10740 ( .A1(n8251), .A2(n8282), .ZN(n11257) );
  OR2_X1 U10741 ( .A1(n8689), .A2(n11257), .ZN(n8253) );
  INV_X1 U10742 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11252) );
  OR2_X1 U10743 ( .A1(n8730), .A2(n11252), .ZN(n8252) );
  NAND4_X1 U10744 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n8252), .ZN(n14035) );
  NAND2_X1 U10745 ( .A1(n8257), .A2(n8256), .ZN(n8261) );
  MUX2_X1 U10746 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8622), .Z(n8258) );
  NAND2_X1 U10747 ( .A1(n8258), .A2(SI_7_), .ZN(n8270) );
  OAI21_X1 U10748 ( .B1(n8258), .B2(SI_7_), .A(n8270), .ZN(n8259) );
  INV_X1 U10749 ( .A(n8259), .ZN(n8260) );
  NAND2_X1 U10750 ( .A1(n8271), .A2(n8262), .ZN(n9900) );
  OR2_X1 U10751 ( .A1(n9900), .A2(n8656), .ZN(n8265) );
  NAND2_X1 U10752 ( .A1(n8277), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8263) );
  XNOR2_X1 U10753 ( .A(n8263), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U10754 ( .A1(n8523), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8522), .B2(
        n10306), .ZN(n8264) );
  NAND2_X1 U10755 ( .A1(n8265), .A2(n8264), .ZN(n11256) );
  MUX2_X1 U10756 ( .A(n14035), .B(n11256), .S(n8795), .Z(n8266) );
  INV_X1 U10757 ( .A(n8266), .ZN(n8268) );
  MUX2_X1 U10758 ( .A(n11256), .B(n14035), .S(n8795), .Z(n8267) );
  NAND2_X1 U10759 ( .A1(n8269), .A2(n8268), .ZN(n8290) );
  NAND2_X1 U10760 ( .A1(n8271), .A2(n8270), .ZN(n8275) );
  MUX2_X1 U10761 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n8622), .Z(n8272) );
  NAND2_X1 U10762 ( .A1(n8272), .A2(SI_8_), .ZN(n8302) );
  OAI21_X1 U10763 ( .B1(n8272), .B2(SI_8_), .A(n8302), .ZN(n8273) );
  INV_X1 U10764 ( .A(n8273), .ZN(n8274) );
  OR2_X1 U10765 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  NAND2_X1 U10766 ( .A1(n8303), .A2(n8276), .ZN(n9988) );
  OR2_X1 U10767 ( .A1(n9988), .A2(n8656), .ZN(n8280) );
  NAND2_X1 U10768 ( .A1(n8278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8310) );
  XNOR2_X1 U10769 ( .A(n8310), .B(P1_IR_REG_8__SCAN_IN), .ZN(n14140) );
  AOI22_X1 U10770 ( .A1(n8523), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8522), .B2(
        n14140), .ZN(n8279) );
  INV_X1 U10771 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n8281) );
  OR2_X1 U10772 ( .A1(n8382), .A2(n8281), .ZN(n8286) );
  NAND2_X1 U10773 ( .A1(n8282), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8296) );
  OR2_X1 U10774 ( .A1(n8282), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10775 ( .A1(n8296), .A2(n8283), .ZN(n11429) );
  OR2_X1 U10776 ( .A1(n8689), .A2(n11429), .ZN(n8285) );
  INV_X1 U10777 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10294) );
  OR2_X1 U10778 ( .A1(n8730), .A2(n10294), .ZN(n8284) );
  OR2_X1 U10779 ( .A1(n11431), .A2(n11627), .ZN(n11341) );
  NAND2_X1 U10780 ( .A1(n11431), .A2(n11627), .ZN(n8288) );
  MUX2_X1 U10781 ( .A(n11341), .B(n8288), .S(n8352), .Z(n8289) );
  NAND3_X1 U10782 ( .A1(n8291), .A2(n8290), .A3(n8289), .ZN(n8294) );
  INV_X1 U10783 ( .A(n11431), .ZN(n8292) );
  MUX2_X1 U10784 ( .A(n11627), .B(n8292), .S(n8352), .Z(n8293) );
  INV_X1 U10785 ( .A(n11627), .ZN(n8767) );
  INV_X1 U10786 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10308) );
  OR2_X1 U10787 ( .A1(n8382), .A2(n10308), .ZN(n8300) );
  NAND2_X1 U10788 ( .A1(n8296), .A2(n8295), .ZN(n8297) );
  NAND2_X1 U10789 ( .A1(n8317), .A2(n8297), .ZN(n11626) );
  OR2_X1 U10790 ( .A1(n8689), .A2(n11626), .ZN(n8299) );
  INV_X1 U10791 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11483) );
  OR2_X1 U10792 ( .A1(n8730), .A2(n11483), .ZN(n8298) );
  MUX2_X1 U10793 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n8622), .Z(n8304) );
  NAND2_X1 U10794 ( .A1(n8304), .A2(SI_9_), .ZN(n8323) );
  OAI21_X1 U10795 ( .B1(n8304), .B2(SI_9_), .A(n8323), .ZN(n8305) );
  INV_X1 U10796 ( .A(n8305), .ZN(n8306) );
  OR2_X1 U10797 ( .A1(n8307), .A2(n8306), .ZN(n8308) );
  INV_X1 U10798 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U10799 ( .A1(n8310), .A2(n8309), .ZN(n8311) );
  NAND2_X1 U10800 ( .A1(n8311), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8348) );
  XNOR2_X1 U10801 ( .A(n8348), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14159) );
  AOI22_X1 U10802 ( .A1(n8523), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8522), .B2(
        n14159), .ZN(n8312) );
  MUX2_X1 U10803 ( .A(n11656), .B(n11621), .S(n8352), .Z(n8315) );
  INV_X1 U10804 ( .A(n11656), .ZN(n11343) );
  MUX2_X1 U10805 ( .A(n11343), .B(n11488), .S(n8795), .Z(n8314) );
  INV_X1 U10806 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10310) );
  OR2_X1 U10807 ( .A1(n8382), .A2(n10310), .ZN(n8321) );
  NAND2_X1 U10808 ( .A1(n8317), .A2(n8316), .ZN(n8318) );
  NAND2_X1 U10809 ( .A1(n8359), .A2(n8318), .ZN(n11658) );
  OR2_X1 U10810 ( .A1(n8689), .A2(n11658), .ZN(n8320) );
  INV_X1 U10811 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10299) );
  OR2_X1 U10812 ( .A1(n8730), .A2(n10299), .ZN(n8319) );
  NAND4_X1 U10813 ( .A1(n8322), .A2(n8321), .A3(n8320), .A4(n8319), .ZN(n14034) );
  MUX2_X1 U10814 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8622), .Z(n8325) );
  NAND2_X1 U10815 ( .A1(n8325), .A2(SI_10_), .ZN(n8344) );
  OAI21_X1 U10816 ( .B1(n8325), .B2(SI_10_), .A(n8344), .ZN(n8341) );
  NAND2_X1 U10817 ( .A1(n10079), .A2(n8758), .ZN(n8330) );
  INV_X1 U10818 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U10819 ( .A1(n8348), .A2(n8326), .ZN(n8327) );
  NAND2_X1 U10820 ( .A1(n8327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8328) );
  XNOR2_X1 U10821 ( .A(n8328), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U10822 ( .A1(n8523), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10324), 
        .B2(n8522), .ZN(n8329) );
  MUX2_X1 U10823 ( .A(n14034), .B(n14792), .S(n8795), .Z(n8333) );
  MUX2_X1 U10824 ( .A(n14034), .B(n14792), .S(n8352), .Z(n8331) );
  NAND2_X1 U10825 ( .A1(n8332), .A2(n8331), .ZN(n8335) );
  INV_X1 U10826 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10317) );
  OR2_X1 U10827 ( .A1(n8382), .A2(n10317), .ZN(n8339) );
  INV_X1 U10828 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8336) );
  XNOR2_X1 U10829 ( .A(n8359), .B(n8336), .ZN(n11763) );
  OR2_X1 U10830 ( .A1(n8689), .A2(n11763), .ZN(n8338) );
  INV_X1 U10831 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11583) );
  OR2_X1 U10832 ( .A1(n8730), .A2(n11583), .ZN(n8337) );
  NAND4_X1 U10833 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(n14033) );
  INV_X1 U10834 ( .A(n8341), .ZN(n8342) );
  MUX2_X1 U10835 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n8622), .Z(n8365) );
  XNOR2_X1 U10836 ( .A(n8365), .B(SI_11_), .ZN(n8368) );
  XNOR2_X1 U10837 ( .A(n8369), .B(n8368), .ZN(n10105) );
  NAND2_X1 U10838 ( .A1(n10105), .A2(n8758), .ZN(n8351) );
  OR2_X1 U10839 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  NAND2_X1 U10840 ( .A1(n8348), .A2(n8347), .ZN(n8370) );
  INV_X1 U10841 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8349) );
  XNOR2_X1 U10842 ( .A(n8370), .B(n8349), .ZN(n10476) );
  AOI22_X1 U10843 ( .A1(n8523), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10476), 
        .B2(n8522), .ZN(n8350) );
  MUX2_X1 U10844 ( .A(n14033), .B(n11768), .S(n8791), .Z(n8354) );
  MUX2_X1 U10845 ( .A(n14033), .B(n11768), .S(n8795), .Z(n8353) );
  INV_X1 U10846 ( .A(n8354), .ZN(n8355) );
  INV_X1 U10847 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8356) );
  OR2_X1 U10848 ( .A1(n8382), .A2(n8356), .ZN(n8363) );
  INV_X1 U10849 ( .A(n8359), .ZN(n8357) );
  AOI21_X1 U10850 ( .B1(n8357), .B2(P1_REG3_REG_11__SCAN_IN), .A(
        P1_REG3_REG_12__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10851 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n8358) );
  OR2_X1 U10852 ( .A1(n8360), .A2(n8383), .ZN(n11742) );
  OR2_X1 U10853 ( .A1(n8689), .A2(n11742), .ZN(n8362) );
  INV_X1 U10854 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10470) );
  OR2_X1 U10855 ( .A1(n8730), .A2(n10470), .ZN(n8361) );
  NAND4_X1 U10856 ( .A1(n8364), .A2(n8363), .A3(n8362), .A4(n8361), .ZN(n14032) );
  INV_X1 U10857 ( .A(n8365), .ZN(n8366) );
  NAND2_X1 U10858 ( .A1(n8366), .A2(n9847), .ZN(n8367) );
  MUX2_X1 U10859 ( .A(n10359), .B(n15054), .S(n8622), .Z(n8393) );
  XNOR2_X1 U10860 ( .A(n8393), .B(SI_12_), .ZN(n8391) );
  NAND2_X1 U10861 ( .A1(n10358), .A2(n8758), .ZN(n8373) );
  NAND2_X1 U10862 ( .A1(n8371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8397) );
  XNOR2_X1 U10863 ( .A(n8397), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U10864 ( .A1(n10657), .A2(n8522), .B1(n8523), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8372) );
  MUX2_X1 U10865 ( .A(n14032), .B(n11889), .S(n8795), .Z(n8377) );
  MUX2_X1 U10866 ( .A(n14032), .B(n11889), .S(n8791), .Z(n8374) );
  NAND2_X1 U10867 ( .A1(n8375), .A2(n8374), .ZN(n8381) );
  INV_X1 U10868 ( .A(n8376), .ZN(n8379) );
  INV_X1 U10869 ( .A(n8377), .ZN(n8378) );
  NAND2_X1 U10870 ( .A1(n8381), .A2(n8380), .ZN(n8403) );
  NAND2_X1 U10871 ( .A1(n8512), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8390) );
  NAND2_X1 U10872 ( .A1(n8383), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8419) );
  OR2_X1 U10873 ( .A1(n8383), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U10874 ( .A1(n8419), .A2(n8384), .ZN(n11949) );
  OR2_X1 U10875 ( .A1(n8689), .A2(n11949), .ZN(n8389) );
  INV_X1 U10876 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8385) );
  OR2_X1 U10877 ( .A1(n8730), .A2(n8385), .ZN(n8388) );
  INV_X1 U10878 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8386) );
  OR2_X1 U10879 ( .A1(n8179), .A2(n8386), .ZN(n8387) );
  NAND4_X1 U10880 ( .A1(n8390), .A2(n8389), .A3(n8388), .A4(n8387), .ZN(n14031) );
  NAND2_X1 U10881 ( .A1(n8393), .A2(n9854), .ZN(n8394) );
  MUX2_X1 U10882 ( .A(n8395), .B(n10448), .S(n8622), .Z(n8406) );
  XNOR2_X1 U10883 ( .A(n8406), .B(SI_13_), .ZN(n8404) );
  NAND2_X1 U10884 ( .A1(n10408), .A2(n8758), .ZN(n8400) );
  INV_X1 U10885 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10886 ( .A1(n8397), .A2(n8396), .ZN(n8398) );
  NAND2_X1 U10887 ( .A1(n8398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8411) );
  XNOR2_X1 U10888 ( .A(n8411), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U10889 ( .A1(n10851), .A2(n8522), .B1(n8523), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8399) );
  MUX2_X1 U10890 ( .A(n14031), .B(n11951), .S(n8791), .Z(n8402) );
  INV_X1 U10891 ( .A(n14031), .ZN(n11873) );
  INV_X1 U10892 ( .A(n11951), .ZN(n11681) );
  MUX2_X1 U10893 ( .A(n11873), .B(n11681), .S(n8795), .Z(n8401) );
  INV_X1 U10894 ( .A(SI_14_), .ZN(n10011) );
  NAND2_X1 U10895 ( .A1(n8452), .A2(n10011), .ZN(n8407) );
  MUX2_X1 U10896 ( .A(n15067), .B(n10638), .S(n8622), .Z(n8446) );
  NAND2_X1 U10897 ( .A1(n8408), .A2(n8446), .ZN(n8409) );
  NAND2_X1 U10898 ( .A1(n8427), .A2(n8409), .ZN(n10637) );
  OR2_X1 U10899 ( .A1(n10637), .A2(n8656), .ZN(n8417) );
  INV_X1 U10900 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10901 ( .A1(n8411), .A2(n8410), .ZN(n8412) );
  NAND2_X1 U10902 ( .A1(n8412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8414) );
  INV_X1 U10903 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8413) );
  OAI22_X1 U10904 ( .A1(n11207), .A2(n8113), .B1(n8157), .B2(n15067), .ZN(
        n8415) );
  INV_X1 U10905 ( .A(n8415), .ZN(n8416) );
  NAND2_X2 U10906 ( .A1(n8417), .A2(n8416), .ZN(n14643) );
  NAND2_X1 U10907 ( .A1(n8512), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8425) );
  INV_X1 U10908 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U10909 ( .A1(n8419), .A2(n8418), .ZN(n8420) );
  NAND2_X1 U10910 ( .A1(n8435), .A2(n8420), .ZN(n14648) );
  OR2_X1 U10911 ( .A1(n8689), .A2(n14648), .ZN(n8424) );
  INV_X1 U10912 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11803) );
  OR2_X1 U10913 ( .A1(n8730), .A2(n11803), .ZN(n8423) );
  INV_X1 U10914 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8421) );
  OR2_X1 U10915 ( .A1(n8179), .A2(n8421), .ZN(n8422) );
  NAND4_X1 U10916 ( .A1(n8425), .A2(n8424), .A3(n8423), .A4(n8422), .ZN(n14030) );
  XNOR2_X1 U10917 ( .A(n14643), .B(n14030), .ZN(n11800) );
  INV_X1 U10918 ( .A(n14643), .ZN(n8442) );
  NAND2_X1 U10919 ( .A1(n8427), .A2(n8426), .ZN(n8428) );
  MUX2_X1 U10920 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n9842), .Z(n8453) );
  XNOR2_X1 U10921 ( .A(n8453), .B(SI_15_), .ZN(n8447) );
  XNOR2_X1 U10922 ( .A(n8428), .B(n8447), .ZN(n10917) );
  NAND2_X1 U10923 ( .A1(n10917), .A2(n8758), .ZN(n8433) );
  OAI21_X1 U10924 ( .B1(n8430), .B2(n8429), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8431) );
  XNOR2_X1 U10925 ( .A(n8431), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U10926 ( .A1(n8523), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8522), 
        .B2(n11849), .ZN(n8432) );
  NAND2_X2 U10927 ( .A1(n8433), .A2(n8432), .ZN(n14663) );
  INV_X1 U10928 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8434) );
  OR2_X1 U10929 ( .A1(n8382), .A2(n8434), .ZN(n8440) );
  INV_X1 U10930 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n14013) );
  AND2_X1 U10931 ( .A1(n8435), .A2(n14013), .ZN(n8436) );
  OR2_X1 U10932 ( .A1(n8436), .A2(n8467), .ZN(n14014) );
  OR2_X1 U10933 ( .A1(n14014), .A2(n8689), .ZN(n8439) );
  INV_X1 U10934 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8437) );
  OR2_X1 U10935 ( .A1(n8730), .A2(n8437), .ZN(n8438) );
  NAND2_X1 U10936 ( .A1(n14663), .A2(n11920), .ZN(n8766) );
  OAI21_X1 U10937 ( .B1(n8442), .B2(n14030), .A(n8766), .ZN(n8443) );
  NAND2_X1 U10938 ( .A1(n8443), .A2(n8795), .ZN(n8444) );
  INV_X1 U10939 ( .A(n14030), .ZN(n11791) );
  OR2_X1 U10940 ( .A1(n14643), .A2(n11791), .ZN(n11784) );
  AOI21_X1 U10941 ( .B1(n6500), .B2(n11784), .A(n8795), .ZN(n8445) );
  NOR2_X1 U10942 ( .A1(n8448), .A2(SI_14_), .ZN(n8451) );
  INV_X1 U10943 ( .A(n8447), .ZN(n8450) );
  NAND2_X1 U10944 ( .A1(n8448), .A2(SI_14_), .ZN(n8449) );
  INV_X1 U10945 ( .A(n8453), .ZN(n8454) );
  NAND2_X1 U10946 ( .A1(n8454), .A2(n10015), .ZN(n8455) );
  MUX2_X1 U10947 ( .A(n10652), .B(n15113), .S(n8622), .Z(n8457) );
  XNOR2_X1 U10948 ( .A(n8457), .B(SI_16_), .ZN(n8475) );
  NAND2_X1 U10949 ( .A1(n8457), .A2(n10077), .ZN(n8458) );
  MUX2_X1 U10950 ( .A(n10835), .B(n10836), .S(n9842), .Z(n8498) );
  XNOR2_X1 U10951 ( .A(n8498), .B(SI_17_), .ZN(n8496) );
  XNOR2_X1 U10952 ( .A(n8497), .B(n8496), .ZN(n10834) );
  NAND2_X1 U10953 ( .A1(n10834), .A2(n8758), .ZN(n8461) );
  NAND2_X1 U10954 ( .A1(n8479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8459) );
  XNOR2_X1 U10955 ( .A(n8459), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14721) );
  AOI22_X1 U10956 ( .A1(n8523), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8522), 
        .B2(n14721), .ZN(n8460) );
  NAND2_X1 U10957 ( .A1(n8469), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8510) );
  OR2_X1 U10958 ( .A1(n8469), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8462) );
  AND2_X1 U10959 ( .A1(n8510), .A2(n8462), .ZN(n14373) );
  NAND2_X1 U10960 ( .A1(n14373), .A2(n8708), .ZN(n8466) );
  NAND2_X1 U10961 ( .A1(n8512), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8465) );
  INV_X1 U10962 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14376) );
  OR2_X1 U10963 ( .A1(n8730), .A2(n14376), .ZN(n8463) );
  XNOR2_X1 U10964 ( .A(n14385), .B(n14350), .ZN(n8485) );
  NOR2_X1 U10965 ( .A1(n8467), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8468) );
  OR2_X1 U10966 ( .A1(n8469), .A2(n8468), .ZN(n14660) );
  INV_X1 U10967 ( .A(n14660), .ZN(n11921) );
  NAND2_X1 U10968 ( .A1(n11921), .A2(n8708), .ZN(n8474) );
  NAND2_X1 U10969 ( .A1(n8512), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8473) );
  INV_X1 U10970 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8470) );
  OR2_X1 U10971 ( .A1(n8179), .A2(n8470), .ZN(n8472) );
  INV_X1 U10972 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14169) );
  OR2_X1 U10973 ( .A1(n8730), .A2(n14169), .ZN(n8471) );
  NAND4_X1 U10974 ( .A1(n8474), .A2(n8473), .A3(n8472), .A4(n8471), .ZN(n14482) );
  INV_X1 U10975 ( .A(n14482), .ZN(n14382) );
  XNOR2_X1 U10976 ( .A(n8476), .B(n8475), .ZN(n10651) );
  NAND2_X1 U10977 ( .A1(n10651), .A2(n8758), .ZN(n8482) );
  NAND2_X1 U10978 ( .A1(n8477), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8478) );
  MUX2_X1 U10979 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8478), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8480) );
  AND2_X1 U10980 ( .A1(n8480), .A2(n8479), .ZN(n14168) );
  AOI22_X1 U10981 ( .A1(n8523), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8522), 
        .B2(n14168), .ZN(n8481) );
  INV_X1 U10982 ( .A(n14654), .ZN(n11924) );
  MUX2_X1 U10983 ( .A(n14382), .B(n11924), .S(n8791), .Z(n8491) );
  OR2_X1 U10984 ( .A1(n14385), .A2(n14350), .ZN(n11967) );
  NAND2_X1 U10985 ( .A1(n14385), .A2(n14350), .ZN(n11966) );
  AND2_X1 U10986 ( .A1(n8791), .A2(n14482), .ZN(n8483) );
  AOI21_X1 U10987 ( .B1(n14654), .B2(n8795), .A(n8483), .ZN(n8484) );
  NAND3_X1 U10988 ( .A1(n11967), .A2(n11966), .A3(n8484), .ZN(n8492) );
  OAI21_X1 U10989 ( .B1(n8485), .B2(n8491), .A(n8492), .ZN(n8486) );
  INV_X1 U10990 ( .A(n14350), .ZN(n14028) );
  AND2_X1 U10991 ( .A1(n8487), .A2(n14028), .ZN(n8489) );
  OAI21_X1 U10992 ( .B1(n14028), .B2(n8795), .A(n14385), .ZN(n8488) );
  OAI21_X1 U10993 ( .B1(n8489), .B2(n14385), .A(n8488), .ZN(n8490) );
  OAI21_X1 U10994 ( .B1(n8492), .B2(n8491), .A(n8490), .ZN(n8493) );
  INV_X1 U10995 ( .A(n8493), .ZN(n8494) );
  NAND2_X1 U10996 ( .A1(n8497), .A2(n8496), .ZN(n8500) );
  NAND2_X1 U10997 ( .A1(n8498), .A2(n10233), .ZN(n8499) );
  MUX2_X1 U10998 ( .A(n11020), .B(n11019), .S(n9842), .Z(n8502) );
  NAND2_X1 U10999 ( .A1(n8503), .A2(n8502), .ZN(n8504) );
  NAND2_X1 U11000 ( .A1(n8521), .A2(n8504), .ZN(n11021) );
  NAND2_X1 U11001 ( .A1(n8505), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8506) );
  XNOR2_X1 U11002 ( .A(n8506), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14184) );
  AOI22_X1 U11003 ( .A1(n8523), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8522), 
        .B2(n14184), .ZN(n8507) );
  AND2_X2 U11004 ( .A1(n8508), .A2(n8507), .ZN(n14476) );
  INV_X1 U11005 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U11006 ( .A1(n8510), .A2(n8509), .ZN(n8511) );
  AND2_X1 U11007 ( .A1(n8527), .A2(n8511), .ZN(n9800) );
  NAND2_X1 U11008 ( .A1(n9800), .A2(n8708), .ZN(n8517) );
  NAND2_X1 U11009 ( .A1(n8512), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8513) );
  AND2_X1 U11010 ( .A1(n8514), .A2(n8513), .ZN(n8516) );
  NAND2_X1 U11011 ( .A1(n8093), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8515) );
  OR2_X1 U11012 ( .A1(n14356), .A2(n14484), .ZN(n11989) );
  MUX2_X1 U11013 ( .A(n13964), .B(n14476), .S(n8795), .Z(n8518) );
  MUX2_X1 U11014 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9842), .Z(n8535) );
  NAND2_X1 U11015 ( .A1(n11235), .A2(n8758), .ZN(n8525) );
  AOI22_X1 U11016 ( .A1(n8523), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14195), 
        .B2(n8522), .ZN(n8524) );
  INV_X1 U11017 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8526) );
  AND2_X1 U11018 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  OR2_X1 U11019 ( .A1(n8528), .A2(n8545), .ZN(n14338) );
  AOI22_X1 U11020 ( .A1(n8512), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n8093), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8530) );
  OAI211_X1 U11021 ( .C1(n14338), .C2(n8689), .A(n8530), .B(n8529), .ZN(n14361) );
  XNOR2_X1 U11022 ( .A(n14470), .B(n14361), .ZN(n14333) );
  NAND2_X1 U11023 ( .A1(n14361), .A2(n8791), .ZN(n8533) );
  OR2_X1 U11024 ( .A1(n14361), .A2(n8791), .ZN(n8532) );
  MUX2_X1 U11025 ( .A(n8533), .B(n8532), .S(n14470), .Z(n8534) );
  NAND2_X1 U11026 ( .A1(n8538), .A2(n10640), .ZN(n8539) );
  INV_X1 U11027 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11539) );
  MUX2_X1 U11028 ( .A(n15074), .B(n11539), .S(n9842), .Z(n8540) );
  NAND2_X1 U11029 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U11030 ( .A1(n8553), .A2(n8542), .ZN(n11538) );
  OR2_X1 U11031 ( .A1(n11538), .A2(n8656), .ZN(n8544) );
  OR2_X1 U11032 ( .A1(n8157), .A2(n15074), .ZN(n8543) );
  OR2_X1 U11033 ( .A1(n8545), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U11034 ( .A1(n8545), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8562) );
  AND2_X1 U11035 ( .A1(n8546), .A2(n8562), .ZN(n14324) );
  NAND2_X1 U11036 ( .A1(n14324), .A2(n8708), .ZN(n8549) );
  NAND2_X1 U11037 ( .A1(n8093), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8547) );
  MUX2_X1 U11038 ( .A(n14322), .B(n13939), .S(n8795), .Z(n8551) );
  MUX2_X1 U11039 ( .A(n14027), .B(n14462), .S(n8795), .Z(n8550) );
  MUX2_X1 U11040 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9842), .Z(n8554) );
  NAND2_X1 U11041 ( .A1(n8554), .A2(SI_21_), .ZN(n8582) );
  OAI21_X1 U11042 ( .B1(n8554), .B2(SI_21_), .A(n8582), .ZN(n8555) );
  INV_X1 U11043 ( .A(n8555), .ZN(n8556) );
  OR2_X1 U11044 ( .A1(n8557), .A2(n8556), .ZN(n8558) );
  NAND2_X1 U11045 ( .A1(n8585), .A2(n8558), .ZN(n11574) );
  OR2_X1 U11046 ( .A1(n11574), .A2(n8656), .ZN(n8560) );
  OR2_X1 U11047 ( .A1(n8157), .A2(n11572), .ZN(n8559) );
  INV_X1 U11048 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8561) );
  OR2_X1 U11049 ( .A1(n8382), .A2(n8561), .ZN(n8566) );
  NAND2_X1 U11050 ( .A1(n8563), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8575) );
  OAI21_X1 U11051 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n8563), .A(n8575), .ZN(
        n14308) );
  OR2_X1 U11052 ( .A1(n8689), .A2(n14308), .ZN(n8565) );
  INV_X1 U11053 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14309) );
  OR2_X1 U11054 ( .A1(n8730), .A2(n14309), .ZN(n8564) );
  NAND4_X1 U11055 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n14326) );
  MUX2_X1 U11056 ( .A(n14455), .B(n14326), .S(n8791), .Z(n8571) );
  MUX2_X1 U11057 ( .A(n14455), .B(n14326), .S(n8795), .Z(n8568) );
  NAND2_X1 U11058 ( .A1(n8569), .A2(n8568), .ZN(n8573) );
  NAND2_X1 U11059 ( .A1(n8573), .A2(n8572), .ZN(n8589) );
  INV_X1 U11060 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8574) );
  OR2_X1 U11061 ( .A1(n8382), .A2(n8574), .ZN(n8579) );
  NAND2_X1 U11062 ( .A1(n8576), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8593) );
  OAI21_X1 U11063 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n8576), .A(n8593), .ZN(
        n14292) );
  OR2_X1 U11064 ( .A1(n8689), .A2(n14292), .ZN(n8578) );
  INV_X1 U11065 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14293) );
  OR2_X1 U11066 ( .A1(n8730), .A2(n14293), .ZN(n8577) );
  NAND4_X1 U11067 ( .A1(n8580), .A2(n8579), .A3(n8578), .A4(n8577), .ZN(n14026) );
  INV_X1 U11068 ( .A(SI_22_), .ZN(n8583) );
  AND2_X1 U11069 ( .A1(n8583), .A2(n8582), .ZN(n8584) );
  OR2_X1 U11070 ( .A1(n9369), .A2(n8622), .ZN(n8587) );
  XNOR2_X1 U11071 ( .A(n8587), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14537) );
  MUX2_X1 U11072 ( .A(n14026), .B(n14449), .S(n8791), .Z(n8590) );
  MUX2_X1 U11073 ( .A(n14026), .B(n14449), .S(n8795), .Z(n8588) );
  INV_X1 U11074 ( .A(n8590), .ZN(n8591) );
  INV_X1 U11075 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8592) );
  OR2_X1 U11076 ( .A1(n8382), .A2(n8592), .ZN(n8597) );
  NAND2_X1 U11077 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n8594), .ZN(n8611) );
  OAI21_X1 U11078 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8594), .A(n8611), .ZN(
        n14273) );
  OR2_X1 U11079 ( .A1(n8689), .A2(n14273), .ZN(n8596) );
  INV_X1 U11080 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14274) );
  OR2_X1 U11081 ( .A1(n8730), .A2(n14274), .ZN(n8595) );
  NAND4_X1 U11082 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n14297) );
  INV_X1 U11083 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8599) );
  MUX2_X1 U11084 ( .A(n8599), .B(n11748), .S(n9842), .Z(n9368) );
  MUX2_X1 U11085 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9842), .Z(n8618) );
  XNOR2_X1 U11086 ( .A(n8618), .B(SI_23_), .ZN(n8601) );
  XNOR2_X1 U11087 ( .A(n8619), .B(n8601), .ZN(n11862) );
  NAND2_X1 U11088 ( .A1(n11862), .A2(n8758), .ZN(n8603) );
  INV_X1 U11089 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11865) );
  OR2_X1 U11090 ( .A1(n8157), .A2(n11865), .ZN(n8602) );
  MUX2_X1 U11091 ( .A(n14297), .B(n14280), .S(n8795), .Z(n8606) );
  MUX2_X1 U11092 ( .A(n14297), .B(n14280), .S(n8791), .Z(n8604) );
  NAND2_X1 U11093 ( .A1(n8605), .A2(n8604), .ZN(n8608) );
  NAND2_X1 U11094 ( .A1(n8608), .A2(n8607), .ZN(n8630) );
  NAND2_X1 U11095 ( .A1(n8512), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8616) );
  INV_X1 U11096 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14505) );
  OR2_X1 U11097 ( .A1(n8179), .A2(n14505), .ZN(n8615) );
  INV_X1 U11098 ( .A(n8611), .ZN(n8609) );
  INV_X1 U11099 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U11100 ( .A1(n8611), .A2(n8610), .ZN(n8612) );
  NAND2_X1 U11101 ( .A1(n8658), .A2(n8612), .ZN(n14246) );
  OR2_X1 U11102 ( .A1(n8689), .A2(n14246), .ZN(n8614) );
  INV_X1 U11103 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14247) );
  OR2_X1 U11104 ( .A1(n8730), .A2(n14247), .ZN(n8613) );
  NAND4_X1 U11105 ( .A1(n8616), .A2(n8615), .A3(n8614), .A4(n8613), .ZN(n14276) );
  INV_X1 U11106 ( .A(n8618), .ZN(n8617) );
  NAND2_X1 U11107 ( .A1(n8620), .A2(n15168), .ZN(n8621) );
  MUX2_X1 U11108 ( .A(n14532), .B(n13804), .S(n8622), .Z(n8623) );
  NAND2_X1 U11109 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  NAND2_X1 U11110 ( .A1(n13802), .A2(n8758), .ZN(n8627) );
  OR2_X1 U11111 ( .A1(n8157), .A2(n14532), .ZN(n8626) );
  MUX2_X1 U11112 ( .A(n14276), .B(n14251), .S(n8795), .Z(n8631) );
  MUX2_X1 U11113 ( .A(n14251), .B(n14276), .S(n8795), .Z(n8628) );
  INV_X1 U11114 ( .A(n8628), .ZN(n8629) );
  NAND2_X1 U11115 ( .A1(n8512), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8637) );
  INV_X1 U11116 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8632) );
  OR2_X1 U11117 ( .A1(n8730), .A2(n8632), .ZN(n8636) );
  INV_X1 U11118 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13953) );
  XNOR2_X1 U11119 ( .A(n8658), .B(n13953), .ZN(n14235) );
  OR2_X1 U11120 ( .A1(n8689), .A2(n14235), .ZN(n8635) );
  INV_X1 U11121 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8633) );
  OR2_X1 U11122 ( .A1(n8179), .A2(n8633), .ZN(n8634) );
  NAND4_X1 U11123 ( .A1(n8637), .A2(n8636), .A3(n8635), .A4(n8634), .ZN(n14255) );
  MUX2_X1 U11124 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9842), .Z(n8648) );
  XNOR2_X1 U11125 ( .A(n8648), .B(SI_25_), .ZN(n8649) );
  XNOR2_X1 U11126 ( .A(n8650), .B(n8649), .ZN(n9411) );
  NAND2_X1 U11127 ( .A1(n9411), .A2(n8758), .ZN(n8641) );
  OR2_X1 U11128 ( .A1(n8157), .A2(n14529), .ZN(n8640) );
  MUX2_X1 U11129 ( .A(n14255), .B(n14425), .S(n8791), .Z(n8642) );
  NAND2_X1 U11130 ( .A1(n8643), .A2(n8642), .ZN(n8647) );
  MUX2_X1 U11131 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n9842), .Z(n8651) );
  NAND2_X1 U11132 ( .A1(n8651), .A2(SI_26_), .ZN(n8677) );
  OAI21_X1 U11133 ( .B1(n8651), .B2(SI_26_), .A(n8677), .ZN(n8652) );
  OR2_X2 U11134 ( .A1(n8653), .A2(n8652), .ZN(n8678) );
  NAND2_X1 U11135 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  NAND2_X1 U11136 ( .A1(n8678), .A2(n8654), .ZN(n14526) );
  OR2_X1 U11137 ( .A1(n8157), .A2(n14525), .ZN(n8655) );
  INV_X1 U11138 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8657) );
  OR2_X1 U11139 ( .A1(n8382), .A2(n8657), .ZN(n8664) );
  INV_X1 U11140 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14007) );
  OAI21_X1 U11141 ( .B1(n8658), .B2(n13953), .A(n14007), .ZN(n8661) );
  INV_X1 U11142 ( .A(n8658), .ZN(n8660) );
  AND2_X1 U11143 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n8659) );
  NAND2_X1 U11144 ( .A1(n8660), .A2(n8659), .ZN(n8671) );
  NAND2_X1 U11145 ( .A1(n8661), .A2(n8671), .ZN(n14222) );
  OR2_X1 U11146 ( .A1(n8689), .A2(n14222), .ZN(n8663) );
  INV_X1 U11147 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14220) );
  OR2_X1 U11148 ( .A1(n8730), .A2(n14220), .ZN(n8662) );
  NAND4_X1 U11149 ( .A1(n8665), .A2(n8664), .A3(n8663), .A4(n8662), .ZN(n14025) );
  MUX2_X1 U11150 ( .A(n14225), .B(n14025), .S(n8795), .Z(n8667) );
  MUX2_X1 U11151 ( .A(n14025), .B(n14225), .S(n8795), .Z(n8666) );
  INV_X1 U11152 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8668) );
  OR2_X1 U11153 ( .A1(n8382), .A2(n8668), .ZN(n8675) );
  INV_X1 U11154 ( .A(n8671), .ZN(n8669) );
  NAND2_X1 U11155 ( .A1(n8669), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8687) );
  INV_X1 U11156 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11157 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  NAND2_X1 U11158 ( .A1(n8687), .A2(n8672), .ZN(n13890) );
  OR2_X1 U11159 ( .A1(n8689), .A2(n13890), .ZN(n8674) );
  INV_X1 U11160 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n12046) );
  OR2_X1 U11161 ( .A1(n8730), .A2(n12046), .ZN(n8673) );
  NAND4_X1 U11162 ( .A1(n8676), .A2(n8675), .A3(n8674), .A4(n8673), .ZN(n14024) );
  NAND2_X2 U11163 ( .A1(n8678), .A2(n8677), .ZN(n8696) );
  MUX2_X1 U11164 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9842), .Z(n8697) );
  XNOR2_X1 U11165 ( .A(n8697), .B(SI_27_), .ZN(n8679) );
  INV_X1 U11166 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14522) );
  OR2_X1 U11167 ( .A1(n8157), .A2(n14522), .ZN(n8680) );
  MUX2_X1 U11168 ( .A(n14024), .B(n14412), .S(n8795), .Z(n8684) );
  NAND2_X1 U11169 ( .A1(n8683), .A2(n8684), .ZN(n8682) );
  MUX2_X1 U11170 ( .A(n14024), .B(n14412), .S(n8791), .Z(n8681) );
  INV_X1 U11171 ( .A(n8684), .ZN(n8685) );
  INV_X1 U11172 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n15056) );
  OR2_X1 U11173 ( .A1(n8382), .A2(n15056), .ZN(n8692) );
  INV_X1 U11174 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13929) );
  NAND2_X1 U11175 ( .A1(n8687), .A2(n13929), .ZN(n8688) );
  NAND2_X1 U11176 ( .A1(n12021), .A2(n8688), .ZN(n13930) );
  OR2_X1 U11177 ( .A1(n8689), .A2(n13930), .ZN(n8691) );
  INV_X1 U11178 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n12004) );
  OR2_X1 U11179 ( .A1(n8730), .A2(n12004), .ZN(n8690) );
  INV_X1 U11180 ( .A(n8697), .ZN(n8694) );
  NAND2_X1 U11181 ( .A1(n8694), .A2(n11664), .ZN(n8695) );
  NAND2_X1 U11182 ( .A1(n8697), .A2(SI_27_), .ZN(n8698) );
  INV_X1 U11183 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11963) );
  INV_X1 U11184 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9628) );
  MUX2_X1 U11185 ( .A(n11963), .B(n9628), .S(n9842), .Z(n8700) );
  INV_X1 U11186 ( .A(SI_28_), .ZN(n11813) );
  NAND2_X1 U11187 ( .A1(n8700), .A2(n11813), .ZN(n8713) );
  INV_X1 U11188 ( .A(n8700), .ZN(n8701) );
  NAND2_X1 U11189 ( .A1(n8701), .A2(SI_28_), .ZN(n8702) );
  NAND2_X1 U11190 ( .A1(n8713), .A2(n8702), .ZN(n8711) );
  NAND2_X1 U11191 ( .A1(n12250), .A2(n8758), .ZN(n8704) );
  OR2_X1 U11192 ( .A1(n8157), .A2(n11963), .ZN(n8703) );
  MUX2_X1 U11193 ( .A(n14401), .B(n13925), .S(n8352), .Z(n8706) );
  INV_X1 U11194 ( .A(n14401), .ZN(n14023) );
  MUX2_X1 U11195 ( .A(n14023), .B(n14407), .S(n8795), .Z(n8705) );
  INV_X1 U11196 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n15060) );
  INV_X1 U11197 ( .A(n12021), .ZN(n8707) );
  AOI22_X1 U11198 ( .A1(n8708), .A2(n8707), .B1(n8093), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n8710) );
  OAI211_X1 U11199 ( .C1(n8382), .C2(n15060), .A(n8710), .B(n8709), .ZN(n14022) );
  INV_X1 U11200 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12032) );
  INV_X1 U11201 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13787) );
  MUX2_X1 U11202 ( .A(n12032), .B(n13787), .S(n9842), .Z(n8720) );
  XNOR2_X1 U11203 ( .A(n8720), .B(SI_29_), .ZN(n8718) );
  NAND2_X1 U11204 ( .A1(n12232), .A2(n8758), .ZN(n8715) );
  OR2_X1 U11205 ( .A1(n8157), .A2(n12032), .ZN(n8714) );
  MUX2_X1 U11206 ( .A(n14404), .B(n14022), .S(n8795), .Z(n8717) );
  INV_X1 U11207 ( .A(SI_29_), .ZN(n13141) );
  NAND2_X1 U11208 ( .A1(n8720), .A2(n13141), .ZN(n8746) );
  MUX2_X1 U11209 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9842), .Z(n8721) );
  NAND2_X1 U11210 ( .A1(n8721), .A2(SI_30_), .ZN(n8749) );
  INV_X1 U11211 ( .A(n8721), .ZN(n8722) );
  INV_X1 U11212 ( .A(SI_30_), .ZN(n15053) );
  NAND2_X1 U11213 ( .A1(n8722), .A2(n15053), .ZN(n8747) );
  AND2_X1 U11214 ( .A1(n8749), .A2(n8747), .ZN(n8723) );
  NAND2_X1 U11215 ( .A1(n12217), .A2(n8758), .ZN(n8726) );
  INV_X1 U11216 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12055) );
  OR2_X1 U11217 ( .A1(n8157), .A2(n12055), .ZN(n8725) );
  INV_X1 U11218 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15070) );
  NAND2_X1 U11219 ( .A1(n8093), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U11220 ( .A1(n8512), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8727) );
  OAI211_X1 U11221 ( .C1(n8179), .C2(n15070), .A(n8728), .B(n8727), .ZN(n14021) );
  INV_X1 U11222 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8729) );
  OR2_X1 U11223 ( .A1(n8382), .A2(n8729), .ZN(n8734) );
  INV_X1 U11224 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14202) );
  OR2_X1 U11225 ( .A1(n8730), .A2(n14202), .ZN(n8733) );
  INV_X1 U11226 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8731) );
  OR2_X1 U11227 ( .A1(n8179), .A2(n8731), .ZN(n8732) );
  INV_X1 U11228 ( .A(n8735), .ZN(n8736) );
  OAI22_X1 U11229 ( .A1(n8791), .A2(n8794), .B1(n9655), .B2(n8736), .ZN(n8737)
         );
  AOI22_X1 U11230 ( .A1(n14210), .A2(n8791), .B1(n14021), .B2(n8737), .ZN(
        n8740) );
  NAND2_X1 U11231 ( .A1(n8739), .A2(n8740), .ZN(n8744) );
  NAND2_X1 U11232 ( .A1(n9655), .A2(n10797), .ZN(n10337) );
  OAI21_X1 U11233 ( .B1(n14204), .B2(n10337), .A(n14021), .ZN(n8738) );
  MUX2_X1 U11234 ( .A(n8738), .B(n14397), .S(n8795), .Z(n8743) );
  INV_X1 U11235 ( .A(n8739), .ZN(n8742) );
  INV_X1 U11236 ( .A(n8740), .ZN(n8741) );
  MUX2_X1 U11237 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9842), .Z(n8745) );
  INV_X1 U11238 ( .A(SI_31_), .ZN(n13130) );
  XNOR2_X1 U11239 ( .A(n8745), .B(n13130), .ZN(n8750) );
  NAND2_X1 U11240 ( .A1(n8750), .A2(n8749), .ZN(n8756) );
  NAND2_X1 U11241 ( .A1(n8747), .A2(n8746), .ZN(n8752) );
  NOR2_X1 U11242 ( .A1(n8752), .A2(n8750), .ZN(n8748) );
  NAND2_X1 U11243 ( .A1(n8757), .A2(n8748), .ZN(n8755) );
  INV_X1 U11244 ( .A(n8750), .ZN(n8753) );
  XNOR2_X1 U11245 ( .A(n8750), .B(n8749), .ZN(n8751) );
  OAI21_X1 U11246 ( .B1(n8753), .B2(n8752), .A(n8751), .ZN(n8754) );
  OAI211_X1 U11247 ( .C1(n8757), .C2(n8756), .A(n8755), .B(n8754), .ZN(n13782)
         );
  NAND2_X1 U11248 ( .A1(n13782), .A2(n8758), .ZN(n8760) );
  INV_X1 U11249 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14516) );
  OR2_X1 U11250 ( .A1(n8157), .A2(n14516), .ZN(n8759) );
  INV_X1 U11251 ( .A(n14536), .ZN(n10336) );
  NAND2_X1 U11252 ( .A1(n10336), .A2(n8138), .ZN(n8761) );
  NAND2_X1 U11253 ( .A1(n10334), .A2(n8761), .ZN(n8762) );
  NAND2_X1 U11254 ( .A1(n11196), .A2(n9655), .ZN(n10803) );
  NAND2_X1 U11255 ( .A1(n8762), .A2(n10803), .ZN(n8793) );
  INV_X1 U11256 ( .A(n8793), .ZN(n8763) );
  NAND2_X1 U11257 ( .A1(n14407), .A2(n14401), .ZN(n12011) );
  OR2_X1 U11258 ( .A1(n14407), .A2(n14401), .ZN(n8764) );
  NAND2_X1 U11259 ( .A1(n12011), .A2(n8764), .ZN(n12002) );
  NAND2_X1 U11260 ( .A1(n14412), .A2(n14005), .ZN(n11977) );
  INV_X1 U11261 ( .A(n14297), .ZN(n13996) );
  XNOR2_X1 U11262 ( .A(n14280), .B(n13996), .ZN(n11974) );
  INV_X1 U11263 ( .A(n14026), .ZN(n14278) );
  XNOR2_X1 U11264 ( .A(n14300), .B(n14278), .ZN(n11994) );
  XNOR2_X1 U11265 ( .A(n14356), .B(n14484), .ZN(n14348) );
  NAND2_X1 U11266 ( .A1(n6500), .A2(n8766), .ZN(n11927) );
  XNOR2_X1 U11267 ( .A(n11768), .B(n11872), .ZN(n11666) );
  NAND2_X1 U11268 ( .A1(n11431), .A2(n8767), .ZN(n8768) );
  NAND2_X1 U11269 ( .A1(n11352), .A2(n8768), .ZN(n11137) );
  INV_X1 U11270 ( .A(n14037), .ZN(n10968) );
  NAND2_X1 U11271 ( .A1(n11268), .A2(n10968), .ZN(n11165) );
  OR2_X1 U11272 ( .A1(n11268), .A2(n10968), .ZN(n8769) );
  INV_X1 U11273 ( .A(n14765), .ZN(n11175) );
  NAND2_X1 U11274 ( .A1(n11175), .A2(n14036), .ZN(n8770) );
  NAND2_X1 U11275 ( .A1(n14765), .A2(n11274), .ZN(n11148) );
  XNOR2_X1 U11276 ( .A(n6651), .B(n10718), .ZN(n11199) );
  NAND4_X1 U11277 ( .A1(n11446), .A2(n10931), .A3(n11199), .A4(n10724), .ZN(
        n8773) );
  XNOR2_X1 U11278 ( .A(n9693), .B(n11132), .ZN(n11093) );
  NOR2_X1 U11279 ( .A1(n8773), .A2(n11093), .ZN(n8774) );
  NAND4_X1 U11280 ( .A1(n11137), .A2(n11272), .A3(n11146), .A4(n8774), .ZN(
        n8776) );
  OR2_X1 U11281 ( .A1(n14792), .A2(n11764), .ZN(n11575) );
  NAND2_X1 U11282 ( .A1(n14792), .A2(n11764), .ZN(n8775) );
  NAND2_X1 U11283 ( .A1(n11575), .A2(n8775), .ZN(n11355) );
  INV_X1 U11284 ( .A(n14035), .ZN(n11149) );
  XNOR2_X1 U11285 ( .A(n11256), .B(n11149), .ZN(n11240) );
  OR4_X1 U11286 ( .A1(n8776), .A2(n11477), .A3(n11355), .A4(n11240), .ZN(n8777) );
  NOR2_X1 U11287 ( .A1(n11666), .A2(n8777), .ZN(n8778) );
  XNOR2_X1 U11288 ( .A(n11951), .B(n14031), .ZN(n11780) );
  XNOR2_X1 U11289 ( .A(n11889), .B(n14032), .ZN(n11735) );
  NAND4_X1 U11290 ( .A1(n11800), .A2(n8778), .A3(n11780), .A4(n11735), .ZN(
        n8779) );
  NOR2_X1 U11291 ( .A1(n11927), .A2(n8779), .ZN(n8780) );
  XNOR2_X1 U11292 ( .A(n14654), .B(n14482), .ZN(n11914) );
  OR2_X1 U11293 ( .A1(n14385), .A2(n14028), .ZN(n11987) );
  NAND2_X1 U11294 ( .A1(n14385), .A2(n14028), .ZN(n11988) );
  NAND2_X1 U11295 ( .A1(n11987), .A2(n11988), .ZN(n14368) );
  NAND4_X1 U11296 ( .A1(n14348), .A2(n8780), .A3(n11914), .A4(n14368), .ZN(
        n8781) );
  NOR2_X1 U11297 ( .A1(n14335), .A2(n8781), .ZN(n8782) );
  XNOR2_X1 U11298 ( .A(n14462), .B(n14027), .ZN(n14320) );
  XNOR2_X1 U11299 ( .A(n14455), .B(n14326), .ZN(n14304) );
  NAND4_X1 U11300 ( .A1(n11994), .A2(n8782), .A3(n14320), .A4(n14304), .ZN(
        n8783) );
  NOR2_X1 U11301 ( .A1(n11974), .A2(n8783), .ZN(n8784) );
  XNOR2_X1 U11302 ( .A(n14425), .B(n14255), .ZN(n14231) );
  NAND4_X1 U11303 ( .A1(n14217), .A2(n8784), .A3(n14231), .A4(n14253), .ZN(
        n8785) );
  XNOR2_X1 U11304 ( .A(n14404), .B(n14022), .ZN(n12016) );
  NAND3_X1 U11305 ( .A1(n8788), .A2(n8787), .A3(n12016), .ZN(n8789) );
  XNOR2_X1 U11306 ( .A(n14195), .B(n8789), .ZN(n8803) );
  NAND2_X1 U11307 ( .A1(n10797), .A2(n11573), .ZN(n8790) );
  INV_X1 U11308 ( .A(n8790), .ZN(n8802) );
  AND2_X1 U11309 ( .A1(n8793), .A2(n8790), .ZN(n8796) );
  NAND2_X1 U11310 ( .A1(n14204), .A2(n8796), .ZN(n8792) );
  NAND2_X1 U11311 ( .A1(n8791), .A2(n14204), .ZN(n8805) );
  MUX2_X1 U11312 ( .A(n8793), .B(n8792), .S(n8805), .Z(n8799) );
  NAND2_X1 U11313 ( .A1(n8795), .A2(n8794), .ZN(n8804) );
  INV_X1 U11314 ( .A(n8796), .ZN(n8807) );
  OAI21_X1 U11315 ( .B1(n14204), .B2(n8807), .A(n8804), .ZN(n8797) );
  OAI21_X1 U11316 ( .B1(n8763), .B2(n8804), .A(n8797), .ZN(n8798) );
  MUX2_X1 U11317 ( .A(n8799), .B(n8798), .S(n14392), .Z(n8800) );
  INV_X1 U11318 ( .A(n8800), .ZN(n8801) );
  INV_X1 U11319 ( .A(n8804), .ZN(n8808) );
  NOR2_X1 U11320 ( .A1(n14392), .A2(n8805), .ZN(n8806) );
  AOI211_X1 U11321 ( .C1(n8808), .C2(n14392), .A(n8807), .B(n8806), .ZN(n8809)
         );
  NAND3_X1 U11322 ( .A1(n8813), .A2(n8812), .A3(n8811), .ZN(n8820) );
  NAND2_X1 U11323 ( .A1(n8815), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8814) );
  MUX2_X1 U11324 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8814), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8818) );
  INV_X1 U11325 ( .A(n8815), .ZN(n8817) );
  NAND2_X1 U11326 ( .A1(n8818), .A2(n8822), .ZN(n9796) );
  INV_X1 U11327 ( .A(n9796), .ZN(n10029) );
  NAND2_X1 U11328 ( .A1(n10029), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11863) );
  NAND2_X1 U11329 ( .A1(n8820), .A2(n8819), .ZN(n8830) );
  INV_X1 U11330 ( .A(n10334), .ZN(n9772) );
  INV_X1 U11331 ( .A(n14055), .ZN(n10031) );
  INV_X1 U11332 ( .A(n14524), .ZN(n14708) );
  NAND2_X1 U11333 ( .A1(n8822), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8823) );
  NAND2_X1 U11334 ( .A1(n8821), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8826) );
  XNOR2_X1 U11335 ( .A(n8826), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U11336 ( .A1(n9789), .A2(n9775), .ZN(n8827) );
  NAND2_X1 U11337 ( .A1(n8138), .A2(n11239), .ZN(n9771) );
  NAND2_X1 U11338 ( .A1(n9772), .A2(n9771), .ZN(n10342) );
  NAND4_X1 U11339 ( .A1(n14483), .A2(n14708), .A3(n10343), .A4(n10342), .ZN(
        n8828) );
  OAI211_X1 U11340 ( .C1(n14536), .C2(n11863), .A(n8828), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8829) );
  NAND2_X1 U11341 ( .A1(n8830), .A2(n8829), .ZN(P1_U3242) );
  OAI21_X1 U11342 ( .B1(n12808), .B2(n12531), .A(n10641), .ZN(n8831) );
  INV_X4 U11343 ( .A(n8835), .ZN(n8907) );
  XNOR2_X1 U11344 ( .A(n13071), .B(n8907), .ZN(n12425) );
  INV_X1 U11345 ( .A(n12425), .ZN(n8896) );
  INV_X2 U11346 ( .A(n8907), .ZN(n8876) );
  XNOR2_X1 U11347 ( .A(n13077), .B(n8876), .ZN(n8832) );
  OAI21_X1 U11348 ( .B1(n12422), .B2(n12697), .A(n12892), .ZN(n8895) );
  NOR3_X1 U11349 ( .A1(n12422), .A2(n12697), .A3(n12892), .ZN(n8894) );
  NOR2_X1 U11350 ( .A1(n8832), .A2(n12903), .ZN(n8893) );
  INV_X2 U11351 ( .A(n8907), .ZN(n10396) );
  NAND3_X1 U11352 ( .A1(n12705), .A2(n8907), .A3(n8834), .ZN(n8837) );
  XNOR2_X1 U11353 ( .A(n8835), .B(n8834), .ZN(n8836) );
  NAND2_X1 U11354 ( .A1(n6618), .A2(n8836), .ZN(n8839) );
  NAND2_X1 U11355 ( .A1(n10399), .A2(n8839), .ZN(n10604) );
  XNOR2_X1 U11356 ( .A(n8907), .B(n10606), .ZN(n8840) );
  XNOR2_X1 U11357 ( .A(n8840), .B(n10402), .ZN(n10605) );
  INV_X1 U11358 ( .A(n8840), .ZN(n8841) );
  NAND2_X1 U11359 ( .A1(n8841), .A2(n10402), .ZN(n8842) );
  XNOR2_X1 U11360 ( .A(n8876), .B(n10584), .ZN(n8843) );
  XNOR2_X1 U11361 ( .A(n8843), .B(n10629), .ZN(n10582) );
  INV_X1 U11362 ( .A(n8843), .ZN(n8844) );
  NAND2_X1 U11363 ( .A1(n10616), .A2(n8844), .ZN(n8845) );
  XNOR2_X1 U11364 ( .A(n8876), .B(n10672), .ZN(n8846) );
  XNOR2_X1 U11365 ( .A(n8846), .B(n10885), .ZN(n10615) );
  NAND2_X1 U11366 ( .A1(n8846), .A2(n10885), .ZN(n8847) );
  XNOR2_X1 U11367 ( .A(n8907), .B(n11011), .ZN(n8848) );
  XNOR2_X1 U11368 ( .A(n8848), .B(n11002), .ZN(n10811) );
  INV_X1 U11369 ( .A(n8848), .ZN(n8849) );
  NAND2_X1 U11370 ( .A1(n8849), .A2(n11002), .ZN(n8850) );
  XNOR2_X1 U11371 ( .A(n8876), .B(n11066), .ZN(n8853) );
  XNOR2_X1 U11372 ( .A(n8853), .B(n11025), .ZN(n11114) );
  INV_X1 U11373 ( .A(n11114), .ZN(n8852) );
  INV_X1 U11374 ( .A(n8853), .ZN(n8854) );
  NAND2_X1 U11375 ( .A1(n12702), .A2(n8854), .ZN(n8855) );
  XNOR2_X1 U11376 ( .A(n12561), .B(n8907), .ZN(n11052) );
  NAND2_X1 U11377 ( .A1(n11053), .A2(n11052), .ZN(n11051) );
  INV_X1 U11378 ( .A(n11052), .ZN(n8856) );
  NAND2_X1 U11379 ( .A1(n8856), .A2(n12701), .ZN(n8857) );
  XNOR2_X1 U11380 ( .A(n10396), .B(n11471), .ZN(n8858) );
  XNOR2_X1 U11381 ( .A(n8858), .B(n11391), .ZN(n12378) );
  NAND2_X1 U11382 ( .A1(n12700), .A2(n8858), .ZN(n8859) );
  XNOR2_X1 U11383 ( .A(n12574), .B(n8876), .ZN(n8861) );
  XNOR2_X1 U11384 ( .A(n8861), .B(n8860), .ZN(n11383) );
  NAND2_X1 U11385 ( .A1(n8861), .A2(n8860), .ZN(n8862) );
  XNOR2_X1 U11386 ( .A(n11498), .B(n8907), .ZN(n8863) );
  XNOR2_X1 U11387 ( .A(n8863), .B(n11390), .ZN(n12359) );
  NAND2_X1 U11388 ( .A1(n8863), .A2(n14590), .ZN(n8864) );
  XNOR2_X1 U11389 ( .A(n11639), .B(n8907), .ZN(n8866) );
  INV_X1 U11390 ( .A(n14576), .ZN(n12362) );
  INV_X1 U11391 ( .A(n8865), .ZN(n8868) );
  INV_X1 U11392 ( .A(n8866), .ZN(n8867) );
  NAND2_X1 U11393 ( .A1(n8868), .A2(n8867), .ZN(n11633) );
  XNOR2_X1 U11394 ( .A(n14585), .B(n10396), .ZN(n11720) );
  AND2_X1 U11395 ( .A1(n11720), .A2(n11818), .ZN(n8870) );
  XNOR2_X1 U11396 ( .A(n14602), .B(n8907), .ZN(n8872) );
  NAND2_X1 U11397 ( .A1(n8872), .A2(n8871), .ZN(n11749) );
  INV_X1 U11398 ( .A(n8872), .ZN(n8873) );
  NAND2_X1 U11399 ( .A1(n8873), .A2(n14577), .ZN(n11750) );
  XNOR2_X1 U11400 ( .A(n12602), .B(n8907), .ZN(n8874) );
  XNOR2_X1 U11401 ( .A(n8874), .B(n12603), .ZN(n11880) );
  NAND2_X1 U11402 ( .A1(n8874), .A2(n12990), .ZN(n8875) );
  XNOR2_X1 U11403 ( .A(n13122), .B(n8907), .ZN(n11905) );
  XNOR2_X1 U11404 ( .A(n13115), .B(n8876), .ZN(n8877) );
  NAND2_X1 U11405 ( .A1(n8877), .A2(n7077), .ZN(n12403) );
  INV_X1 U11406 ( .A(n8877), .ZN(n8878) );
  NAND2_X1 U11407 ( .A1(n8878), .A2(n12991), .ZN(n12404) );
  XNOR2_X1 U11408 ( .A(n13109), .B(n8907), .ZN(n8879) );
  XNOR2_X1 U11409 ( .A(n8879), .B(n12955), .ZN(n12414) );
  NAND2_X1 U11410 ( .A1(n8879), .A2(n12981), .ZN(n8880) );
  XNOR2_X1 U11411 ( .A(n13032), .B(n8907), .ZN(n8881) );
  XNOR2_X1 U11412 ( .A(n8881), .B(n12941), .ZN(n12451) );
  NAND2_X1 U11413 ( .A1(n8881), .A2(n12969), .ZN(n8882) );
  XNOR2_X1 U11414 ( .A(n13098), .B(n8907), .ZN(n8883) );
  XNOR2_X1 U11415 ( .A(n8883), .B(n12926), .ZN(n12371) );
  INV_X1 U11416 ( .A(n8883), .ZN(n8884) );
  NAND2_X1 U11417 ( .A1(n8884), .A2(n12926), .ZN(n8885) );
  XNOR2_X1 U11418 ( .A(n12932), .B(n8907), .ZN(n8886) );
  XNOR2_X1 U11419 ( .A(n8886), .B(n12940), .ZN(n12434) );
  NAND2_X1 U11420 ( .A1(n8886), .A2(n12698), .ZN(n8887) );
  XNOR2_X1 U11421 ( .A(n13021), .B(n8907), .ZN(n8888) );
  XNOR2_X1 U11422 ( .A(n8888), .B(n12902), .ZN(n12388) );
  NAND2_X1 U11423 ( .A1(n12389), .A2(n12388), .ZN(n12387) );
  NAND2_X1 U11424 ( .A1(n8888), .A2(n12927), .ZN(n8889) );
  XNOR2_X1 U11425 ( .A(n13082), .B(n10396), .ZN(n8890) );
  INV_X1 U11426 ( .A(n8890), .ZN(n8891) );
  XNOR2_X1 U11427 ( .A(n13008), .B(n8907), .ZN(n8897) );
  XNOR2_X1 U11428 ( .A(n8897), .B(n12881), .ZN(n12396) );
  XNOR2_X1 U11429 ( .A(n13060), .B(n8907), .ZN(n8898) );
  XNOR2_X1 U11430 ( .A(n8898), .B(n8900), .ZN(n12462) );
  INV_X1 U11431 ( .A(n8898), .ZN(n8899) );
  XNOR2_X1 U11432 ( .A(n12662), .B(n8907), .ZN(n8901) );
  XNOR2_X1 U11433 ( .A(n8901), .B(n12696), .ZN(n12345) );
  NAND2_X1 U11434 ( .A1(n14522), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8903) );
  XNOR2_X1 U11435 ( .A(n9628), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8904) );
  XNOR2_X1 U11436 ( .A(n9627), .B(n8904), .ZN(n11811) );
  NAND2_X1 U11437 ( .A1(n11811), .A2(n12486), .ZN(n8906) );
  OR2_X1 U11438 ( .A1(n12487), .A2(n11813), .ZN(n8905) );
  NAND2_X1 U11439 ( .A1(n13054), .A2(n12349), .ZN(n12522) );
  XNOR2_X1 U11440 ( .A(n12663), .B(n8907), .ZN(n8908) );
  XNOR2_X1 U11441 ( .A(n8909), .B(n8908), .ZN(n8914) );
  NAND4_X1 U11442 ( .A1(n8918), .A2(n8910), .A3(n15026), .A4(n8916), .ZN(n8913) );
  OR2_X1 U11443 ( .A1(n8911), .A2(n8935), .ZN(n8912) );
  NAND2_X1 U11444 ( .A1(n8914), .A2(n12449), .ZN(n8945) );
  INV_X1 U11445 ( .A(n13054), .ZN(n9625) );
  OR2_X1 U11446 ( .A1(n8918), .A2(n12675), .ZN(n8915) );
  INV_X1 U11447 ( .A(n8916), .ZN(n8917) );
  OR2_X1 U11448 ( .A1(n8918), .A2(n8917), .ZN(n8923) );
  INV_X1 U11449 ( .A(n8920), .ZN(n12686) );
  NAND3_X1 U11450 ( .A1(n8935), .A2(n8921), .A3(n12686), .ZN(n8922) );
  NAND4_X1 U11451 ( .A1(n8923), .A2(n9654), .A3(n8922), .A4(n10351), .ZN(n8924) );
  NAND2_X1 U11452 ( .A1(n8924), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8928) );
  INV_X1 U11453 ( .A(n8935), .ZN(n8925) );
  OR2_X1 U11454 ( .A1(n12689), .A2(n8925), .ZN(n8926) );
  OR2_X1 U11455 ( .A1(n10130), .A2(P3_U3151), .ZN(n12693) );
  AND2_X1 U11456 ( .A1(n8926), .A2(n12693), .ZN(n8927) );
  INV_X1 U11457 ( .A(n8929), .ZN(n12818) );
  NAND2_X1 U11458 ( .A1(n8930), .A2(n12818), .ZN(n12477) );
  NAND2_X1 U11459 ( .A1(n6447), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U11460 ( .A1(n8931), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8933) );
  NAND2_X1 U11461 ( .A1(n6449), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8932) );
  OR2_X1 U11462 ( .A1(n12689), .A2(n8935), .ZN(n8938) );
  AOI22_X1 U11463 ( .A1(n6439), .A2(n12696), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8940) );
  OAI21_X1 U11464 ( .B1(n12837), .B2(n12455), .A(n8940), .ZN(n8941) );
  AOI21_X1 U11465 ( .B1(n12841), .B2(n12464), .A(n8941), .ZN(n8942) );
  INV_X1 U11466 ( .A(n8943), .ZN(n8944) );
  NAND2_X1 U11467 ( .A1(n8945), .A2(n8944), .ZN(P3_U3160) );
  NAND2_X1 U11468 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9087) );
  INV_X1 U11469 ( .A(n9087), .ZN(n8946) );
  NAND2_X1 U11470 ( .A1(n8946), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9107) );
  INV_X1 U11471 ( .A(n9107), .ZN(n8947) );
  NAND2_X1 U11472 ( .A1(n8947), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9124) );
  INV_X1 U11473 ( .A(n9124), .ZN(n8948) );
  NAND2_X1 U11474 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n8949) );
  INV_X1 U11475 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9229) );
  INV_X1 U11476 ( .A(n9284), .ZN(n8953) );
  NAND2_X1 U11477 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n8955) );
  INV_X1 U11478 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13238) );
  INV_X1 U11479 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13218) );
  INV_X1 U11480 ( .A(n9415), .ZN(n8958) );
  NAND2_X1 U11481 ( .A1(n8958), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9417) );
  INV_X1 U11482 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13257) );
  NAND2_X1 U11483 ( .A1(n9417), .A2(n13257), .ZN(n8959) );
  NAND2_X1 U11484 ( .A1(n9435), .A2(n8959), .ZN(n13459) );
  INV_X1 U11485 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9101) );
  INV_X1 U11486 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8961) );
  NOR2_X1 U11487 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n8965) );
  NOR2_X1 U11488 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .ZN(n8964) );
  NOR2_X1 U11489 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n8963) );
  NOR2_X1 U11490 ( .A1(n8999), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U11491 ( .A1(n9479), .A2(n8970), .ZN(n9455) );
  NOR3_X1 U11492 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .A3(P2_IR_REG_26__SCAN_IN), .ZN(n8971) );
  INV_X1 U11493 ( .A(n8971), .ZN(n8972) );
  INV_X1 U11494 ( .A(n9013), .ZN(n8973) );
  NAND2_X1 U11495 ( .A1(n8973), .A2(n9010), .ZN(n8977) );
  INV_X1 U11496 ( .A(n8977), .ZN(n8975) );
  NAND2_X1 U11497 ( .A1(n8975), .A2(n8974), .ZN(n13783) );
  OR2_X1 U11498 ( .A1(n13459), .A2(n9492), .ZN(n8985) );
  INV_X1 U11499 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13458) );
  INV_X1 U11500 ( .A(n8980), .ZN(n12053) );
  NAND2_X1 U11501 ( .A1(n12236), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U11502 ( .A1(n6647), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8981) );
  OAI211_X1 U11503 ( .C1(n13458), .C2(n12239), .A(n8982), .B(n8981), .ZN(n8983) );
  INV_X1 U11504 ( .A(n8983), .ZN(n8984) );
  NOR2_X1 U11505 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8989) );
  INV_X1 U11506 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8988) );
  INV_X1 U11507 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8987) );
  NAND4_X1 U11508 ( .A1(n8989), .A2(n8988), .A3(n8987), .A4(n8986), .ZN(n8990)
         );
  NOR2_X2 U11509 ( .A1(n9280), .A2(n8990), .ZN(n8994) );
  INV_X1 U11510 ( .A(n8994), .ZN(n8991) );
  INV_X1 U11511 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U11512 ( .A1(n8994), .A2(n8993), .ZN(n8995) );
  INV_X1 U11513 ( .A(n8999), .ZN(n9001) );
  NAND4_X1 U11514 ( .A1(n8998), .A2(n9003), .A3(n9002), .A4(n9057), .ZN(n9295)
         );
  NAND2_X1 U11515 ( .A1(n9005), .A2(n9004), .ZN(n9008) );
  OAI21_X1 U11516 ( .B1(n9008), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9007) );
  XNOR2_X1 U11517 ( .A(n9007), .B(n9006), .ZN(n10089) );
  XNOR2_X2 U11518 ( .A(n9009), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13330) );
  NAND2_X1 U11519 ( .A1(n13472), .A2(n9321), .ZN(n9429) );
  INV_X1 U11520 ( .A(n9429), .ZN(n9432) );
  BUF_X4 U11521 ( .A(n9033), .Z(n9862) );
  NAND2_X4 U11522 ( .A1(n9862), .A2(n9842), .ZN(n9038) );
  OR2_X1 U11523 ( .A1(n14526), .A2(n9038), .ZN(n9016) );
  NAND2_X1 U11524 ( .A1(n12251), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9015) );
  XNOR2_X1 U11525 ( .A(n13681), .B(n13164), .ZN(n9431) );
  NAND2_X1 U11526 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9017) );
  MUX2_X1 U11527 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9017), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9020) );
  INV_X1 U11528 ( .A(n9018), .ZN(n9019) );
  INV_X1 U11529 ( .A(n9952), .ZN(n9962) );
  NAND2_X1 U11530 ( .A1(n6460), .A2(n9962), .ZN(n9021) );
  NAND2_X1 U11531 ( .A1(n9026), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U11532 ( .A1(n9027), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U11533 ( .A1(n9045), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U11534 ( .A1(n6734), .A2(n9321), .ZN(n9035) );
  XNOR2_X1 U11535 ( .A(n10435), .B(n9035), .ZN(n10019) );
  NAND2_X1 U11536 ( .A1(n9045), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U11537 ( .A1(n12235), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9030) );
  NAND2_X1 U11538 ( .A1(n9026), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U11539 ( .A1(n9027), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11540 ( .A1(n9842), .A2(SI_0_), .ZN(n9032) );
  XNOR2_X1 U11541 ( .A(n9032), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13806) );
  NAND2_X1 U11542 ( .A1(n12064), .A2(n12059), .ZN(n10518) );
  OR2_X1 U11543 ( .A1(n10518), .A2(n9395), .ZN(n10083) );
  INV_X1 U11544 ( .A(n12059), .ZN(n12063) );
  NAND2_X1 U11545 ( .A1(n9331), .A2(n12063), .ZN(n9034) );
  AND2_X1 U11546 ( .A1(n10083), .A2(n9034), .ZN(n10020) );
  NAND2_X1 U11547 ( .A1(n10019), .A2(n10020), .ZN(n10436) );
  INV_X1 U11548 ( .A(n10435), .ZN(n9036) );
  NAND2_X1 U11549 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  NAND2_X1 U11550 ( .A1(n10436), .A2(n9037), .ZN(n9050) );
  NOR2_X1 U11551 ( .A1(n9844), .A2(n9038), .ZN(n9044) );
  INV_X1 U11552 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13784) );
  NOR2_X1 U11553 ( .A1(n9018), .A2(n13784), .ZN(n9039) );
  MUX2_X1 U11554 ( .A(n13784), .B(n9039), .S(P2_IR_REG_2__SCAN_IN), .Z(n9040)
         );
  INV_X1 U11555 ( .A(n9040), .ZN(n9042) );
  INV_X1 U11556 ( .A(n9057), .ZN(n9041) );
  NAND2_X1 U11557 ( .A1(n9042), .A2(n9041), .ZN(n14819) );
  OAI22_X1 U11558 ( .A1(n9244), .A2(n9843), .B1(n9862), .B2(n14819), .ZN(n9043) );
  XNOR2_X1 U11559 ( .A(n13164), .B(n12073), .ZN(n9051) );
  NAND2_X1 U11560 ( .A1(n9026), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11561 ( .A1(n9027), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11562 ( .A1(n9045), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U11563 ( .A1(n13295), .A2(n9255), .ZN(n9052) );
  XNOR2_X1 U11564 ( .A(n9051), .B(n9052), .ZN(n10437) );
  NAND2_X1 U11565 ( .A1(n9050), .A2(n10437), .ZN(n10443) );
  INV_X1 U11566 ( .A(n9051), .ZN(n9053) );
  NAND2_X1 U11567 ( .A1(n9053), .A2(n9052), .ZN(n9054) );
  NAND2_X1 U11568 ( .A1(n10443), .A2(n9054), .ZN(n10376) );
  OR2_X1 U11569 ( .A1(n9896), .A2(n9038), .ZN(n9061) );
  NOR2_X1 U11570 ( .A1(n9057), .A2(n13784), .ZN(n9055) );
  MUX2_X1 U11571 ( .A(n13784), .B(n9055), .S(P2_IR_REG_3__SCAN_IN), .Z(n9059)
         );
  NAND2_X1 U11572 ( .A1(n9057), .A2(n9056), .ZN(n9071) );
  INV_X1 U11573 ( .A(n9071), .ZN(n9058) );
  AOI22_X1 U11574 ( .A1(n12251), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6461), 
        .B2(n9883), .ZN(n9060) );
  XNOR2_X1 U11575 ( .A(n12087), .B(n9331), .ZN(n9066) );
  INV_X1 U11576 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9884) );
  OR2_X1 U11577 ( .A1(n12239), .A2(n9884), .ZN(n9065) );
  OR2_X1 U11578 ( .A1(n9492), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9064) );
  INV_X1 U11579 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9062) );
  NOR2_X1 U11580 ( .A1(n12088), .A2(n9395), .ZN(n9067) );
  NAND2_X1 U11581 ( .A1(n9066), .A2(n9067), .ZN(n9079) );
  INV_X1 U11582 ( .A(n9066), .ZN(n10386) );
  INV_X1 U11583 ( .A(n9067), .ZN(n9068) );
  NAND2_X1 U11584 ( .A1(n10386), .A2(n9068), .ZN(n9069) );
  NAND2_X1 U11585 ( .A1(n9079), .A2(n9069), .ZN(n10375) );
  NAND2_X1 U11586 ( .A1(n9839), .A2(n12249), .ZN(n9074) );
  NAND2_X1 U11587 ( .A1(n9071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9070) );
  MUX2_X1 U11588 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9070), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9072) );
  AND2_X1 U11589 ( .A1(n9072), .A2(n9098), .ZN(n9966) );
  AOI22_X1 U11590 ( .A1(n12251), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6461), 
        .B2(n9966), .ZN(n9073) );
  NAND2_X1 U11591 ( .A1(n9074), .A2(n9073), .ZN(n12095) );
  XNOR2_X1 U11592 ( .A(n12095), .B(n13164), .ZN(n9081) );
  NAND2_X1 U11593 ( .A1(n9045), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U11594 ( .A1(n12235), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9077) );
  OAI21_X1 U11595 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9087), .ZN(n10698) );
  OR2_X1 U11596 ( .A1(n9492), .A2(n10698), .ZN(n9076) );
  NAND2_X1 U11597 ( .A1(n9027), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9075) );
  NAND4_X1 U11598 ( .A1(n9078), .A2(n9077), .A3(n9076), .A4(n9075), .ZN(n13293) );
  NAND2_X1 U11599 ( .A1(n13293), .A2(n9255), .ZN(n9082) );
  XNOR2_X1 U11600 ( .A(n9081), .B(n9082), .ZN(n10387) );
  AND2_X1 U11601 ( .A1(n10387), .A2(n9079), .ZN(n9080) );
  INV_X1 U11602 ( .A(n9081), .ZN(n10364) );
  NAND2_X1 U11603 ( .A1(n9849), .A2(n12249), .ZN(n9085) );
  NAND2_X1 U11604 ( .A1(n9098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9083) );
  XNOR2_X1 U11605 ( .A(n9083), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U11606 ( .A1(n12251), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6461), 
        .B2(n9973), .ZN(n9084) );
  XNOR2_X1 U11607 ( .A(n12102), .B(n13164), .ZN(n9094) );
  INV_X2 U11608 ( .A(n12220), .ZN(n12236) );
  NAND2_X1 U11609 ( .A1(n12236), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U11610 ( .A1(n12235), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9091) );
  INV_X1 U11611 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U11612 ( .A1(n9087), .A2(n9086), .ZN(n9088) );
  NAND2_X1 U11613 ( .A1(n9107), .A2(n9088), .ZN(n10755) );
  OR2_X1 U11614 ( .A1(n9492), .A2(n10755), .ZN(n9090) );
  NAND2_X1 U11615 ( .A1(n9027), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9089) );
  NAND4_X1 U11616 ( .A1(n9092), .A2(n9091), .A3(n9090), .A4(n9089), .ZN(n13292) );
  NAND2_X1 U11617 ( .A1(n13292), .A2(n9255), .ZN(n9095) );
  XNOR2_X1 U11618 ( .A(n9094), .B(n9095), .ZN(n10363) );
  INV_X1 U11619 ( .A(n9094), .ZN(n9096) );
  NAND2_X1 U11620 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  INV_X1 U11621 ( .A(n9102), .ZN(n9099) );
  NAND2_X1 U11622 ( .A1(n9099), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9100) );
  MUX2_X1 U11623 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9100), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n9103) );
  NAND2_X1 U11624 ( .A1(n9102), .A2(n9101), .ZN(n9119) );
  AND2_X1 U11625 ( .A1(n9103), .A2(n9119), .ZN(n9999) );
  AOI22_X1 U11626 ( .A1(n12251), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6461), 
        .B2(n9999), .ZN(n9104) );
  XNOR2_X1 U11627 ( .A(n12109), .B(n9331), .ZN(n9113) );
  NAND2_X1 U11628 ( .A1(n12236), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9112) );
  INV_X1 U11629 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10000) );
  INV_X1 U11630 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U11631 ( .A1(n9107), .A2(n9106), .ZN(n9108) );
  NAND2_X1 U11632 ( .A1(n9124), .A2(n9108), .ZN(n10818) );
  OR2_X1 U11633 ( .A1(n9492), .A2(n10818), .ZN(n9110) );
  INV_X1 U11634 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10772) );
  OR2_X1 U11635 ( .A1(n12239), .A2(n10772), .ZN(n9109) );
  AND4_X2 U11636 ( .A1(n9112), .A2(n9111), .A3(n9110), .A4(n9109), .ZN(n12108)
         );
  NOR2_X1 U11637 ( .A1(n12108), .A2(n9395), .ZN(n9114) );
  NAND2_X1 U11638 ( .A1(n9113), .A2(n9114), .ZN(n9117) );
  INV_X1 U11639 ( .A(n9113), .ZN(n10644) );
  INV_X1 U11640 ( .A(n9114), .ZN(n9115) );
  NAND2_X1 U11641 ( .A1(n10644), .A2(n9115), .ZN(n9116) );
  NAND2_X1 U11642 ( .A1(n9117), .A2(n9116), .ZN(n10822) );
  NAND2_X1 U11643 ( .A1(n9119), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9118) );
  MUX2_X1 U11644 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9118), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n9120) );
  AND2_X1 U11645 ( .A1(n9120), .A2(n9137), .ZN(n10002) );
  AOI22_X1 U11646 ( .A1(n12251), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6461), 
        .B2(n10002), .ZN(n9121) );
  XNOR2_X1 U11647 ( .A(n12115), .B(n13164), .ZN(n9130) );
  NAND2_X1 U11648 ( .A1(n12236), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U11649 ( .A1(n12235), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9128) );
  INV_X1 U11650 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9123) );
  NAND2_X1 U11651 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  NAND2_X1 U11652 ( .A1(n9156), .A2(n9125), .ZN(n10788) );
  OR2_X1 U11653 ( .A1(n9492), .A2(n10788), .ZN(n9127) );
  NAND2_X1 U11654 ( .A1(n9027), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9126) );
  NAND4_X1 U11655 ( .A1(n9129), .A2(n9128), .A3(n9127), .A4(n9126), .ZN(n13290) );
  AND2_X1 U11656 ( .A1(n13290), .A2(n9255), .ZN(n9131) );
  NAND2_X1 U11657 ( .A1(n9130), .A2(n9131), .ZN(n9147) );
  INV_X1 U11658 ( .A(n9130), .ZN(n10870) );
  INV_X1 U11659 ( .A(n9131), .ZN(n9132) );
  NAND2_X1 U11660 ( .A1(n10870), .A2(n9132), .ZN(n9133) );
  AND2_X1 U11661 ( .A1(n9147), .A2(n9133), .ZN(n10642) );
  NAND2_X1 U11662 ( .A1(n9134), .A2(n10642), .ZN(n10869) );
  OR2_X1 U11663 ( .A1(n9988), .A2(n9038), .ZN(n9141) );
  NAND2_X1 U11664 ( .A1(n9137), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9136) );
  MUX2_X1 U11665 ( .A(n9136), .B(P2_IR_REG_31__SCAN_IN), .S(n9135), .Z(n9138)
         );
  NAND2_X1 U11666 ( .A1(n9138), .A2(n9167), .ZN(n10064) );
  OAI22_X1 U11667 ( .A1(n9244), .A2(n10166), .B1(n10064), .B2(n9862), .ZN(
        n9139) );
  INV_X1 U11668 ( .A(n9139), .ZN(n9140) );
  AND2_X2 U11669 ( .A1(n9141), .A2(n9140), .ZN(n14897) );
  XNOR2_X1 U11670 ( .A(n14897), .B(n9331), .ZN(n10974) );
  NAND2_X1 U11671 ( .A1(n12236), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9146) );
  INV_X1 U11672 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9142) );
  OR2_X1 U11673 ( .A1(n12218), .A2(n9142), .ZN(n9145) );
  INV_X1 U11674 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9155) );
  XNOR2_X1 U11675 ( .A(n9156), .B(n9155), .ZN(n10991) );
  OR2_X1 U11676 ( .A1(n9492), .A2(n10991), .ZN(n9144) );
  INV_X1 U11677 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10992) );
  OR2_X1 U11678 ( .A1(n12239), .A2(n10992), .ZN(n9143) );
  NAND2_X1 U11679 ( .A1(n13289), .A2(n9255), .ZN(n9148) );
  XNOR2_X1 U11680 ( .A(n10974), .B(n9148), .ZN(n10879) );
  NAND3_X1 U11681 ( .A1(n10869), .A2(n9147), .A3(n10879), .ZN(n10873) );
  INV_X1 U11682 ( .A(n10974), .ZN(n9149) );
  NAND2_X1 U11683 ( .A1(n9149), .A2(n9148), .ZN(n9150) );
  NAND2_X1 U11684 ( .A1(n10873), .A2(n9150), .ZN(n9162) );
  OR2_X1 U11685 ( .A1(n10014), .A2(n9038), .ZN(n9153) );
  NAND2_X1 U11686 ( .A1(n9167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9151) );
  XNOR2_X1 U11687 ( .A(n9151), .B(P2_IR_REG_9__SCAN_IN), .ZN(n14853) );
  AOI22_X1 U11688 ( .A1(n12251), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n14853), 
        .B2(n6461), .ZN(n9152) );
  NAND2_X2 U11689 ( .A1(n9153), .A2(n9152), .ZN(n12130) );
  XNOR2_X1 U11690 ( .A(n12130), .B(n13164), .ZN(n9163) );
  NAND2_X1 U11691 ( .A1(n6647), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11692 ( .A1(n12236), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9160) );
  INV_X1 U11693 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9154) );
  OAI21_X1 U11694 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9157) );
  NAND2_X1 U11695 ( .A1(n9157), .A2(n9172), .ZN(n11045) );
  OR2_X1 U11696 ( .A1(n9492), .A2(n11045), .ZN(n9159) );
  NAND2_X1 U11697 ( .A1(n9027), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9158) );
  NAND4_X1 U11698 ( .A1(n9161), .A2(n9160), .A3(n9159), .A4(n9158), .ZN(n13288) );
  NAND2_X1 U11699 ( .A1(n13288), .A2(n9255), .ZN(n9164) );
  XNOR2_X1 U11700 ( .A(n9163), .B(n9164), .ZN(n10975) );
  NAND2_X1 U11701 ( .A1(n9162), .A2(n10975), .ZN(n10981) );
  INV_X1 U11702 ( .A(n9163), .ZN(n9165) );
  NAND2_X1 U11703 ( .A1(n9165), .A2(n9164), .ZN(n9166) );
  NAND2_X1 U11704 ( .A1(n10079), .A2(n12249), .ZN(n9171) );
  INV_X1 U11705 ( .A(n9185), .ZN(n9168) );
  NAND2_X1 U11706 ( .A1(n9168), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9169) );
  XNOR2_X1 U11707 ( .A(n9169), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U11708 ( .A1(n10260), .A2(n6461), .B1(n12251), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n9170) );
  XNOR2_X1 U11709 ( .A(n13655), .B(n9331), .ZN(n9179) );
  NAND2_X1 U11710 ( .A1(n12236), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U11711 ( .A1(n6647), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9176) );
  INV_X1 U11712 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U11713 ( .A1(n9172), .A2(n11081), .ZN(n9173) );
  NAND2_X1 U11714 ( .A1(n9195), .A2(n9173), .ZN(n13652) );
  OR2_X1 U11715 ( .A1(n9492), .A2(n13652), .ZN(n9175) );
  NAND2_X1 U11716 ( .A1(n9027), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9174) );
  NAND4_X1 U11717 ( .A1(n9177), .A2(n9176), .A3(n9175), .A4(n9174), .ZN(n13287) );
  NAND2_X1 U11718 ( .A1(n13287), .A2(n9255), .ZN(n9180) );
  XNOR2_X1 U11719 ( .A(n9179), .B(n9180), .ZN(n11077) );
  INV_X1 U11720 ( .A(n11077), .ZN(n9178) );
  INV_X1 U11721 ( .A(n9179), .ZN(n9182) );
  INV_X1 U11722 ( .A(n9180), .ZN(n9181) );
  NAND2_X1 U11723 ( .A1(n9182), .A2(n9181), .ZN(n9183) );
  NAND2_X1 U11724 ( .A1(n10105), .A2(n12249), .ZN(n9192) );
  INV_X1 U11725 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9184) );
  INV_X1 U11726 ( .A(n9189), .ZN(n9186) );
  NAND2_X1 U11727 ( .A1(n9186), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9187) );
  MUX2_X1 U11728 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9187), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n9190) );
  INV_X1 U11729 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9188) );
  INV_X1 U11730 ( .A(n9208), .ZN(n9205) );
  AOI22_X1 U11731 ( .A1(n10597), .A2(n6461), .B1(n12251), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n9191) );
  XNOR2_X1 U11732 ( .A(n14908), .B(n9331), .ZN(n9204) );
  INV_X1 U11733 ( .A(n9204), .ZN(n9202) );
  NAND2_X1 U11734 ( .A1(n12236), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9200) );
  INV_X1 U11735 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9193) );
  OR2_X1 U11736 ( .A1(n12218), .A2(n9193), .ZN(n9199) );
  NAND2_X1 U11737 ( .A1(n9195), .A2(n9194), .ZN(n9196) );
  NAND2_X1 U11738 ( .A1(n9214), .A2(n9196), .ZN(n11372) );
  OR2_X1 U11739 ( .A1(n9492), .A2(n11372), .ZN(n9198) );
  INV_X1 U11740 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11373) );
  OR2_X1 U11741 ( .A1(n12239), .A2(n11373), .ZN(n9197) );
  NOR2_X1 U11742 ( .A1(n12141), .A2(n9395), .ZN(n9203) );
  INV_X1 U11743 ( .A(n9203), .ZN(n9201) );
  AND2_X1 U11744 ( .A1(n9204), .A2(n9203), .ZN(n11180) );
  NAND2_X1 U11745 ( .A1(n10358), .A2(n12249), .ZN(n9212) );
  NAND2_X1 U11746 ( .A1(n9205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9206) );
  MUX2_X1 U11747 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9206), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9209) );
  INV_X1 U11748 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U11749 ( .A1(n9208), .A2(n9207), .ZN(n9241) );
  NAND2_X1 U11750 ( .A1(n9209), .A2(n9241), .ZN(n10684) );
  OAI22_X1 U11751 ( .A1(n10684), .A2(n9862), .B1(n9244), .B2(n15054), .ZN(
        n9210) );
  INV_X1 U11752 ( .A(n9210), .ZN(n9211) );
  XNOR2_X1 U11753 ( .A(n14631), .B(n13164), .ZN(n9220) );
  NAND2_X1 U11754 ( .A1(n12236), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9219) );
  INV_X1 U11755 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9213) );
  OR2_X1 U11756 ( .A1(n12218), .A2(n9213), .ZN(n9218) );
  INV_X1 U11757 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10594) );
  NAND2_X1 U11758 ( .A1(n9214), .A2(n10594), .ZN(n9215) );
  NAND2_X1 U11759 ( .A1(n9230), .A2(n9215), .ZN(n11511) );
  OR2_X1 U11760 ( .A1(n9492), .A2(n11511), .ZN(n9217) );
  INV_X1 U11761 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11512) );
  OR2_X1 U11762 ( .A1(n12239), .A2(n11512), .ZN(n9216) );
  NAND2_X1 U11763 ( .A1(n13285), .A2(n9255), .ZN(n9221) );
  NAND2_X1 U11764 ( .A1(n9220), .A2(n9221), .ZN(n9225) );
  INV_X1 U11765 ( .A(n9220), .ZN(n9223) );
  INV_X1 U11766 ( .A(n9221), .ZN(n9222) );
  NAND2_X1 U11767 ( .A1(n9223), .A2(n9222), .ZN(n9224) );
  AND2_X1 U11768 ( .A1(n9225), .A2(n9224), .ZN(n11300) );
  NAND2_X1 U11769 ( .A1(n11298), .A2(n9225), .ZN(n11435) );
  NAND2_X1 U11770 ( .A1(n10408), .A2(n12249), .ZN(n9228) );
  NAND2_X1 U11771 ( .A1(n9241), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9226) );
  AOI22_X1 U11772 ( .A1(n11122), .A2(n6461), .B1(n12251), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n9227) );
  XNOR2_X1 U11773 ( .A(n12157), .B(n9331), .ZN(n9236) );
  NAND2_X1 U11774 ( .A1(n6647), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9235) );
  NAND2_X1 U11775 ( .A1(n12236), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U11776 ( .A1(n9230), .A2(n9229), .ZN(n9231) );
  NAND2_X1 U11777 ( .A1(n9249), .A2(n9231), .ZN(n11436) );
  OR2_X1 U11778 ( .A1(n9492), .A2(n11436), .ZN(n9233) );
  NAND2_X1 U11779 ( .A1(n9027), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9232) );
  NAND4_X1 U11780 ( .A1(n9235), .A2(n9234), .A3(n9233), .A4(n9232), .ZN(n13284) );
  NAND2_X1 U11781 ( .A1(n13284), .A2(n9255), .ZN(n9237) );
  XNOR2_X1 U11782 ( .A(n9236), .B(n9237), .ZN(n11434) );
  INV_X1 U11783 ( .A(n9236), .ZN(n9239) );
  INV_X1 U11784 ( .A(n9237), .ZN(n9238) );
  NAND2_X1 U11785 ( .A1(n9239), .A2(n9238), .ZN(n9240) );
  OAI21_X1 U11786 ( .B1(n9241), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9243) );
  INV_X1 U11787 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n9242) );
  OAI22_X1 U11788 ( .A1(n11524), .A2(n9862), .B1(n9244), .B2(n10638), .ZN(
        n9245) );
  INV_X1 U11789 ( .A(n9245), .ZN(n9246) );
  XNOR2_X1 U11790 ( .A(n14620), .B(n9331), .ZN(n9256) );
  NAND2_X1 U11791 ( .A1(n6647), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U11792 ( .A1(n9249), .A2(n9248), .ZN(n9250) );
  AND2_X1 U11793 ( .A1(n9271), .A2(n9250), .ZN(n11614) );
  NAND2_X1 U11794 ( .A1(n9026), .A2(n11614), .ZN(n9253) );
  NAND2_X1 U11795 ( .A1(n9027), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11796 ( .A1(n12236), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9251) );
  NAND4_X1 U11797 ( .A1(n9254), .A2(n9253), .A3(n9252), .A4(n9251), .ZN(n13388) );
  NAND2_X1 U11798 ( .A1(n13388), .A2(n9255), .ZN(n9257) );
  NAND2_X1 U11799 ( .A1(n9256), .A2(n9257), .ZN(n9262) );
  INV_X1 U11800 ( .A(n9256), .ZN(n9259) );
  INV_X1 U11801 ( .A(n9257), .ZN(n9258) );
  NAND2_X1 U11802 ( .A1(n9259), .A2(n9258), .ZN(n9260) );
  NAND2_X1 U11803 ( .A1(n9262), .A2(n9260), .ZN(n11613) );
  NAND2_X1 U11804 ( .A1(n10917), .A2(n12249), .ZN(n9267) );
  NAND2_X1 U11805 ( .A1(n9456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9264) );
  MUX2_X1 U11806 ( .A(n9264), .B(P2_IR_REG_31__SCAN_IN), .S(n9263), .Z(n9265)
         );
  NAND2_X1 U11807 ( .A1(n9265), .A2(n9280), .ZN(n11602) );
  INV_X1 U11808 ( .A(n11602), .ZN(n11596) );
  AOI22_X1 U11809 ( .A1(n12251), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6461), 
        .B2(n11596), .ZN(n9266) );
  XNOR2_X1 U11810 ( .A(n13781), .B(n9331), .ZN(n9276) );
  NAND2_X1 U11811 ( .A1(n6647), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U11812 ( .A1(n12236), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9268) );
  AND2_X1 U11813 ( .A1(n9269), .A2(n9268), .ZN(n9275) );
  INV_X1 U11814 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11815 ( .A1(n9271), .A2(n9270), .ZN(n9272) );
  NAND2_X1 U11816 ( .A1(n9284), .A2(n9272), .ZN(n13637) );
  OR2_X1 U11817 ( .A1(n13637), .A2(n9492), .ZN(n9274) );
  NAND2_X1 U11818 ( .A1(n9027), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9273) );
  NOR2_X1 U11819 ( .A1(n13389), .A2(n9395), .ZN(n13271) );
  INV_X1 U11820 ( .A(n9276), .ZN(n9277) );
  NOR2_X1 U11821 ( .A1(n9278), .A2(n9277), .ZN(n9279) );
  NAND2_X1 U11822 ( .A1(n10651), .A2(n12249), .ZN(n9283) );
  NAND2_X1 U11823 ( .A1(n9280), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9281) );
  XNOR2_X1 U11824 ( .A(n9281), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U11825 ( .A1(n12251), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6461), 
        .B2(n11832), .ZN(n9282) );
  XNOR2_X1 U11826 ( .A(n13390), .B(n13164), .ZN(n9289) );
  INV_X1 U11827 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U11828 ( .A1(n9284), .A2(n13198), .ZN(n9285) );
  NAND2_X1 U11829 ( .A1(n9299), .A2(n9285), .ZN(n13618) );
  OR2_X1 U11830 ( .A1(n13618), .A2(n9492), .ZN(n9288) );
  AOI22_X1 U11831 ( .A1(n9027), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n6647), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n9287) );
  NAND2_X1 U11832 ( .A1(n12236), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9286) );
  OR2_X1 U11833 ( .A1(n13633), .A2(n9395), .ZN(n9290) );
  NAND2_X1 U11834 ( .A1(n9289), .A2(n9290), .ZN(n9294) );
  INV_X1 U11835 ( .A(n9289), .ZN(n9292) );
  INV_X1 U11836 ( .A(n9290), .ZN(n9291) );
  NAND2_X1 U11837 ( .A1(n9292), .A2(n9291), .ZN(n9293) );
  AND2_X1 U11838 ( .A1(n9294), .A2(n9293), .ZN(n13194) );
  NAND2_X1 U11839 ( .A1(n10834), .A2(n12249), .ZN(n9298) );
  NAND2_X1 U11840 ( .A1(n9295), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9296) );
  XNOR2_X1 U11841 ( .A(n9296), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U11842 ( .A1(n12251), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6461), 
        .B2(n13313), .ZN(n9297) );
  XNOR2_X1 U11843 ( .A(n13604), .B(n13164), .ZN(n9304) );
  NAND2_X1 U11844 ( .A1(n9299), .A2(n11828), .ZN(n9300) );
  AND2_X1 U11845 ( .A1(n9314), .A2(n9300), .ZN(n13601) );
  NAND2_X1 U11846 ( .A1(n13601), .A2(n9026), .ZN(n9303) );
  AOI22_X1 U11847 ( .A1(n12236), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n6647), 
        .B2(P2_REG1_REG_17__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U11848 ( .A1(n9027), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9301) );
  OR2_X1 U11849 ( .A1(n13393), .A2(n9395), .ZN(n9305) );
  NAND2_X1 U11850 ( .A1(n9304), .A2(n9305), .ZN(n9309) );
  INV_X1 U11851 ( .A(n9304), .ZN(n9307) );
  INV_X1 U11852 ( .A(n9305), .ZN(n9306) );
  NAND2_X1 U11853 ( .A1(n9307), .A2(n9306), .ZN(n9308) );
  AND2_X1 U11854 ( .A1(n9309), .A2(n9308), .ZN(n13206) );
  OR2_X1 U11855 ( .A1(n11021), .A2(n9038), .ZN(n9313) );
  NAND2_X1 U11856 ( .A1(n9310), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9311) );
  XNOR2_X1 U11857 ( .A(n9311), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14864) );
  AOI22_X1 U11858 ( .A1(n12251), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6461), 
        .B2(n14864), .ZN(n9312) );
  XNOR2_X1 U11859 ( .A(n13593), .B(n13164), .ZN(n9322) );
  INV_X1 U11860 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13248) );
  NAND2_X1 U11861 ( .A1(n9314), .A2(n13248), .ZN(n9315) );
  NAND2_X1 U11862 ( .A1(n9341), .A2(n9315), .ZN(n13589) );
  OR2_X1 U11863 ( .A1(n13589), .A2(n9492), .ZN(n9320) );
  INV_X1 U11864 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n14861) );
  NAND2_X1 U11865 ( .A1(n6647), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11866 ( .A1(n12236), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9316) );
  OAI211_X1 U11867 ( .C1(n12239), .C2(n14861), .A(n9317), .B(n9316), .ZN(n9318) );
  INV_X1 U11868 ( .A(n9318), .ZN(n9319) );
  NAND2_X1 U11869 ( .A1(n13359), .A2(n9255), .ZN(n9323) );
  XNOR2_X1 U11870 ( .A(n9322), .B(n9323), .ZN(n13245) );
  INV_X1 U11871 ( .A(n9322), .ZN(n9325) );
  INV_X1 U11872 ( .A(n9323), .ZN(n9324) );
  NAND2_X1 U11873 ( .A1(n9325), .A2(n9324), .ZN(n9326) );
  NAND2_X1 U11874 ( .A1(n11235), .A2(n12249), .ZN(n9328) );
  AOI22_X1 U11875 ( .A1(n12251), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6461), 
        .B2(n13330), .ZN(n9327) );
  XNOR2_X1 U11876 ( .A(n13578), .B(n9331), .ZN(n13151) );
  NAND2_X1 U11877 ( .A1(n12251), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9329) );
  XNOR2_X1 U11878 ( .A(n13715), .B(n9331), .ZN(n9349) );
  INV_X1 U11879 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9333) );
  INV_X1 U11880 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9332) );
  OAI21_X1 U11881 ( .B1(n9341), .B2(n9333), .A(n9332), .ZN(n9334) );
  AND2_X1 U11882 ( .A1(n9334), .A2(n9354), .ZN(n13562) );
  NAND2_X1 U11883 ( .A1(n13562), .A2(n9026), .ZN(n9340) );
  INV_X1 U11884 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U11885 ( .A1(n12236), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11886 ( .A1(n6647), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9335) );
  OAI211_X1 U11887 ( .C1(n9337), .C2(n12239), .A(n9336), .B(n9335), .ZN(n9338)
         );
  INV_X1 U11888 ( .A(n9338), .ZN(n9339) );
  NAND2_X1 U11889 ( .A1(n9340), .A2(n9339), .ZN(n13543) );
  NAND2_X1 U11890 ( .A1(n13543), .A2(n9255), .ZN(n9348) );
  XNOR2_X1 U11891 ( .A(n9349), .B(n9348), .ZN(n13229) );
  XNOR2_X1 U11892 ( .A(n9341), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n13576) );
  NAND2_X1 U11893 ( .A1(n13576), .A2(n9026), .ZN(n9346) );
  INV_X1 U11894 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U11895 ( .A1(n12236), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U11896 ( .A1(n9027), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9342) );
  OAI211_X1 U11897 ( .C1(n12218), .C2(n13324), .A(n9343), .B(n9342), .ZN(n9344) );
  INV_X1 U11898 ( .A(n9344), .ZN(n9345) );
  NOR2_X1 U11899 ( .A1(n13247), .A2(n9395), .ZN(n13152) );
  NAND2_X1 U11900 ( .A1(n9349), .A2(n9348), .ZN(n9350) );
  OR2_X1 U11901 ( .A1(n11574), .A2(n9038), .ZN(n9352) );
  NAND2_X1 U11902 ( .A1(n12251), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9351) );
  XNOR2_X1 U11903 ( .A(n13552), .B(n13164), .ZN(n9363) );
  INV_X1 U11904 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U11905 ( .A1(n9354), .A2(n9353), .ZN(n9355) );
  NAND2_X1 U11906 ( .A1(n9373), .A2(n9355), .ZN(n13549) );
  OR2_X1 U11907 ( .A1(n13549), .A2(n9492), .ZN(n9361) );
  INV_X1 U11908 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11909 ( .A1(n12236), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U11910 ( .A1(n6647), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9356) );
  OAI211_X1 U11911 ( .C1(n9358), .C2(n12239), .A(n9357), .B(n9356), .ZN(n9359)
         );
  INV_X1 U11912 ( .A(n9359), .ZN(n9360) );
  NAND2_X1 U11913 ( .A1(n13524), .A2(n9255), .ZN(n9364) );
  XNOR2_X1 U11914 ( .A(n9363), .B(n9364), .ZN(n13175) );
  INV_X1 U11915 ( .A(n13175), .ZN(n9362) );
  INV_X1 U11916 ( .A(n9363), .ZN(n9366) );
  INV_X1 U11917 ( .A(n9364), .ZN(n9365) );
  NAND2_X1 U11918 ( .A1(n9366), .A2(n9365), .ZN(n9367) );
  NAND2_X1 U11919 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  NAND2_X1 U11920 ( .A1(n12251), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9372) );
  XNOR2_X1 U11921 ( .A(n13526), .B(n13164), .ZN(n9380) );
  NAND2_X1 U11922 ( .A1(n9373), .A2(n13238), .ZN(n9374) );
  AND2_X1 U11923 ( .A1(n9387), .A2(n9374), .ZN(n13530) );
  NAND2_X1 U11924 ( .A1(n13530), .A2(n9026), .ZN(n9379) );
  INV_X1 U11925 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13532) );
  NAND2_X1 U11926 ( .A1(n12236), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11927 ( .A1(n6647), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9375) );
  OAI211_X1 U11928 ( .C1(n13532), .C2(n12239), .A(n9376), .B(n9375), .ZN(n9377) );
  INV_X1 U11929 ( .A(n9377), .ZN(n9378) );
  OR2_X1 U11930 ( .A1(n13233), .A2(n9395), .ZN(n13234) );
  INV_X1 U11931 ( .A(n9380), .ZN(n9381) );
  NOR2_X1 U11932 ( .A1(n9382), .A2(n9381), .ZN(n9383) );
  AOI21_X1 U11933 ( .B1(n13235), .B2(n13234), .A(n9383), .ZN(n9398) );
  NAND2_X1 U11934 ( .A1(n11862), .A2(n12249), .ZN(n9385) );
  NAND2_X1 U11935 ( .A1(n12251), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9384) );
  XNOR2_X1 U11936 ( .A(n13698), .B(n13164), .ZN(n9397) );
  INV_X1 U11937 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U11938 ( .A1(n9387), .A2(n9386), .ZN(n9388) );
  NAND2_X1 U11939 ( .A1(n9401), .A2(n9388), .ZN(n13145) );
  OR2_X1 U11940 ( .A1(n13145), .A2(n9492), .ZN(n9394) );
  INV_X1 U11941 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9391) );
  NAND2_X1 U11942 ( .A1(n12236), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U11943 ( .A1(n6647), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9389) );
  OAI211_X1 U11944 ( .C1(n9391), .C2(n12239), .A(n9390), .B(n9389), .ZN(n9392)
         );
  INV_X1 U11945 ( .A(n9392), .ZN(n9393) );
  NOR2_X1 U11946 ( .A1(n13406), .A2(n9395), .ZN(n9396) );
  NAND2_X1 U11947 ( .A1(n13802), .A2(n12249), .ZN(n9400) );
  NAND2_X1 U11948 ( .A1(n12251), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9399) );
  XNOR2_X1 U11949 ( .A(n13692), .B(n13164), .ZN(n13184) );
  NAND2_X1 U11950 ( .A1(n9401), .A2(n13218), .ZN(n9402) );
  AND2_X1 U11951 ( .A1(n9415), .A2(n9402), .ZN(n13497) );
  NAND2_X1 U11952 ( .A1(n13497), .A2(n9026), .ZN(n9408) );
  INV_X1 U11953 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U11954 ( .A1(n12236), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9404) );
  NAND2_X1 U11955 ( .A1(n6647), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9403) );
  OAI211_X1 U11956 ( .C1(n9405), .C2(n12239), .A(n9404), .B(n9403), .ZN(n9406)
         );
  INV_X1 U11957 ( .A(n9406), .ZN(n9407) );
  NAND2_X1 U11958 ( .A1(n9408), .A2(n9407), .ZN(n13408) );
  AND2_X1 U11959 ( .A1(n13408), .A2(n9255), .ZN(n9409) );
  NAND2_X1 U11960 ( .A1(n13184), .A2(n9409), .ZN(n9410) );
  OAI21_X1 U11961 ( .B1(n13184), .B2(n9409), .A(n9410), .ZN(n13214) );
  INV_X1 U11962 ( .A(n9410), .ZN(n9428) );
  NAND2_X1 U11963 ( .A1(n9411), .A2(n12249), .ZN(n9413) );
  NAND2_X1 U11964 ( .A1(n12251), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9412) );
  XNOR2_X1 U11965 ( .A(n13763), .B(n13164), .ZN(n9424) );
  INV_X1 U11966 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11967 ( .A1(n9415), .A2(n9414), .ZN(n9416) );
  NAND2_X1 U11968 ( .A1(n9417), .A2(n9416), .ZN(n13187) );
  OR2_X1 U11969 ( .A1(n13187), .A2(n9492), .ZN(n9423) );
  INV_X1 U11970 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9420) );
  NAND2_X1 U11971 ( .A1(n6647), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9419) );
  NAND2_X1 U11972 ( .A1(n12236), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9418) );
  OAI211_X1 U11973 ( .C1(n9420), .C2(n12239), .A(n9419), .B(n9418), .ZN(n9421)
         );
  INV_X1 U11974 ( .A(n9421), .ZN(n9422) );
  NAND2_X1 U11975 ( .A1(n9423), .A2(n9422), .ZN(n13455) );
  AND2_X1 U11976 ( .A1(n13455), .A2(n9321), .ZN(n9425) );
  NAND2_X1 U11977 ( .A1(n9424), .A2(n9425), .ZN(n9430) );
  INV_X1 U11978 ( .A(n9424), .ZN(n13263) );
  INV_X1 U11979 ( .A(n9425), .ZN(n9426) );
  NAND2_X1 U11980 ( .A1(n13263), .A2(n9426), .ZN(n9427) );
  AND2_X1 U11981 ( .A1(n9430), .A2(n9427), .ZN(n13183) );
  XNOR2_X1 U11982 ( .A(n9431), .B(n9429), .ZN(n13264) );
  NAND2_X1 U11983 ( .A1(n13794), .A2(n12249), .ZN(n9434) );
  NAND2_X1 U11984 ( .A1(n12251), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9433) );
  XNOR2_X1 U11985 ( .A(n13446), .B(n13164), .ZN(n9443) );
  INV_X1 U11986 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U11987 ( .A1(n9435), .A2(n9507), .ZN(n9436) );
  NAND2_X1 U11988 ( .A1(n9502), .A2(n9026), .ZN(n9441) );
  INV_X1 U11989 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13439) );
  NAND2_X1 U11990 ( .A1(n12236), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9438) );
  NAND2_X1 U11991 ( .A1(n6647), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9437) );
  OAI211_X1 U11992 ( .C1(n13439), .C2(n12239), .A(n9438), .B(n9437), .ZN(n9439) );
  INV_X1 U11993 ( .A(n9439), .ZN(n9440) );
  AND2_X1 U11994 ( .A1(n13456), .A2(n9321), .ZN(n9442) );
  NAND2_X1 U11995 ( .A1(n9443), .A2(n9442), .ZN(n13161) );
  OAI21_X1 U11996 ( .B1(n9443), .B2(n9442), .A(n13161), .ZN(n9444) );
  NOR4_X1 U11997 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9454) );
  NOR4_X1 U11998 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9449) );
  NOR4_X1 U11999 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9448) );
  NOR4_X1 U12000 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9447) );
  NOR4_X1 U12001 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9446) );
  NAND4_X1 U12002 ( .A1(n9449), .A2(n9448), .A3(n9447), .A4(n9446), .ZN(n9450)
         );
  NOR4_X1 U12003 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n9451), .A4(n9450), .ZN(n9453) );
  NOR4_X1 U12004 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9452) );
  NAND3_X1 U12005 ( .A1(n9454), .A2(n9453), .A3(n9452), .ZN(n9471) );
  NAND2_X1 U12006 ( .A1(n9464), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9461) );
  MUX2_X1 U12007 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9461), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9462) );
  NAND2_X1 U12008 ( .A1(n9467), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9463) );
  MUX2_X1 U12009 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9463), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9465) );
  NAND2_X1 U12010 ( .A1(n9482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9466) );
  MUX2_X1 U12011 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9466), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9468) );
  NAND2_X1 U12012 ( .A1(n9468), .A2(n9467), .ZN(n13805) );
  XNOR2_X1 U12013 ( .A(P2_B_REG_SCAN_IN), .B(n13805), .ZN(n9469) );
  NAND2_X1 U12014 ( .A1(n13799), .A2(n9469), .ZN(n9470) );
  AND2_X1 U12015 ( .A1(n9471), .A2(n14873), .ZN(n10102) );
  INV_X1 U12016 ( .A(n10102), .ZN(n10519) );
  INV_X1 U12017 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14879) );
  NAND2_X1 U12018 ( .A1(n14873), .A2(n14879), .ZN(n9473) );
  INV_X1 U12019 ( .A(n9478), .ZN(n13798) );
  NAND2_X1 U12020 ( .A1(n13798), .A2(n13799), .ZN(n9472) );
  NAND2_X1 U12021 ( .A1(n9473), .A2(n9472), .ZN(n14880) );
  INV_X1 U12022 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14876) );
  NAND2_X1 U12023 ( .A1(n14873), .A2(n14876), .ZN(n9475) );
  NAND2_X1 U12024 ( .A1(n13798), .A2(n13805), .ZN(n9474) );
  NAND2_X1 U12025 ( .A1(n9475), .A2(n9474), .ZN(n14877) );
  NOR2_X1 U12026 ( .A1(n14880), .A2(n14877), .ZN(n9476) );
  NAND2_X1 U12027 ( .A1(n10519), .A2(n9476), .ZN(n9503) );
  NOR2_X1 U12028 ( .A1(n13799), .A2(n13805), .ZN(n9477) );
  INV_X1 U12029 ( .A(n9479), .ZN(n9480) );
  OAI21_X1 U12030 ( .B1(n9295), .B2(n9480), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9481) );
  MUX2_X1 U12031 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9481), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n9483) );
  NAND2_X1 U12032 ( .A1(n9483), .A2(n9482), .ZN(n11836) );
  AND2_X1 U12033 ( .A1(n9866), .A2(n11836), .ZN(n9504) );
  INV_X1 U12034 ( .A(n14881), .ZN(n14878) );
  NOR2_X1 U12035 ( .A1(n9503), .A2(n14878), .ZN(n9498) );
  NAND2_X1 U12036 ( .A1(n12331), .A2(n12334), .ZN(n12285) );
  NOR2_X1 U12037 ( .A1(n14889), .A2(n9861), .ZN(n9484) );
  INV_X1 U12038 ( .A(n12331), .ZN(n12295) );
  NAND2_X1 U12039 ( .A1(n9498), .A2(n15201), .ZN(n9488) );
  NAND2_X1 U12040 ( .A1(n13639), .A2(n13330), .ZN(n10463) );
  INV_X1 U12041 ( .A(n10463), .ZN(n9487) );
  INV_X1 U12042 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13169) );
  INV_X1 U12043 ( .A(n13383), .ZN(n9491) );
  NAND2_X1 U12044 ( .A1(n9489), .A2(n13169), .ZN(n9490) );
  NAND2_X1 U12045 ( .A1(n9491), .A2(n9490), .ZN(n13423) );
  INV_X1 U12046 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13427) );
  NAND2_X1 U12047 ( .A1(n12236), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9494) );
  NAND2_X1 U12048 ( .A1(n6647), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9493) );
  OAI211_X1 U12049 ( .C1(n13427), .C2(n12239), .A(n9494), .B(n9493), .ZN(n9495) );
  INV_X1 U12050 ( .A(n9495), .ZN(n9496) );
  INV_X1 U12051 ( .A(n12285), .ZN(n12340) );
  NAND2_X1 U12052 ( .A1(n9498), .A2(n12340), .ZN(n13199) );
  INV_X1 U12053 ( .A(n13199), .ZN(n13251) );
  AND2_X1 U12054 ( .A1(n13251), .A2(n13544), .ZN(n13261) );
  INV_X1 U12055 ( .A(n13472), .ZN(n13435) );
  INV_X1 U12056 ( .A(n9500), .ZN(n9501) );
  NOR2_X1 U12057 ( .A1(n13435), .A2(n13277), .ZN(n9509) );
  INV_X1 U12058 ( .A(n9502), .ZN(n13440) );
  NAND2_X1 U12059 ( .A1(n9503), .A2(n10463), .ZN(n10018) );
  NAND2_X1 U12060 ( .A1(n9861), .A2(n12285), .ZN(n10017) );
  AND2_X1 U12061 ( .A1(n9504), .A2(n10017), .ZN(n9505) );
  NAND2_X1 U12062 ( .A1(n10018), .A2(n9505), .ZN(n9506) );
  OAI22_X1 U12063 ( .A1(n13440), .A2(n13276), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9507), .ZN(n9508) );
  AOI211_X1 U12064 ( .C1(n13379), .C2(n13261), .A(n9509), .B(n9508), .ZN(n9510) );
  INV_X1 U12065 ( .A(n9511), .ZN(n9512) );
  INV_X1 U12066 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14692) );
  INV_X1 U12067 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10664) );
  INV_X1 U12068 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n9537) );
  XNOR2_X1 U12069 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9546) );
  INV_X1 U12070 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n9535) );
  INV_X1 U12071 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10322) );
  XOR2_X1 U12072 ( .A(n9535), .B(n10322), .Z(n9548) );
  INV_X1 U12073 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9531) );
  XNOR2_X1 U12074 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9585) );
  INV_X1 U12075 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n9514) );
  XOR2_X1 U12076 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n9562) );
  NOR2_X1 U12077 ( .A1(n9516), .A2(n9517), .ZN(n9519) );
  NOR2_X1 U12078 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n9554), .ZN(n9518) );
  NOR2_X1 U12079 ( .A1(n9520), .A2(n15131), .ZN(n9522) );
  NOR2_X1 U12080 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14123), .ZN(n9524) );
  NOR2_X1 U12081 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9525), .ZN(n9527) );
  XNOR2_X1 U12082 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n9525), .ZN(n9578) );
  XOR2_X1 U12083 ( .A(n9529), .B(n14138), .Z(n9552) );
  NAND2_X1 U12084 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n9532), .ZN(n9550) );
  NAND2_X1 U12085 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n9550), .ZN(n9533) );
  NAND2_X1 U12086 ( .A1(n9549), .A2(n9533), .ZN(n9547) );
  NAND2_X1 U12087 ( .A1(n9546), .A2(n9545), .ZN(n9536) );
  INV_X1 U12088 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14968) );
  NAND2_X1 U12089 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14968), .ZN(n9538) );
  INV_X1 U12090 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10859) );
  NAND2_X1 U12091 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n10859), .ZN(n9539) );
  INV_X1 U12092 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n11714) );
  INV_X1 U12093 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14560) );
  NAND2_X1 U12094 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14560), .ZN(n9541) );
  INV_X1 U12095 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9540) );
  AOI22_X1 U12096 ( .A1(n9601), .A2(n9541), .B1(P3_ADDR_REG_15__SCAN_IN), .B2(
        n9540), .ZN(n9606) );
  XOR2_X1 U12097 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(P3_ADDR_REG_16__SCAN_IN), 
        .Z(n9542) );
  XNOR2_X1 U12098 ( .A(n9606), .B(n9542), .ZN(n14690) );
  INV_X1 U12099 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14681) );
  XNOR2_X1 U12100 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9544) );
  XNOR2_X1 U12101 ( .A(n9544), .B(n9543), .ZN(n14680) );
  XNOR2_X1 U12102 ( .A(n9546), .B(n9545), .ZN(n9598) );
  XOR2_X1 U12103 ( .A(n9548), .B(n9547), .Z(n9593) );
  INV_X1 U12104 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14946) );
  NAND2_X1 U12105 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  XNOR2_X1 U12106 ( .A(n14946), .B(n9551), .ZN(n9591) );
  XOR2_X1 U12107 ( .A(n9553), .B(n9552), .Z(n9583) );
  NAND2_X1 U12108 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9555), .ZN(n9568) );
  INV_X1 U12109 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15127) );
  XNOR2_X1 U12110 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n9556) );
  XOR2_X1 U12111 ( .A(n9557), .B(n9556), .Z(n9559) );
  OR2_X1 U12112 ( .A1(n15127), .A2(n9559), .ZN(n9561) );
  AOI21_X1 U12113 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n9558), .A(n9557), .ZN(
        n15218) );
  INV_X1 U12114 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15217) );
  NOR2_X1 U12115 ( .A1(n15218), .A2(n15217), .ZN(n15223) );
  XNOR2_X1 U12116 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9559), .ZN(n15222) );
  NAND2_X1 U12117 ( .A1(n15223), .A2(n15222), .ZN(n9560) );
  NAND2_X1 U12118 ( .A1(n9561), .A2(n9560), .ZN(n14545) );
  XNOR2_X1 U12119 ( .A(n6564), .B(n9562), .ZN(n14544) );
  NOR2_X1 U12120 ( .A1(n14545), .A2(n14544), .ZN(n9563) );
  INV_X1 U12121 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14827) );
  NAND2_X1 U12122 ( .A1(n14545), .A2(n14544), .ZN(n14543) );
  OAI21_X1 U12123 ( .B1(n9563), .B2(n14827), .A(n14543), .ZN(n9566) );
  XNOR2_X1 U12124 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n9564), .ZN(n9565) );
  NAND2_X1 U12125 ( .A1(n9568), .A2(n9567), .ZN(n9571) );
  XNOR2_X1 U12126 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9569), .ZN(n9570) );
  NOR2_X1 U12127 ( .A1(n9571), .A2(n9570), .ZN(n9573) );
  XNOR2_X1 U12128 ( .A(n9571), .B(n9570), .ZN(n15216) );
  NOR2_X1 U12129 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15216), .ZN(n9572) );
  NAND2_X1 U12130 ( .A1(n9574), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9577) );
  XOR2_X1 U12131 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), .Z(
        n9575) );
  XNOR2_X1 U12132 ( .A(n9576), .B(n9575), .ZN(n14547) );
  XNOR2_X1 U12133 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9578), .ZN(n15220) );
  NAND2_X1 U12134 ( .A1(n15219), .A2(n15220), .ZN(n9581) );
  NAND2_X1 U12135 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9579), .ZN(n9580) );
  XNOR2_X1 U12136 ( .A(n9585), .B(n9584), .ZN(n9587) );
  NAND2_X1 U12137 ( .A1(n9586), .A2(n9587), .ZN(n9589) );
  NAND2_X1 U12138 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n14550), .ZN(n9588) );
  NAND2_X1 U12139 ( .A1(n9591), .A2(n9590), .ZN(n9592) );
  NAND2_X1 U12140 ( .A1(n9593), .A2(n9594), .ZN(n9596) );
  NAND2_X1 U12141 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n14677), .ZN(n9595) );
  NAND2_X1 U12142 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  XNOR2_X1 U12143 ( .A(n9598), .B(n9597), .ZN(n14678) );
  XOR2_X1 U12144 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n9599) );
  XNOR2_X1 U12145 ( .A(n9600), .B(n9599), .ZN(n14685) );
  XNOR2_X1 U12146 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n9602) );
  XOR2_X1 U12147 ( .A(n9602), .B(n9601), .Z(n9604) );
  INV_X1 U12148 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n9608) );
  INV_X1 U12149 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n9607) );
  OR2_X1 U12150 ( .A1(n9607), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9605) );
  AOI22_X1 U12151 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n9607), .B1(n9606), .B2(
        n9605), .ZN(n9612) );
  XNOR2_X1 U12152 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9612), .ZN(n9613) );
  XOR2_X1 U12153 ( .A(n9608), .B(n9613), .Z(n14554) );
  INV_X1 U12154 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U12155 ( .A1(n14553), .A2(n14554), .ZN(n14552) );
  INV_X1 U12156 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U12157 ( .A1(n9612), .A2(n9611), .ZN(n9615) );
  NAND2_X1 U12158 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n9613), .ZN(n9614) );
  NAND2_X1 U12159 ( .A1(n9615), .A2(n9614), .ZN(n9619) );
  INV_X1 U12160 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12775) );
  NOR2_X1 U12161 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n12775), .ZN(n9616) );
  AOI21_X1 U12162 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n12775), .A(n9616), .ZN(
        n9620) );
  XNOR2_X1 U12163 ( .A(n9619), .B(n9620), .ZN(n9617) );
  NAND2_X1 U12164 ( .A1(n9620), .A2(n9619), .ZN(n9621) );
  OAI21_X1 U12165 ( .B1(n12775), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9621), .ZN(
        n9622) );
  INV_X1 U12166 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9643) );
  OR2_X1 U12167 ( .A1(n12662), .A2(n12696), .ZN(n12831) );
  AND2_X1 U12168 ( .A1(n12663), .A2(n12831), .ZN(n9624) );
  AND2_X1 U12169 ( .A1(n11963), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9626) );
  XNOR2_X1 U12170 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12029) );
  XNOR2_X1 U12171 ( .A(n12031), .B(n12029), .ZN(n13137) );
  NAND2_X1 U12172 ( .A1(n13137), .A2(n12486), .ZN(n9631) );
  NAND2_X1 U12173 ( .A1(n9629), .A2(SI_29_), .ZN(n9630) );
  NAND2_X1 U12174 ( .A1(n9631), .A2(n9630), .ZN(n9641) );
  NAND2_X1 U12175 ( .A1(n9641), .A2(n12837), .ZN(n12668) );
  XNOR2_X1 U12176 ( .A(n9632), .B(n12515), .ZN(n9640) );
  INV_X1 U12177 ( .A(P3_B_REG_SCAN_IN), .ZN(n9633) );
  NOR2_X1 U12178 ( .A1(n6710), .A2(n9633), .ZN(n9634) );
  OR2_X1 U12179 ( .A1(n12958), .A2(n9634), .ZN(n12816) );
  NAND2_X1 U12180 ( .A1(n6449), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U12181 ( .A1(n6447), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U12182 ( .A1(n8931), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9635) );
  OAI22_X1 U12183 ( .A1(n12349), .A2(n12956), .B1(n12816), .B2(n12493), .ZN(
        n9638) );
  INV_X1 U12184 ( .A(n9641), .ZN(n9642) );
  NOR2_X1 U12185 ( .A1(n12822), .A2(n12826), .ZN(n9649) );
  MUX2_X1 U12186 ( .A(n9643), .B(n9649), .S(n15051), .Z(n9648) );
  INV_X1 U12187 ( .A(n12659), .ZN(n9644) );
  AND2_X1 U12188 ( .A1(n12662), .A2(n12857), .ZN(n12520) );
  INV_X1 U12189 ( .A(n9646), .ZN(n12521) );
  XNOR2_X1 U12190 ( .A(n12677), .B(n12515), .ZN(n12829) );
  NAND2_X1 U12191 ( .A1(n9648), .A2(n9647), .ZN(P3_U3488) );
  INV_X1 U12192 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9650) );
  MUX2_X1 U12193 ( .A(n9650), .B(n9649), .S(n15039), .Z(n9652) );
  INV_X1 U12194 ( .A(n15032), .ZN(n14603) );
  NAND2_X1 U12195 ( .A1(n9652), .A2(n9651), .ZN(P3_U3456) );
  NAND2_X1 U12196 ( .A1(n11836), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9653) );
  INV_X2 U12197 ( .A(n9684), .ZN(n13880) );
  INV_X2 U12198 ( .A(n13880), .ZN(n13923) );
  AND2_X2 U12199 ( .A1(n14355), .A2(n13876), .ZN(n9680) );
  OAI22_X1 U12200 ( .A1(n14476), .A2(n13923), .B1(n13964), .B2(n13920), .ZN(
        n13818) );
  OAI22_X1 U12201 ( .A1(n14476), .A2(n13924), .B1(n13964), .B2(n13923), .ZN(
        n9659) );
  XNOR2_X1 U12202 ( .A(n9659), .B(n13921), .ZN(n13819) );
  XOR2_X1 U12203 ( .A(n13818), .B(n13819), .Z(n9769) );
  AND2_X1 U12204 ( .A1(n9680), .A2(n14034), .ZN(n9660) );
  AOI21_X1 U12205 ( .B1(n14792), .B2(n13868), .A(n9660), .ZN(n9723) );
  INV_X2 U12206 ( .A(n9684), .ZN(n13829) );
  AOI22_X1 U12207 ( .A1(n14792), .A2(n6456), .B1(n13829), .B2(n14034), .ZN(
        n9661) );
  XNOR2_X1 U12208 ( .A(n9661), .B(n13921), .ZN(n9722) );
  NAND2_X1 U12209 ( .A1(n9680), .A2(n14038), .ZN(n9663) );
  NAND2_X1 U12210 ( .A1(n14694), .A2(n13880), .ZN(n9662) );
  NAND2_X1 U12211 ( .A1(n9663), .A2(n9662), .ZN(n9692) );
  NAND2_X1 U12212 ( .A1(n14038), .A2(n13880), .ZN(n9665) );
  NAND2_X1 U12213 ( .A1(n6456), .A2(n14694), .ZN(n9664) );
  NAND2_X1 U12214 ( .A1(n9665), .A2(n9664), .ZN(n9666) );
  XNOR2_X1 U12215 ( .A(n9666), .B(n13921), .ZN(n9691) );
  NAND2_X1 U12216 ( .A1(n6651), .A2(n13880), .ZN(n9670) );
  AOI21_X1 U12217 ( .B1(n10718), .B2(n6456), .A(n9668), .ZN(n9669) );
  NAND2_X1 U12218 ( .A1(n9670), .A2(n9669), .ZN(n10121) );
  NAND2_X1 U12219 ( .A1(n9680), .A2(n6651), .ZN(n9674) );
  OAI21_X1 U12220 ( .B1(n13865), .B2(n10121), .A(n10120), .ZN(n10412) );
  NAND2_X1 U12221 ( .A1(n9679), .A2(n9675), .ZN(n9677) );
  INV_X1 U12222 ( .A(n11449), .ZN(n14738) );
  NAND2_X1 U12223 ( .A1(n14738), .A2(n6456), .ZN(n9676) );
  NAND2_X1 U12224 ( .A1(n9677), .A2(n9676), .ZN(n9678) );
  XNOR2_X1 U12225 ( .A(n9681), .B(n9682), .ZN(n10411) );
  INV_X1 U12226 ( .A(n9681), .ZN(n9683) );
  AOI22_X1 U12227 ( .A1(n9680), .A2(n14740), .B1(n13829), .B2(n10727), .ZN(
        n9688) );
  NAND2_X1 U12228 ( .A1(n14740), .A2(n13880), .ZN(n9686) );
  NAND2_X1 U12229 ( .A1(n6456), .A2(n10727), .ZN(n9685) );
  NAND2_X1 U12230 ( .A1(n9686), .A2(n9685), .ZN(n9687) );
  XOR2_X1 U12231 ( .A(n9688), .B(n9690), .Z(n10487) );
  INV_X1 U12232 ( .A(n9688), .ZN(n9689) );
  OAI22_X1 U12233 ( .A1(n10488), .A2(n10487), .B1(n9690), .B2(n9689), .ZN(
        n14700) );
  XNOR2_X1 U12234 ( .A(n9691), .B(n9692), .ZN(n14701) );
  AOI22_X1 U12235 ( .A1(n9693), .A2(n9680), .B1(n13829), .B2(n11143), .ZN(
        n9695) );
  OAI22_X1 U12236 ( .A1(n11273), .A2(n13923), .B1(n11132), .B2(n13924), .ZN(
        n9694) );
  XNOR2_X1 U12237 ( .A(n9694), .B(n13921), .ZN(n10965) );
  INV_X1 U12238 ( .A(n11268), .ZN(n14761) );
  OAI22_X1 U12239 ( .A1(n14761), .A2(n13924), .B1(n10968), .B2(n13923), .ZN(
        n9696) );
  XOR2_X1 U12240 ( .A(n13921), .B(n9696), .Z(n10954) );
  INV_X1 U12241 ( .A(n10954), .ZN(n9699) );
  NAND2_X1 U12242 ( .A1(n11268), .A2(n13880), .ZN(n9698) );
  NAND2_X1 U12243 ( .A1(n9680), .A2(n14037), .ZN(n9697) );
  NAND2_X1 U12244 ( .A1(n9698), .A2(n9697), .ZN(n9700) );
  NOR2_X1 U12245 ( .A1(n9699), .A2(n9700), .ZN(n9701) );
  INV_X1 U12246 ( .A(n9700), .ZN(n10953) );
  OAI22_X1 U12247 ( .A1(n11175), .A2(n13923), .B1(n11274), .B2(n13920), .ZN(
        n9706) );
  NAND2_X1 U12248 ( .A1(n14765), .A2(n6456), .ZN(n9703) );
  NAND2_X1 U12249 ( .A1(n14036), .A2(n13880), .ZN(n9702) );
  NAND2_X1 U12250 ( .A1(n9703), .A2(n9702), .ZN(n9704) );
  XNOR2_X1 U12251 ( .A(n9704), .B(n13921), .ZN(n9705) );
  XOR2_X1 U12252 ( .A(n9706), .B(n9705), .Z(n11069) );
  AOI22_X1 U12253 ( .A1(n11256), .A2(n6456), .B1(n13829), .B2(n14035), .ZN(
        n9707) );
  XNOR2_X1 U12254 ( .A(n9707), .B(n13921), .ZN(n9709) );
  AND2_X1 U12255 ( .A1(n9680), .A2(n14035), .ZN(n9708) );
  AOI21_X1 U12256 ( .B1(n11256), .B2(n13829), .A(n9708), .ZN(n9710) );
  XNOR2_X1 U12257 ( .A(n9709), .B(n9710), .ZN(n11187) );
  NAND2_X1 U12258 ( .A1(n11431), .A2(n6456), .ZN(n9712) );
  OR2_X1 U12259 ( .A1(n11627), .A2(n13923), .ZN(n9711) );
  NAND2_X1 U12260 ( .A1(n9712), .A2(n9711), .ZN(n9713) );
  XNOR2_X1 U12261 ( .A(n9713), .B(n13865), .ZN(n9716) );
  NOR2_X1 U12262 ( .A1(n11627), .A2(n13920), .ZN(n9714) );
  AOI21_X1 U12263 ( .B1(n11431), .B2(n13829), .A(n9714), .ZN(n9715) );
  NAND2_X1 U12264 ( .A1(n9716), .A2(n9715), .ZN(n9717) );
  OAI21_X1 U12265 ( .B1(n9716), .B2(n9715), .A(n9717), .ZN(n11425) );
  OAI22_X1 U12266 ( .A1(n11621), .A2(n13923), .B1(n11656), .B2(n13920), .ZN(
        n9720) );
  XNOR2_X1 U12267 ( .A(n9719), .B(n9720), .ZN(n11623) );
  OAI22_X1 U12268 ( .A1(n11621), .A2(n13924), .B1(n11656), .B2(n13923), .ZN(
        n9718) );
  XOR2_X1 U12269 ( .A(n13921), .B(n9718), .Z(n11624) );
  NAND2_X1 U12270 ( .A1(n11623), .A2(n11624), .ZN(n11622) );
  XOR2_X1 U12271 ( .A(n9723), .B(n9722), .Z(n11653) );
  INV_X1 U12272 ( .A(n9719), .ZN(n9721) );
  OR2_X1 U12273 ( .A1(n9721), .A2(n9720), .ZN(n11650) );
  OAI22_X1 U12274 ( .A1(n14669), .A2(n13924), .B1(n11872), .B2(n13923), .ZN(
        n9724) );
  XNOR2_X1 U12275 ( .A(n9724), .B(n13921), .ZN(n9726) );
  OAI22_X1 U12276 ( .A1(n14669), .A2(n13923), .B1(n11872), .B2(n13920), .ZN(
        n9725) );
  XNOR2_X1 U12277 ( .A(n9726), .B(n9725), .ZN(n11761) );
  NOR2_X1 U12278 ( .A1(n9726), .A2(n9725), .ZN(n11868) );
  NAND2_X1 U12279 ( .A1(n11889), .A2(n6456), .ZN(n9728) );
  NAND2_X1 U12280 ( .A1(n14032), .A2(n13880), .ZN(n9727) );
  NAND2_X1 U12281 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  XNOR2_X1 U12282 ( .A(n9729), .B(n13865), .ZN(n9731) );
  AND2_X1 U12283 ( .A1(n9680), .A2(n14032), .ZN(n9730) );
  AOI21_X1 U12284 ( .B1(n11889), .B2(n13829), .A(n9730), .ZN(n9732) );
  XNOR2_X1 U12285 ( .A(n9731), .B(n9732), .ZN(n11867) );
  INV_X1 U12286 ( .A(n9731), .ZN(n9734) );
  INV_X1 U12287 ( .A(n9732), .ZN(n9733) );
  AND2_X1 U12288 ( .A1(n9680), .A2(n14031), .ZN(n9735) );
  AOI21_X1 U12289 ( .B1(n11951), .B2(n13829), .A(n9735), .ZN(n9739) );
  OAI22_X1 U12290 ( .A1(n11681), .A2(n13924), .B1(n11873), .B2(n13923), .ZN(
        n9736) );
  XNOR2_X1 U12291 ( .A(n9736), .B(n13921), .ZN(n9737) );
  XOR2_X1 U12292 ( .A(n9739), .B(n9737), .Z(n11944) );
  INV_X1 U12293 ( .A(n9737), .ZN(n9738) );
  OAI22_X1 U12294 ( .A1(n11945), .A2(n11944), .B1(n9739), .B2(n9738), .ZN(
        n14641) );
  NAND2_X1 U12295 ( .A1(n14643), .A2(n6456), .ZN(n9741) );
  NAND2_X1 U12296 ( .A1(n14030), .A2(n13880), .ZN(n9740) );
  NAND2_X1 U12297 ( .A1(n9741), .A2(n9740), .ZN(n9742) );
  XNOR2_X1 U12298 ( .A(n9742), .B(n13865), .ZN(n9745) );
  AND2_X1 U12299 ( .A1(n9680), .A2(n14030), .ZN(n9743) );
  AOI21_X1 U12300 ( .B1(n14643), .B2(n13829), .A(n9743), .ZN(n9744) );
  NAND2_X1 U12301 ( .A1(n9745), .A2(n9744), .ZN(n9746) );
  OAI21_X1 U12302 ( .B1(n9745), .B2(n9744), .A(n9746), .ZN(n14640) );
  NAND2_X1 U12303 ( .A1(n14663), .A2(n6456), .ZN(n9748) );
  NAND2_X1 U12304 ( .A1(n14029), .A2(n13880), .ZN(n9747) );
  NAND2_X1 U12305 ( .A1(n9748), .A2(n9747), .ZN(n9749) );
  XNOR2_X1 U12306 ( .A(n9749), .B(n13865), .ZN(n9750) );
  AOI22_X1 U12307 ( .A1(n14663), .A2(n13868), .B1(n9680), .B2(n14029), .ZN(
        n14011) );
  NAND2_X1 U12308 ( .A1(n14654), .A2(n6456), .ZN(n9752) );
  NAND2_X1 U12309 ( .A1(n14482), .A2(n13868), .ZN(n9751) );
  NAND2_X1 U12310 ( .A1(n9752), .A2(n9751), .ZN(n9753) );
  XNOR2_X1 U12311 ( .A(n9753), .B(n13865), .ZN(n9756) );
  AND2_X1 U12312 ( .A1(n9680), .A2(n14482), .ZN(n9754) );
  AOI21_X1 U12313 ( .B1(n14654), .B2(n13829), .A(n9754), .ZN(n9755) );
  NAND2_X1 U12314 ( .A1(n9756), .A2(n9755), .ZN(n13958) );
  OAI21_X1 U12315 ( .B1(n9756), .B2(n9755), .A(n13958), .ZN(n14651) );
  NAND2_X1 U12316 ( .A1(n14385), .A2(n6456), .ZN(n9760) );
  OR2_X1 U12317 ( .A1(n14350), .A2(n13923), .ZN(n9759) );
  NAND2_X1 U12318 ( .A1(n9760), .A2(n9759), .ZN(n9761) );
  XNOR2_X1 U12319 ( .A(n9761), .B(n13865), .ZN(n9764) );
  NOR2_X1 U12320 ( .A1(n14350), .A2(n13920), .ZN(n9762) );
  AOI21_X1 U12321 ( .B1(n14385), .B2(n13880), .A(n9762), .ZN(n9763) );
  NAND2_X1 U12322 ( .A1(n9764), .A2(n9763), .ZN(n9767) );
  OR2_X1 U12323 ( .A1(n9764), .A2(n9763), .ZN(n9765) );
  AND2_X1 U12324 ( .A1(n9767), .A2(n9765), .ZN(n13959) );
  OAI21_X1 U12325 ( .B1(n9769), .B2(n9768), .A(n13909), .ZN(n9793) );
  NOR2_X1 U12326 ( .A1(n14793), .A2(n9772), .ZN(n9792) );
  INV_X1 U12327 ( .A(n9775), .ZN(n14531) );
  NAND3_X1 U12328 ( .A1(n14535), .A2(P1_B_REG_SCAN_IN), .A3(n14531), .ZN(n9773) );
  OR2_X1 U12329 ( .A1(n9789), .A2(n9775), .ZN(n9904) );
  OAI21_X1 U12330 ( .B1(n10714), .B2(P1_D_REG_1__SCAN_IN), .A(n9904), .ZN(
        n10341) );
  INV_X1 U12331 ( .A(n10343), .ZN(n9776) );
  NOR2_X1 U12332 ( .A1(n10341), .A2(n9776), .ZN(n9801) );
  INV_X1 U12333 ( .A(n10714), .ZN(n9788) );
  NOR4_X1 U12334 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9780) );
  NOR4_X1 U12335 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9779) );
  NOR4_X1 U12336 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9778) );
  NOR4_X1 U12337 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9777) );
  NAND4_X1 U12338 ( .A1(n9780), .A2(n9779), .A3(n9778), .A4(n9777), .ZN(n9786)
         );
  NOR2_X1 U12339 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .ZN(
        n9784) );
  NOR4_X1 U12340 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9783) );
  NOR4_X1 U12341 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9782) );
  NOR4_X1 U12342 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n9781) );
  NAND4_X1 U12343 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(n9785)
         );
  NOR2_X1 U12344 ( .A1(n9786), .A2(n9785), .ZN(n10713) );
  NAND2_X1 U12345 ( .A1(n10713), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U12346 ( .A1(n9788), .A2(n9787), .ZN(n9790) );
  INV_X1 U12347 ( .A(n9789), .ZN(n14527) );
  NAND2_X1 U12348 ( .A1(n14535), .A2(n14527), .ZN(n10712) );
  NAND2_X1 U12349 ( .A1(n9790), .A2(n10712), .ZN(n10345) );
  INV_X1 U12350 ( .A(n10345), .ZN(n9802) );
  NAND2_X1 U12351 ( .A1(n9801), .A2(n9802), .ZN(n9795) );
  INV_X1 U12352 ( .A(n9795), .ZN(n9791) );
  AND2_X1 U12353 ( .A1(n9793), .A2(n14655), .ZN(n9806) );
  AND2_X1 U12354 ( .A1(n11196), .A2(n10343), .ZN(n9794) );
  NAND2_X1 U12355 ( .A1(n9795), .A2(n14374), .ZN(n14697) );
  NOR2_X1 U12356 ( .A1(n14476), .A2(n14015), .ZN(n9805) );
  NAND2_X1 U12357 ( .A1(n9770), .A2(n11196), .ZN(n10344) );
  OAI21_X1 U12358 ( .B1(n10345), .B2(n10341), .A(n10344), .ZN(n9798) );
  NAND4_X1 U12359 ( .A1(n9798), .A2(n10342), .A3(n9797), .A4(n9796), .ZN(n9799) );
  INV_X1 U12360 ( .A(n9800), .ZN(n14358) );
  NAND2_X1 U12361 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11847)
         );
  OAI21_X1 U12362 ( .B1(n14707), .B2(n14358), .A(n11847), .ZN(n9804) );
  INV_X1 U12363 ( .A(n14361), .ZN(n14475) );
  AND2_X1 U12364 ( .A1(n9801), .A2(n10342), .ZN(n10795) );
  NOR2_X2 U12365 ( .A1(n10334), .A2(n10031), .ZN(n14739) );
  NAND2_X1 U12366 ( .A1(n14704), .A2(n14739), .ZN(n13975) );
  NAND2_X1 U12367 ( .A1(n14704), .A2(n14483), .ZN(n13974) );
  OAI22_X1 U12368 ( .A1(n14475), .A2(n13975), .B1(n14350), .B2(n13974), .ZN(
        n9803) );
  INV_X2 U12369 ( .A(n10409), .ZN(n14528) );
  INV_X2 U12370 ( .A(n11861), .ZN(n14534) );
  OAI222_X1 U12371 ( .A1(n14528), .A2(n8100), .B1(n14534), .B2(n9903), .C1(
        P1_U3086), .C2(n10042), .ZN(P1_U3354) );
  OAI222_X1 U12372 ( .A1(n14528), .A2(n9807), .B1(n14534), .B2(n9844), .C1(
        P1_U3086), .C2(n14057), .ZN(P1_U3353) );
  NOR2_X1 U12373 ( .A1(n9842), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13134) );
  INV_X1 U12374 ( .A(n9808), .ZN(n9810) );
  NAND2_X2 U12375 ( .A1(n9842), .A2(P3_U3151), .ZN(n13142) );
  INV_X1 U12376 ( .A(SI_5_), .ZN(n9809) );
  OAI222_X1 U12377 ( .A1(n10243), .A2(P3_U3151), .B1(n13140), .B2(n9810), .C1(
        n13142), .C2(n9809), .ZN(P3_U3290) );
  INV_X1 U12378 ( .A(n14074), .ZN(n9812) );
  OAI222_X1 U12379 ( .A1(P1_U3086), .A2(n9812), .B1(n14534), .B2(n9896), .C1(
        n9811), .C2(n14528), .ZN(P1_U3352) );
  OAI222_X1 U12380 ( .A1(n13140), .A2(n9814), .B1(n13142), .B2(n9813), .C1(
        n10908), .C2(P3_U3151), .ZN(P3_U3287) );
  OAI222_X1 U12381 ( .A1(n10552), .A2(P3_U3151), .B1(n13140), .B2(n9816), .C1(
        n9815), .C2(n13142), .ZN(P3_U3289) );
  OAI222_X1 U12382 ( .A1(n10142), .A2(P3_U3151), .B1(n13140), .B2(n9818), .C1(
        n9817), .C2(n13142), .ZN(P3_U3295) );
  INV_X1 U12383 ( .A(n9819), .ZN(n9821) );
  INV_X1 U12384 ( .A(SI_4_), .ZN(n9820) );
  OAI222_X1 U12385 ( .A1(n13140), .A2(n9821), .B1(n13142), .B2(n9820), .C1(
        n10240), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12386 ( .A(n9822), .ZN(n9824) );
  INV_X1 U12387 ( .A(SI_7_), .ZN(n9823) );
  OAI222_X1 U12388 ( .A1(n13140), .A2(n9824), .B1(n13142), .B2(n9823), .C1(
        P3_U3151), .C2(n14932), .ZN(P3_U3288) );
  OAI222_X1 U12389 ( .A1(P3_U3151), .A2(n10145), .B1(n13142), .B2(n6719), .C1(
        n13140), .C2(n9825), .ZN(P3_U3294) );
  INV_X1 U12390 ( .A(n9826), .ZN(n9828) );
  INV_X1 U12391 ( .A(SI_2_), .ZN(n9827) );
  OAI222_X1 U12392 ( .A1(n13140), .A2(n9828), .B1(n13142), .B2(n9827), .C1(
        n6453), .C2(P3_U3151), .ZN(P3_U3293) );
  INV_X1 U12393 ( .A(n9829), .ZN(n9831) );
  INV_X1 U12394 ( .A(SI_3_), .ZN(n9830) );
  OAI222_X1 U12395 ( .A1(n10185), .A2(P3_U3151), .B1(n13140), .B2(n9831), .C1(
        n9830), .C2(n13142), .ZN(P3_U3292) );
  OAI222_X1 U12396 ( .A1(n13140), .A2(n9833), .B1(n13142), .B2(n9832), .C1(
        n10898), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12397 ( .A1(n13140), .A2(n9835), .B1(n13142), .B2(n9834), .C1(
        n14944), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12398 ( .A(n13127), .ZN(n9838) );
  INV_X1 U12399 ( .A(n10348), .ZN(n9836) );
  NAND2_X1 U12400 ( .A1(n9836), .A2(n9838), .ZN(n9837) );
  OAI21_X1 U12401 ( .B1(n15111), .B2(n9838), .A(n9837), .ZN(P3_U3377) );
  INV_X1 U12402 ( .A(n14093), .ZN(n9841) );
  INV_X1 U12403 ( .A(n9839), .ZN(n9845) );
  OAI222_X1 U12404 ( .A1(P1_U3086), .A2(n9841), .B1(n14534), .B2(n9845), .C1(
        n9840), .C2(n14528), .ZN(P1_U3351) );
  NAND2_X2 U12405 ( .A1(n9842), .A2(P2_U3088), .ZN(n13800) );
  NAND2_X2 U12406 ( .A1(n9014), .A2(P2_U3088), .ZN(n13803) );
  OAI222_X1 U12407 ( .A1(P2_U3088), .A2(n14819), .B1(n13800), .B2(n9844), .C1(
        n9843), .C2(n13803), .ZN(P2_U3325) );
  INV_X1 U12408 ( .A(n9966), .ZN(n9976) );
  OAI222_X1 U12409 ( .A1(P2_U3088), .A2(n9976), .B1(n13800), .B2(n9845), .C1(
        n10162), .C2(n13803), .ZN(P2_U3323) );
  INV_X1 U12410 ( .A(n11413), .ZN(n9846) );
  OAI222_X1 U12411 ( .A1(n13140), .A2(n9848), .B1(n13142), .B2(n9847), .C1(
        n9846), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12412 ( .A(n14109), .ZN(n9851) );
  INV_X1 U12413 ( .A(n9849), .ZN(n9859) );
  OAI222_X1 U12414 ( .A1(n9851), .A2(P1_U3086), .B1(n14534), .B2(n9859), .C1(
        n9850), .C2(n14528), .ZN(P1_U3350) );
  INV_X1 U12415 ( .A(n14125), .ZN(n9853) );
  OAI222_X1 U12416 ( .A1(P1_U3086), .A2(n9853), .B1(n14534), .B2(n9898), .C1(
        n9852), .C2(n14528), .ZN(P1_U3349) );
  INV_X1 U12417 ( .A(n11416), .ZN(n11703) );
  OAI222_X1 U12418 ( .A1(n13140), .A2(n9855), .B1(n11703), .B2(P3_U3151), .C1(
        n9854), .C2(n13142), .ZN(P3_U3283) );
  NAND2_X1 U12419 ( .A1(n10343), .A2(n10714), .ZN(n14736) );
  INV_X1 U12420 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9858) );
  INV_X1 U12421 ( .A(n10712), .ZN(n9856) );
  AOI22_X1 U12422 ( .A1(n14736), .A2(n9858), .B1(n9857), .B2(n9856), .ZN(
        P1_U3445) );
  INV_X1 U12423 ( .A(n9973), .ZN(n9998) );
  OAI222_X1 U12424 ( .A1(n13803), .A2(n9860), .B1(n13800), .B2(n9859), .C1(
        P2_U3088), .C2(n9998), .ZN(P2_U3322) );
  INV_X1 U12425 ( .A(n11836), .ZN(n9865) );
  NAND2_X1 U12426 ( .A1(n9861), .A2(n11836), .ZN(n9863) );
  NAND2_X1 U12427 ( .A1(n9863), .A2(n9862), .ZN(n9864) );
  OAI21_X1 U12428 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(n9886) );
  NAND2_X1 U12429 ( .A1(n9886), .A2(n9500), .ZN(n14836) );
  OR2_X1 U12430 ( .A1(n14836), .A2(P2_U3088), .ZN(n14820) );
  INV_X1 U12431 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9867) );
  MUX2_X1 U12432 ( .A(n9867), .B(P2_REG1_REG_2__SCAN_IN), .S(n14819), .Z(
        n14823) );
  INV_X1 U12433 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9953) );
  MUX2_X1 U12434 ( .A(n9953), .B(P2_REG1_REG_1__SCAN_IN), .S(n9952), .Z(n9869)
         );
  AND2_X1 U12435 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9868) );
  NAND2_X1 U12436 ( .A1(n9869), .A2(n9868), .ZN(n9957) );
  OAI21_X1 U12437 ( .B1(n9953), .B2(n9952), .A(n9957), .ZN(n14824) );
  NAND2_X1 U12438 ( .A1(n14823), .A2(n14824), .ZN(n14822) );
  INV_X1 U12439 ( .A(n14819), .ZN(n9870) );
  NAND2_X1 U12440 ( .A1(n9870), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9941) );
  INV_X1 U12441 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n15178) );
  MUX2_X1 U12442 ( .A(n15178), .B(P2_REG1_REG_3__SCAN_IN), .S(n9883), .Z(n9942) );
  AOI21_X1 U12443 ( .B1(n14822), .B2(n9941), .A(n9942), .ZN(n9944) );
  INV_X1 U12444 ( .A(n9883), .ZN(n9948) );
  NOR2_X1 U12445 ( .A1(n9948), .A2(n15178), .ZN(n9876) );
  INV_X1 U12446 ( .A(n9876), .ZN(n9872) );
  MUX2_X1 U12447 ( .A(n9874), .B(P2_REG1_REG_4__SCAN_IN), .S(n9966), .Z(n9871)
         );
  NAND2_X1 U12448 ( .A1(n9872), .A2(n9871), .ZN(n9877) );
  OR2_X1 U12449 ( .A1(n9500), .A2(P2_U3088), .ZN(n13792) );
  INV_X1 U12450 ( .A(n13795), .ZN(n12341) );
  NOR2_X1 U12451 ( .A1(n13792), .A2(n12341), .ZN(n9873) );
  INV_X1 U12452 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9874) );
  MUX2_X1 U12453 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9874), .S(n9966), .Z(n9875)
         );
  OAI21_X1 U12454 ( .B1(n9944), .B2(n9876), .A(n9875), .ZN(n9969) );
  OAI211_X1 U12455 ( .C1(n9944), .C2(n9877), .A(n14868), .B(n9969), .ZN(n9878)
         );
  OAI21_X1 U12456 ( .B1(n7124), .B2(n14857), .A(n9878), .ZN(n9892) );
  INV_X1 U12457 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9879) );
  MUX2_X1 U12458 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9879), .S(n9966), .Z(n9888)
         );
  INV_X1 U12459 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9882) );
  MUX2_X1 U12460 ( .A(n9882), .B(P2_REG2_REG_2__SCAN_IN), .S(n14819), .Z(
        n14816) );
  INV_X1 U12461 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9880) );
  MUX2_X1 U12462 ( .A(n9880), .B(P2_REG2_REG_1__SCAN_IN), .S(n9952), .Z(n9951)
         );
  AND2_X1 U12463 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9950) );
  NAND2_X1 U12464 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  NAND2_X1 U12465 ( .A1(n9962), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U12466 ( .A1(n9949), .A2(n9881), .ZN(n14815) );
  NAND2_X1 U12467 ( .A1(n14816), .A2(n14815), .ZN(n14814) );
  OAI21_X1 U12468 ( .B1(n9882), .B2(n14819), .A(n14814), .ZN(n9937) );
  MUX2_X1 U12469 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9884), .S(n9883), .Z(n9938)
         );
  NOR2_X1 U12470 ( .A1(n13792), .A2(n13795), .ZN(n9885) );
  NAND2_X1 U12471 ( .A1(n9887), .A2(n9888), .ZN(n9975) );
  OAI211_X1 U12472 ( .C1(n9888), .C2(n9887), .A(n14865), .B(n9975), .ZN(n9889)
         );
  INV_X1 U12473 ( .A(n9889), .ZN(n9891) );
  AND2_X1 U12474 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9890) );
  NOR3_X1 U12475 ( .A1(n9892), .A2(n9891), .A3(n9890), .ZN(n9893) );
  OAI21_X1 U12476 ( .B1(n9976), .B2(n14820), .A(n9893), .ZN(P2_U3218) );
  INV_X1 U12477 ( .A(n13803), .ZN(n13790) );
  NAND2_X1 U12478 ( .A1(n13790), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U12479 ( .A1(n10002), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14835) );
  OAI211_X1 U12480 ( .C1(n9900), .C2(n13800), .A(n9894), .B(n14835), .ZN(
        P2_U3320) );
  OAI222_X1 U12481 ( .A1(P2_U3088), .A2(n9948), .B1(n13800), .B2(n9896), .C1(
        n9895), .C2(n13803), .ZN(P2_U3324) );
  INV_X1 U12482 ( .A(n9999), .ZN(n13298) );
  OAI222_X1 U12483 ( .A1(P2_U3088), .A2(n13298), .B1(n13800), .B2(n9898), .C1(
        n9897), .C2(n13803), .ZN(P2_U3321) );
  INV_X1 U12484 ( .A(n10306), .ZN(n9901) );
  OAI222_X1 U12485 ( .A1(P1_U3086), .A2(n9901), .B1(n14534), .B2(n9900), .C1(
        n9899), .C2(n14528), .ZN(P1_U3348) );
  OAI222_X1 U12486 ( .A1(P2_U3088), .A2(n9952), .B1(n13800), .B2(n9903), .C1(
        n9902), .C2(n13803), .ZN(P2_U3326) );
  INV_X1 U12487 ( .A(n14736), .ZN(n14735) );
  OAI22_X1 U12488 ( .A1(n14735), .A2(P1_D_REG_1__SCAN_IN), .B1(n9905), .B2(
        n9904), .ZN(n9906) );
  INV_X1 U12489 ( .A(n9906), .ZN(P1_U3446) );
  NOR2_X1 U12490 ( .A1(n13127), .A2(n9907), .ZN(n9910) );
  CLKBUF_X1 U12491 ( .A(n9910), .Z(n9934) );
  INV_X1 U12492 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U12493 ( .A1(n9934), .A2(n9908), .ZN(P3_U3254) );
  INV_X1 U12494 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9909) );
  NOR2_X1 U12495 ( .A1(n9934), .A2(n9909), .ZN(P3_U3263) );
  INV_X1 U12496 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9911) );
  NOR2_X1 U12497 ( .A1(n9934), .A2(n9911), .ZN(P3_U3262) );
  INV_X1 U12498 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U12499 ( .A1(n9910), .A2(n9912), .ZN(P3_U3243) );
  INV_X1 U12500 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9913) );
  NOR2_X1 U12501 ( .A1(n9910), .A2(n9913), .ZN(P3_U3240) );
  INV_X1 U12502 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n15186) );
  NOR2_X1 U12503 ( .A1(n9910), .A2(n15186), .ZN(P3_U3241) );
  INV_X1 U12504 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9914) );
  NOR2_X1 U12505 ( .A1(n9934), .A2(n9914), .ZN(P3_U3255) );
  INV_X1 U12506 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9915) );
  NOR2_X1 U12507 ( .A1(n9910), .A2(n9915), .ZN(P3_U3244) );
  INV_X1 U12508 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9916) );
  NOR2_X1 U12509 ( .A1(n9934), .A2(n9916), .ZN(P3_U3261) );
  INV_X1 U12510 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U12511 ( .A1(n9910), .A2(n9917), .ZN(P3_U3260) );
  INV_X1 U12512 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U12513 ( .A1(n9934), .A2(n9918), .ZN(P3_U3259) );
  INV_X1 U12514 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9919) );
  NOR2_X1 U12515 ( .A1(n9910), .A2(n9919), .ZN(P3_U3258) );
  INV_X1 U12516 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U12517 ( .A1(n9934), .A2(n9920), .ZN(P3_U3257) );
  INV_X1 U12518 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9921) );
  NOR2_X1 U12519 ( .A1(n9934), .A2(n9921), .ZN(P3_U3256) );
  INV_X1 U12520 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9922) );
  NOR2_X1 U12521 ( .A1(n9934), .A2(n9922), .ZN(P3_U3247) );
  INV_X1 U12522 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9923) );
  NOR2_X1 U12523 ( .A1(n9910), .A2(n9923), .ZN(P3_U3236) );
  INV_X1 U12524 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9924) );
  NOR2_X1 U12525 ( .A1(n9934), .A2(n9924), .ZN(P3_U3253) );
  INV_X1 U12526 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U12527 ( .A1(n9934), .A2(n9925), .ZN(P3_U3252) );
  INV_X1 U12528 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9926) );
  NOR2_X1 U12529 ( .A1(n9934), .A2(n9926), .ZN(P3_U3251) );
  INV_X1 U12530 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n15129) );
  NOR2_X1 U12531 ( .A1(n9910), .A2(n15129), .ZN(P3_U3245) );
  INV_X1 U12532 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n15124) );
  NOR2_X1 U12533 ( .A1(n9934), .A2(n15124), .ZN(P3_U3249) );
  INV_X1 U12534 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9927) );
  NOR2_X1 U12535 ( .A1(n9934), .A2(n9927), .ZN(P3_U3248) );
  INV_X1 U12536 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U12537 ( .A1(n9910), .A2(n9928), .ZN(P3_U3239) );
  INV_X1 U12538 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9929) );
  NOR2_X1 U12539 ( .A1(n9934), .A2(n9929), .ZN(P3_U3246) );
  INV_X1 U12540 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9930) );
  NOR2_X1 U12541 ( .A1(n9910), .A2(n9930), .ZN(P3_U3237) );
  INV_X1 U12542 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9931) );
  NOR2_X1 U12543 ( .A1(n9910), .A2(n9931), .ZN(P3_U3238) );
  INV_X1 U12544 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U12545 ( .A1(n9934), .A2(n9932), .ZN(P3_U3235) );
  INV_X1 U12546 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9933) );
  NOR2_X1 U12547 ( .A1(n9934), .A2(n9933), .ZN(P3_U3242) );
  INV_X1 U12548 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n15172) );
  NOR2_X1 U12549 ( .A1(n9934), .A2(n15172), .ZN(P3_U3250) );
  INV_X1 U12550 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9935) );
  NOR2_X1 U12551 ( .A1(n9934), .A2(n9935), .ZN(P3_U3234) );
  INV_X1 U12552 ( .A(n14857), .ZN(n14859) );
  OAI211_X1 U12553 ( .C1(n9938), .C2(n9937), .A(n14865), .B(n9936), .ZN(n9940)
         );
  INV_X1 U12554 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10377) );
  OR2_X1 U12555 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10377), .ZN(n9939) );
  NAND2_X1 U12556 ( .A1(n9940), .A2(n9939), .ZN(n9946) );
  INV_X1 U12557 ( .A(n14868), .ZN(n13328) );
  AND3_X1 U12558 ( .A1(n9942), .A2(n14822), .A3(n9941), .ZN(n9943) );
  NOR3_X1 U12559 ( .A1(n13328), .A2(n9944), .A3(n9943), .ZN(n9945) );
  AOI211_X1 U12560 ( .C1(n14859), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n9946), .B(
        n9945), .ZN(n9947) );
  OAI21_X1 U12561 ( .B1(n9948), .B2(n14820), .A(n9947), .ZN(P2_U3217) );
  INV_X1 U12562 ( .A(n14820), .ZN(n14863) );
  INV_X1 U12563 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10705) );
  OAI211_X1 U12564 ( .C1(n9951), .C2(n9950), .A(n14865), .B(n9949), .ZN(n9959)
         );
  INV_X1 U12565 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14916) );
  INV_X1 U12566 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9955) );
  MUX2_X1 U12567 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9953), .S(n9952), .Z(n9954)
         );
  OAI21_X1 U12568 ( .B1(n14916), .B2(n9955), .A(n9954), .ZN(n9956) );
  NAND3_X1 U12569 ( .A1(n14868), .A2(n9957), .A3(n9956), .ZN(n9958) );
  OAI211_X1 U12570 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10705), .A(n9959), .B(
        n9958), .ZN(n9961) );
  NOR2_X1 U12571 ( .A1(n15127), .A2(n14857), .ZN(n9960) );
  AOI211_X1 U12572 ( .C1(n14863), .C2(n9962), .A(n9961), .B(n9960), .ZN(n9963)
         );
  INV_X1 U12573 ( .A(n9963), .ZN(P2_U3215) );
  INV_X1 U12574 ( .A(n11695), .ZN(n14965) );
  OAI222_X1 U12575 ( .A1(n13140), .A2(n9965), .B1(n14965), .B2(P3_U3151), .C1(
        n9964), .C2(n13142), .ZN(P3_U3282) );
  NAND2_X1 U12576 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10366) );
  INV_X1 U12577 ( .A(n10366), .ZN(n9972) );
  NAND2_X1 U12578 ( .A1(n9966), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9968) );
  INV_X1 U12579 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9997) );
  MUX2_X1 U12580 ( .A(n9997), .B(P2_REG1_REG_5__SCAN_IN), .S(n9973), .Z(n9967)
         );
  AOI21_X1 U12581 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n13306) );
  AND3_X1 U12582 ( .A1(n9969), .A2(n9968), .A3(n9967), .ZN(n9970) );
  NOR3_X1 U12583 ( .A1(n13328), .A2(n13306), .A3(n9970), .ZN(n9971) );
  AOI211_X1 U12584 ( .C1(n14859), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n9972), .B(
        n9971), .ZN(n9980) );
  INV_X1 U12585 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9974) );
  MUX2_X1 U12586 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9974), .S(n9973), .Z(n9978)
         );
  OAI21_X1 U12587 ( .B1(n9976), .B2(n9879), .A(n9975), .ZN(n9977) );
  NAND2_X1 U12588 ( .A1(n9977), .A2(n9978), .ZN(n9993) );
  OAI211_X1 U12589 ( .C1(n9978), .C2(n9977), .A(n14865), .B(n9993), .ZN(n9979)
         );
  OAI211_X1 U12590 ( .C1(n14820), .C2(n9998), .A(n9980), .B(n9979), .ZN(
        P2_U3219) );
  INV_X1 U12591 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U12592 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14865), .B1(n14868), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n9984) );
  INV_X1 U12593 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10528) );
  NAND2_X1 U12594 ( .A1(n14865), .A2(n10528), .ZN(n9982) );
  NAND2_X1 U12595 ( .A1(n14868), .A2(n14916), .ZN(n9981) );
  AND3_X1 U12596 ( .A1(n14820), .A2(n9982), .A3(n9981), .ZN(n9983) );
  MUX2_X1 U12597 ( .A(n9984), .B(n9983), .S(P2_IR_REG_0__SCAN_IN), .Z(n9986)
         );
  NAND2_X1 U12598 ( .A1(n14859), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n9985) );
  OAI211_X1 U12599 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10527), .A(n9986), .B(
        n9985), .ZN(P2_U3214) );
  INV_X1 U12600 ( .A(n14140), .ZN(n10307) );
  OAI222_X1 U12601 ( .A1(P1_U3086), .A2(n10307), .B1(n14534), .B2(n9988), .C1(
        n9987), .C2(n14528), .ZN(P1_U3347) );
  OAI222_X1 U12602 ( .A1(P2_U3088), .A2(n10064), .B1(n13800), .B2(n9988), .C1(
        n10166), .C2(n13803), .ZN(P2_U3319) );
  INV_X1 U12603 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n9990) );
  NAND2_X1 U12604 ( .A1(n10616), .A2(P3_U3897), .ZN(n9989) );
  OAI21_X1 U12605 ( .B1(P3_U3897), .B2(n9990), .A(n9989), .ZN(P3_U3494) );
  INV_X1 U12606 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n9992) );
  NAND2_X1 U12607 ( .A1(n12991), .A2(P3_U3897), .ZN(n9991) );
  OAI21_X1 U12608 ( .B1(P3_U3897), .B2(n9992), .A(n9991), .ZN(P3_U3507) );
  OAI21_X1 U12609 ( .B1(n9974), .B2(n9998), .A(n9993), .ZN(n13303) );
  MUX2_X1 U12610 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10772), .S(n9999), .Z(
        n13302) );
  INV_X1 U12611 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9994) );
  MUX2_X1 U12612 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9994), .S(n10002), .Z(
        n14831) );
  AND2_X1 U12613 ( .A1(n14830), .A2(n14831), .ZN(n14828) );
  MUX2_X1 U12614 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10992), .S(n10064), .Z(
        n9995) );
  AOI211_X1 U12615 ( .C1(n9996), .C2(n9995), .A(n11825), .B(n14849), .ZN(
        n10010) );
  NOR2_X1 U12616 ( .A1(n9998), .A2(n9997), .ZN(n13305) );
  MUX2_X1 U12617 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10000), .S(n9999), .Z(
        n13304) );
  OAI21_X1 U12618 ( .B1(n13306), .B2(n13305), .A(n13304), .ZN(n13308) );
  OAI21_X1 U12619 ( .B1(n10000), .B2(n13298), .A(n13308), .ZN(n14840) );
  INV_X1 U12620 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10001) );
  MUX2_X1 U12621 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10001), .S(n10002), .Z(
        n14839) );
  NAND2_X1 U12622 ( .A1(n14840), .A2(n14839), .ZN(n14838) );
  NAND2_X1 U12623 ( .A1(n10002), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10004) );
  MUX2_X1 U12624 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9142), .S(n10064), .Z(
        n10003) );
  AOI21_X1 U12625 ( .B1(n14838), .B2(n10004), .A(n10003), .ZN(n10065) );
  AND3_X1 U12626 ( .A1(n14838), .A2(n10004), .A3(n10003), .ZN(n10005) );
  NOR3_X1 U12627 ( .A1(n10065), .A2(n10005), .A3(n13328), .ZN(n10009) );
  NAND2_X1 U12628 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10874) );
  INV_X1 U12629 ( .A(n10874), .ZN(n10006) );
  AOI21_X1 U12630 ( .B1(n14859), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n10006), .ZN(
        n10007) );
  OAI21_X1 U12631 ( .B1(n10064), .B2(n14820), .A(n10007), .ZN(n10008) );
  OR3_X1 U12632 ( .A1(n10010), .A2(n10009), .A3(n10008), .ZN(P2_U3222) );
  INV_X1 U12633 ( .A(n11698), .ZN(n11700) );
  OAI222_X1 U12634 ( .A1(n13140), .A2(n10012), .B1(n13142), .B2(n10011), .C1(
        n11700), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12635 ( .A(n14853), .ZN(n10060) );
  OAI222_X1 U12636 ( .A1(P2_U3088), .A2(n10060), .B1(n13800), .B2(n10014), 
        .C1(n10164), .C2(n13803), .ZN(P2_U3318) );
  INV_X1 U12637 ( .A(n14159), .ZN(n10309) );
  OAI222_X1 U12638 ( .A1(P1_U3086), .A2(n10309), .B1(n14534), .B2(n10014), 
        .C1(n10013), .C2(n14528), .ZN(P1_U3346) );
  OAI222_X1 U12639 ( .A1(n13140), .A2(n10016), .B1(n14559), .B2(P3_U3151), 
        .C1(n10015), .C2(n13142), .ZN(P3_U3280) );
  INV_X1 U12640 ( .A(n12076), .ZN(n10706) );
  INV_X1 U12641 ( .A(n13295), .ZN(n10452) );
  OAI22_X1 U12642 ( .A1(n10517), .A2(n13630), .B1(n10452), .B2(n13632), .ZN(
        n10096) );
  NAND2_X1 U12643 ( .A1(n14881), .A2(n10017), .ZN(n10465) );
  INV_X1 U12644 ( .A(n10465), .ZN(n10521) );
  AND2_X1 U12645 ( .A1(n10018), .A2(n10521), .ZN(n10433) );
  INV_X1 U12646 ( .A(n10433), .ZN(n10085) );
  AOI22_X1 U12647 ( .A1(n13251), .A2(n10096), .B1(n10085), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10023) );
  OAI21_X1 U12648 ( .B1(n10020), .B2(n10019), .A(n10436), .ZN(n10021) );
  NAND2_X1 U12649 ( .A1(n10021), .A2(n9485), .ZN(n10022) );
  OAI211_X1 U12650 ( .C1(n10706), .C2(n13258), .A(n10023), .B(n10022), .ZN(
        P2_U3194) );
  INV_X1 U12651 ( .A(n10042), .ZN(n14044) );
  INV_X1 U12652 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14803) );
  MUX2_X1 U12653 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n14803), .S(n10042), .Z(
        n14041) );
  NAND2_X1 U12654 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14042) );
  NOR2_X1 U12655 ( .A1(n14041), .A2(n14042), .ZN(n14040) );
  AOI21_X1 U12656 ( .B1(n14044), .B2(P1_REG1_REG_1__SCAN_IN), .A(n14040), .ZN(
        n14064) );
  INV_X1 U12657 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10733) );
  MUX2_X1 U12658 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10733), .S(n14057), .Z(
        n14063) );
  NOR2_X1 U12659 ( .A1(n14064), .A2(n14063), .ZN(n14079) );
  NOR2_X1 U12660 ( .A1(n14057), .A2(n10733), .ZN(n14075) );
  INV_X1 U12661 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10024) );
  MUX2_X1 U12662 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10024), .S(n14074), .Z(
        n10025) );
  NAND2_X1 U12663 ( .A1(n14074), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14089) );
  MUX2_X1 U12664 ( .A(n8181), .B(P1_REG1_REG_4__SCAN_IN), .S(n14093), .Z(
        n14088) );
  AOI21_X1 U12665 ( .B1(n14090), .B2(n14089), .A(n14088), .ZN(n14087) );
  AOI21_X1 U12666 ( .B1(n14093), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14087), .ZN(
        n14106) );
  MUX2_X1 U12667 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n8211), .S(n14109), .Z(
        n14107) );
  OAI21_X1 U12668 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n14109), .A(n14105), .ZN(
        n14117) );
  MUX2_X1 U12669 ( .A(n14118), .B(P1_REG1_REG_6__SCAN_IN), .S(n14125), .Z(
        n10026) );
  OR2_X1 U12670 ( .A1(n14117), .A2(n10026), .ZN(n14119) );
  NAND2_X1 U12671 ( .A1(n14125), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10028) );
  MUX2_X1 U12672 ( .A(n8248), .B(P1_REG1_REG_7__SCAN_IN), .S(n10306), .Z(
        n10027) );
  NAND3_X1 U12673 ( .A1(n14119), .A2(n10028), .A3(n10027), .ZN(n10030) );
  OAI21_X1 U12674 ( .B1(n10334), .B2(n10029), .A(n8113), .ZN(n10034) );
  NOR2_X1 U12675 ( .A1(n10343), .A2(n8819), .ZN(n10032) );
  OR2_X1 U12676 ( .A1(n10034), .A2(n10032), .ZN(n14718) );
  NOR2_X2 U12677 ( .A1(n14718), .A2(n14708), .ZN(n14194) );
  NAND2_X1 U12678 ( .A1(n10030), .A2(n14194), .ZN(n10059) );
  NOR2_X2 U12679 ( .A1(n14718), .A2(n10031), .ZN(n14722) );
  INV_X1 U12680 ( .A(n10032), .ZN(n10033) );
  AND2_X1 U12681 ( .A1(n10034), .A2(n10033), .ZN(n14733) );
  OR2_X1 U12682 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8249), .ZN(n11189) );
  OAI21_X1 U12683 ( .B1(n14199), .B2(n15108), .A(n11189), .ZN(n10035) );
  AOI21_X1 U12684 ( .B1(n10306), .B2(n14722), .A(n10035), .ZN(n10058) );
  INV_X1 U12685 ( .A(n14718), .ZN(n10037) );
  NOR2_X1 U12686 ( .A1(n14055), .A2(n14524), .ZN(n10036) );
  NAND2_X1 U12687 ( .A1(n10037), .A2(n10036), .ZN(n14190) );
  MUX2_X1 U12688 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10038), .S(n14074), .Z(
        n10044) );
  MUX2_X1 U12689 ( .A(n10039), .B(P1_REG2_REG_2__SCAN_IN), .S(n14057), .Z(
        n14062) );
  MUX2_X1 U12690 ( .A(n10040), .B(P1_REG2_REG_1__SCAN_IN), .S(n10042), .Z(
        n14046) );
  AND2_X1 U12691 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10041) );
  NAND2_X1 U12692 ( .A1(n14046), .A2(n10041), .ZN(n14045) );
  OAI21_X1 U12693 ( .B1(n10040), .B2(n10042), .A(n14045), .ZN(n14061) );
  NAND2_X1 U12694 ( .A1(n14062), .A2(n14061), .ZN(n14070) );
  OR2_X1 U12695 ( .A1(n14057), .A2(n10039), .ZN(n14069) );
  NAND2_X1 U12696 ( .A1(n14070), .A2(n14069), .ZN(n10043) );
  NAND2_X1 U12697 ( .A1(n10044), .A2(n10043), .ZN(n14095) );
  NAND2_X1 U12698 ( .A1(n14074), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14094) );
  NAND2_X1 U12699 ( .A1(n14095), .A2(n14094), .ZN(n10046) );
  MUX2_X1 U12700 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11097), .S(n14093), .Z(
        n10045) );
  NAND2_X1 U12701 ( .A1(n10046), .A2(n10045), .ZN(n14112) );
  NAND2_X1 U12702 ( .A1(n14093), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U12703 ( .A1(n14112), .A2(n14111), .ZN(n10049) );
  MUX2_X1 U12704 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10047), .S(n14109), .Z(
        n10048) );
  NAND2_X1 U12705 ( .A1(n10049), .A2(n10048), .ZN(n14128) );
  NAND2_X1 U12706 ( .A1(n14109), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14126) );
  NAND2_X1 U12707 ( .A1(n14128), .A2(n14126), .ZN(n10051) );
  MUX2_X1 U12708 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11172), .S(n14125), .Z(
        n10050) );
  NAND2_X1 U12709 ( .A1(n10051), .A2(n10050), .ZN(n14130) );
  NAND2_X1 U12710 ( .A1(n14125), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U12711 ( .A1(n14130), .A2(n10055), .ZN(n10053) );
  MUX2_X1 U12712 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11252), .S(n10306), .Z(
        n10052) );
  NAND2_X1 U12713 ( .A1(n10053), .A2(n10052), .ZN(n14143) );
  MUX2_X1 U12714 ( .A(n11252), .B(P1_REG2_REG_7__SCAN_IN), .S(n10306), .Z(
        n10054) );
  NAND3_X1 U12715 ( .A1(n14130), .A2(n10055), .A3(n10054), .ZN(n10056) );
  NAND3_X1 U12716 ( .A1(n14724), .A2(n14143), .A3(n10056), .ZN(n10057) );
  OAI211_X1 U12717 ( .C1(n10305), .C2(n10059), .A(n10058), .B(n10057), .ZN(
        P1_U3250) );
  NOR2_X1 U12718 ( .A1(n14733), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12719 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11046) );
  NOR2_X1 U12720 ( .A1(n10064), .A2(n10992), .ZN(n14848) );
  XNOR2_X1 U12721 ( .A(n14853), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n14847) );
  AOI21_X1 U12722 ( .B1(n10060), .B2(n11046), .A(n14846), .ZN(n10063) );
  INV_X1 U12723 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10061) );
  MUX2_X1 U12724 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10061), .S(n10260), .Z(
        n10062) );
  NAND2_X1 U12725 ( .A1(n10063), .A2(n10062), .ZN(n10254) );
  OAI211_X1 U12726 ( .C1(n10063), .C2(n10062), .A(n10254), .B(n14865), .ZN(
        n10076) );
  INV_X1 U12727 ( .A(n10064), .ZN(n10066) );
  AOI21_X1 U12728 ( .B1(n10066), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10065), .ZN(
        n14845) );
  INV_X1 U12729 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10067) );
  MUX2_X1 U12730 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10067), .S(n14853), .Z(
        n14844) );
  NAND2_X1 U12731 ( .A1(n14845), .A2(n14844), .ZN(n14843) );
  OAI21_X1 U12732 ( .B1(n14853), .B2(P2_REG1_REG_9__SCAN_IN), .A(n14843), .ZN(
        n10070) );
  INV_X1 U12733 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10068) );
  MUX2_X1 U12734 ( .A(n10068), .B(P2_REG1_REG_10__SCAN_IN), .S(n10260), .Z(
        n10069) );
  AOI21_X1 U12735 ( .B1(n10070), .B2(n10069), .A(n13328), .ZN(n10074) );
  OR2_X1 U12736 ( .A1(n10070), .A2(n10069), .ZN(n10263) );
  INV_X1 U12737 ( .A(n10260), .ZN(n10255) );
  NOR2_X1 U12738 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11081), .ZN(n10071) );
  AOI21_X1 U12739 ( .B1(n14859), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10071), 
        .ZN(n10072) );
  OAI21_X1 U12740 ( .B1(n10255), .B2(n14820), .A(n10072), .ZN(n10073) );
  AOI21_X1 U12741 ( .B1(n10074), .B2(n10263), .A(n10073), .ZN(n10075) );
  NAND2_X1 U12742 ( .A1(n10076), .A2(n10075), .ZN(P2_U3224) );
  INV_X1 U12743 ( .A(n12740), .ZN(n12733) );
  OAI222_X1 U12744 ( .A1(n13140), .A2(n10078), .B1(n12733), .B2(P3_U3151), 
        .C1(n10077), .C2(n13142), .ZN(P3_U3279) );
  INV_X1 U12745 ( .A(n10324), .ZN(n10319) );
  INV_X1 U12746 ( .A(n10079), .ZN(n10081) );
  OAI222_X1 U12747 ( .A1(n10319), .A2(P1_U3086), .B1(n14534), .B2(n10081), 
        .C1(n10080), .C2(n14528), .ZN(P1_U3345) );
  OAI222_X1 U12748 ( .A1(n13803), .A2(n10082), .B1(n13800), .B2(n10081), .C1(
        P2_U3088), .C2(n10255), .ZN(P2_U3317) );
  INV_X1 U12749 ( .A(n6734), .ZN(n10524) );
  NAND2_X1 U12750 ( .A1(n9485), .A2(n9321), .ZN(n13262) );
  OAI22_X1 U12751 ( .A1(n13262), .A2(n10517), .B1(n12063), .B2(n13272), .ZN(
        n10084) );
  NAND2_X1 U12752 ( .A1(n10084), .A2(n10083), .ZN(n10087) );
  AOI22_X1 U12753 ( .A1(n13281), .A2(n12059), .B1(n10085), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10086) );
  OAI211_X1 U12754 ( .C1(n10524), .C2(n13278), .A(n10087), .B(n10086), .ZN(
        P2_U3204) );
  INV_X1 U12755 ( .A(n10518), .ZN(n10091) );
  INV_X1 U12756 ( .A(n10111), .ZN(n10090) );
  AOI21_X1 U12757 ( .B1(n10091), .B2(n12297), .A(n10090), .ZN(n10711) );
  INV_X1 U12758 ( .A(n10711), .ZN(n10099) );
  NAND2_X1 U12759 ( .A1(n6761), .A2(n12059), .ZN(n10092) );
  NAND2_X1 U12760 ( .A1(n10092), .A2(n13639), .ZN(n10093) );
  NOR2_X1 U12761 ( .A1(n10113), .A2(n10093), .ZN(n10708) );
  NOR2_X1 U12762 ( .A1(n12064), .A2(n12063), .ZN(n10094) );
  OAI21_X1 U12763 ( .B1(n10094), .B2(n12297), .A(n10116), .ZN(n10097) );
  NAND2_X1 U12764 ( .A1(n12343), .A2(n13330), .ZN(n12229) );
  OR2_X1 U12765 ( .A1(n12329), .A2(n12331), .ZN(n10095) );
  AOI21_X1 U12766 ( .B1(n10097), .B2(n13635), .A(n10096), .ZN(n10704) );
  INV_X1 U12767 ( .A(n10704), .ZN(n10098) );
  AOI211_X1 U12768 ( .C1(n14623), .C2(n10099), .A(n10708), .B(n10098), .ZN(
        n10570) );
  INV_X1 U12769 ( .A(n14877), .ZN(n10100) );
  NAND2_X1 U12770 ( .A1(n10100), .A2(n10463), .ZN(n10101) );
  NOR2_X1 U12771 ( .A1(n10101), .A2(n10465), .ZN(n10103) );
  INV_X1 U12772 ( .A(n14880), .ZN(n10520) );
  NOR2_X1 U12773 ( .A1(n10520), .A2(n10102), .ZN(n10467) );
  NAND2_X1 U12774 ( .A1(n14922), .A2(n14889), .ZN(n13749) );
  AOI22_X1 U12775 ( .A1(n13742), .A2(n6761), .B1(n14920), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10104) );
  OAI21_X1 U12776 ( .B1(n10570), .B2(n14920), .A(n10104), .ZN(P2_U3500) );
  INV_X1 U12777 ( .A(n10105), .ZN(n10108) );
  INV_X1 U12778 ( .A(n10476), .ZN(n10106) );
  OAI222_X1 U12779 ( .A1(n14528), .A2(n10107), .B1(n14534), .B2(n10108), .C1(
        P1_U3086), .C2(n10106), .ZN(P1_U3344) );
  INV_X1 U12780 ( .A(n10597), .ZN(n10590) );
  OAI222_X1 U12781 ( .A1(n13803), .A2(n10109), .B1(n13800), .B2(n10108), .C1(
        P2_U3088), .C2(n10590), .ZN(P2_U3316) );
  OR2_X1 U12782 ( .A1(n6734), .A2(n6761), .ZN(n10110) );
  NAND2_X1 U12783 ( .A1(n10111), .A2(n10110), .ZN(n10112) );
  INV_X1 U12784 ( .A(n12296), .ZN(n10117) );
  NAND2_X1 U12785 ( .A1(n10112), .A2(n10117), .ZN(n10419) );
  OAI21_X1 U12786 ( .B1(n10112), .B2(n10117), .A(n10419), .ZN(n10734) );
  OAI21_X1 U12787 ( .B1(n10113), .B2(n10736), .A(n13639), .ZN(n10114) );
  NOR2_X1 U12788 ( .A1(n10114), .A2(n10457), .ZN(n10739) );
  OR2_X1 U12789 ( .A1(n6734), .A2(n10706), .ZN(n10115) );
  XNOR2_X1 U12790 ( .A(n10117), .B(n10423), .ZN(n10118) );
  INV_X1 U12791 ( .A(n13635), .ZN(n11543) );
  AOI22_X1 U12792 ( .A1(n13294), .A2(n13544), .B1(n13542), .B2(n6734), .ZN(
        n10434) );
  OAI21_X1 U12793 ( .B1(n10118), .B2(n11543), .A(n10434), .ZN(n10740) );
  AOI211_X1 U12794 ( .C1(n14623), .C2(n10734), .A(n10739), .B(n10740), .ZN(
        n10578) );
  AOI22_X1 U12795 ( .A1(n13742), .A2(n12073), .B1(n14920), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10119) );
  OAI21_X1 U12796 ( .B1(n10578), .B2(n14920), .A(n10119), .ZN(P2_U3501) );
  INV_X1 U12797 ( .A(n6450), .ZN(n11203) );
  OAI21_X1 U12798 ( .B1(n10122), .B2(n10121), .A(n10120), .ZN(n14052) );
  NAND2_X1 U12799 ( .A1(n14052), .A2(n14655), .ZN(n10124) );
  NAND2_X1 U12800 ( .A1(n14697), .A2(n10342), .ZN(n10489) );
  AOI22_X1 U12801 ( .A1(n14653), .A2(n10718), .B1(n10489), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10123) );
  OAI211_X1 U12802 ( .C1(n11203), .C2(n13975), .A(n10124), .B(n10123), .ZN(
        P1_U3232) );
  MUX2_X1 U12803 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n11411), .Z(n10168) );
  XNOR2_X1 U12804 ( .A(n10168), .B(n6454), .ZN(n10169) );
  MUX2_X1 U12805 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n7491), .Z(n10126) );
  XOR2_X1 U12806 ( .A(n10145), .B(n10126), .Z(n10199) );
  INV_X1 U12807 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10125) );
  INV_X1 U12808 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10159) );
  MUX2_X1 U12809 ( .A(n10125), .B(n10159), .S(n7491), .Z(n12707) );
  AND2_X1 U12810 ( .A1(n12707), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n12712) );
  INV_X1 U12811 ( .A(n10145), .ZN(n10211) );
  INV_X1 U12812 ( .A(n10126), .ZN(n10127) );
  XOR2_X1 U12813 ( .A(n10170), .B(n10169), .Z(n10155) );
  INV_X1 U12814 ( .A(n6454), .ZN(n10153) );
  AOI21_X1 U12815 ( .B1(n6458), .B2(n10130), .A(n10129), .ZN(n10132) );
  NAND2_X1 U12816 ( .A1(n10131), .A2(n12693), .ZN(n10133) );
  NAND2_X1 U12817 ( .A1(n10132), .A2(n10133), .ZN(n10141) );
  MUX2_X1 U12818 ( .A(n12706), .B(n10141), .S(n6710), .Z(n14966) );
  INV_X1 U12819 ( .A(n10132), .ZN(n10134) );
  AOI22_X1 U12820 ( .A1(n14923), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10151) );
  INV_X1 U12821 ( .A(n14983), .ZN(n12710) );
  INV_X1 U12822 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10136) );
  AND2_X1 U12823 ( .A1(n10142), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n12711) );
  NAND2_X1 U12824 ( .A1(n7521), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10137) );
  OAI21_X1 U12825 ( .B1(n10145), .B2(n12711), .A(n10137), .ZN(n10202) );
  INV_X1 U12826 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15001) );
  OR2_X1 U12827 ( .A1(n10202), .A2(n15001), .ZN(n10200) );
  NAND2_X1 U12828 ( .A1(n10200), .A2(n10137), .ZN(n10138) );
  NAND2_X1 U12829 ( .A1(n10139), .A2(n10138), .ZN(n10174) );
  OAI21_X1 U12830 ( .B1(n10139), .B2(n10138), .A(n10174), .ZN(n10140) );
  NAND2_X1 U12831 ( .A1(n12710), .A2(n10140), .ZN(n10150) );
  INV_X1 U12832 ( .A(n14977), .ZN(n12709) );
  INV_X1 U12833 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15042) );
  NAND2_X1 U12834 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10142), .ZN(n10143) );
  INV_X1 U12835 ( .A(n10143), .ZN(n10144) );
  OAI21_X1 U12836 ( .B1(n10145), .B2(n10144), .A(n7448), .ZN(n10203) );
  INV_X1 U12837 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15040) );
  NAND2_X1 U12838 ( .A1(n10205), .A2(n7448), .ZN(n10146) );
  OAI21_X1 U12839 ( .B1(n10147), .B2(n10146), .A(n10184), .ZN(n10148) );
  NAND2_X1 U12840 ( .A1(n12709), .A2(n10148), .ZN(n10149) );
  NAND3_X1 U12841 ( .A1(n10151), .A2(n10150), .A3(n10149), .ZN(n10152) );
  AOI21_X1 U12842 ( .B1(n10153), .B2(n14954), .A(n10152), .ZN(n10154) );
  OAI21_X1 U12843 ( .B1(n10155), .B2(n14975), .A(n10154), .ZN(P3_U3184) );
  AND2_X1 U12844 ( .A1(n6657), .A2(n12529), .ZN(n12525) );
  NOR2_X1 U12845 ( .A1(n14985), .A2(n12525), .ZN(n12497) );
  OR3_X1 U12846 ( .A1(n12497), .A2(n15015), .A3(n10156), .ZN(n10158) );
  OR2_X1 U12847 ( .A1(n6618), .A2(n12958), .ZN(n10157) );
  NAND2_X1 U12848 ( .A1(n10158), .A2(n10157), .ZN(n10446) );
  NOR2_X1 U12849 ( .A1(n15051), .A2(n10159), .ZN(n10160) );
  AOI21_X1 U12850 ( .B1(n10446), .B2(n15051), .A(n10160), .ZN(n10161) );
  OAI21_X1 U12851 ( .B1(n12529), .B2(n13027), .A(n10161), .ZN(P3_U3459) );
  MUX2_X1 U12852 ( .A(n10162), .B(n11273), .S(P1_U4016), .Z(n10163) );
  INV_X1 U12853 ( .A(n10163), .ZN(P1_U3564) );
  MUX2_X1 U12854 ( .A(n10164), .B(n11656), .S(P1_U4016), .Z(n10165) );
  INV_X1 U12855 ( .A(n10165), .ZN(P1_U3569) );
  MUX2_X1 U12856 ( .A(n10166), .B(n11627), .S(P1_U4016), .Z(n10167) );
  INV_X1 U12857 ( .A(n10167), .ZN(P1_U3568) );
  MUX2_X1 U12858 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12799), .Z(n10234) );
  XNOR2_X1 U12859 ( .A(n10234), .B(n10240), .ZN(n10235) );
  OAI22_X1 U12860 ( .A1(n10170), .A2(n10169), .B1(n10168), .B2(n6453), .ZN(
        n10214) );
  MUX2_X1 U12861 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n11411), .Z(n10171) );
  XOR2_X1 U12862 ( .A(n10185), .B(n10171), .Z(n10215) );
  INV_X1 U12863 ( .A(n10185), .ZN(n10228) );
  INV_X1 U12864 ( .A(n10171), .ZN(n10172) );
  AOI22_X1 U12865 ( .A1(n10214), .A2(n10215), .B1(n10228), .B2(n10172), .ZN(
        n10236) );
  XOR2_X1 U12866 ( .A(n10236), .B(n10235), .Z(n10198) );
  NAND2_X1 U12867 ( .A1(n6453), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10173) );
  NAND2_X1 U12868 ( .A1(n10174), .A2(n10173), .ZN(n10175) );
  NAND2_X1 U12869 ( .A1(n10175), .A2(n10185), .ZN(n10179) );
  OAI21_X1 U12870 ( .B1(n10175), .B2(n10185), .A(n10179), .ZN(n10218) );
  INV_X1 U12871 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10827) );
  INV_X1 U12872 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10176) );
  MUX2_X1 U12873 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10176), .S(n10240), .Z(
        n10178) );
  INV_X1 U12874 ( .A(n10178), .ZN(n10180) );
  NAND3_X1 U12875 ( .A1(n10216), .A2(n10180), .A3(n10179), .ZN(n10181) );
  NAND2_X1 U12876 ( .A1(n10237), .A2(n10181), .ZN(n10196) );
  NAND2_X1 U12877 ( .A1(n6454), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10183) );
  OAI21_X1 U12878 ( .B1(n10186), .B2(n10185), .A(n10189), .ZN(n10220) );
  INV_X1 U12879 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U12880 ( .A1(n10222), .A2(n10189), .ZN(n10187) );
  INV_X1 U12881 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10671) );
  MUX2_X1 U12882 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10671), .S(n10240), .Z(
        n10188) );
  NAND2_X1 U12883 ( .A1(n10187), .A2(n10188), .ZN(n10242) );
  INV_X1 U12884 ( .A(n10188), .ZN(n10190) );
  NAND3_X1 U12885 ( .A1(n10222), .A2(n10190), .A3(n10189), .ZN(n10191) );
  AND2_X1 U12886 ( .A1(n10242), .A2(n10191), .ZN(n10193) );
  NAND2_X1 U12887 ( .A1(n14923), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U12888 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10617) );
  OAI211_X1 U12889 ( .C1(n14977), .C2(n10193), .A(n10192), .B(n10617), .ZN(
        n10195) );
  NOR2_X1 U12890 ( .A1(n14966), .A2(n10240), .ZN(n10194) );
  AOI211_X1 U12891 ( .C1(n12710), .C2(n10196), .A(n10195), .B(n10194), .ZN(
        n10197) );
  OAI21_X1 U12892 ( .B1(n10198), .B2(n14975), .A(n10197), .ZN(P3_U3186) );
  XOR2_X1 U12893 ( .A(n12712), .B(n10199), .Z(n10213) );
  INV_X1 U12894 ( .A(n10200), .ZN(n10201) );
  AOI21_X1 U12895 ( .B1(n15001), .B2(n10202), .A(n10201), .ZN(n10209) );
  AOI22_X1 U12896 ( .A1(n14923), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10208) );
  NAND2_X1 U12897 ( .A1(n10203), .A2(n15040), .ZN(n10204) );
  NAND2_X1 U12898 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  NAND2_X1 U12899 ( .A1(n12709), .A2(n10206), .ZN(n10207) );
  OAI211_X1 U12900 ( .C1(n10209), .C2(n14983), .A(n10208), .B(n10207), .ZN(
        n10210) );
  AOI21_X1 U12901 ( .B1(n10211), .B2(n14954), .A(n10210), .ZN(n10212) );
  OAI21_X1 U12902 ( .B1(n14975), .B2(n10213), .A(n10212), .ZN(P3_U3183) );
  XOR2_X1 U12903 ( .A(n10214), .B(n10215), .Z(n10230) );
  INV_X1 U12904 ( .A(n10216), .ZN(n10217) );
  AOI21_X1 U12905 ( .B1(n10827), .B2(n10218), .A(n10217), .ZN(n10226) );
  AND2_X1 U12906 ( .A1(P3_U3151), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n10583) );
  AOI21_X1 U12907 ( .B1(n14923), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10583), .ZN(
        n10225) );
  NAND2_X1 U12908 ( .A1(n10220), .A2(n10219), .ZN(n10221) );
  NAND2_X1 U12909 ( .A1(n10222), .A2(n10221), .ZN(n10223) );
  NAND2_X1 U12910 ( .A1(n12709), .A2(n10223), .ZN(n10224) );
  OAI211_X1 U12911 ( .C1(n10226), .C2(n14983), .A(n10225), .B(n10224), .ZN(
        n10227) );
  AOI21_X1 U12912 ( .B1(n10228), .B2(n14954), .A(n10227), .ZN(n10229) );
  OAI21_X1 U12913 ( .B1(n10230), .B2(n14975), .A(n10229), .ZN(P3_U3185) );
  INV_X1 U12914 ( .A(n10231), .ZN(n10232) );
  OAI222_X1 U12915 ( .A1(n13142), .A2(n10233), .B1(n13140), .B2(n10232), .C1(
        P3_U3151), .C2(n12778), .ZN(P3_U3278) );
  MUX2_X1 U12916 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12799), .Z(n10271) );
  XOR2_X1 U12917 ( .A(n10243), .B(n10271), .Z(n10273) );
  OAI22_X1 U12918 ( .A1(n10236), .A2(n10235), .B1(n10234), .B2(n10240), .ZN(
        n10274) );
  XOR2_X1 U12919 ( .A(n10274), .B(n10273), .Z(n10253) );
  INV_X1 U12920 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10890) );
  NAND2_X1 U12921 ( .A1(n10238), .A2(n10890), .ZN(n10239) );
  AOI21_X1 U12922 ( .B1(n10281), .B2(n10239), .A(n14983), .ZN(n10251) );
  INV_X1 U12923 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10247) );
  NAND2_X1 U12924 ( .A1(n10240), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10241) );
  NAND2_X1 U12925 ( .A1(n10244), .A2(n10243), .ZN(n10285) );
  INV_X1 U12926 ( .A(n10287), .ZN(n10245) );
  AOI21_X1 U12927 ( .B1(n10247), .B2(n10246), .A(n10245), .ZN(n10249) );
  OR2_X1 U12928 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7559), .ZN(n10812) );
  NAND2_X1 U12929 ( .A1(n14923), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10248) );
  OAI211_X1 U12930 ( .C1(n10249), .C2(n14977), .A(n10812), .B(n10248), .ZN(
        n10250) );
  AOI211_X1 U12931 ( .C1(n14954), .C2(n6715), .A(n10251), .B(n10250), .ZN(
        n10252) );
  OAI21_X1 U12932 ( .B1(n10253), .B2(n14975), .A(n10252), .ZN(P3_U3187) );
  MUX2_X1 U12933 ( .A(n11373), .B(P2_REG2_REG_11__SCAN_IN), .S(n10597), .Z(
        n10257) );
  OAI21_X1 U12934 ( .B1(n10255), .B2(n10061), .A(n10254), .ZN(n10256) );
  AOI21_X1 U12935 ( .B1(n10257), .B2(n10256), .A(n10589), .ZN(n10268) );
  AND2_X1 U12936 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10259) );
  NOR2_X1 U12937 ( .A1(n10590), .A2(n14820), .ZN(n10258) );
  AOI211_X1 U12938 ( .C1(n14859), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n10259), 
        .B(n10258), .ZN(n10267) );
  NAND2_X1 U12939 ( .A1(n10260), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10262) );
  MUX2_X1 U12940 ( .A(n9193), .B(P2_REG1_REG_11__SCAN_IN), .S(n10597), .Z(
        n10261) );
  AOI21_X1 U12941 ( .B1(n10263), .B2(n10262), .A(n10261), .ZN(n10596) );
  INV_X1 U12942 ( .A(n10596), .ZN(n10265) );
  NAND3_X1 U12943 ( .A1(n10263), .A2(n10262), .A3(n10261), .ZN(n10264) );
  NAND3_X1 U12944 ( .A1(n10265), .A2(n14868), .A3(n10264), .ZN(n10266) );
  OAI211_X1 U12945 ( .C1(n10268), .C2(n11825), .A(n10267), .B(n10266), .ZN(
        P2_U3225) );
  INV_X1 U12946 ( .A(n12802), .ZN(n12788) );
  OAI222_X1 U12947 ( .A1(n13140), .A2(n10270), .B1(n13142), .B2(n10269), .C1(
        n12788), .C2(P3_U3151), .ZN(P3_U3277) );
  MUX2_X1 U12948 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12799), .Z(n10534) );
  XNOR2_X1 U12949 ( .A(n10534), .B(n10552), .ZN(n10535) );
  INV_X1 U12950 ( .A(n10271), .ZN(n10272) );
  XOR2_X1 U12951 ( .A(n10536), .B(n10535), .Z(n10293) );
  INV_X1 U12952 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15132) );
  NOR2_X1 U12953 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15132), .ZN(n11107) );
  AOI21_X1 U12954 ( .B1(n14923), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11107), .ZN(
        n10275) );
  OAI21_X1 U12955 ( .B1(n14966), .B2(n10552), .A(n10275), .ZN(n10291) );
  NAND2_X1 U12956 ( .A1(n10281), .A2(n10279), .ZN(n10277) );
  INV_X1 U12957 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10276) );
  MUX2_X1 U12958 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n10276), .S(n10552), .Z(
        n10278) );
  NAND2_X1 U12959 ( .A1(n10277), .A2(n10278), .ZN(n10542) );
  INV_X1 U12960 ( .A(n10278), .ZN(n10280) );
  NAND3_X1 U12961 ( .A1(n10281), .A2(n10280), .A3(n10279), .ZN(n10282) );
  AOI21_X1 U12962 ( .B1(n10542), .B2(n10282), .A(n14983), .ZN(n10290) );
  NAND2_X1 U12963 ( .A1(n10287), .A2(n10285), .ZN(n10283) );
  INV_X1 U12964 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15084) );
  MUX2_X1 U12965 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n15084), .S(n10552), .Z(
        n10284) );
  INV_X1 U12966 ( .A(n10284), .ZN(n10286) );
  NAND3_X1 U12967 ( .A1(n10287), .A2(n10286), .A3(n10285), .ZN(n10288) );
  AOI21_X1 U12968 ( .B1(n10554), .B2(n10288), .A(n14977), .ZN(n10289) );
  NOR3_X1 U12969 ( .A1(n10291), .A2(n10290), .A3(n10289), .ZN(n10292) );
  OAI21_X1 U12970 ( .B1(n10293), .B2(n14975), .A(n10292), .ZN(P3_U3188) );
  INV_X1 U12971 ( .A(n14722), .ZN(n11859) );
  NAND2_X1 U12972 ( .A1(n10306), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n14142) );
  NAND2_X1 U12973 ( .A1(n14143), .A2(n14142), .ZN(n10296) );
  MUX2_X1 U12974 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10294), .S(n14140), .Z(
        n10295) );
  NAND2_X1 U12975 ( .A1(n10296), .A2(n10295), .ZN(n14156) );
  NAND2_X1 U12976 ( .A1(n14140), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n14155) );
  NAND2_X1 U12977 ( .A1(n14156), .A2(n14155), .ZN(n10298) );
  MUX2_X1 U12978 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11483), .S(n14159), .Z(
        n10297) );
  NAND2_X1 U12979 ( .A1(n10298), .A2(n10297), .ZN(n14158) );
  NAND2_X1 U12980 ( .A1(n14159), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U12981 ( .A1(n14158), .A2(n10303), .ZN(n10301) );
  MUX2_X1 U12982 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10299), .S(n10324), .Z(
        n10300) );
  NAND2_X1 U12983 ( .A1(n10301), .A2(n10300), .ZN(n10329) );
  MUX2_X1 U12984 ( .A(n10299), .B(P1_REG2_REG_10__SCAN_IN), .S(n10324), .Z(
        n10302) );
  NAND3_X1 U12985 ( .A1(n14158), .A2(n10303), .A3(n10302), .ZN(n10304) );
  NAND3_X1 U12986 ( .A1(n10329), .A2(n14724), .A3(n10304), .ZN(n10316) );
  NAND2_X1 U12987 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11657)
         );
  AOI21_X1 U12988 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10306), .A(n10305), .ZN(
        n14134) );
  MUX2_X1 U12989 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n8281), .S(n14140), .Z(
        n14135) );
  NAND2_X1 U12990 ( .A1(n14134), .A2(n14135), .ZN(n14150) );
  NAND2_X1 U12991 ( .A1(n10307), .A2(n8281), .ZN(n14148) );
  MUX2_X1 U12992 ( .A(n10308), .B(P1_REG1_REG_9__SCAN_IN), .S(n14159), .Z(
        n14149) );
  AOI21_X1 U12993 ( .B1(n14150), .B2(n14148), .A(n14149), .ZN(n14152) );
  MUX2_X1 U12994 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10310), .S(n10324), .Z(
        n10311) );
  NAND2_X1 U12995 ( .A1(n10312), .A2(n10311), .ZN(n10318) );
  OAI211_X1 U12996 ( .C1(n10312), .C2(n10311), .A(n14194), .B(n10318), .ZN(
        n10313) );
  NAND2_X1 U12997 ( .A1(n11657), .A2(n10313), .ZN(n10314) );
  AOI21_X1 U12998 ( .B1(n14733), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10314), 
        .ZN(n10315) );
  OAI211_X1 U12999 ( .C1(n11859), .C2(n10319), .A(n10316), .B(n10315), .ZN(
        P1_U3253) );
  MUX2_X1 U13000 ( .A(n10317), .B(P1_REG1_REG_11__SCAN_IN), .S(n10476), .Z(
        n10321) );
  OAI21_X1 U13001 ( .B1(n10310), .B2(n10319), .A(n10318), .ZN(n10320) );
  AOI21_X1 U13002 ( .B1(n10321), .B2(n10320), .A(n10479), .ZN(n10333) );
  NAND2_X1 U13003 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11762)
         );
  OAI21_X1 U13004 ( .B1(n14199), .B2(n10322), .A(n11762), .ZN(n10323) );
  AOI21_X1 U13005 ( .B1(n14722), .B2(n10476), .A(n10323), .ZN(n10332) );
  NAND2_X1 U13006 ( .A1(n10324), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10328) );
  NAND2_X1 U13007 ( .A1(n10329), .A2(n10328), .ZN(n10326) );
  MUX2_X1 U13008 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11583), .S(n10476), .Z(
        n10325) );
  NAND2_X1 U13009 ( .A1(n10326), .A2(n10325), .ZN(n10472) );
  MUX2_X1 U13010 ( .A(n11583), .B(P1_REG2_REG_11__SCAN_IN), .S(n10476), .Z(
        n10327) );
  NAND3_X1 U13011 ( .A1(n10329), .A2(n10328), .A3(n10327), .ZN(n10330) );
  NAND3_X1 U13012 ( .A1(n10472), .A2(n14724), .A3(n10330), .ZN(n10331) );
  OAI211_X1 U13013 ( .C1(n10333), .C2(n14729), .A(n10332), .B(n10331), .ZN(
        P1_U3254) );
  NAND2_X1 U13014 ( .A1(n10718), .A2(n9770), .ZN(n11195) );
  INV_X1 U13015 ( .A(n11195), .ZN(n10340) );
  AND2_X1 U13016 ( .A1(n10334), .A2(n11239), .ZN(n10335) );
  NAND2_X1 U13017 ( .A1(n13921), .A2(n10335), .ZN(n11278) );
  NAND2_X1 U13018 ( .A1(n10336), .A2(n11196), .ZN(n14430) );
  NAND2_X1 U13019 ( .A1(n14536), .A2(n14195), .ZN(n10338) );
  AOI21_X1 U13020 ( .B1(n14753), .B2(n14795), .A(n11199), .ZN(n10339) );
  AOI211_X1 U13021 ( .C1(n14739), .C2(n6450), .A(n10340), .B(n10339), .ZN(
        n14737) );
  NAND4_X1 U13022 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10717) );
  NAND2_X1 U13023 ( .A1(n14811), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10346) );
  OAI21_X1 U13024 ( .B1(n14737), .B2(n14811), .A(n10346), .ZN(P1_U3528) );
  INV_X1 U13025 ( .A(n10347), .ZN(n13128) );
  NAND2_X1 U13026 ( .A1(n10350), .A2(n10348), .ZN(n10349) );
  OAI21_X1 U13027 ( .B1(n10350), .B2(n13128), .A(n10349), .ZN(n10352) );
  NAND3_X1 U13028 ( .A1(n10353), .A2(n10352), .A3(n10351), .ZN(n10355) );
  MUX2_X1 U13029 ( .A(n10446), .B(P3_REG2_REG_0__SCAN_IN), .S(n15004), .Z(
        n10357) );
  OR2_X1 U13030 ( .A1(n10355), .A2(n12675), .ZN(n11500) );
  NOR2_X2 U13031 ( .A1(n11500), .A2(n15026), .ZN(n12994) );
  INV_X1 U13032 ( .A(n12994), .ZN(n12847) );
  INV_X1 U13033 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10394) );
  OAI22_X1 U13034 ( .A1(n12847), .A2(n12529), .B1(n14580), .B2(n10394), .ZN(
        n10356) );
  OR2_X1 U13035 ( .A1(n10357), .A2(n10356), .ZN(P3_U3233) );
  INV_X1 U13036 ( .A(n10358), .ZN(n10360) );
  OAI222_X1 U13037 ( .A1(P2_U3088), .A2(n10684), .B1(n13800), .B2(n10360), 
        .C1(n15054), .C2(n13803), .ZN(P2_U3315) );
  INV_X1 U13038 ( .A(n10657), .ZN(n10361) );
  OAI222_X1 U13039 ( .A1(P1_U3086), .A2(n10361), .B1(n14534), .B2(n10360), 
        .C1(n10359), .C2(n14528), .ZN(P1_U3343) );
  OAI22_X1 U13040 ( .A1(n13262), .A2(n12096), .B1(n10364), .B2(n13272), .ZN(
        n10365) );
  NAND3_X1 U13041 ( .A1(n10362), .A2(n7331), .A3(n10365), .ZN(n10371) );
  OAI21_X1 U13042 ( .B1(n13276), .B2(n10755), .A(n10366), .ZN(n10367) );
  INV_X1 U13043 ( .A(n10367), .ZN(n10370) );
  INV_X1 U13044 ( .A(n13277), .ZN(n13265) );
  AOI22_X1 U13045 ( .A1(n13265), .A2(n13293), .B1(n13261), .B2(n13291), .ZN(
        n10369) );
  NAND2_X1 U13046 ( .A1(n13281), .A2(n12102), .ZN(n10368) );
  AND4_X1 U13047 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        n10372) );
  OAI21_X1 U13048 ( .B1(n10373), .B2(n13272), .A(n10372), .ZN(P2_U3199) );
  INV_X1 U13049 ( .A(n10382), .ZN(n10374) );
  AOI211_X1 U13050 ( .C1(n10376), .C2(n10375), .A(n13272), .B(n10374), .ZN(
        n10381) );
  INV_X1 U13051 ( .A(n12087), .ZN(n15202) );
  AOI22_X1 U13052 ( .A1(n13261), .A2(n13293), .B1(n15202), .B2(n13281), .ZN(
        n10379) );
  AOI22_X1 U13053 ( .A1(n13240), .A2(n10377), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10378) );
  OAI211_X1 U13054 ( .C1(n10452), .C2(n13277), .A(n10379), .B(n10378), .ZN(
        n10380) );
  OR2_X1 U13055 ( .A1(n10381), .A2(n10380), .ZN(P2_U3190) );
  OAI21_X1 U13056 ( .B1(n10387), .B2(n10382), .A(n10362), .ZN(n10390) );
  AOI22_X1 U13057 ( .A1(n13294), .A2(n13542), .B1(n13544), .B2(n13292), .ZN(
        n10430) );
  INV_X1 U13058 ( .A(n10430), .ZN(n10383) );
  AOI22_X1 U13059 ( .A1(n13251), .A2(n10383), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10385) );
  NAND2_X1 U13060 ( .A1(n13281), .A2(n12095), .ZN(n10384) );
  OAI211_X1 U13061 ( .C1(n13276), .C2(n10698), .A(n10385), .B(n10384), .ZN(
        n10389) );
  NOR4_X1 U13062 ( .A1(n10387), .A2(n13262), .A3(n10386), .A4(n12088), .ZN(
        n10388) );
  AOI211_X1 U13063 ( .C1(n9485), .C2(n10390), .A(n10389), .B(n10388), .ZN(
        n10391) );
  INV_X1 U13064 ( .A(n10391), .ZN(P2_U3202) );
  INV_X1 U13065 ( .A(n12464), .ZN(n12438) );
  NAND2_X1 U13066 ( .A1(n12438), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10609) );
  INV_X1 U13067 ( .A(n10609), .ZN(n10407) );
  INV_X1 U13068 ( .A(n12449), .ZN(n12471) );
  OAI22_X1 U13069 ( .A1(n12497), .A2(n12471), .B1(n12529), .B2(n12459), .ZN(
        n10392) );
  AOI21_X1 U13070 ( .B1(n12463), .B2(n12705), .A(n10392), .ZN(n10393) );
  OAI21_X1 U13071 ( .B1(n10407), .B2(n10394), .A(n10393), .ZN(P3_U3172) );
  INV_X1 U13072 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10406) );
  INV_X1 U13073 ( .A(n14985), .ZN(n10397) );
  NAND3_X1 U13074 ( .A1(n10397), .A2(n6779), .A3(n10396), .ZN(n10398) );
  OAI211_X1 U13075 ( .C1(n10400), .C2(n14990), .A(n10399), .B(n10398), .ZN(
        n10401) );
  NAND2_X1 U13076 ( .A1(n10401), .A2(n12449), .ZN(n10405) );
  OAI22_X1 U13077 ( .A1(n12455), .A2(n10402), .B1(n12459), .B2(n7939), .ZN(
        n10403) );
  AOI21_X1 U13078 ( .B1(n6439), .B2(n6657), .A(n10403), .ZN(n10404) );
  OAI211_X1 U13079 ( .C1(n10407), .C2(n10406), .A(n10405), .B(n10404), .ZN(
        P3_U3162) );
  INV_X1 U13080 ( .A(n10408), .ZN(n10449) );
  AOI22_X1 U13081 ( .A1(n10851), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10409), .ZN(n10410) );
  OAI21_X1 U13082 ( .B1(n10449), .B2(n14534), .A(n10410), .ZN(P1_U3342) );
  XOR2_X1 U13083 ( .A(n10412), .B(n10411), .Z(n10415) );
  AOI22_X1 U13084 ( .A1(n14653), .A2(n14738), .B1(n10489), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10414) );
  INV_X1 U13085 ( .A(n13975), .ZN(n10490) );
  INV_X1 U13086 ( .A(n13974), .ZN(n10491) );
  AOI22_X1 U13087 ( .A1(n10490), .A2(n14740), .B1(n10491), .B2(n6651), .ZN(
        n10413) );
  OAI211_X1 U13088 ( .C1(n10415), .C2(n14699), .A(n10414), .B(n10413), .ZN(
        P1_U3222) );
  OAI222_X1 U13089 ( .A1(n12808), .A2(P3_U3151), .B1(n13142), .B2(n10417), 
        .C1(n13140), .C2(n10416), .ZN(P3_U3276) );
  OR2_X1 U13090 ( .A1(n13295), .A2(n12073), .ZN(n10418) );
  NAND2_X1 U13091 ( .A1(n10419), .A2(n10418), .ZN(n10451) );
  XNOR2_X2 U13092 ( .A(n12087), .B(n13294), .ZN(n12298) );
  NAND2_X1 U13093 ( .A1(n12088), .A2(n12087), .ZN(n10420) );
  XNOR2_X1 U13094 ( .A(n12095), .B(n13293), .ZN(n12301) );
  INV_X1 U13095 ( .A(n12301), .ZN(n10429) );
  OAI21_X1 U13096 ( .B1(n10421), .B2(n10429), .A(n10745), .ZN(n10693) );
  AOI21_X1 U13097 ( .B1(n10458), .B2(n12095), .A(n13620), .ZN(n10422) );
  AND2_X1 U13098 ( .A1(n10422), .A2(n10754), .ZN(n10700) );
  INV_X1 U13099 ( .A(n12298), .ZN(n10426) );
  NAND2_X1 U13100 ( .A1(n10423), .A2(n12296), .ZN(n10425) );
  OR2_X1 U13101 ( .A1(n10736), .A2(n13295), .ZN(n10424) );
  NAND2_X1 U13102 ( .A1(n15202), .A2(n12088), .ZN(n10427) );
  XNOR2_X1 U13103 ( .A(n10747), .B(n10429), .ZN(n10431) );
  OAI21_X1 U13104 ( .B1(n10431), .B2(n11543), .A(n10430), .ZN(n10696) );
  AOI211_X1 U13105 ( .C1(n14623), .C2(n10693), .A(n10700), .B(n10696), .ZN(
        n10574) );
  AOI22_X1 U13106 ( .A1(n13742), .A2(n12095), .B1(n14920), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n10432) );
  OAI21_X1 U13107 ( .B1(n10574), .B2(n14920), .A(n10432), .ZN(P2_U3503) );
  INV_X1 U13108 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10735) );
  OAI22_X1 U13109 ( .A1(n13199), .A2(n10434), .B1(n10433), .B2(n10735), .ZN(
        n10441) );
  INV_X1 U13110 ( .A(n13262), .ZN(n13270) );
  AOI22_X1 U13111 ( .A1(n13270), .A2(n6734), .B1(n9485), .B2(n10435), .ZN(
        n10439) );
  INV_X1 U13112 ( .A(n10436), .ZN(n10438) );
  NOR3_X1 U13113 ( .A1(n10439), .A2(n10438), .A3(n10437), .ZN(n10440) );
  AOI211_X1 U13114 ( .C1(n12073), .C2(n13281), .A(n10441), .B(n10440), .ZN(
        n10442) );
  OAI21_X1 U13115 ( .B1(n10443), .B2(n13272), .A(n10442), .ZN(P2_U3209) );
  INV_X1 U13116 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10444) );
  NOR2_X1 U13117 ( .A1(n15039), .A2(n10444), .ZN(n10445) );
  AOI21_X1 U13118 ( .B1(n15039), .B2(n10446), .A(n10445), .ZN(n10447) );
  OAI21_X1 U13119 ( .B1(n12529), .B2(n13097), .A(n10447), .ZN(P3_U3390) );
  INV_X1 U13120 ( .A(n11122), .ZN(n10690) );
  OAI222_X1 U13121 ( .A1(P2_U3088), .A2(n10690), .B1(n13800), .B2(n10449), 
        .C1(n10448), .C2(n13803), .ZN(P2_U3314) );
  OAI21_X1 U13122 ( .B1(n10451), .B2(n12298), .A(n10450), .ZN(n15208) );
  INV_X1 U13123 ( .A(n15208), .ZN(n10461) );
  INV_X1 U13124 ( .A(n10088), .ZN(n14912) );
  OAI22_X1 U13125 ( .A1(n12096), .A2(n13632), .B1(n10452), .B2(n13630), .ZN(
        n10456) );
  XNOR2_X1 U13126 ( .A(n12298), .B(n10453), .ZN(n10454) );
  NOR2_X1 U13127 ( .A1(n10454), .A2(n11543), .ZN(n10455) );
  AOI211_X1 U13128 ( .C1(n14912), .C2(n15208), .A(n10456), .B(n10455), .ZN(
        n15205) );
  INV_X1 U13129 ( .A(n10457), .ZN(n10459) );
  AOI21_X1 U13130 ( .B1(n15202), .B2(n10459), .A(n6921), .ZN(n15199) );
  AOI22_X1 U13131 ( .A1(n15199), .A2(n13639), .B1(n14889), .B2(n15202), .ZN(
        n10460) );
  OAI211_X1 U13132 ( .C1(n10461), .C2(n14903), .A(n15205), .B(n10460), .ZN(
        n10468) );
  NAND2_X1 U13133 ( .A1(n10468), .A2(n14922), .ZN(n10462) );
  OAI21_X1 U13134 ( .B1(n14922), .B2(n15178), .A(n10462), .ZN(P2_U3502) );
  NAND2_X1 U13135 ( .A1(n14877), .A2(n10463), .ZN(n10464) );
  NOR2_X1 U13136 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  NAND2_X1 U13137 ( .A1(n10468), .A2(n14915), .ZN(n10469) );
  OAI21_X1 U13138 ( .B1(n14915), .B2(n9062), .A(n10469), .ZN(P2_U3439) );
  MUX2_X1 U13139 ( .A(n10470), .B(P1_REG2_REG_12__SCAN_IN), .S(n10657), .Z(
        n10475) );
  NAND2_X1 U13140 ( .A1(n10476), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10471) );
  NAND2_X1 U13141 ( .A1(n10472), .A2(n10471), .ZN(n10474) );
  OR2_X1 U13142 ( .A1(n10474), .A2(n10475), .ZN(n10659) );
  INV_X1 U13143 ( .A(n10659), .ZN(n10473) );
  AOI21_X1 U13144 ( .B1(n10475), .B2(n10474), .A(n10473), .ZN(n10486) );
  NOR2_X1 U13145 ( .A1(n10476), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10477) );
  MUX2_X1 U13146 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n8356), .S(n10657), .Z(
        n10478) );
  OAI21_X1 U13147 ( .B1(n10479), .B2(n10477), .A(n10478), .ZN(n10654) );
  INV_X1 U13148 ( .A(n10654), .ZN(n10481) );
  NOR3_X1 U13149 ( .A1(n10479), .A2(n10478), .A3(n10477), .ZN(n10480) );
  OAI21_X1 U13150 ( .B1(n10481), .B2(n10480), .A(n14194), .ZN(n10485) );
  INV_X1 U13151 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10482) );
  NAND2_X1 U13152 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n11871)
         );
  OAI21_X1 U13153 ( .B1(n14199), .B2(n10482), .A(n11871), .ZN(n10483) );
  AOI21_X1 U13154 ( .B1(n10657), .B2(n14722), .A(n10483), .ZN(n10484) );
  OAI211_X1 U13155 ( .C1(n10486), .C2(n14190), .A(n10485), .B(n10484), .ZN(
        P1_U3255) );
  XOR2_X1 U13156 ( .A(n10488), .B(n10487), .Z(n10494) );
  AOI22_X1 U13157 ( .A1(n14653), .A2(n10727), .B1(n10489), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13158 ( .A1(n10491), .A2(n6450), .B1(n10490), .B2(n14038), .ZN(
        n10492) );
  OAI211_X1 U13159 ( .C1(n10494), .C2(n14699), .A(n10493), .B(n10492), .ZN(
        P1_U3237) );
  OAI21_X1 U13160 ( .B1(n10496), .B2(n12495), .A(n10495), .ZN(n10831) );
  OAI211_X1 U13161 ( .C1(n10498), .C2(n7944), .A(n14991), .B(n10497), .ZN(
        n10500) );
  AOI22_X1 U13162 ( .A1(n14987), .A2(n14989), .B1(n12704), .B2(n14988), .ZN(
        n10499) );
  NAND2_X1 U13163 ( .A1(n10500), .A2(n10499), .ZN(n10826) );
  AOI21_X1 U13164 ( .B1(n15032), .B2(n10831), .A(n10826), .ZN(n10505) );
  AOI22_X1 U13165 ( .A1(n8048), .A2(n10584), .B1(n15049), .B2(
        P3_REG1_REG_3__SCAN_IN), .ZN(n10501) );
  OAI21_X1 U13166 ( .B1(n10505), .B2(n15049), .A(n10501), .ZN(P3_U3462) );
  INV_X1 U13167 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10502) );
  OAI22_X1 U13168 ( .A1(n10828), .A2(n13097), .B1(n15039), .B2(n10502), .ZN(
        n10503) );
  INV_X1 U13169 ( .A(n10503), .ZN(n10504) );
  OAI21_X1 U13170 ( .B1(n10505), .B2(n15037), .A(n10504), .ZN(P3_U3399) );
  OAI21_X1 U13171 ( .B1(n10507), .B2(n12534), .A(n10506), .ZN(n15012) );
  INV_X1 U13172 ( .A(n15012), .ZN(n10516) );
  NOR2_X1 U13173 ( .A1(n14996), .A2(n10849), .ZN(n10622) );
  INV_X1 U13174 ( .A(n10622), .ZN(n10508) );
  NOR2_X1 U13175 ( .A1(n15004), .A2(n10508), .ZN(n14999) );
  INV_X1 U13176 ( .A(n14999), .ZN(n11474) );
  NAND2_X1 U13177 ( .A1(n10606), .A2(n15015), .ZN(n15009) );
  NOR2_X1 U13178 ( .A1(n15009), .A2(n12675), .ZN(n10513) );
  XNOR2_X1 U13179 ( .A(n10509), .B(n12534), .ZN(n10512) );
  OAI22_X1 U13180 ( .A1(n6618), .A2(n12956), .B1(n10629), .B2(n12958), .ZN(
        n10510) );
  AOI21_X1 U13181 ( .B1(n15012), .B2(n15029), .A(n10510), .ZN(n10511) );
  OAI21_X1 U13182 ( .B1(n12954), .B2(n10512), .A(n10511), .ZN(n15010) );
  AOI211_X1 U13183 ( .C1(n14998), .C2(P3_REG3_REG_2__SCAN_IN), .A(n10513), .B(
        n15010), .ZN(n10514) );
  MUX2_X1 U13184 ( .A(n10136), .B(n10514), .S(n15002), .Z(n10515) );
  OAI21_X1 U13185 ( .B1(n10516), .B2(n11474), .A(n10515), .ZN(P3_U3231) );
  NAND2_X1 U13186 ( .A1(n10518), .A2(n12062), .ZN(n14882) );
  NAND4_X1 U13187 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n14877), .ZN(
        n10522) );
  OR2_X1 U13188 ( .A1(n12286), .A2(n12334), .ZN(n10694) );
  INV_X1 U13189 ( .A(n10694), .ZN(n15209) );
  NAND2_X1 U13190 ( .A1(n15210), .A2(n15209), .ZN(n11518) );
  OAI21_X1 U13191 ( .B1(n13649), .B2(n12331), .A(n13641), .ZN(n10526) );
  AND2_X1 U13192 ( .A1(n12059), .A2(n10523), .ZN(n14884) );
  NOR2_X1 U13193 ( .A1(n14912), .A2(n13635), .ZN(n10525) );
  OAI22_X1 U13194 ( .A1(n14882), .A2(n10525), .B1(n10524), .B2(n13632), .ZN(
        n14883) );
  AOI22_X1 U13195 ( .A1(n10526), .A2(n14884), .B1(n15210), .B2(n14883), .ZN(
        n10531) );
  OAI22_X1 U13196 ( .A1(n15210), .A2(n10528), .B1(n10527), .B2(n13651), .ZN(
        n10529) );
  INV_X1 U13197 ( .A(n10529), .ZN(n10530) );
  OAI211_X1 U13198 ( .C1(n14882), .C2(n11518), .A(n10531), .B(n10530), .ZN(
        P2_U3265) );
  INV_X1 U13199 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10533) );
  INV_X1 U13200 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10532) );
  MUX2_X1 U13201 ( .A(n10533), .B(n10532), .S(n12799), .Z(n10902) );
  XNOR2_X1 U13202 ( .A(n10902), .B(n10908), .ZN(n10540) );
  MUX2_X1 U13203 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12799), .Z(n10537) );
  OR2_X1 U13204 ( .A1(n10537), .A2(n14932), .ZN(n10538) );
  OAI22_X1 U13205 ( .A1(n10536), .A2(n10535), .B1(n10534), .B2(n10552), .ZN(
        n14926) );
  XOR2_X1 U13206 ( .A(n14932), .B(n10537), .Z(n14925) );
  NAND2_X1 U13207 ( .A1(n14926), .A2(n14925), .ZN(n14924) );
  NAND2_X1 U13208 ( .A1(n10538), .A2(n14924), .ZN(n10539) );
  NAND2_X1 U13209 ( .A1(n10540), .A2(n10539), .ZN(n10903) );
  OAI21_X1 U13210 ( .B1(n10540), .B2(n10539), .A(n10903), .ZN(n10565) );
  NAND2_X1 U13211 ( .A1(n10552), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10541) );
  INV_X1 U13212 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n14928) );
  INV_X1 U13213 ( .A(n10545), .ZN(n10543) );
  MUX2_X1 U13214 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n10533), .S(n10908), .Z(
        n10547) );
  INV_X1 U13215 ( .A(n10547), .ZN(n10549) );
  INV_X1 U13216 ( .A(n10910), .ZN(n10548) );
  AOI21_X1 U13217 ( .B1(n10550), .B2(n10549), .A(n10548), .ZN(n10563) );
  NOR2_X1 U13218 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10551), .ZN(n12380) );
  MUX2_X1 U13219 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n10532), .S(n10908), .Z(
        n10557) );
  NAND2_X1 U13220 ( .A1(n10552), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10553) );
  NAND2_X1 U13221 ( .A1(n10554), .A2(n10553), .ZN(n10555) );
  INV_X1 U13222 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15044) );
  INV_X1 U13223 ( .A(n10557), .ZN(n10559) );
  NAND2_X1 U13224 ( .A1(n10559), .A2(n10558), .ZN(n10560) );
  AOI21_X1 U13225 ( .B1(n10896), .B2(n10560), .A(n14977), .ZN(n10561) );
  AOI211_X1 U13226 ( .C1(n14923), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n12380), .B(
        n10561), .ZN(n10562) );
  OAI21_X1 U13227 ( .B1(n10563), .B2(n14983), .A(n10562), .ZN(n10564) );
  AOI21_X1 U13228 ( .B1(n14936), .B2(n10565), .A(n10564), .ZN(n10566) );
  OAI21_X1 U13229 ( .B1(n10908), .B2(n14966), .A(n10566), .ZN(P3_U3190) );
  INV_X1 U13230 ( .A(n14915), .ZN(n14913) );
  NAND2_X1 U13231 ( .A1(n14915), .A2(n14889), .ZN(n13780) );
  INV_X1 U13232 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10567) );
  OAI22_X1 U13233 ( .A1(n13780), .A2(n10706), .B1(n14915), .B2(n10567), .ZN(
        n10568) );
  INV_X1 U13234 ( .A(n10568), .ZN(n10569) );
  OAI21_X1 U13235 ( .B1(n10570), .B2(n14913), .A(n10569), .ZN(P2_U3433) );
  INV_X1 U13236 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10571) );
  OAI22_X1 U13237 ( .A1(n13780), .A2(n12097), .B1(n14915), .B2(n10571), .ZN(
        n10572) );
  INV_X1 U13238 ( .A(n10572), .ZN(n10573) );
  OAI21_X1 U13239 ( .B1(n10574), .B2(n14913), .A(n10573), .ZN(P2_U3442) );
  INV_X1 U13240 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10575) );
  OAI22_X1 U13241 ( .A1(n13780), .A2(n10736), .B1(n14915), .B2(n10575), .ZN(
        n10576) );
  INV_X1 U13242 ( .A(n10576), .ZN(n10577) );
  OAI21_X1 U13243 ( .B1(n10578), .B2(n14913), .A(n10577), .ZN(P2_U3436) );
  INV_X1 U13244 ( .A(n10579), .ZN(n10580) );
  AOI211_X1 U13245 ( .C1(n10582), .C2(n10581), .A(n12471), .B(n10580), .ZN(
        n10588) );
  AOI22_X1 U13246 ( .A1(n6439), .A2(n14989), .B1(n12463), .B2(n12704), .ZN(
        n10586) );
  INV_X1 U13247 ( .A(n12459), .ZN(n12469) );
  AOI21_X1 U13248 ( .B1(n12469), .B2(n10584), .A(n10583), .ZN(n10585) );
  OAI211_X1 U13249 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12438), .A(n10586), .B(
        n10585), .ZN(n10587) );
  OR2_X1 U13250 ( .A1(n10588), .A2(n10587), .ZN(P3_U3158) );
  MUX2_X1 U13251 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11512), .S(n10684), .Z(
        n10593) );
  AOI21_X1 U13252 ( .B1(n10590), .B2(n11373), .A(n10589), .ZN(n10592) );
  INV_X1 U13253 ( .A(n10679), .ZN(n10591) );
  AOI21_X1 U13254 ( .B1(n10593), .B2(n10592), .A(n10591), .ZN(n10603) );
  NOR2_X1 U13255 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10594), .ZN(n11303) );
  NOR2_X1 U13256 ( .A1(n14820), .A2(n10684), .ZN(n10595) );
  AOI211_X1 U13257 ( .C1(n14859), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n11303), 
        .B(n10595), .ZN(n10602) );
  AOI21_X1 U13258 ( .B1(n10597), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10596), 
        .ZN(n10599) );
  MUX2_X1 U13259 ( .A(n9213), .B(P2_REG1_REG_12__SCAN_IN), .S(n10684), .Z(
        n10598) );
  NOR2_X1 U13260 ( .A1(n10599), .A2(n10598), .ZN(n10600) );
  AND2_X1 U13261 ( .A1(n10599), .A2(n10598), .ZN(n10683) );
  OAI21_X1 U13262 ( .B1(n10600), .B2(n10683), .A(n14868), .ZN(n10601) );
  OAI211_X1 U13263 ( .C1(n10603), .C2(n11825), .A(n10602), .B(n10601), .ZN(
        P2_U3226) );
  XOR2_X1 U13264 ( .A(n10604), .B(n10605), .Z(n10611) );
  INV_X1 U13265 ( .A(n6439), .ZN(n12467) );
  AOI22_X1 U13266 ( .A1(n12463), .A2(n10616), .B1(n12469), .B2(n10606), .ZN(
        n10607) );
  OAI21_X1 U13267 ( .B1(n12467), .B2(n6618), .A(n10607), .ZN(n10608) );
  AOI21_X1 U13268 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10609), .A(n10608), .ZN(
        n10610) );
  OAI21_X1 U13269 ( .B1(n10611), .B2(n12471), .A(n10610), .ZN(P3_U3177) );
  INV_X1 U13270 ( .A(n10612), .ZN(n10613) );
  AOI21_X1 U13271 ( .B1(n10615), .B2(n10614), .A(n10613), .ZN(n10621) );
  AOI22_X1 U13272 ( .A1(n6439), .A2(n10616), .B1(n12463), .B2(n12703), .ZN(
        n10618) );
  OAI211_X1 U13273 ( .C1(n12459), .C2(n10675), .A(n10618), .B(n10617), .ZN(
        n10619) );
  AOI21_X1 U13274 ( .B1(n10633), .B2(n12464), .A(n10619), .ZN(n10620) );
  OAI21_X1 U13275 ( .B1(n10621), .B2(n12471), .A(n10620), .ZN(P3_U3170) );
  NOR2_X1 U13276 ( .A1(n15029), .A2(n10622), .ZN(n10623) );
  OAI21_X1 U13277 ( .B1(n10625), .B2(n12547), .A(n10624), .ZN(n10670) );
  INV_X1 U13278 ( .A(n10670), .ZN(n10636) );
  OAI211_X1 U13279 ( .C1(n10628), .C2(n10627), .A(n10626), .B(n14991), .ZN(
        n10632) );
  OAI22_X1 U13280 ( .A1(n11002), .A2(n12958), .B1(n10629), .B2(n12956), .ZN(
        n10630) );
  INV_X1 U13281 ( .A(n10630), .ZN(n10631) );
  AND2_X1 U13282 ( .A1(n10632), .A2(n10631), .ZN(n10668) );
  MUX2_X1 U13283 ( .A(n10176), .B(n10668), .S(n15002), .Z(n10635) );
  AOI22_X1 U13284 ( .A1(n12994), .A2(n10672), .B1(n14998), .B2(n10633), .ZN(
        n10634) );
  OAI211_X1 U13285 ( .C1(n12997), .C2(n10636), .A(n10635), .B(n10634), .ZN(
        P3_U3229) );
  OAI222_X1 U13286 ( .A1(P1_U3086), .A2(n11207), .B1(n14534), .B2(n10637), 
        .C1(n15067), .C2(n14528), .ZN(P1_U3341) );
  OAI222_X1 U13287 ( .A1(n13803), .A2(n10638), .B1(n13800), .B2(n10637), .C1(
        n11524), .C2(P2_U3088), .ZN(P2_U3313) );
  OAI222_X1 U13288 ( .A1(n10641), .A2(P3_U3151), .B1(n13142), .B2(n10640), 
        .C1(n13140), .C2(n10639), .ZN(P3_U3275) );
  INV_X1 U13289 ( .A(n12115), .ZN(n12117) );
  INV_X1 U13290 ( .A(n10642), .ZN(n10643) );
  AOI21_X1 U13291 ( .B1(n10819), .B2(n10643), .A(n13272), .ZN(n10646) );
  NOR3_X1 U13292 ( .A1(n10644), .A2(n12108), .A3(n13262), .ZN(n10645) );
  OAI21_X1 U13293 ( .B1(n10646), .B2(n10645), .A(n10869), .ZN(n10650) );
  INV_X1 U13294 ( .A(n10788), .ZN(n10648) );
  AND2_X1 U13295 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14832) );
  OAI22_X1 U13296 ( .A1(n13278), .A2(n12123), .B1(n12108), .B2(n13277), .ZN(
        n10647) );
  AOI211_X1 U13297 ( .C1(n13240), .C2(n10648), .A(n14832), .B(n10647), .ZN(
        n10649) );
  OAI211_X1 U13298 ( .C1(n12117), .C2(n13258), .A(n10650), .B(n10649), .ZN(
        P2_U3185) );
  INV_X1 U13299 ( .A(n14168), .ZN(n11853) );
  INV_X1 U13300 ( .A(n10651), .ZN(n10653) );
  OAI222_X1 U13301 ( .A1(P1_U3086), .A2(n11853), .B1(n14534), .B2(n10653), 
        .C1(n10652), .C2(n14528), .ZN(P1_U3339) );
  INV_X1 U13302 ( .A(n11832), .ZN(n11609) );
  OAI222_X1 U13303 ( .A1(n13803), .A2(n15113), .B1(n13800), .B2(n10653), .C1(
        n11609), .C2(P2_U3088), .ZN(P2_U3311) );
  OAI21_X1 U13304 ( .B1(n10657), .B2(P1_REG1_REG_12__SCAN_IN), .A(n10654), 
        .ZN(n10656) );
  INV_X1 U13305 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11779) );
  MUX2_X1 U13306 ( .A(n11779), .B(P1_REG1_REG_13__SCAN_IN), .S(n10851), .Z(
        n10655) );
  AOI211_X1 U13307 ( .C1(n10656), .C2(n10655), .A(n14729), .B(n10850), .ZN(
        n10667) );
  OR2_X1 U13308 ( .A1(n10657), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10658) );
  NAND2_X1 U13309 ( .A1(n10659), .A2(n10658), .ZN(n10662) );
  MUX2_X1 U13310 ( .A(n8385), .B(P1_REG2_REG_13__SCAN_IN), .S(n10851), .Z(
        n10661) );
  INV_X1 U13311 ( .A(n10853), .ZN(n10660) );
  AOI211_X1 U13312 ( .C1(n10662), .C2(n10661), .A(n14190), .B(n10660), .ZN(
        n10666) );
  NAND2_X1 U13313 ( .A1(n14722), .A2(n10851), .ZN(n10663) );
  NAND2_X1 U13314 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11947)
         );
  OAI211_X1 U13315 ( .C1(n10664), .C2(n14199), .A(n10663), .B(n11947), .ZN(
        n10665) );
  OR3_X1 U13316 ( .A1(n10667), .A2(n10666), .A3(n10665), .ZN(P1_U3256) );
  INV_X1 U13317 ( .A(n10668), .ZN(n10669) );
  AOI21_X1 U13318 ( .B1(n15032), .B2(n10670), .A(n10669), .ZN(n10678) );
  AOI22_X1 U13319 ( .A1(n8048), .A2(n10672), .B1(n15049), .B2(
        P3_REG1_REG_4__SCAN_IN), .ZN(n10673) );
  OAI21_X1 U13320 ( .B1(n10678), .B2(n15049), .A(n10673), .ZN(P3_U3463) );
  INV_X1 U13321 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10674) );
  OAI22_X1 U13322 ( .A1(n10675), .A2(n13097), .B1(n15039), .B2(n10674), .ZN(
        n10676) );
  INV_X1 U13323 ( .A(n10676), .ZN(n10677) );
  OAI21_X1 U13324 ( .B1(n10678), .B2(n15037), .A(n10677), .ZN(P3_U3402) );
  XNOR2_X1 U13325 ( .A(n11122), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n10682) );
  INV_X1 U13326 ( .A(n10684), .ZN(n10680) );
  NOR2_X1 U13327 ( .A1(n10681), .A2(n10682), .ZN(n11119) );
  AOI211_X1 U13328 ( .C1(n10682), .C2(n10681), .A(n11825), .B(n11119), .ZN(
        n10692) );
  AOI21_X1 U13329 ( .B1(n9213), .B2(n10684), .A(n10683), .ZN(n10687) );
  INV_X1 U13330 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10685) );
  MUX2_X1 U13331 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n10685), .S(n11122), .Z(
        n10686) );
  NAND2_X1 U13332 ( .A1(n10687), .A2(n10686), .ZN(n11125) );
  OAI211_X1 U13333 ( .C1(n10687), .C2(n10686), .A(n11125), .B(n14868), .ZN(
        n10689) );
  AND2_X1 U13334 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n11438) );
  AOI21_X1 U13335 ( .B1(n14859), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n11438), 
        .ZN(n10688) );
  OAI211_X1 U13336 ( .C1(n14820), .C2(n10690), .A(n10689), .B(n10688), .ZN(
        n10691) );
  OR2_X1 U13337 ( .A1(n10692), .A2(n10691), .ZN(P2_U3227) );
  INV_X1 U13338 ( .A(n10693), .ZN(n10703) );
  NAND2_X1 U13339 ( .A1(n10088), .A2(n10694), .ZN(n10695) );
  INV_X1 U13340 ( .A(n10696), .ZN(n10697) );
  MUX2_X1 U13341 ( .A(n9879), .B(n10697), .S(n15210), .Z(n10702) );
  OAI22_X1 U13342 ( .A1(n13603), .A2(n12097), .B1(n10698), .B2(n13651), .ZN(
        n10699) );
  AOI21_X1 U13343 ( .B1(n13658), .B2(n10700), .A(n10699), .ZN(n10701) );
  OAI211_X1 U13344 ( .C1(n10703), .C2(n13627), .A(n10702), .B(n10701), .ZN(
        P2_U3261) );
  MUX2_X1 U13345 ( .A(n9880), .B(n10704), .S(n15210), .Z(n10710) );
  OAI22_X1 U13346 ( .A1(n13603), .A2(n10706), .B1(n10705), .B2(n13651), .ZN(
        n10707) );
  AOI21_X1 U13347 ( .B1(n13658), .B2(n10708), .A(n10707), .ZN(n10709) );
  OAI211_X1 U13348 ( .C1(n10711), .C2(n13627), .A(n10710), .B(n10709), .ZN(
        P2_U3264) );
  OAI21_X1 U13349 ( .B1(n10714), .B2(P1_D_REG_0__SCAN_IN), .A(n10712), .ZN(
        n10716) );
  OR2_X1 U13350 ( .A1(n10714), .A2(n10713), .ZN(n10715) );
  NAND2_X1 U13351 ( .A1(n10716), .A2(n10715), .ZN(n10793) );
  NAND2_X1 U13352 ( .A1(n14039), .A2(n10718), .ZN(n11442) );
  NAND2_X1 U13353 ( .A1(n10719), .A2(n11442), .ZN(n11445) );
  OR2_X1 U13354 ( .A1(n9679), .A2(n14738), .ZN(n10720) );
  INV_X1 U13355 ( .A(n10724), .ZN(n10721) );
  NAND2_X1 U13356 ( .A1(n10722), .A2(n10721), .ZN(n10922) );
  OAI21_X1 U13357 ( .B1(n10722), .B2(n10721), .A(n10922), .ZN(n10806) );
  INV_X1 U13358 ( .A(n10806), .ZN(n10729) );
  INV_X1 U13359 ( .A(n10723), .ZN(n10725) );
  OAI21_X1 U13360 ( .B1(n10725), .B2(n10724), .A(n10930), .ZN(n10726) );
  AOI222_X1 U13361 ( .A1(n14489), .A2(n10726), .B1(n14038), .B2(n14739), .C1(
        n6450), .C2(n14483), .ZN(n10809) );
  AOI211_X1 U13362 ( .C1(n10727), .C2(n11447), .A(n14355), .B(n10926), .ZN(
        n10802) );
  AOI21_X1 U13363 ( .B1(n14793), .B2(n10727), .A(n10802), .ZN(n10728) );
  OAI211_X1 U13364 ( .C1(n14753), .C2(n10729), .A(n10809), .B(n10728), .ZN(
        n10731) );
  NAND2_X1 U13365 ( .A1(n10731), .A2(n14802), .ZN(n10730) );
  OAI21_X1 U13366 ( .B1(n14802), .B2(n8119), .A(n10730), .ZN(P1_U3465) );
  NAND2_X1 U13367 ( .A1(n10731), .A2(n14813), .ZN(n10732) );
  OAI21_X1 U13368 ( .B1(n14813), .B2(n10733), .A(n10732), .ZN(P1_U3530) );
  INV_X1 U13369 ( .A(n10734), .ZN(n10743) );
  OAI22_X1 U13370 ( .A1(n15210), .A2(n9882), .B1(n10735), .B2(n13651), .ZN(
        n10738) );
  NOR2_X1 U13371 ( .A1(n13603), .A2(n10736), .ZN(n10737) );
  AOI211_X1 U13372 ( .C1(n10739), .C2(n13658), .A(n10738), .B(n10737), .ZN(
        n10742) );
  NAND2_X1 U13373 ( .A1(n10740), .A2(n15210), .ZN(n10741) );
  OAI211_X1 U13374 ( .C1(n13627), .C2(n10743), .A(n10742), .B(n10741), .ZN(
        P2_U3263) );
  NAND2_X1 U13375 ( .A1(n12097), .A2(n12096), .ZN(n10744) );
  XNOR2_X1 U13376 ( .A(n12102), .B(n13292), .ZN(n12300) );
  OAI21_X1 U13377 ( .B1(n10746), .B2(n10750), .A(n10761), .ZN(n10841) );
  INV_X1 U13378 ( .A(n10841), .ZN(n10759) );
  OAI22_X1 U13379 ( .A1(n12096), .A2(n13630), .B1(n12108), .B2(n13632), .ZN(
        n10753) );
  NAND2_X1 U13380 ( .A1(n10747), .A2(n12301), .ZN(n10749) );
  NAND2_X1 U13381 ( .A1(n12095), .A2(n12096), .ZN(n10748) );
  XNOR2_X1 U13382 ( .A(n10764), .B(n10750), .ZN(n10751) );
  NOR2_X1 U13383 ( .A1(n10751), .A2(n11543), .ZN(n10752) );
  AOI211_X1 U13384 ( .C1(n14912), .C2(n10841), .A(n10753), .B(n10752), .ZN(
        n10838) );
  MUX2_X1 U13385 ( .A(n9974), .B(n10838), .S(n15210), .Z(n10758) );
  AOI211_X1 U13386 ( .C1(n12102), .C2(n10754), .A(n13620), .B(n10773), .ZN(
        n10840) );
  INV_X1 U13387 ( .A(n12102), .ZN(n12105) );
  OAI22_X1 U13388 ( .A1(n12105), .A2(n13603), .B1(n13651), .B2(n10755), .ZN(
        n10756) );
  AOI21_X1 U13389 ( .B1(n10840), .B2(n13658), .A(n10756), .ZN(n10757) );
  OAI211_X1 U13390 ( .C1(n10759), .C2(n11518), .A(n10758), .B(n10757), .ZN(
        P2_U3260) );
  OR2_X1 U13391 ( .A1(n12102), .A2(n13292), .ZN(n10760) );
  INV_X1 U13392 ( .A(n12303), .ZN(n10766) );
  OAI21_X1 U13393 ( .B1(n10762), .B2(n10766), .A(n10780), .ZN(n10771) );
  INV_X1 U13394 ( .A(n10771), .ZN(n14892) );
  INV_X1 U13395 ( .A(n13292), .ZN(n12104) );
  OAI22_X1 U13396 ( .A1(n12116), .A2(n13632), .B1(n12104), .B2(n13630), .ZN(
        n10770) );
  AND2_X1 U13397 ( .A1(n12102), .A2(n12104), .ZN(n10763) );
  OR2_X1 U13398 ( .A1(n12102), .A2(n12104), .ZN(n10765) );
  NAND2_X1 U13399 ( .A1(n10767), .A2(n10766), .ZN(n10768) );
  AOI21_X1 U13400 ( .B1(n10783), .B2(n10768), .A(n11543), .ZN(n10769) );
  AOI211_X1 U13401 ( .C1(n14912), .C2(n10771), .A(n10770), .B(n10769), .ZN(
        n14891) );
  MUX2_X1 U13402 ( .A(n10772), .B(n14891), .S(n15210), .Z(n10778) );
  INV_X1 U13403 ( .A(n10773), .ZN(n10775) );
  INV_X1 U13404 ( .A(n10787), .ZN(n10774) );
  AOI211_X1 U13405 ( .C1(n14888), .C2(n10775), .A(n13620), .B(n10774), .ZN(
        n14887) );
  OAI22_X1 U13406 ( .A1(n12109), .A2(n13603), .B1(n13651), .B2(n10818), .ZN(
        n10776) );
  AOI21_X1 U13407 ( .B1(n14887), .B2(n13658), .A(n10776), .ZN(n10777) );
  OAI211_X1 U13408 ( .C1(n14892), .C2(n11518), .A(n10778), .B(n10777), .ZN(
        P2_U3259) );
  NAND2_X1 U13409 ( .A1(n12109), .A2(n12108), .ZN(n10779) );
  OAI21_X1 U13410 ( .B1(n10781), .B2(n12305), .A(n10983), .ZN(n10944) );
  INV_X1 U13411 ( .A(n10944), .ZN(n10792) );
  NAND2_X1 U13412 ( .A1(n14888), .A2(n12108), .ZN(n10782) );
  AOI21_X1 U13413 ( .B1(n10784), .B2(n12305), .A(n11543), .ZN(n10786) );
  OAI22_X1 U13414 ( .A1(n12123), .A2(n13632), .B1(n12108), .B2(n13630), .ZN(
        n10785) );
  AOI21_X1 U13415 ( .B1(n10786), .B2(n10987), .A(n10785), .ZN(n10941) );
  MUX2_X1 U13416 ( .A(n10941), .B(n9994), .S(n13649), .Z(n10791) );
  AOI211_X1 U13417 ( .C1(n12115), .C2(n10787), .A(n13620), .B(n7445), .ZN(
        n10943) );
  OAI22_X1 U13418 ( .A1(n12117), .A2(n13603), .B1(n13651), .B2(n10788), .ZN(
        n10789) );
  AOI21_X1 U13419 ( .B1(n10943), .B2(n13658), .A(n10789), .ZN(n10790) );
  OAI211_X1 U13420 ( .C1(n10792), .C2(n13627), .A(n10791), .B(n10790), .ZN(
        P2_U3258) );
  INV_X1 U13421 ( .A(n10793), .ZN(n10794) );
  NAND2_X1 U13422 ( .A1(n10795), .A2(n10794), .ZN(n12022) );
  INV_X2 U13423 ( .A(n14377), .ZN(n14325) );
  OAI22_X1 U13424 ( .A1(n14377), .A2(n10039), .B1(n10796), .B2(n14374), .ZN(
        n10801) );
  AND2_X1 U13425 ( .A1(n9770), .A2(n10797), .ZN(n10798) );
  NOR2_X1 U13426 ( .A1(n14364), .A2(n10799), .ZN(n10800) );
  AOI211_X1 U13427 ( .C1(n10802), .C2(n14357), .A(n10801), .B(n10800), .ZN(
        n10808) );
  INV_X1 U13428 ( .A(n10803), .ZN(n10804) );
  NAND2_X1 U13429 ( .A1(n14377), .A2(n10804), .ZN(n14262) );
  NAND2_X1 U13430 ( .A1(n14377), .A2(n14254), .ZN(n10805) );
  NAND2_X1 U13431 ( .A1(n10806), .A2(n14337), .ZN(n10807) );
  OAI211_X1 U13432 ( .C1(n10809), .C2(n14325), .A(n10808), .B(n10807), .ZN(
        P1_U3291) );
  XOR2_X1 U13433 ( .A(n10810), .B(n10811), .Z(n10816) );
  AOI22_X1 U13434 ( .A1(n6439), .A2(n12704), .B1(n12463), .B2(n12702), .ZN(
        n10813) );
  OAI211_X1 U13435 ( .C1(n12459), .C2(n11014), .A(n10813), .B(n10812), .ZN(
        n10814) );
  AOI21_X1 U13436 ( .B1(n10888), .B2(n12464), .A(n10814), .ZN(n10815) );
  OAI21_X1 U13437 ( .B1(n10816), .B2(n12471), .A(n10815), .ZN(P3_U3167) );
  AOI22_X1 U13438 ( .A1(n13265), .A2(n13292), .B1(n13261), .B2(n13290), .ZN(
        n10817) );
  NAND2_X1 U13439 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13297) );
  OAI211_X1 U13440 ( .C1(n10818), .C2(n13276), .A(n10817), .B(n13297), .ZN(
        n10824) );
  INV_X1 U13441 ( .A(n10819), .ZN(n10820) );
  AOI211_X1 U13442 ( .C1(n10822), .C2(n10821), .A(n13272), .B(n10820), .ZN(
        n10823) );
  AOI211_X1 U13443 ( .C1(n14888), .C2(n13281), .A(n10824), .B(n10823), .ZN(
        n10825) );
  INV_X1 U13444 ( .A(n10825), .ZN(P2_U3211) );
  INV_X1 U13445 ( .A(n10826), .ZN(n10833) );
  OAI22_X1 U13446 ( .A1(n15002), .A2(n10827), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n14580), .ZN(n10830) );
  NOR2_X1 U13447 ( .A1(n12847), .A2(n10828), .ZN(n10829) );
  AOI211_X1 U13448 ( .C1(n10831), .C2(n14599), .A(n10830), .B(n10829), .ZN(
        n10832) );
  OAI21_X1 U13449 ( .B1(n10833), .B2(n15004), .A(n10832), .ZN(P3_U3230) );
  INV_X1 U13450 ( .A(n14721), .ZN(n11854) );
  INV_X1 U13451 ( .A(n10834), .ZN(n10837) );
  OAI222_X1 U13452 ( .A1(P1_U3086), .A2(n11854), .B1(n14534), .B2(n10837), 
        .C1(n10835), .C2(n14528), .ZN(P1_U3338) );
  INV_X1 U13453 ( .A(n13313), .ZN(n13318) );
  OAI222_X1 U13454 ( .A1(P2_U3088), .A2(n13318), .B1(n13800), .B2(n10837), 
        .C1(n10836), .C2(n13803), .ZN(P2_U3310) );
  INV_X1 U13455 ( .A(n10838), .ZN(n10839) );
  AOI211_X1 U13456 ( .C1(n14901), .C2(n10841), .A(n10840), .B(n10839), .ZN(
        n10846) );
  AOI22_X1 U13457 ( .A1(n13742), .A2(n12102), .B1(n14920), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10842) );
  OAI21_X1 U13458 ( .B1(n10846), .B2(n14920), .A(n10842), .ZN(P2_U3504) );
  INV_X1 U13459 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10843) );
  OAI22_X1 U13460 ( .A1(n12105), .A2(n13780), .B1(n14915), .B2(n10843), .ZN(
        n10844) );
  INV_X1 U13461 ( .A(n10844), .ZN(n10845) );
  OAI21_X1 U13462 ( .B1(n10846), .B2(n14913), .A(n10845), .ZN(P2_U3445) );
  OAI222_X1 U13463 ( .A1(n10849), .A2(P3_U3151), .B1(n13142), .B2(n10848), 
        .C1(n13140), .C2(n10847), .ZN(P3_U3274) );
  AOI21_X1 U13464 ( .B1(n10851), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10850), 
        .ZN(n10864) );
  INV_X1 U13465 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11904) );
  NOR3_X1 U13466 ( .A1(n10864), .A2(n11904), .A3(n14729), .ZN(n10855) );
  NAND2_X1 U13467 ( .A1(n10851), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U13468 ( .A1(n10853), .A2(n10852), .ZN(n10858) );
  NOR3_X1 U13469 ( .A1(n10858), .A2(P1_REG2_REG_14__SCAN_IN), .A3(n14190), 
        .ZN(n10854) );
  NOR3_X1 U13470 ( .A1(n10855), .A2(n14722), .A3(n10854), .ZN(n10868) );
  AOI21_X1 U13471 ( .B1(n11207), .B2(P1_REG2_REG_14__SCAN_IN), .A(n10858), 
        .ZN(n10856) );
  NOR2_X1 U13472 ( .A1(n10856), .A2(n14190), .ZN(n10861) );
  MUX2_X1 U13473 ( .A(n11803), .B(P1_REG2_REG_14__SCAN_IN), .S(n11207), .Z(
        n10857) );
  NAND2_X1 U13474 ( .A1(n10858), .A2(n10857), .ZN(n11206) );
  NAND2_X1 U13475 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14646)
         );
  OAI21_X1 U13476 ( .B1(n14199), .B2(n10859), .A(n14646), .ZN(n10860) );
  AOI21_X1 U13477 ( .B1(n10861), .B2(n11206), .A(n10860), .ZN(n10867) );
  INV_X1 U13478 ( .A(n11207), .ZN(n10862) );
  NOR3_X1 U13479 ( .A1(n10864), .A2(P1_REG1_REG_14__SCAN_IN), .A3(n10862), 
        .ZN(n10865) );
  MUX2_X1 U13480 ( .A(n11904), .B(P1_REG1_REG_14__SCAN_IN), .S(n11207), .Z(
        n10863) );
  OAI21_X1 U13481 ( .B1(n10865), .B2(n11204), .A(n14194), .ZN(n10866) );
  OAI211_X1 U13482 ( .C1(n10868), .C2(n11207), .A(n10867), .B(n10866), .ZN(
        P1_U3257) );
  INV_X1 U13483 ( .A(n10869), .ZN(n10872) );
  NOR3_X1 U13484 ( .A1(n10870), .A2(n12116), .A3(n13262), .ZN(n10871) );
  AOI21_X1 U13485 ( .B1(n10872), .B2(n9485), .A(n10871), .ZN(n10880) );
  INV_X1 U13486 ( .A(n10873), .ZN(n10977) );
  NOR2_X1 U13487 ( .A1(n14897), .A2(n13258), .ZN(n10877) );
  AOI22_X1 U13488 ( .A1(n13265), .A2(n13290), .B1(n13261), .B2(n13288), .ZN(
        n10875) );
  OAI211_X1 U13489 ( .C1(n10991), .C2(n13276), .A(n10875), .B(n10874), .ZN(
        n10876) );
  AOI211_X1 U13490 ( .C1(n10977), .C2(n9485), .A(n10877), .B(n10876), .ZN(
        n10878) );
  OAI21_X1 U13491 ( .B1(n10880), .B2(n10879), .A(n10878), .ZN(P2_U3193) );
  INV_X1 U13492 ( .A(n10881), .ZN(n10882) );
  AOI21_X1 U13493 ( .B1(n12552), .B2(n10883), .A(n10882), .ZN(n10884) );
  OAI222_X1 U13494 ( .A1(n12958), .A2(n11025), .B1(n12956), .B2(n10885), .C1(
        n12954), .C2(n10884), .ZN(n11009) );
  INV_X1 U13495 ( .A(n11009), .ZN(n10894) );
  OAI21_X1 U13496 ( .B1(n10887), .B2(n12552), .A(n10886), .ZN(n11010) );
  NOR2_X1 U13497 ( .A1(n12847), .A2(n11014), .ZN(n10892) );
  INV_X1 U13498 ( .A(n10888), .ZN(n10889) );
  OAI22_X1 U13499 ( .A1(n15002), .A2(n10890), .B1(n10889), .B2(n14580), .ZN(
        n10891) );
  AOI211_X1 U13500 ( .C1(n11010), .C2(n14599), .A(n10892), .B(n10891), .ZN(
        n10893) );
  OAI21_X1 U13501 ( .B1(n10894), .B2(n15004), .A(n10893), .ZN(P3_U3228) );
  INV_X1 U13502 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15047) );
  NAND2_X1 U13503 ( .A1(n10908), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10895) );
  AOI21_X1 U13504 ( .B1(n15047), .B2(n10897), .A(n11331), .ZN(n10916) );
  MUX2_X1 U13505 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12799), .Z(n10899) );
  NAND2_X1 U13506 ( .A1(n10898), .A2(n10899), .ZN(n11317) );
  INV_X1 U13507 ( .A(n10899), .ZN(n10900) );
  NAND2_X1 U13508 ( .A1(n10900), .A2(n11330), .ZN(n11315) );
  NAND2_X1 U13509 ( .A1(n11317), .A2(n11315), .ZN(n10905) );
  INV_X1 U13510 ( .A(n10908), .ZN(n10901) );
  NAND2_X1 U13511 ( .A1(n10902), .A2(n10901), .ZN(n10904) );
  XNOR2_X1 U13512 ( .A(n10905), .B(n11318), .ZN(n10907) );
  NAND2_X1 U13513 ( .A1(n14923), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n10906) );
  NAND2_X1 U13514 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11384) );
  OAI211_X1 U13515 ( .C1(n14975), .C2(n10907), .A(n10906), .B(n11384), .ZN(
        n10914) );
  INV_X1 U13516 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U13517 ( .A1(n10908), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10909) );
  AOI21_X1 U13518 ( .B1(n11397), .B2(n10911), .A(n11307), .ZN(n10912) );
  NOR2_X1 U13519 ( .A1(n10912), .A2(n14983), .ZN(n10913) );
  AOI211_X1 U13520 ( .C1(n14954), .C2(n11330), .A(n10914), .B(n10913), .ZN(
        n10915) );
  OAI21_X1 U13521 ( .B1(n10916), .B2(n14977), .A(n10915), .ZN(P3_U3191) );
  INV_X1 U13522 ( .A(n11849), .ZN(n11208) );
  INV_X1 U13523 ( .A(n10917), .ZN(n10919) );
  OAI222_X1 U13524 ( .A1(n11208), .A2(P1_U3086), .B1(n14534), .B2(n10919), 
        .C1(n10918), .C2(n14528), .ZN(P1_U3340) );
  OAI222_X1 U13525 ( .A1(n13803), .A2(n10920), .B1(n13800), .B2(n10919), .C1(
        P2_U3088), .C2(n11602), .ZN(P2_U3312) );
  INV_X1 U13526 ( .A(n14262), .ZN(n12049) );
  NAND2_X1 U13527 ( .A1(n10922), .A2(n10921), .ZN(n10924) );
  INV_X1 U13528 ( .A(n10931), .ZN(n10923) );
  NAND2_X1 U13529 ( .A1(n10924), .A2(n10923), .ZN(n11087) );
  OR2_X1 U13530 ( .A1(n10924), .A2(n10923), .ZN(n10925) );
  NAND2_X1 U13531 ( .A1(n11087), .A2(n10925), .ZN(n14751) );
  INV_X1 U13532 ( .A(n11098), .ZN(n11099) );
  OAI211_X1 U13533 ( .C1(n10927), .C2(n10926), .A(n11099), .B(n14370), .ZN(
        n14748) );
  INV_X1 U13534 ( .A(n14374), .ZN(n14323) );
  INV_X1 U13535 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14073) );
  AOI22_X1 U13536 ( .A1(n14384), .A2(n14694), .B1(n14323), .B2(n14073), .ZN(
        n10928) );
  OAI21_X1 U13537 ( .B1(n14387), .B2(n14748), .A(n10928), .ZN(n10939) );
  NAND2_X1 U13538 ( .A1(n14751), .A2(n14254), .ZN(n10937) );
  NAND2_X1 U13539 ( .A1(n10932), .A2(n10931), .ZN(n11092) );
  OAI21_X1 U13540 ( .B1(n10932), .B2(n10931), .A(n11092), .ZN(n10935) );
  OR2_X1 U13541 ( .A1(n11273), .A2(n14474), .ZN(n10934) );
  NAND2_X1 U13542 ( .A1(n14740), .A2(n14483), .ZN(n10933) );
  NAND2_X1 U13543 ( .A1(n10934), .A2(n10933), .ZN(n14703) );
  AOI21_X1 U13544 ( .B1(n10935), .B2(n14489), .A(n14703), .ZN(n10936) );
  NAND2_X1 U13545 ( .A1(n10937), .A2(n10936), .ZN(n14749) );
  MUX2_X1 U13546 ( .A(n14749), .B(P1_REG2_REG_3__SCAN_IN), .S(n14325), .Z(
        n10938) );
  AOI211_X1 U13547 ( .C1(n12049), .C2(n14751), .A(n10939), .B(n10938), .ZN(
        n10940) );
  INV_X1 U13548 ( .A(n10940), .ZN(P1_U3290) );
  INV_X1 U13549 ( .A(n10941), .ZN(n10942) );
  AOI211_X1 U13550 ( .C1(n14623), .C2(n10944), .A(n10943), .B(n10942), .ZN(
        n10949) );
  INV_X1 U13551 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10945) );
  OAI22_X1 U13552 ( .A1(n12117), .A2(n13780), .B1(n14915), .B2(n10945), .ZN(
        n10946) );
  INV_X1 U13553 ( .A(n10946), .ZN(n10947) );
  OAI21_X1 U13554 ( .B1(n10949), .B2(n14913), .A(n10947), .ZN(P2_U3451) );
  AOI22_X1 U13555 ( .A1(n12115), .A2(n13742), .B1(n14920), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10948) );
  OAI21_X1 U13556 ( .B1(n10949), .B2(n14920), .A(n10948), .ZN(P2_U3506) );
  INV_X1 U13557 ( .A(n10950), .ZN(n10952) );
  OAI22_X1 U13558 ( .A1(n12690), .A2(P3_U3151), .B1(SI_22_), .B2(n13142), .ZN(
        n10951) );
  AOI21_X1 U13559 ( .B1(n10952), .B2(n13134), .A(n10951), .ZN(P3_U3273) );
  XNOR2_X1 U13560 ( .A(n10954), .B(n10953), .ZN(n10955) );
  XNOR2_X1 U13561 ( .A(n10956), .B(n10955), .ZN(n10961) );
  INV_X1 U13562 ( .A(n11267), .ZN(n10957) );
  NAND2_X1 U13563 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14102) );
  OAI21_X1 U13564 ( .B1(n14707), .B2(n10957), .A(n14102), .ZN(n10959) );
  OAI22_X1 U13565 ( .A1(n11274), .A2(n13975), .B1(n13974), .B2(n11273), .ZN(
        n10958) );
  AOI211_X1 U13566 ( .C1(n14653), .C2(n11268), .A(n10959), .B(n10958), .ZN(
        n10960) );
  OAI21_X1 U13567 ( .B1(n10961), .B2(n14699), .A(n10960), .ZN(P1_U3227) );
  INV_X1 U13568 ( .A(n10962), .ZN(n10963) );
  NOR2_X1 U13569 ( .A1(n10964), .A2(n10963), .ZN(n10966) );
  XNOR2_X1 U13570 ( .A(n10966), .B(n10965), .ZN(n10972) );
  NOR2_X1 U13571 ( .A1(n11132), .A2(n14775), .ZN(n14756) );
  NAND2_X1 U13572 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14084) );
  OAI21_X1 U13573 ( .B1(n14707), .B2(n11100), .A(n14084), .ZN(n10970) );
  INV_X1 U13574 ( .A(n14038), .ZN(n10967) );
  OAI22_X1 U13575 ( .A1(n10968), .A2(n13975), .B1(n13974), .B2(n10967), .ZN(
        n10969) );
  AOI211_X1 U13576 ( .C1(n14756), .C2(n14697), .A(n10970), .B(n10969), .ZN(
        n10971) );
  OAI21_X1 U13577 ( .B1(n10972), .B2(n14699), .A(n10971), .ZN(P1_U3230) );
  AOI22_X1 U13578 ( .A1(n13265), .A2(n13289), .B1(n13261), .B2(n13287), .ZN(
        n10973) );
  NAND2_X1 U13579 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14855) );
  OAI211_X1 U13580 ( .C1(n11045), .C2(n13276), .A(n10973), .B(n14855), .ZN(
        n10979) );
  AOI22_X1 U13581 ( .A1(n10974), .A2(n9485), .B1(n13270), .B2(n13289), .ZN(
        n10976) );
  NOR3_X1 U13582 ( .A1(n10977), .A2(n10976), .A3(n10975), .ZN(n10978) );
  AOI211_X1 U13583 ( .C1(n12130), .C2(n13281), .A(n10979), .B(n10978), .ZN(
        n10980) );
  OAI21_X1 U13584 ( .B1(n10981), .B2(n13272), .A(n10980), .ZN(P2_U3203) );
  OR2_X1 U13585 ( .A1(n12115), .A2(n13290), .ZN(n10982) );
  INV_X1 U13586 ( .A(n14897), .ZN(n10995) );
  NAND2_X1 U13587 ( .A1(n10984), .A2(n12307), .ZN(n10985) );
  NAND2_X1 U13588 ( .A1(n11037), .A2(n10985), .ZN(n14895) );
  OR2_X1 U13589 ( .A1(n12115), .A2(n12116), .ZN(n10986) );
  XOR2_X1 U13590 ( .A(n11038), .B(n12307), .Z(n10989) );
  INV_X1 U13591 ( .A(n13288), .ZN(n12131) );
  OAI22_X1 U13592 ( .A1(n12116), .A2(n13630), .B1(n12131), .B2(n13632), .ZN(
        n10988) );
  AOI21_X1 U13593 ( .B1(n10989), .B2(n13635), .A(n10988), .ZN(n10990) );
  OAI21_X1 U13594 ( .B1(n10088), .B2(n14895), .A(n10990), .ZN(n14898) );
  NAND2_X1 U13595 ( .A1(n14898), .A2(n15210), .ZN(n10997) );
  INV_X1 U13596 ( .A(n13603), .ZN(n13654) );
  OAI22_X1 U13597 ( .A1(n15210), .A2(n10992), .B1(n10991), .B2(n13651), .ZN(
        n10994) );
  NAND2_X1 U13598 ( .A1(n14897), .A2(n7445), .ZN(n11044) );
  OAI211_X1 U13599 ( .C1(n14897), .C2(n7445), .A(n13639), .B(n11044), .ZN(
        n14896) );
  NOR2_X1 U13600 ( .A1(n14896), .A2(n13641), .ZN(n10993) );
  AOI211_X1 U13601 ( .C1(n13654), .C2(n10995), .A(n10994), .B(n10993), .ZN(
        n10996) );
  OAI211_X1 U13602 ( .C1(n14895), .C2(n11518), .A(n10997), .B(n10996), .ZN(
        P2_U3257) );
  OAI21_X1 U13603 ( .B1(n10999), .B2(n12498), .A(n10998), .ZN(n11062) );
  INV_X1 U13604 ( .A(n11062), .ZN(n11008) );
  AOI21_X1 U13605 ( .B1(n11000), .B2(n12498), .A(n12954), .ZN(n11005) );
  OAI22_X1 U13606 ( .A1(n11002), .A2(n12956), .B1(n11001), .B2(n12958), .ZN(
        n11003) );
  AOI21_X1 U13607 ( .B1(n11005), .B2(n11004), .A(n11003), .ZN(n11060) );
  MUX2_X1 U13608 ( .A(n11060), .B(n10276), .S(n15004), .Z(n11007) );
  AOI22_X1 U13609 ( .A1(n12994), .A2(n11066), .B1(n14998), .B2(n11117), .ZN(
        n11006) );
  OAI211_X1 U13610 ( .C1(n12997), .C2(n11008), .A(n11007), .B(n11006), .ZN(
        P3_U3227) );
  AOI21_X1 U13611 ( .B1(n15032), .B2(n11010), .A(n11009), .ZN(n11017) );
  AOI22_X1 U13612 ( .A1(n8048), .A2(n11011), .B1(n15049), .B2(
        P3_REG1_REG_5__SCAN_IN), .ZN(n11012) );
  OAI21_X1 U13613 ( .B1(n11017), .B2(n15049), .A(n11012), .ZN(P3_U3464) );
  INV_X1 U13614 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11013) );
  OAI22_X1 U13615 ( .A1(n11014), .A2(n13097), .B1(n15039), .B2(n11013), .ZN(
        n11015) );
  INV_X1 U13616 ( .A(n11015), .ZN(n11016) );
  OAI21_X1 U13617 ( .B1(n11017), .B2(n15037), .A(n11016), .ZN(P3_U3405) );
  NAND2_X1 U13618 ( .A1(n12706), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11018) );
  OAI21_X1 U13619 ( .B1(n12837), .B2(n12706), .A(n11018), .ZN(P3_U3520) );
  INV_X1 U13620 ( .A(n14864), .ZN(n13321) );
  OAI222_X1 U13621 ( .A1(n13803), .A2(n11019), .B1(n13800), .B2(n11021), .C1(
        n13321), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13622 ( .A(n14184), .ZN(n11860) );
  OAI222_X1 U13623 ( .A1(P1_U3086), .A2(n11860), .B1(n14534), .B2(n11021), 
        .C1(n11020), .C2(n14528), .ZN(P1_U3337) );
  NAND2_X1 U13624 ( .A1(n12706), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11022) );
  OAI21_X1 U13625 ( .B1(n12349), .B2(n12706), .A(n11022), .ZN(P3_U3519) );
  OAI211_X1 U13626 ( .C1(n11024), .C2(n12561), .A(n11023), .B(n14991), .ZN(
        n11028) );
  OAI22_X1 U13627 ( .A1(n11025), .A2(n12956), .B1(n11391), .B2(n12958), .ZN(
        n11026) );
  INV_X1 U13628 ( .A(n11026), .ZN(n11027) );
  AND2_X1 U13629 ( .A1(n11028), .A2(n11027), .ZN(n15018) );
  OR2_X1 U13630 ( .A1(n11029), .A2(n12502), .ZN(n11030) );
  NAND2_X1 U13631 ( .A1(n11031), .A2(n11030), .ZN(n15016) );
  NOR2_X1 U13632 ( .A1(n12847), .A2(n11055), .ZN(n11034) );
  INV_X1 U13633 ( .A(n11057), .ZN(n11032) );
  OAI22_X1 U13634 ( .A1(n15002), .A2(n14928), .B1(n11032), .B2(n14580), .ZN(
        n11033) );
  AOI211_X1 U13635 ( .C1(n15016), .C2(n14599), .A(n11034), .B(n11033), .ZN(
        n11035) );
  OAI21_X1 U13636 ( .B1(n15018), .B2(n15004), .A(n11035), .ZN(P3_U3226) );
  OR2_X1 U13637 ( .A1(n14897), .A2(n12123), .ZN(n11036) );
  NAND2_X1 U13638 ( .A1(n11037), .A2(n11036), .ZN(n11284) );
  XNOR2_X1 U13639 ( .A(n12130), .B(n13288), .ZN(n12306) );
  XNOR2_X1 U13640 ( .A(n11284), .B(n11283), .ZN(n11226) );
  NAND2_X1 U13641 ( .A1(n11038), .A2(n12307), .ZN(n11040) );
  NAND2_X1 U13642 ( .A1(n14897), .A2(n13289), .ZN(n11039) );
  XNOR2_X1 U13643 ( .A(n6743), .B(n11283), .ZN(n11042) );
  INV_X1 U13644 ( .A(n13287), .ZN(n11366) );
  OAI22_X1 U13645 ( .A1(n11366), .A2(n13632), .B1(n12123), .B2(n13630), .ZN(
        n11041) );
  AOI21_X1 U13646 ( .B1(n11042), .B2(n13635), .A(n11041), .ZN(n11043) );
  OAI21_X1 U13647 ( .B1(n11226), .B2(n10088), .A(n11043), .ZN(n11227) );
  NAND2_X1 U13648 ( .A1(n11227), .A2(n15210), .ZN(n11050) );
  AOI211_X1 U13649 ( .C1(n12130), .C2(n11044), .A(n13620), .B(n6701), .ZN(
        n11228) );
  INV_X1 U13650 ( .A(n12130), .ZN(n12132) );
  NOR2_X1 U13651 ( .A1(n12132), .A2(n13603), .ZN(n11048) );
  OAI22_X1 U13652 ( .A1(n15210), .A2(n11046), .B1(n11045), .B2(n13651), .ZN(
        n11047) );
  AOI211_X1 U13653 ( .C1(n11228), .C2(n13658), .A(n11048), .B(n11047), .ZN(
        n11049) );
  OAI211_X1 U13654 ( .C1(n11226), .C2(n11518), .A(n11050), .B(n11049), .ZN(
        P2_U3256) );
  OAI211_X1 U13655 ( .C1(n11053), .C2(n11052), .A(n11051), .B(n12449), .ZN(
        n11059) );
  AOI22_X1 U13656 ( .A1(n6439), .A2(n12702), .B1(n12463), .B2(n12700), .ZN(
        n11054) );
  NAND2_X1 U13657 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_U3151), .ZN(n14938) );
  OAI211_X1 U13658 ( .C1(n11055), .C2(n12459), .A(n11054), .B(n14938), .ZN(
        n11056) );
  AOI21_X1 U13659 ( .B1(n11057), .B2(n12464), .A(n11056), .ZN(n11058) );
  NAND2_X1 U13660 ( .A1(n11059), .A2(n11058), .ZN(P3_U3153) );
  INV_X1 U13661 ( .A(n11060), .ZN(n11061) );
  AOI21_X1 U13662 ( .B1(n15032), .B2(n11062), .A(n11061), .ZN(n11068) );
  INV_X1 U13663 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11063) );
  OAI22_X1 U13664 ( .A1(n11110), .A2(n13097), .B1(n15039), .B2(n11063), .ZN(
        n11064) );
  INV_X1 U13665 ( .A(n11064), .ZN(n11065) );
  OAI21_X1 U13666 ( .B1(n11068), .B2(n15037), .A(n11065), .ZN(P3_U3408) );
  AOI22_X1 U13667 ( .A1(n8048), .A2(n11066), .B1(n15049), .B2(
        P3_REG1_REG_6__SCAN_IN), .ZN(n11067) );
  OAI21_X1 U13668 ( .B1(n11068), .B2(n15049), .A(n11067), .ZN(P3_U3465) );
  XNOR2_X1 U13669 ( .A(n11070), .B(n11069), .ZN(n11076) );
  NAND2_X1 U13670 ( .A1(n14037), .A2(n14483), .ZN(n11072) );
  NAND2_X1 U13671 ( .A1(n14035), .A2(n14739), .ZN(n11071) );
  NAND2_X1 U13672 ( .A1(n11072), .A2(n11071), .ZN(n11168) );
  NAND2_X1 U13673 ( .A1(n14704), .A2(n11168), .ZN(n11073) );
  NAND2_X1 U13674 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14122) );
  OAI211_X1 U13675 ( .C1(n14707), .C2(n11174), .A(n11073), .B(n14122), .ZN(
        n11074) );
  AOI21_X1 U13676 ( .B1(n14653), .B2(n14765), .A(n11074), .ZN(n11075) );
  OAI21_X1 U13677 ( .B1(n11076), .B2(n14699), .A(n11075), .ZN(P1_U3239) );
  AOI21_X1 U13678 ( .B1(n11078), .B2(n11077), .A(n13272), .ZN(n11080) );
  NAND2_X1 U13679 ( .A1(n11080), .A2(n11079), .ZN(n11085) );
  INV_X1 U13680 ( .A(n13652), .ZN(n11083) );
  INV_X1 U13681 ( .A(n12141), .ZN(n13286) );
  AOI22_X1 U13682 ( .A1(n13286), .A2(n13544), .B1(n13542), .B2(n13288), .ZN(
        n11291) );
  OAI22_X1 U13683 ( .A1(n13199), .A2(n11291), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11081), .ZN(n11082) );
  AOI21_X1 U13684 ( .B1(n11083), .B2(n13240), .A(n11082), .ZN(n11084) );
  OAI211_X1 U13685 ( .C1(n6700), .C2(n13258), .A(n11085), .B(n11084), .ZN(
        P2_U3189) );
  OR2_X1 U13686 ( .A1(n14038), .A2(n14694), .ZN(n11086) );
  NAND2_X1 U13687 ( .A1(n11087), .A2(n11086), .ZN(n11088) );
  NAND2_X1 U13688 ( .A1(n11088), .A2(n11093), .ZN(n11134) );
  OAI21_X1 U13689 ( .B1(n11088), .B2(n11093), .A(n11134), .ZN(n11089) );
  INV_X1 U13690 ( .A(n11089), .ZN(n14754) );
  INV_X1 U13691 ( .A(n11090), .ZN(n11091) );
  NAND2_X1 U13692 ( .A1(n11092), .A2(n11091), .ZN(n11095) );
  INV_X1 U13693 ( .A(n11093), .ZN(n11094) );
  NAND2_X1 U13694 ( .A1(n11095), .A2(n11094), .ZN(n11145) );
  OAI21_X1 U13695 ( .B1(n11095), .B2(n11094), .A(n11145), .ZN(n11096) );
  AOI222_X1 U13696 ( .A1(n14489), .A2(n11096), .B1(n14037), .B2(n14739), .C1(
        n14038), .C2(n14483), .ZN(n14752) );
  MUX2_X1 U13697 ( .A(n11097), .B(n14752), .S(n14377), .Z(n11103) );
  AND2_X1 U13698 ( .A1(n11098), .A2(n11132), .ZN(n11266) );
  AOI211_X1 U13699 ( .C1(n11143), .C2(n11099), .A(n14355), .B(n11266), .ZN(
        n14755) );
  OAI22_X1 U13700 ( .A1(n14364), .A2(n11132), .B1(n14374), .B2(n11100), .ZN(
        n11101) );
  AOI21_X1 U13701 ( .B1(n14755), .B2(n14357), .A(n11101), .ZN(n11102) );
  OAI211_X1 U13702 ( .C1(n14391), .C2(n14754), .A(n11103), .B(n11102), .ZN(
        P1_U3289) );
  NAND2_X1 U13703 ( .A1(n11104), .A2(n13134), .ZN(n11105) );
  OAI211_X1 U13704 ( .C1(n11106), .C2(n13142), .A(n11105), .B(n12693), .ZN(
        P3_U3272) );
  AOI22_X1 U13705 ( .A1(n6439), .A2(n12703), .B1(n12463), .B2(n12701), .ZN(
        n11109) );
  INV_X1 U13706 ( .A(n11107), .ZN(n11108) );
  OAI211_X1 U13707 ( .C1(n11110), .C2(n12459), .A(n11109), .B(n11108), .ZN(
        n11116) );
  INV_X1 U13708 ( .A(n11111), .ZN(n11112) );
  AOI211_X1 U13709 ( .C1(n11114), .C2(n11113), .A(n12471), .B(n11112), .ZN(
        n11115) );
  AOI211_X1 U13710 ( .C1(n11117), .C2(n12464), .A(n11116), .B(n11115), .ZN(
        n11118) );
  INV_X1 U13711 ( .A(n11118), .ZN(P3_U3179) );
  XNOR2_X1 U13712 ( .A(n11525), .B(n11524), .ZN(n11121) );
  INV_X1 U13713 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11120) );
  NOR2_X1 U13714 ( .A1(n11120), .A2(n11121), .ZN(n11526) );
  AOI211_X1 U13715 ( .C1(n11121), .C2(n11120), .A(n11526), .B(n11825), .ZN(
        n11131) );
  NAND2_X1 U13716 ( .A1(n11122), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11124) );
  INV_X1 U13717 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14628) );
  MUX2_X1 U13718 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14628), .S(n11524), .Z(
        n11123) );
  AOI21_X1 U13719 ( .B1(n11125), .B2(n11124), .A(n11123), .ZN(n11519) );
  AND3_X1 U13720 ( .A1(n11125), .A2(n11124), .A3(n11123), .ZN(n11126) );
  NOR3_X1 U13721 ( .A1(n11519), .A2(n11126), .A3(n13328), .ZN(n11130) );
  NAND2_X1 U13722 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11615)
         );
  INV_X1 U13723 ( .A(n11615), .ZN(n11127) );
  AOI21_X1 U13724 ( .B1(n14859), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n11127), 
        .ZN(n11128) );
  OAI21_X1 U13725 ( .B1(n11524), .B2(n14820), .A(n11128), .ZN(n11129) );
  OR3_X1 U13726 ( .A1(n11131), .A2(n11130), .A3(n11129), .ZN(P2_U3228) );
  NAND2_X1 U13727 ( .A1(n11273), .A2(n11132), .ZN(n11133) );
  NAND2_X1 U13728 ( .A1(n11134), .A2(n11133), .ZN(n11264) );
  INV_X1 U13729 ( .A(n11272), .ZN(n11263) );
  NAND2_X1 U13730 ( .A1(n11264), .A2(n11263), .ZN(n11262) );
  OR2_X1 U13731 ( .A1(n11268), .A2(n14037), .ZN(n11135) );
  OR2_X1 U13732 ( .A1(n11256), .A2(n14035), .ZN(n11136) );
  NAND2_X1 U13733 ( .A1(n11243), .A2(n11136), .ZN(n11138) );
  NAND2_X1 U13734 ( .A1(n11138), .A2(n11152), .ZN(n11353) );
  OAI21_X1 U13735 ( .B1(n11138), .B2(n11152), .A(n11353), .ZN(n11217) );
  INV_X1 U13736 ( .A(n11217), .ZN(n11160) );
  OAI22_X1 U13737 ( .A1(n14377), .A2(n10294), .B1(n11429), .B2(n14374), .ZN(
        n11142) );
  NAND2_X1 U13738 ( .A1(n11266), .A2(n14761), .ZN(n11265) );
  OR2_X1 U13739 ( .A1(n11253), .A2(n11256), .ZN(n11254) );
  NAND2_X1 U13740 ( .A1(n11254), .A2(n11431), .ZN(n11139) );
  NAND2_X1 U13741 ( .A1(n11139), .A2(n14370), .ZN(n11140) );
  OR2_X1 U13742 ( .A1(n11140), .A2(n11484), .ZN(n11218) );
  NOR2_X1 U13743 ( .A1(n11218), .A2(n14387), .ZN(n11141) );
  AOI211_X1 U13744 ( .C1(n14384), .C2(n11431), .A(n11142), .B(n11141), .ZN(
        n11159) );
  NAND2_X1 U13745 ( .A1(n11273), .A2(n11143), .ZN(n11144) );
  NAND2_X1 U13746 ( .A1(n11270), .A2(n11165), .ZN(n11147) );
  NAND2_X1 U13747 ( .A1(n11147), .A2(n11146), .ZN(n11167) );
  INV_X1 U13748 ( .A(n11240), .ZN(n11245) );
  NAND2_X1 U13749 ( .A1(n11246), .A2(n11245), .ZN(n11244) );
  NAND2_X1 U13750 ( .A1(n11256), .A2(n11149), .ZN(n11150) );
  NAND2_X1 U13751 ( .A1(n11244), .A2(n11150), .ZN(n11151) );
  AOI21_X1 U13752 ( .B1(n11151), .B2(n11152), .A(n14795), .ZN(n11154) );
  INV_X1 U13753 ( .A(n11151), .ZN(n11153) );
  NAND2_X1 U13754 ( .A1(n11154), .A2(n11342), .ZN(n11219) );
  INV_X1 U13755 ( .A(n11219), .ZN(n11157) );
  OR2_X1 U13756 ( .A1(n11656), .A2(n14474), .ZN(n11156) );
  NAND2_X1 U13757 ( .A1(n14035), .A2(n14483), .ZN(n11155) );
  NAND2_X1 U13758 ( .A1(n11156), .A2(n11155), .ZN(n11427) );
  OAI21_X1 U13759 ( .B1(n11157), .B2(n11427), .A(n14377), .ZN(n11158) );
  OAI211_X1 U13760 ( .C1(n11160), .C2(n14391), .A(n11159), .B(n11158), .ZN(
        P1_U3285) );
  OR2_X1 U13761 ( .A1(n11161), .A2(n11164), .ZN(n11162) );
  NAND2_X1 U13762 ( .A1(n11163), .A2(n11162), .ZN(n14769) );
  INV_X1 U13763 ( .A(n14769), .ZN(n11179) );
  NAND2_X1 U13764 ( .A1(n14769), .A2(n14254), .ZN(n11171) );
  NAND3_X1 U13765 ( .A1(n11270), .A2(n11165), .A3(n11164), .ZN(n11166) );
  NAND2_X1 U13766 ( .A1(n11167), .A2(n11166), .ZN(n11169) );
  AOI21_X1 U13767 ( .B1(n11169), .B2(n14489), .A(n11168), .ZN(n11170) );
  AND2_X1 U13768 ( .A1(n11171), .A2(n11170), .ZN(n14771) );
  MUX2_X1 U13769 ( .A(n11172), .B(n14771), .S(n14377), .Z(n11178) );
  AOI21_X1 U13770 ( .B1(n11265), .B2(n14765), .A(n14355), .ZN(n11173) );
  AND2_X1 U13771 ( .A1(n11173), .A2(n11253), .ZN(n14767) );
  OAI22_X1 U13772 ( .A1(n14364), .A2(n11175), .B1(n14374), .B2(n11174), .ZN(
        n11176) );
  AOI21_X1 U13773 ( .B1(n14767), .B2(n14357), .A(n11176), .ZN(n11177) );
  OAI211_X1 U13774 ( .C1(n11179), .C2(n14262), .A(n11178), .B(n11177), .ZN(
        P1_U3287) );
  NOR2_X1 U13775 ( .A1(n6599), .A2(n11180), .ZN(n11181) );
  XNOR2_X1 U13776 ( .A(n11182), .B(n11181), .ZN(n11186) );
  INV_X1 U13777 ( .A(n14908), .ZN(n11375) );
  OAI22_X1 U13778 ( .A1(n11366), .A2(n13630), .B1(n12150), .B2(n13632), .ZN(
        n11368) );
  AOI22_X1 U13779 ( .A1(n13251), .A2(n11368), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11183) );
  OAI21_X1 U13780 ( .B1(n11372), .B2(n13276), .A(n11183), .ZN(n11184) );
  AOI21_X1 U13781 ( .B1(n11375), .B2(n13281), .A(n11184), .ZN(n11185) );
  OAI21_X1 U13782 ( .B1(n11186), .B2(n13272), .A(n11185), .ZN(P2_U3208) );
  XNOR2_X1 U13783 ( .A(n11188), .B(n11187), .ZN(n11193) );
  OAI21_X1 U13784 ( .B1(n14707), .B2(n11257), .A(n11189), .ZN(n11191) );
  OAI22_X1 U13785 ( .A1(n11274), .A2(n13974), .B1(n13975), .B2(n11627), .ZN(
        n11190) );
  AOI211_X1 U13786 ( .C1(n14653), .C2(n11256), .A(n11191), .B(n11190), .ZN(
        n11192) );
  OAI21_X1 U13787 ( .B1(n11193), .B2(n14699), .A(n11192), .ZN(P1_U3213) );
  AND2_X1 U13788 ( .A1(n14377), .A2(n14739), .ZN(n14379) );
  INV_X1 U13789 ( .A(n14379), .ZN(n11457) );
  NOR2_X1 U13790 ( .A1(n14374), .A2(n11194), .ZN(n11198) );
  NOR3_X1 U13791 ( .A1(n14325), .A2(n11196), .A3(n11195), .ZN(n11197) );
  AOI211_X1 U13792 ( .C1(n14325), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11198), .B(
        n11197), .ZN(n11202) );
  NAND2_X1 U13793 ( .A1(n14377), .A2(n14489), .ZN(n14346) );
  INV_X1 U13794 ( .A(n14346), .ZN(n14389) );
  INV_X1 U13795 ( .A(n11199), .ZN(n11200) );
  OAI21_X1 U13796 ( .B1(n14337), .B2(n14389), .A(n11200), .ZN(n11201) );
  OAI211_X1 U13797 ( .C1(n11203), .C2(n11457), .A(n11202), .B(n11201), .ZN(
        P1_U3293) );
  XNOR2_X1 U13798 ( .A(n11849), .B(n11839), .ZN(n11205) );
  NOR2_X1 U13799 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n11205), .ZN(n11840) );
  AOI21_X1 U13800 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n11205), .A(n11840), 
        .ZN(n11216) );
  OAI21_X1 U13801 ( .B1(n11803), .B2(n11207), .A(n11206), .ZN(n11848) );
  XOR2_X1 U13802 ( .A(n11208), .B(n11848), .Z(n11209) );
  NOR2_X1 U13803 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11209), .ZN(n11850) );
  AOI21_X1 U13804 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11209), .A(n11850), 
        .ZN(n11213) );
  NOR2_X1 U13805 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14013), .ZN(n11210) );
  AOI21_X1 U13806 ( .B1(n14733), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n11210), 
        .ZN(n11212) );
  NAND2_X1 U13807 ( .A1(n14722), .A2(n11849), .ZN(n11211) );
  OAI211_X1 U13808 ( .C1(n11213), .C2(n14190), .A(n11212), .B(n11211), .ZN(
        n11214) );
  INV_X1 U13809 ( .A(n11214), .ZN(n11215) );
  OAI21_X1 U13810 ( .B1(n11216), .B2(n14729), .A(n11215), .ZN(P1_U3258) );
  NAND2_X1 U13811 ( .A1(n11217), .A2(n14799), .ZN(n11221) );
  AOI21_X1 U13812 ( .B1(n11431), .B2(n14793), .A(n11427), .ZN(n11220) );
  NAND4_X1 U13813 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11223) );
  NAND2_X1 U13814 ( .A1(n11223), .A2(n14813), .ZN(n11222) );
  OAI21_X1 U13815 ( .B1(n14813), .B2(n8281), .A(n11222), .ZN(P1_U3536) );
  INV_X1 U13816 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11225) );
  NAND2_X1 U13817 ( .A1(n11223), .A2(n14802), .ZN(n11224) );
  OAI21_X1 U13818 ( .B1(n14802), .B2(n11225), .A(n11224), .ZN(P1_U3483) );
  INV_X1 U13819 ( .A(n11226), .ZN(n11229) );
  AOI211_X1 U13820 ( .C1(n14901), .C2(n11229), .A(n11228), .B(n11227), .ZN(
        n11234) );
  AOI22_X1 U13821 ( .A1(n12130), .A2(n13742), .B1(n14920), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11230) );
  OAI21_X1 U13822 ( .B1(n11234), .B2(n14920), .A(n11230), .ZN(P2_U3508) );
  INV_X1 U13823 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11231) );
  OAI22_X1 U13824 ( .A1(n12132), .A2(n13780), .B1(n14915), .B2(n11231), .ZN(
        n11232) );
  INV_X1 U13825 ( .A(n11232), .ZN(n11233) );
  OAI21_X1 U13826 ( .B1(n11234), .B2(n14913), .A(n11233), .ZN(P2_U3457) );
  INV_X1 U13827 ( .A(n11235), .ZN(n11238) );
  OAI222_X1 U13828 ( .A1(n13803), .A2(n11236), .B1(n13800), .B2(n11238), .C1(
        n12334), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13829 ( .A1(P1_U3086), .A2(n11239), .B1(n14534), .B2(n11238), 
        .C1(n11237), .C2(n14528), .ZN(P1_U3336) );
  OR2_X1 U13830 ( .A1(n11241), .A2(n11240), .ZN(n11242) );
  NAND2_X1 U13831 ( .A1(n11243), .A2(n11242), .ZN(n14778) );
  INV_X1 U13832 ( .A(n14778), .ZN(n11261) );
  NAND2_X1 U13833 ( .A1(n14778), .A2(n14254), .ZN(n11251) );
  OAI21_X1 U13834 ( .B1(n11246), .B2(n11245), .A(n11244), .ZN(n11249) );
  NAND2_X1 U13835 ( .A1(n14036), .A2(n14483), .ZN(n11247) );
  OAI21_X1 U13836 ( .B1(n11627), .B2(n14474), .A(n11247), .ZN(n11248) );
  AOI21_X1 U13837 ( .B1(n11249), .B2(n14489), .A(n11248), .ZN(n11250) );
  AND2_X1 U13838 ( .A1(n11251), .A2(n11250), .ZN(n14780) );
  MUX2_X1 U13839 ( .A(n11252), .B(n14780), .S(n14377), .Z(n11260) );
  AOI21_X1 U13840 ( .B1(n11253), .B2(n11256), .A(n14355), .ZN(n11255) );
  AND2_X1 U13841 ( .A1(n11255), .A2(n11254), .ZN(n14773) );
  INV_X1 U13842 ( .A(n11256), .ZN(n14776) );
  OAI22_X1 U13843 ( .A1(n14776), .A2(n14364), .B1(n14374), .B2(n11257), .ZN(
        n11258) );
  AOI21_X1 U13844 ( .B1(n14773), .B2(n14357), .A(n11258), .ZN(n11259) );
  OAI211_X1 U13845 ( .C1(n11261), .C2(n14262), .A(n11260), .B(n11259), .ZN(
        P1_U3286) );
  OAI21_X1 U13846 ( .B1(n11264), .B2(n11263), .A(n11262), .ZN(n14764) );
  OAI211_X1 U13847 ( .C1(n11266), .C2(n14761), .A(n14370), .B(n11265), .ZN(
        n14760) );
  AOI22_X1 U13848 ( .A1(n14384), .A2(n11268), .B1(n11267), .B2(n14323), .ZN(
        n11269) );
  OAI21_X1 U13849 ( .B1(n14760), .B2(n14387), .A(n11269), .ZN(n11281) );
  INV_X1 U13850 ( .A(n14764), .ZN(n11279) );
  OAI21_X1 U13851 ( .B1(n11272), .B2(n11271), .A(n11270), .ZN(n11276) );
  OAI22_X1 U13852 ( .A1(n11274), .A2(n14474), .B1(n11273), .B2(n14400), .ZN(
        n11275) );
  AOI21_X1 U13853 ( .B1(n11276), .B2(n14489), .A(n11275), .ZN(n11277) );
  OAI21_X1 U13854 ( .B1(n11279), .B2(n11278), .A(n11277), .ZN(n14762) );
  MUX2_X1 U13855 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n14762), .S(n14377), .Z(
        n11280) );
  AOI211_X1 U13856 ( .C1(n12049), .C2(n14764), .A(n11281), .B(n11280), .ZN(
        n11282) );
  INV_X1 U13857 ( .A(n11282), .ZN(P1_U3288) );
  NAND2_X1 U13858 ( .A1(n11284), .A2(n11283), .ZN(n11286) );
  NAND2_X1 U13859 ( .A1(n12130), .A2(n13288), .ZN(n11285) );
  XNOR2_X1 U13860 ( .A(n13655), .B(n13287), .ZN(n12309) );
  XNOR2_X1 U13861 ( .A(n11363), .B(n12309), .ZN(n13657) );
  NAND2_X1 U13862 ( .A1(n13655), .A2(n11287), .ZN(n11288) );
  NAND2_X1 U13863 ( .A1(n11288), .A2(n13639), .ZN(n11289) );
  NOR2_X1 U13864 ( .A1(n11370), .A2(n11289), .ZN(n13659) );
  INV_X1 U13865 ( .A(n12309), .ZN(n11362) );
  OAI211_X1 U13866 ( .C1(n6594), .C2(n12309), .A(n13635), .B(n11367), .ZN(
        n11292) );
  NAND2_X1 U13867 ( .A1(n11292), .A2(n11291), .ZN(n13650) );
  AOI211_X1 U13868 ( .C1(n14623), .C2(n13657), .A(n13659), .B(n13650), .ZN(
        n11297) );
  AOI22_X1 U13869 ( .A1(n13655), .A2(n13742), .B1(n14920), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11293) );
  OAI21_X1 U13870 ( .B1(n11297), .B2(n14920), .A(n11293), .ZN(P2_U3509) );
  INV_X1 U13871 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11294) );
  NOR2_X1 U13872 ( .A1(n14915), .A2(n11294), .ZN(n11295) );
  AOI21_X1 U13873 ( .B1(n13655), .B2(n6641), .A(n11295), .ZN(n11296) );
  OAI21_X1 U13874 ( .B1(n11297), .B2(n14913), .A(n11296), .ZN(P2_U3460) );
  OAI21_X1 U13875 ( .B1(n11300), .B2(n11299), .A(n11298), .ZN(n11301) );
  NAND2_X1 U13876 ( .A1(n11301), .A2(n9485), .ZN(n11306) );
  INV_X1 U13877 ( .A(n11511), .ZN(n11304) );
  INV_X1 U13878 ( .A(n13284), .ZN(n12158) );
  OAI22_X1 U13879 ( .A1(n13278), .A2(n12158), .B1(n12141), .B2(n13277), .ZN(
        n11302) );
  AOI211_X1 U13880 ( .C1(n13240), .C2(n11304), .A(n11303), .B(n11302), .ZN(
        n11305) );
  OAI211_X1 U13881 ( .C1(n14631), .C2(n13258), .A(n11306), .B(n11305), .ZN(
        P2_U3196) );
  INV_X1 U13882 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11311) );
  NOR2_X1 U13883 ( .A1(n11330), .A2(n6575), .ZN(n11308) );
  INV_X1 U13884 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11309) );
  MUX2_X1 U13885 ( .A(n11309), .B(P3_REG2_REG_10__SCAN_IN), .S(n14944), .Z(
        n14942) );
  AOI21_X1 U13886 ( .B1(n11311), .B2(n11310), .A(n11414), .ZN(n11340) );
  INV_X1 U13887 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11312) );
  MUX2_X1 U13888 ( .A(n11311), .B(n11312), .S(n12799), .Z(n11313) );
  AND2_X1 U13889 ( .A1(n11413), .A2(n11313), .ZN(n11410) );
  NOR2_X1 U13890 ( .A1(n11413), .A2(n11313), .ZN(n11314) );
  OR2_X1 U13891 ( .A1(n11410), .A2(n11314), .ZN(n11324) );
  MUX2_X1 U13892 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12799), .Z(n11319) );
  OR2_X1 U13893 ( .A1(n11319), .A2(n14944), .ZN(n11321) );
  INV_X1 U13894 ( .A(n11321), .ZN(n11322) );
  INV_X1 U13895 ( .A(n11315), .ZN(n11316) );
  NAND2_X1 U13896 ( .A1(n14944), .A2(n11319), .ZN(n11320) );
  NAND2_X1 U13897 ( .A1(n11321), .A2(n11320), .ZN(n14956) );
  NOR2_X1 U13898 ( .A1(n14957), .A2(n14956), .ZN(n14955) );
  NOR2_X1 U13899 ( .A1(n11322), .A2(n14955), .ZN(n11323) );
  NOR2_X1 U13900 ( .A1(n11323), .A2(n11324), .ZN(n11409) );
  AOI21_X1 U13901 ( .B1(n11324), .B2(n11323), .A(n11409), .ZN(n11328) );
  NAND2_X1 U13902 ( .A1(n14923), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11327) );
  INV_X1 U13903 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11325) );
  NOR2_X1 U13904 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11325), .ZN(n11635) );
  INV_X1 U13905 ( .A(n11635), .ZN(n11326) );
  OAI211_X1 U13906 ( .C1(n11328), .C2(n14975), .A(n11327), .B(n11326), .ZN(
        n11338) );
  NOR2_X1 U13907 ( .A1(n11330), .A2(n11329), .ZN(n11332) );
  INV_X1 U13908 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11333) );
  MUX2_X1 U13909 ( .A(n11333), .B(P3_REG1_REG_10__SCAN_IN), .S(n14944), .Z(
        n14947) );
  NAND2_X1 U13910 ( .A1(n14944), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11334) );
  XNOR2_X1 U13911 ( .A(n11413), .B(n11402), .ZN(n11335) );
  NOR2_X1 U13912 ( .A1(n11312), .A2(n11335), .ZN(n11403) );
  AOI21_X1 U13913 ( .B1(n11312), .B2(n11335), .A(n11403), .ZN(n11336) );
  NOR2_X1 U13914 ( .A1(n11336), .A2(n14977), .ZN(n11337) );
  AOI211_X1 U13915 ( .C1(n14954), .C2(n11413), .A(n11338), .B(n11337), .ZN(
        n11339) );
  OAI21_X1 U13916 ( .B1(n11340), .B2(n14983), .A(n11339), .ZN(P3_U3193) );
  OAI21_X1 U13917 ( .B1(n11346), .B2(n11345), .A(n11576), .ZN(n14796) );
  NAND2_X1 U13918 ( .A1(n14377), .A2(n14483), .ZN(n14381) );
  INV_X1 U13919 ( .A(n11658), .ZN(n11347) );
  AOI22_X1 U13920 ( .A1(n14325), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11347), 
        .B2(n14323), .ZN(n11348) );
  OAI21_X1 U13921 ( .B1(n11656), .B2(n14381), .A(n11348), .ZN(n11351) );
  AOI211_X1 U13922 ( .C1(n14792), .C2(n11485), .A(n14355), .B(n6598), .ZN(
        n14790) );
  INV_X1 U13923 ( .A(n14790), .ZN(n11349) );
  NAND2_X1 U13924 ( .A1(n14033), .A2(n14739), .ZN(n11655) );
  AOI21_X1 U13925 ( .B1(n11349), .B2(n11655), .A(n14387), .ZN(n11350) );
  AOI211_X1 U13926 ( .C1(n14384), .C2(n14792), .A(n11351), .B(n11350), .ZN(
        n11358) );
  NAND2_X1 U13927 ( .A1(n11621), .A2(n11656), .ZN(n11354) );
  OAI21_X1 U13928 ( .B1(n11356), .B2(n11355), .A(n11581), .ZN(n14798) );
  NAND2_X1 U13929 ( .A1(n14798), .A2(n14337), .ZN(n11357) );
  OAI211_X1 U13930 ( .C1(n14796), .C2(n14346), .A(n11358), .B(n11357), .ZN(
        P1_U3283) );
  INV_X1 U13931 ( .A(n11359), .ZN(n11360) );
  OAI222_X1 U13932 ( .A1(P3_U3151), .A2(n11361), .B1(n13140), .B2(n11360), 
        .C1(n15168), .C2(n13142), .ZN(P3_U3271) );
  XNOR2_X1 U13933 ( .A(n11375), .B(n12141), .ZN(n12311) );
  NAND2_X1 U13934 ( .A1(n11363), .A2(n11362), .ZN(n11365) );
  NAND2_X1 U13935 ( .A1(n13655), .A2(n13287), .ZN(n11364) );
  XOR2_X1 U13936 ( .A(n11504), .B(n12311), .Z(n14911) );
  INV_X1 U13937 ( .A(n14911), .ZN(n14904) );
  OAI21_X1 U13938 ( .B1(n6591), .B2(n7046), .A(n11507), .ZN(n11369) );
  AOI21_X1 U13939 ( .B1(n11369), .B2(n13635), .A(n11368), .ZN(n14906) );
  INV_X1 U13940 ( .A(n14906), .ZN(n11378) );
  NOR2_X1 U13941 ( .A1(n14908), .A2(n11370), .ZN(n11371) );
  OR3_X1 U13942 ( .A1(n11513), .A2(n11371), .A3(n13620), .ZN(n14905) );
  OAI22_X1 U13943 ( .A1(n15210), .A2(n11373), .B1(n11372), .B2(n13651), .ZN(
        n11374) );
  AOI21_X1 U13944 ( .B1(n11375), .B2(n13654), .A(n11374), .ZN(n11376) );
  OAI21_X1 U13945 ( .B1(n14905), .B2(n13641), .A(n11376), .ZN(n11377) );
  AOI21_X1 U13946 ( .B1(n11378), .B2(n15210), .A(n11377), .ZN(n11379) );
  OAI21_X1 U13947 ( .B1(n13627), .B2(n14904), .A(n11379), .ZN(P2_U3254) );
  INV_X1 U13948 ( .A(n11380), .ZN(n11381) );
  AOI21_X1 U13949 ( .B1(n11383), .B2(n11382), .A(n11381), .ZN(n11388) );
  AOI22_X1 U13950 ( .A1(n6439), .A2(n12700), .B1(n12463), .B2(n14590), .ZN(
        n11385) );
  OAI211_X1 U13951 ( .C1(n12459), .C2(n15027), .A(n11385), .B(n11384), .ZN(
        n11386) );
  AOI21_X1 U13952 ( .B1(n11395), .B2(n12464), .A(n11386), .ZN(n11387) );
  OAI21_X1 U13953 ( .B1(n11388), .B2(n12471), .A(n11387), .ZN(P3_U3171) );
  AOI21_X1 U13954 ( .B1(n11389), .B2(n12572), .A(n12954), .ZN(n11394) );
  OAI22_X1 U13955 ( .A1(n11391), .A2(n12956), .B1(n11390), .B2(n12958), .ZN(
        n11392) );
  AOI21_X1 U13956 ( .B1(n11394), .B2(n11393), .A(n11392), .ZN(n15025) );
  INV_X1 U13957 ( .A(n11395), .ZN(n11396) );
  OAI22_X1 U13958 ( .A1(n15002), .A2(n11397), .B1(n11396), .B2(n14580), .ZN(
        n11398) );
  AOI21_X1 U13959 ( .B1(n12574), .B2(n12994), .A(n11398), .ZN(n11401) );
  XNOR2_X1 U13960 ( .A(n11399), .B(n12572), .ZN(n15030) );
  NAND2_X1 U13961 ( .A1(n15030), .A2(n14599), .ZN(n11400) );
  OAI211_X1 U13962 ( .C1(n15025), .C2(n15004), .A(n11401), .B(n11400), .ZN(
        P3_U3224) );
  NOR2_X1 U13963 ( .A1(n11413), .A2(n11402), .ZN(n11404) );
  INV_X1 U13964 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11405) );
  MUX2_X1 U13965 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n11405), .S(n11416), .Z(
        n11407) );
  INV_X1 U13966 ( .A(n11685), .ZN(n11406) );
  AOI21_X1 U13967 ( .B1(n11408), .B2(n11407), .A(n11406), .ZN(n11424) );
  MUX2_X1 U13968 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12799), .Z(n11704) );
  XOR2_X1 U13969 ( .A(n11416), .B(n11704), .Z(n11705) );
  XNOR2_X1 U13970 ( .A(n11707), .B(n11705), .ZN(n11422) );
  NOR2_X1 U13971 ( .A1(n11413), .A2(n11412), .ZN(n11415) );
  INV_X1 U13972 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11417) );
  MUX2_X1 U13973 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n11417), .S(n11416), .Z(
        n11691) );
  XNOR2_X1 U13974 ( .A(n11692), .B(n11691), .ZN(n11418) );
  NAND2_X1 U13975 ( .A1(n12710), .A2(n11418), .ZN(n11420) );
  AND2_X1 U13976 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11723) );
  AOI21_X1 U13977 ( .B1(n14923), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11723), 
        .ZN(n11419) );
  OAI211_X1 U13978 ( .C1(n14966), .C2(n11703), .A(n11420), .B(n11419), .ZN(
        n11421) );
  AOI21_X1 U13979 ( .B1(n14936), .B2(n11422), .A(n11421), .ZN(n11423) );
  OAI21_X1 U13980 ( .B1(n11424), .B2(n14977), .A(n11423), .ZN(P3_U3194) );
  AOI21_X1 U13981 ( .B1(n11426), .B2(n11425), .A(n6600), .ZN(n11433) );
  NAND2_X1 U13982 ( .A1(n11427), .A2(n14704), .ZN(n11428) );
  NAND2_X1 U13983 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n14137) );
  OAI211_X1 U13984 ( .C1(n14707), .C2(n11429), .A(n11428), .B(n14137), .ZN(
        n11430) );
  AOI21_X1 U13985 ( .B1(n11431), .B2(n14653), .A(n11430), .ZN(n11432) );
  OAI21_X1 U13986 ( .B1(n11433), .B2(n14699), .A(n11432), .ZN(P1_U3221) );
  XNOR2_X1 U13987 ( .A(n11435), .B(n11434), .ZN(n11441) );
  INV_X1 U13988 ( .A(n11436), .ZN(n11550) );
  INV_X1 U13989 ( .A(n13388), .ZN(n13631) );
  OAI22_X1 U13990 ( .A1(n13278), .A2(n13631), .B1(n12150), .B2(n13277), .ZN(
        n11437) );
  AOI211_X1 U13991 ( .C1(n13240), .C2(n11550), .A(n11438), .B(n11437), .ZN(
        n11440) );
  NAND2_X1 U13992 ( .A1(n12157), .A2(n13281), .ZN(n11439) );
  OAI211_X1 U13993 ( .C1(n11441), .C2(n13272), .A(n11440), .B(n11439), .ZN(
        P2_U3206) );
  INV_X1 U13994 ( .A(n11442), .ZN(n11443) );
  NAND2_X1 U13995 ( .A1(n11446), .A2(n11443), .ZN(n11444) );
  NAND2_X1 U13996 ( .A1(n11445), .A2(n11444), .ZN(n14744) );
  NAND2_X1 U13997 ( .A1(n14744), .A2(n14254), .ZN(n11454) );
  AOI21_X1 U13998 ( .B1(n11446), .B2(n6651), .A(n14795), .ZN(n11452) );
  OAI21_X1 U13999 ( .B1(n11449), .B2(n11448), .A(n11447), .ZN(n11456) );
  XNOR2_X1 U14000 ( .A(n11456), .B(n6450), .ZN(n11450) );
  AND2_X1 U14001 ( .A1(n11450), .A2(n14489), .ZN(n11451) );
  OAI22_X1 U14002 ( .A1(n11452), .A2(n14483), .B1(n11451), .B2(n6651), .ZN(
        n11453) );
  AND2_X1 U14003 ( .A1(n11454), .A2(n11453), .ZN(n14746) );
  OAI22_X1 U14004 ( .A1(n14377), .A2(n10040), .B1(n11455), .B2(n14374), .ZN(
        n11460) );
  INV_X1 U14005 ( .A(n14740), .ZN(n11458) );
  OR2_X1 U14006 ( .A1(n11456), .A2(n14355), .ZN(n14741) );
  OAI22_X1 U14007 ( .A1(n11458), .A2(n11457), .B1(n14387), .B2(n14741), .ZN(
        n11459) );
  AOI211_X1 U14008 ( .C1(n14384), .C2(n14738), .A(n11460), .B(n11459), .ZN(
        n11462) );
  NAND2_X1 U14009 ( .A1(n14744), .A2(n12049), .ZN(n11461) );
  OAI211_X1 U14010 ( .C1(n14325), .C2(n14746), .A(n11462), .B(n11461), .ZN(
        P1_U3292) );
  OAI222_X1 U14011 ( .A1(n8138), .A2(P1_U3086), .B1(n14534), .B2(n11538), .C1(
        n15074), .C2(n14528), .ZN(P1_U3335) );
  XNOR2_X1 U14012 ( .A(n11463), .B(n11465), .ZN(n15019) );
  OAI21_X1 U14013 ( .B1(n6711), .B2(n11465), .A(n11464), .ZN(n11467) );
  NAND2_X1 U14014 ( .A1(n11467), .A2(n14991), .ZN(n11469) );
  AOI22_X1 U14015 ( .A1(n12701), .A2(n14987), .B1(n14988), .B2(n12699), .ZN(
        n11468) );
  OAI211_X1 U14016 ( .C1(n14995), .C2(n15019), .A(n11469), .B(n11468), .ZN(
        n15020) );
  MUX2_X1 U14017 ( .A(n15020), .B(P3_REG2_REG_8__SCAN_IN), .S(n15004), .Z(
        n11470) );
  INV_X1 U14018 ( .A(n11470), .ZN(n11473) );
  INV_X1 U14019 ( .A(n11500), .ZN(n14598) );
  NOR2_X1 U14020 ( .A1(n11471), .A2(n15026), .ZN(n15021) );
  AOI22_X1 U14021 ( .A1(n14598), .A2(n15021), .B1(n14998), .B2(n12382), .ZN(
        n11472) );
  OAI211_X1 U14022 ( .C1(n15019), .C2(n11474), .A(n11473), .B(n11472), .ZN(
        P3_U3225) );
  OAI21_X1 U14023 ( .B1(n11476), .B2(n11477), .A(n11475), .ZN(n14786) );
  INV_X1 U14024 ( .A(n14786), .ZN(n11492) );
  OAI22_X1 U14025 ( .A1(n11764), .A2(n14474), .B1(n11627), .B2(n14400), .ZN(
        n11482) );
  NAND2_X1 U14026 ( .A1(n11478), .A2(n11477), .ZN(n11479) );
  AOI21_X1 U14027 ( .B1(n11480), .B2(n11479), .A(n14795), .ZN(n11481) );
  AOI211_X1 U14028 ( .C1(n14254), .C2(n14786), .A(n11482), .B(n11481), .ZN(
        n14788) );
  MUX2_X1 U14029 ( .A(n11483), .B(n14788), .S(n14377), .Z(n11491) );
  INV_X1 U14030 ( .A(n11484), .ZN(n11487) );
  INV_X1 U14031 ( .A(n11485), .ZN(n11486) );
  AOI211_X1 U14032 ( .C1(n11488), .C2(n11487), .A(n14355), .B(n11486), .ZN(
        n14783) );
  OAI22_X1 U14033 ( .A1(n11621), .A2(n14364), .B1(n11626), .B2(n14374), .ZN(
        n11489) );
  AOI21_X1 U14034 ( .B1(n14783), .B2(n14357), .A(n11489), .ZN(n11490) );
  OAI211_X1 U14035 ( .C1(n11492), .C2(n14262), .A(n11491), .B(n11490), .ZN(
        P1_U3284) );
  OAI211_X1 U14036 ( .C1(n11494), .C2(n12577), .A(n11493), .B(n14991), .ZN(
        n11496) );
  AOI22_X1 U14037 ( .A1(n14987), .A2(n12699), .B1(n14576), .B2(n14988), .ZN(
        n11495) );
  AND2_X1 U14038 ( .A1(n11496), .A2(n11495), .ZN(n15036) );
  INV_X1 U14039 ( .A(n12577), .ZN(n12501) );
  XNOR2_X1 U14040 ( .A(n11497), .B(n12501), .ZN(n15033) );
  NAND2_X1 U14041 ( .A1(n11498), .A2(n15015), .ZN(n15035) );
  AOI22_X1 U14042 ( .A1(n15004), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n14998), 
        .B2(n12364), .ZN(n11499) );
  OAI21_X1 U14043 ( .B1(n11500), .B2(n15035), .A(n11499), .ZN(n11501) );
  AOI21_X1 U14044 ( .B1(n15033), .B2(n14599), .A(n11501), .ZN(n11502) );
  OAI21_X1 U14045 ( .B1(n15036), .B2(n15004), .A(n11502), .ZN(P3_U3223) );
  NOR2_X1 U14046 ( .A1(n14908), .A2(n12141), .ZN(n11503) );
  NAND2_X1 U14047 ( .A1(n14908), .A2(n12141), .ZN(n11505) );
  XNOR2_X1 U14048 ( .A(n11540), .B(n13285), .ZN(n12313) );
  XNOR2_X1 U14049 ( .A(n11546), .B(n12313), .ZN(n14629) );
  OR2_X1 U14050 ( .A1(n14908), .A2(n13286), .ZN(n11506) );
  XNOR2_X1 U14051 ( .A(n11542), .B(n12313), .ZN(n11509) );
  OAI22_X1 U14052 ( .A1(n12158), .A2(n13632), .B1(n12141), .B2(n13630), .ZN(
        n11508) );
  AOI21_X1 U14053 ( .B1(n11509), .B2(n13635), .A(n11508), .ZN(n11510) );
  OAI21_X1 U14054 ( .B1(n14629), .B2(n10088), .A(n11510), .ZN(n14632) );
  NAND2_X1 U14055 ( .A1(n14632), .A2(n15210), .ZN(n11517) );
  OAI22_X1 U14056 ( .A1(n15210), .A2(n11512), .B1(n11511), .B2(n13651), .ZN(
        n11515) );
  OAI211_X1 U14057 ( .C1(n14631), .C2(n11513), .A(n13639), .B(n11549), .ZN(
        n14630) );
  NOR2_X1 U14058 ( .A1(n14630), .A2(n13641), .ZN(n11514) );
  AOI211_X1 U14059 ( .C1(n13654), .C2(n11540), .A(n11515), .B(n11514), .ZN(
        n11516) );
  OAI211_X1 U14060 ( .C1(n14629), .C2(n11518), .A(n11517), .B(n11516), .ZN(
        P2_U3253) );
  INV_X1 U14061 ( .A(n11524), .ZN(n11520) );
  AOI21_X1 U14062 ( .B1(n11520), .B2(P2_REG1_REG_14__SCAN_IN), .A(n11519), 
        .ZN(n11603) );
  INV_X1 U14063 ( .A(n11603), .ZN(n11521) );
  XNOR2_X1 U14064 ( .A(n11521), .B(n11596), .ZN(n11601) );
  XNOR2_X1 U14065 ( .A(n11601), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n11532) );
  NOR2_X1 U14066 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9270), .ZN(n11522) );
  AOI21_X1 U14067 ( .B1(n14859), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n11522), 
        .ZN(n11523) );
  OAI21_X1 U14068 ( .B1(n11602), .B2(n14820), .A(n11523), .ZN(n11531) );
  INV_X1 U14069 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11529) );
  NOR2_X1 U14070 ( .A1(n11525), .A2(n11524), .ZN(n11527) );
  XNOR2_X1 U14071 ( .A(n11593), .B(n11602), .ZN(n11528) );
  AOI211_X1 U14072 ( .C1(n11529), .C2(n11528), .A(n11825), .B(n11594), .ZN(
        n11530) );
  AOI211_X1 U14073 ( .C1(n14868), .C2(n11532), .A(n11531), .B(n11530), .ZN(
        n11533) );
  INV_X1 U14074 ( .A(n11533), .ZN(P2_U3229) );
  INV_X1 U14075 ( .A(n11534), .ZN(n11537) );
  INV_X1 U14076 ( .A(SI_25_), .ZN(n11535) );
  OAI222_X1 U14077 ( .A1(n13140), .A2(n11537), .B1(P3_U3151), .B2(n11536), 
        .C1(n11535), .C2(n13142), .ZN(P3_U3270) );
  OAI222_X1 U14078 ( .A1(n13803), .A2(n11539), .B1(P2_U3088), .B2(n12331), 
        .C1(n13800), .C2(n11538), .ZN(P2_U3307) );
  NOR2_X1 U14079 ( .A1(n14631), .A2(n13285), .ZN(n11541) );
  XNOR2_X1 U14080 ( .A(n12157), .B(n13284), .ZN(n12312) );
  XNOR2_X1 U14081 ( .A(n11556), .B(n12312), .ZN(n11544) );
  OAI222_X1 U14082 ( .A1(n13632), .A2(n13631), .B1(n13630), .B2(n12150), .C1(
        n11544), .C2(n11543), .ZN(n11642) );
  INV_X1 U14083 ( .A(n11642), .ZN(n11555) );
  AND2_X1 U14084 ( .A1(n14631), .A2(n12150), .ZN(n11545) );
  OR2_X1 U14085 ( .A1(n14631), .A2(n12150), .ZN(n11547) );
  XNOR2_X1 U14086 ( .A(n11564), .B(n12312), .ZN(n11644) );
  INV_X1 U14087 ( .A(n12157), .ZN(n12159) );
  INV_X1 U14088 ( .A(n11566), .ZN(n11548) );
  AOI211_X1 U14089 ( .C1(n12157), .C2(n11549), .A(n13620), .B(n11548), .ZN(
        n11643) );
  NAND2_X1 U14090 ( .A1(n11643), .A2(n13658), .ZN(n11552) );
  INV_X1 U14091 ( .A(n13651), .ZN(n15200) );
  AOI22_X1 U14092 ( .A1(n13649), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11550), 
        .B2(n15200), .ZN(n11551) );
  OAI211_X1 U14093 ( .C1(n12159), .C2(n13603), .A(n11552), .B(n11551), .ZN(
        n11553) );
  AOI21_X1 U14094 ( .B1(n13656), .B2(n11644), .A(n11553), .ZN(n11554) );
  OAI21_X1 U14095 ( .B1(n11555), .B2(n13649), .A(n11554), .ZN(P2_U3252) );
  OR2_X1 U14096 ( .A1(n12157), .A2(n12158), .ZN(n11557) );
  NAND2_X1 U14097 ( .A1(n14620), .A2(n13631), .ZN(n13348) );
  OR2_X1 U14098 ( .A1(n14620), .A2(n13631), .ZN(n11558) );
  NAND2_X1 U14099 ( .A1(n11559), .A2(n11565), .ZN(n11560) );
  NAND2_X1 U14100 ( .A1(n13349), .A2(n11560), .ZN(n11562) );
  OAI22_X1 U14101 ( .A1(n13389), .A2(n13632), .B1(n12158), .B2(n13630), .ZN(
        n11561) );
  AOI21_X1 U14102 ( .B1(n11562), .B2(n13635), .A(n11561), .ZN(n14627) );
  AND2_X1 U14103 ( .A1(n12157), .A2(n13284), .ZN(n11563) );
  XNOR2_X1 U14104 ( .A(n13387), .B(n11565), .ZN(n14624) );
  AND2_X1 U14105 ( .A1(n14620), .A2(n11566), .ZN(n11567) );
  OR3_X1 U14106 ( .A1(n13640), .A2(n11567), .A3(n13620), .ZN(n14622) );
  AOI22_X1 U14107 ( .A1(n13649), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11614), 
        .B2(n15200), .ZN(n11569) );
  NAND2_X1 U14108 ( .A1(n14620), .A2(n13654), .ZN(n11568) );
  OAI211_X1 U14109 ( .C1(n14622), .C2(n13641), .A(n11569), .B(n11568), .ZN(
        n11570) );
  AOI21_X1 U14110 ( .B1(n14624), .B2(n13656), .A(n11570), .ZN(n11571) );
  OAI21_X1 U14111 ( .B1(n14627), .B2(n13649), .A(n11571), .ZN(P2_U3251) );
  OAI222_X1 U14112 ( .A1(n11573), .A2(P1_U3086), .B1(n14534), .B2(n11574), 
        .C1(n11572), .C2(n14528), .ZN(P1_U3334) );
  OAI222_X1 U14113 ( .A1(n13803), .A2(n15180), .B1(P2_U3088), .B2(n12329), 
        .C1(n13800), .C2(n11574), .ZN(P2_U3306) );
  XNOR2_X1 U14114 ( .A(n11668), .B(n11666), .ZN(n11577) );
  NAND2_X1 U14115 ( .A1(n11577), .A2(n14489), .ZN(n11579) );
  AOI22_X1 U14116 ( .A1(n14483), .A2(n14034), .B1(n14032), .B2(n14739), .ZN(
        n11578) );
  NAND2_X1 U14117 ( .A1(n11579), .A2(n11578), .ZN(n14670) );
  INV_X1 U14118 ( .A(n14670), .ZN(n11588) );
  OR2_X1 U14119 ( .A1(n14792), .A2(n14034), .ZN(n11580) );
  OAI21_X1 U14120 ( .B1(n11582), .B2(n11666), .A(n11672), .ZN(n14672) );
  OAI211_X1 U14121 ( .C1(n14669), .C2(n6598), .A(n14370), .B(n11741), .ZN(
        n14668) );
  OAI22_X1 U14122 ( .A1(n14377), .A2(n11583), .B1(n11763), .B2(n14374), .ZN(
        n11584) );
  AOI21_X1 U14123 ( .B1(n11768), .B2(n14384), .A(n11584), .ZN(n11585) );
  OAI21_X1 U14124 ( .B1(n14668), .B2(n14387), .A(n11585), .ZN(n11586) );
  AOI21_X1 U14125 ( .B1(n14672), .B2(n14337), .A(n11586), .ZN(n11587) );
  OAI21_X1 U14126 ( .B1(n11588), .B2(n14325), .A(n11587), .ZN(P1_U3282) );
  INV_X1 U14127 ( .A(n11589), .ZN(n11590) );
  OAI222_X1 U14128 ( .A1(n11592), .A2(P3_U3151), .B1(n13142), .B2(n11591), 
        .C1(n13140), .C2(n11590), .ZN(P3_U3269) );
  INV_X1 U14129 ( .A(n11593), .ZN(n11595) );
  NAND2_X1 U14130 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n11832), .ZN(n11597) );
  OAI21_X1 U14131 ( .B1(n11832), .B2(P2_REG2_REG_16__SCAN_IN), .A(n11597), 
        .ZN(n11598) );
  NOR2_X1 U14132 ( .A1(n11599), .A2(n11598), .ZN(n11824) );
  AOI211_X1 U14133 ( .C1(n11599), .C2(n11598), .A(n11824), .B(n11825), .ZN(
        n11611) );
  INV_X1 U14134 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11600) );
  OAI22_X1 U14135 ( .A1(n11603), .A2(n11602), .B1(n11601), .B2(n11600), .ZN(
        n11605) );
  XOR2_X1 U14136 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n11832), .Z(n11604) );
  NAND2_X1 U14137 ( .A1(n11604), .A2(n11605), .ZN(n11830) );
  OAI211_X1 U14138 ( .C1(n11605), .C2(n11604), .A(n14868), .B(n11830), .ZN(
        n11608) );
  NOR2_X1 U14139 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13198), .ZN(n11606) );
  AOI21_X1 U14140 ( .B1(n14859), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11606), 
        .ZN(n11607) );
  OAI211_X1 U14141 ( .C1(n14820), .C2(n11609), .A(n11608), .B(n11607), .ZN(
        n11610) );
  OR2_X1 U14142 ( .A1(n11611), .A2(n11610), .ZN(P2_U3230) );
  AOI21_X1 U14143 ( .B1(n11613), .B2(n11612), .A(n6601), .ZN(n11620) );
  INV_X1 U14144 ( .A(n11614), .ZN(n11617) );
  AOI22_X1 U14145 ( .A1(n13265), .A2(n13284), .B1(n13261), .B2(n13350), .ZN(
        n11616) );
  OAI211_X1 U14146 ( .C1(n11617), .C2(n13276), .A(n11616), .B(n11615), .ZN(
        n11618) );
  AOI21_X1 U14147 ( .B1(n14620), .B2(n13281), .A(n11618), .ZN(n11619) );
  OAI21_X1 U14148 ( .B1(n11620), .B2(n13272), .A(n11619), .ZN(P2_U3187) );
  INV_X1 U14149 ( .A(n14697), .ZN(n13908) );
  OR2_X1 U14150 ( .A1(n11621), .A2(n14775), .ZN(n14782) );
  OAI21_X1 U14151 ( .B1(n11624), .B2(n11623), .A(n11651), .ZN(n11625) );
  NAND2_X1 U14152 ( .A1(n11625), .A2(n14655), .ZN(n11631) );
  INV_X1 U14153 ( .A(n14707), .ZN(n13982) );
  INV_X1 U14154 ( .A(n11626), .ZN(n11629) );
  AND2_X1 U14155 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14153) );
  OAI22_X1 U14156 ( .A1(n11764), .A2(n13975), .B1(n13974), .B2(n11627), .ZN(
        n11628) );
  AOI211_X1 U14157 ( .C1(n13982), .C2(n11629), .A(n14153), .B(n11628), .ZN(
        n11630) );
  OAI211_X1 U14158 ( .C1(n13908), .C2(n14782), .A(n11631), .B(n11630), .ZN(
        P1_U3231) );
  NAND2_X1 U14159 ( .A1(n11633), .A2(n11632), .ZN(n11634) );
  XNOR2_X1 U14160 ( .A(n11634), .B(n12362), .ZN(n11641) );
  AOI21_X1 U14161 ( .B1(n6439), .B2(n14590), .A(n11635), .ZN(n11637) );
  NAND2_X1 U14162 ( .A1(n12464), .A2(n14593), .ZN(n11636) );
  OAI211_X1 U14163 ( .C1(n11818), .C2(n12455), .A(n11637), .B(n11636), .ZN(
        n11638) );
  AOI21_X1 U14164 ( .B1(n11639), .B2(n12469), .A(n11638), .ZN(n11640) );
  OAI21_X1 U14165 ( .B1(n11641), .B2(n12471), .A(n11640), .ZN(P3_U3176) );
  AOI211_X1 U14166 ( .C1(n14623), .C2(n11644), .A(n11643), .B(n11642), .ZN(
        n11649) );
  INV_X1 U14167 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11645) );
  OAI22_X1 U14168 ( .A1(n12159), .A2(n13780), .B1(n14915), .B2(n11645), .ZN(
        n11646) );
  INV_X1 U14169 ( .A(n11646), .ZN(n11647) );
  OAI21_X1 U14170 ( .B1(n11649), .B2(n14913), .A(n11647), .ZN(P2_U3469) );
  AOI22_X1 U14171 ( .A1(n12157), .A2(n13742), .B1(n14920), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n11648) );
  OAI21_X1 U14172 ( .B1(n11649), .B2(n14920), .A(n11648), .ZN(P2_U3512) );
  INV_X1 U14173 ( .A(n14792), .ZN(n11662) );
  AND2_X1 U14174 ( .A1(n11651), .A2(n11650), .ZN(n11654) );
  OAI211_X1 U14175 ( .C1(n11654), .C2(n11653), .A(n14655), .B(n11652), .ZN(
        n11661) );
  OAI21_X1 U14176 ( .B1(n11656), .B2(n14400), .A(n11655), .ZN(n14791) );
  OAI21_X1 U14177 ( .B1(n14707), .B2(n11658), .A(n11657), .ZN(n11659) );
  AOI21_X1 U14178 ( .B1(n14704), .B2(n14791), .A(n11659), .ZN(n11660) );
  OAI211_X1 U14179 ( .C1(n11662), .C2(n14015), .A(n11661), .B(n11660), .ZN(
        P1_U3217) );
  INV_X1 U14180 ( .A(n11663), .ZN(n11665) );
  OAI222_X1 U14181 ( .A1(n7491), .A2(P3_U3151), .B1(n13140), .B2(n11665), .C1(
        n11664), .C2(n13142), .ZN(P3_U3268) );
  INV_X1 U14182 ( .A(n11666), .ZN(n11667) );
  NAND2_X1 U14183 ( .A1(n11736), .A2(n11735), .ZN(n11670) );
  INV_X1 U14184 ( .A(n14032), .ZN(n11765) );
  OR2_X1 U14185 ( .A1(n11889), .A2(n11765), .ZN(n11669) );
  NAND2_X1 U14186 ( .A1(n11670), .A2(n11669), .ZN(n11781) );
  INV_X1 U14187 ( .A(n11780), .ZN(n11674) );
  XNOR2_X1 U14188 ( .A(n11781), .B(n11674), .ZN(n11671) );
  OAI22_X1 U14189 ( .A1(n11791), .A2(n14474), .B1(n11765), .B2(n14400), .ZN(
        n11946) );
  AOI21_X1 U14190 ( .B1(n11671), .B2(n14489), .A(n11946), .ZN(n11774) );
  INV_X1 U14191 ( .A(n11735), .ZN(n11733) );
  NAND2_X1 U14192 ( .A1(n11734), .A2(n11733), .ZN(n11732) );
  OR2_X1 U14193 ( .A1(n11889), .A2(n14032), .ZN(n11673) );
  NAND2_X1 U14194 ( .A1(n11732), .A2(n11673), .ZN(n11675) );
  OAI21_X1 U14195 ( .B1(n11675), .B2(n11674), .A(n11787), .ZN(n11771) );
  INV_X1 U14196 ( .A(n11677), .ZN(n11740) );
  INV_X1 U14197 ( .A(n11805), .ZN(n11676) );
  AOI21_X1 U14198 ( .B1(n11951), .B2(n11677), .A(n11676), .ZN(n11772) );
  NAND3_X1 U14199 ( .A1(n11772), .A2(n14370), .A3(n14357), .ZN(n11680) );
  INV_X1 U14200 ( .A(n11949), .ZN(n11678) );
  AOI22_X1 U14201 ( .A1(n14325), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n11678), 
        .B2(n14323), .ZN(n11679) );
  OAI211_X1 U14202 ( .C1(n11681), .C2(n14364), .A(n11680), .B(n11679), .ZN(
        n11682) );
  AOI21_X1 U14203 ( .B1(n11771), .B2(n14337), .A(n11682), .ZN(n11683) );
  OAI21_X1 U14204 ( .B1(n14325), .B2(n11774), .A(n11683), .ZN(P1_U3280) );
  NAND2_X1 U14205 ( .A1(n11703), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n11684) );
  NOR2_X1 U14206 ( .A1(n11695), .A2(n11686), .ZN(n11687) );
  INV_X1 U14207 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14971) );
  NAND2_X1 U14208 ( .A1(n11700), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12723) );
  INV_X1 U14209 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U14210 ( .A1(n11698), .A2(n11941), .ZN(n11688) );
  NAND2_X1 U14211 ( .A1(n12723), .A2(n11688), .ZN(n11701) );
  INV_X1 U14212 ( .A(n12717), .ZN(n11689) );
  AOI21_X1 U14213 ( .B1(n11690), .B2(n11701), .A(n11689), .ZN(n11719) );
  NAND2_X1 U14214 ( .A1(n11703), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n11693) );
  INV_X1 U14215 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14964) );
  NAND2_X1 U14216 ( .A1(n11700), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12736) );
  INV_X1 U14217 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11697) );
  NAND2_X1 U14218 ( .A1(n11698), .A2(n11697), .ZN(n11699) );
  NAND2_X1 U14219 ( .A1(n12736), .A2(n11699), .ZN(n12734) );
  XNOR2_X1 U14220 ( .A(n12735), .B(n12734), .ZN(n11717) );
  NOR2_X1 U14221 ( .A1(n14966), .A2(n11700), .ZN(n11716) );
  INV_X1 U14222 ( .A(n14923), .ZN(n14967) );
  MUX2_X1 U14223 ( .A(n12734), .B(n11701), .S(n12799), .Z(n11710) );
  MUX2_X1 U14224 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12799), .Z(n11702) );
  NOR2_X1 U14225 ( .A1(n11702), .A2(n14965), .ZN(n11711) );
  XNOR2_X1 U14226 ( .A(n11702), .B(n14965), .ZN(n14974) );
  NAND2_X1 U14227 ( .A1(n11704), .A2(n11703), .ZN(n11709) );
  INV_X1 U14228 ( .A(n11705), .ZN(n11706) );
  NAND2_X1 U14229 ( .A1(n11707), .A2(n11706), .ZN(n11708) );
  NAND2_X1 U14230 ( .A1(n11709), .A2(n11708), .ZN(n14973) );
  NOR2_X1 U14231 ( .A1(n14974), .A2(n14973), .ZN(n14972) );
  OR3_X2 U14232 ( .A1(n11710), .A2(n11711), .A3(n14972), .ZN(n12725) );
  OAI21_X1 U14233 ( .B1(n11711), .B2(n14972), .A(n11710), .ZN(n11712) );
  NAND3_X1 U14234 ( .A1(n14936), .A2(n12725), .A3(n11712), .ZN(n11713) );
  NAND2_X1 U14235 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n11882)
         );
  OAI211_X1 U14236 ( .C1(n14967), .C2(n11714), .A(n11713), .B(n11882), .ZN(
        n11715) );
  AOI211_X1 U14237 ( .C1(n12710), .C2(n11717), .A(n11716), .B(n11715), .ZN(
        n11718) );
  OAI21_X1 U14238 ( .B1(n11719), .B2(n14977), .A(n11718), .ZN(P3_U3196) );
  XNOR2_X1 U14239 ( .A(n11720), .B(n14591), .ZN(n11721) );
  XNOR2_X1 U14240 ( .A(n11722), .B(n11721), .ZN(n11730) );
  NAND2_X1 U14241 ( .A1(n14585), .A2(n12469), .ZN(n11728) );
  AOI21_X1 U14242 ( .B1(n6439), .B2(n14576), .A(n11723), .ZN(n11727) );
  NAND2_X1 U14243 ( .A1(n12464), .A2(n11724), .ZN(n11726) );
  NAND2_X1 U14244 ( .A1(n12463), .A2(n14577), .ZN(n11725) );
  NAND4_X1 U14245 ( .A1(n11728), .A2(n11727), .A3(n11726), .A4(n11725), .ZN(
        n11729) );
  AOI21_X1 U14246 ( .B1(n11730), .B2(n12449), .A(n11729), .ZN(n11731) );
  INV_X1 U14247 ( .A(n11731), .ZN(P3_U3164) );
  OAI21_X1 U14248 ( .B1(n11734), .B2(n11733), .A(n11732), .ZN(n11887) );
  OAI22_X1 U14249 ( .A1(n11872), .A2(n14400), .B1(n11873), .B2(n14474), .ZN(
        n11739) );
  XNOR2_X1 U14250 ( .A(n11736), .B(n11735), .ZN(n11737) );
  NOR2_X1 U14251 ( .A1(n11737), .A2(n14795), .ZN(n11738) );
  AOI211_X1 U14252 ( .C1(n14254), .C2(n11887), .A(n11739), .B(n11738), .ZN(
        n11891) );
  AOI211_X1 U14253 ( .C1(n11889), .C2(n11741), .A(n14355), .B(n11740), .ZN(
        n11888) );
  NAND2_X1 U14254 ( .A1(n11888), .A2(n14357), .ZN(n11744) );
  INV_X1 U14255 ( .A(n11742), .ZN(n11876) );
  AOI22_X1 U14256 ( .A1(n14325), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11876), 
        .B2(n14323), .ZN(n11743) );
  OAI211_X1 U14257 ( .C1(n6855), .C2(n14364), .A(n11744), .B(n11743), .ZN(
        n11745) );
  AOI21_X1 U14258 ( .B1(n11887), .B2(n12049), .A(n11745), .ZN(n11746) );
  OAI21_X1 U14259 ( .B1(n11891), .B2(n14325), .A(n11746), .ZN(P1_U3281) );
  OAI222_X1 U14260 ( .A1(n13803), .A2(n11748), .B1(P2_U3088), .B2(n6756), .C1(
        n13800), .C2(n11747), .ZN(P2_U3305) );
  NAND2_X1 U14261 ( .A1(n11750), .A2(n11749), .ZN(n11752) );
  XOR2_X1 U14262 ( .A(n11752), .B(n11751), .Z(n11759) );
  INV_X1 U14263 ( .A(n11753), .ZN(n11819) );
  NOR2_X1 U14264 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11754), .ZN(n14981) );
  NOR2_X1 U14265 ( .A1(n12455), .A2(n12603), .ZN(n11755) );
  AOI211_X1 U14266 ( .C1(n6439), .C2(n14591), .A(n14981), .B(n11755), .ZN(
        n11756) );
  OAI21_X1 U14267 ( .B1(n11819), .B2(n12438), .A(n11756), .ZN(n11757) );
  AOI21_X1 U14268 ( .B1(n11821), .B2(n12469), .A(n11757), .ZN(n11758) );
  OAI21_X1 U14269 ( .B1(n11759), .B2(n12471), .A(n11758), .ZN(P3_U3174) );
  AOI21_X1 U14270 ( .B1(n11761), .B2(n11760), .A(n6590), .ZN(n11770) );
  OAI21_X1 U14271 ( .B1(n14707), .B2(n11763), .A(n11762), .ZN(n11767) );
  OAI22_X1 U14272 ( .A1(n11765), .A2(n13975), .B1(n13974), .B2(n11764), .ZN(
        n11766) );
  AOI211_X1 U14273 ( .C1(n11768), .C2(n14653), .A(n11767), .B(n11766), .ZN(
        n11769) );
  OAI21_X1 U14274 ( .B1(n11770), .B2(n14699), .A(n11769), .ZN(P1_U3236) );
  INV_X1 U14275 ( .A(n11771), .ZN(n11775) );
  AOI22_X1 U14276 ( .A1(n11772), .A2(n14370), .B1(n14793), .B2(n11951), .ZN(
        n11773) );
  OAI211_X1 U14277 ( .C1(n11775), .C2(n14753), .A(n11774), .B(n11773), .ZN(
        n11777) );
  NAND2_X1 U14278 ( .A1(n11777), .A2(n14802), .ZN(n11776) );
  OAI21_X1 U14279 ( .B1(n14802), .B2(n8386), .A(n11776), .ZN(P1_U3498) );
  NAND2_X1 U14280 ( .A1(n11777), .A2(n14813), .ZN(n11778) );
  OAI21_X1 U14281 ( .B1(n14813), .B2(n11779), .A(n11778), .ZN(P1_U3541) );
  NAND2_X1 U14282 ( .A1(n11781), .A2(n11780), .ZN(n11783) );
  OR2_X1 U14283 ( .A1(n11951), .A2(n11873), .ZN(n11782) );
  NAND2_X1 U14284 ( .A1(n11783), .A2(n11782), .ZN(n11798) );
  NAND2_X1 U14285 ( .A1(n11798), .A2(n11800), .ZN(n11785) );
  NAND2_X1 U14286 ( .A1(n11785), .A2(n11784), .ZN(n11915) );
  XNOR2_X1 U14287 ( .A(n11915), .B(n7120), .ZN(n14665) );
  OR2_X1 U14288 ( .A1(n11951), .A2(n14031), .ZN(n11786) );
  NAND2_X1 U14289 ( .A1(n14643), .A2(n14030), .ZN(n11789) );
  XNOR2_X1 U14290 ( .A(n11926), .B(n7120), .ZN(n14667) );
  NAND2_X1 U14291 ( .A1(n14667), .A2(n14337), .ZN(n11797) );
  INV_X1 U14292 ( .A(n11919), .ZN(n11790) );
  AOI211_X1 U14293 ( .C1(n14663), .C2(n6587), .A(n14355), .B(n11790), .ZN(
        n14661) );
  OAI22_X1 U14294 ( .A1(n14382), .A2(n14474), .B1(n11791), .B2(n14400), .ZN(
        n14662) );
  INV_X1 U14295 ( .A(n14662), .ZN(n11792) );
  OAI22_X1 U14296 ( .A1(n11792), .A2(n14325), .B1(n14014), .B2(n14374), .ZN(
        n11793) );
  AOI21_X1 U14297 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14325), .A(n11793), 
        .ZN(n11794) );
  OAI21_X1 U14298 ( .B1(n14016), .B2(n14364), .A(n11794), .ZN(n11795) );
  AOI21_X1 U14299 ( .B1(n14661), .B2(n14357), .A(n11795), .ZN(n11796) );
  OAI211_X1 U14300 ( .C1(n14665), .C2(n14346), .A(n11797), .B(n11796), .ZN(
        P1_U3278) );
  XOR2_X1 U14301 ( .A(n11800), .B(n11798), .Z(n11799) );
  OAI22_X1 U14302 ( .A1(n11873), .A2(n14400), .B1(n11920), .B2(n14474), .ZN(
        n14645) );
  AOI21_X1 U14303 ( .B1(n11799), .B2(n14489), .A(n14645), .ZN(n11899) );
  OAI21_X1 U14304 ( .B1(n11802), .B2(n11788), .A(n11801), .ZN(n11900) );
  OAI22_X1 U14305 ( .A1(n14377), .A2(n11803), .B1(n14648), .B2(n14374), .ZN(
        n11804) );
  AOI21_X1 U14306 ( .B1(n14643), .B2(n14384), .A(n11804), .ZN(n11808) );
  AOI21_X1 U14307 ( .B1(n14643), .B2(n11805), .A(n14355), .ZN(n11806) );
  AND2_X1 U14308 ( .A1(n11806), .A2(n6587), .ZN(n11897) );
  NAND2_X1 U14309 ( .A1(n11897), .A2(n14357), .ZN(n11807) );
  OAI211_X1 U14310 ( .C1(n11900), .C2(n14391), .A(n11808), .B(n11807), .ZN(
        n11809) );
  INV_X1 U14311 ( .A(n11809), .ZN(n11810) );
  OAI21_X1 U14312 ( .B1(n14325), .B2(n11899), .A(n11810), .ZN(P1_U3279) );
  INV_X1 U14313 ( .A(n11811), .ZN(n11812) );
  OAI222_X1 U14314 ( .A1(P3_U3151), .A2(n6710), .B1(n13142), .B2(n11813), .C1(
        n13140), .C2(n11812), .ZN(P3_U3267) );
  INV_X1 U14315 ( .A(n12594), .ZN(n11814) );
  XNOR2_X1 U14316 ( .A(n11815), .B(n12506), .ZN(n14604) );
  XNOR2_X1 U14317 ( .A(n11816), .B(n12506), .ZN(n11817) );
  OAI222_X1 U14318 ( .A1(n12956), .A2(n11818), .B1(n12958), .B2(n12603), .C1(
        n11817), .C2(n12954), .ZN(n14606) );
  NAND2_X1 U14319 ( .A1(n14606), .A2(n15002), .ZN(n11823) );
  OAI22_X1 U14320 ( .A1(n15002), .A2(n14964), .B1(n11819), .B2(n14580), .ZN(
        n11820) );
  AOI21_X1 U14321 ( .B1(n11821), .B2(n12994), .A(n11820), .ZN(n11822) );
  OAI211_X1 U14322 ( .C1(n12997), .C2(n14604), .A(n11823), .B(n11822), .ZN(
        P3_U3220) );
  AOI21_X1 U14323 ( .B1(n11832), .B2(P2_REG2_REG_16__SCAN_IN), .A(n11824), 
        .ZN(n11827) );
  XNOR2_X1 U14324 ( .A(n13313), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n11826) );
  NOR2_X1 U14325 ( .A1(n11827), .A2(n11826), .ZN(n13312) );
  AOI211_X1 U14326 ( .C1(n11827), .C2(n11826), .A(n13312), .B(n11825), .ZN(
        n11829) );
  NOR2_X1 U14327 ( .A1(n11828), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13210) );
  NOR2_X1 U14328 ( .A1(n11829), .A2(n13210), .ZN(n11835) );
  XNOR2_X1 U14329 ( .A(n13313), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n13319) );
  INV_X1 U14330 ( .A(n11830), .ZN(n11831) );
  AOI21_X1 U14331 ( .B1(n11832), .B2(P2_REG1_REG_16__SCAN_IN), .A(n11831), 
        .ZN(n13320) );
  XOR2_X1 U14332 ( .A(n13319), .B(n13320), .Z(n11833) );
  AOI22_X1 U14333 ( .A1(n14859), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(n14868), 
        .B2(n11833), .ZN(n11834) );
  OAI211_X1 U14334 ( .C1(n13318), .C2(n14820), .A(n11835), .B(n11834), .ZN(
        P2_U3231) );
  INV_X1 U14335 ( .A(n11862), .ZN(n11838) );
  AOI21_X1 U14336 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n13790), .A(n12339), 
        .ZN(n11837) );
  OAI21_X1 U14337 ( .B1(n11838), .B2(n13800), .A(n11837), .ZN(P2_U3304) );
  NOR2_X1 U14338 ( .A1(n11849), .A2(n11839), .ZN(n11841) );
  INV_X1 U14339 ( .A(n14165), .ZN(n11843) );
  XNOR2_X1 U14340 ( .A(n14168), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14164) );
  INV_X1 U14341 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11842) );
  OAI22_X1 U14342 ( .A1(n11843), .A2(n14164), .B1(n11842), .B2(n11853), .ZN(
        n14720) );
  INV_X1 U14343 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11844) );
  XNOR2_X1 U14344 ( .A(n14721), .B(n11844), .ZN(n14719) );
  XNOR2_X1 U14345 ( .A(n14176), .B(n14184), .ZN(n11845) );
  NAND2_X1 U14346 ( .A1(n11845), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14178) );
  OAI211_X1 U14347 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11845), .A(n14194), 
        .B(n14178), .ZN(n11846) );
  NAND2_X1 U14348 ( .A1(n11847), .A2(n11846), .ZN(n11857) );
  XOR2_X1 U14349 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n14721), .Z(n14725) );
  NOR2_X1 U14350 ( .A1(n11849), .A2(n11848), .ZN(n11851) );
  NOR2_X1 U14351 ( .A1(n11851), .A2(n11850), .ZN(n14172) );
  NAND2_X1 U14352 ( .A1(n14168), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11852) );
  OAI211_X1 U14353 ( .C1(n14168), .C2(P1_REG2_REG_16__SCAN_IN), .A(n14172), 
        .B(n11852), .ZN(n14170) );
  OAI21_X1 U14354 ( .B1(n11853), .B2(n14169), .A(n14170), .ZN(n14726) );
  NAND2_X1 U14355 ( .A1(n14725), .A2(n14726), .ZN(n14723) );
  OAI21_X1 U14356 ( .B1(n11854), .B2(n14376), .A(n14723), .ZN(n14185) );
  XNOR2_X1 U14357 ( .A(n14185), .B(n14184), .ZN(n14182) );
  INV_X1 U14358 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14359) );
  XNOR2_X1 U14359 ( .A(n14182), .B(n14359), .ZN(n11855) );
  NOR2_X1 U14360 ( .A1(n14190), .A2(n11855), .ZN(n11856) );
  AOI211_X1 U14361 ( .C1(n14733), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n11857), 
        .B(n11856), .ZN(n11858) );
  OAI21_X1 U14362 ( .B1(n11860), .B2(n11859), .A(n11858), .ZN(P1_U3261) );
  NAND2_X1 U14363 ( .A1(n11862), .A2(n11861), .ZN(n11864) );
  OAI211_X1 U14364 ( .C1(n11865), .C2(n14528), .A(n11864), .B(n11863), .ZN(
        P1_U3332) );
  INV_X1 U14365 ( .A(n11866), .ZN(n11870) );
  OAI21_X1 U14366 ( .B1(n6590), .B2(n11868), .A(n11867), .ZN(n11869) );
  NAND3_X1 U14367 ( .A1(n11870), .A2(n14655), .A3(n11869), .ZN(n11878) );
  INV_X1 U14368 ( .A(n11871), .ZN(n11875) );
  OAI22_X1 U14369 ( .A1(n11873), .A2(n13975), .B1(n13974), .B2(n11872), .ZN(
        n11874) );
  AOI211_X1 U14370 ( .C1(n11876), .C2(n13982), .A(n11875), .B(n11874), .ZN(
        n11877) );
  OAI211_X1 U14371 ( .C1(n6855), .C2(n14015), .A(n11878), .B(n11877), .ZN(
        P1_U3224) );
  INV_X1 U14372 ( .A(n12602), .ZN(n12601) );
  OAI211_X1 U14373 ( .C1(n11881), .C2(n11880), .A(n11879), .B(n12449), .ZN(
        n11886) );
  NAND2_X1 U14374 ( .A1(n6439), .A2(n14577), .ZN(n11883) );
  OAI211_X1 U14375 ( .C1(n12409), .C2(n12455), .A(n11883), .B(n11882), .ZN(
        n11884) );
  AOI21_X1 U14376 ( .B1(n11958), .B2(n12464), .A(n11884), .ZN(n11885) );
  OAI211_X1 U14377 ( .C1(n12601), .C2(n12459), .A(n11886), .B(n11885), .ZN(
        P3_U3155) );
  INV_X1 U14378 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11894) );
  INV_X1 U14379 ( .A(n11887), .ZN(n11892) );
  AOI21_X1 U14380 ( .B1(n14793), .B2(n11889), .A(n11888), .ZN(n11890) );
  OAI211_X1 U14381 ( .C1(n11892), .C2(n14430), .A(n11891), .B(n11890), .ZN(
        n11895) );
  NAND2_X1 U14382 ( .A1(n11895), .A2(n14802), .ZN(n11893) );
  OAI21_X1 U14383 ( .B1(n14802), .B2(n11894), .A(n11893), .ZN(P1_U3495) );
  NAND2_X1 U14384 ( .A1(n11895), .A2(n14813), .ZN(n11896) );
  OAI21_X1 U14385 ( .B1(n14813), .B2(n8356), .A(n11896), .ZN(P1_U3540) );
  AOI21_X1 U14386 ( .B1(n14793), .B2(n14643), .A(n11897), .ZN(n11898) );
  OAI211_X1 U14387 ( .C1(n11900), .C2(n14753), .A(n11899), .B(n11898), .ZN(
        n11902) );
  NAND2_X1 U14388 ( .A1(n11902), .A2(n14802), .ZN(n11901) );
  OAI21_X1 U14389 ( .B1(n14802), .B2(n8421), .A(n11901), .ZN(P1_U3501) );
  NAND2_X1 U14390 ( .A1(n11902), .A2(n14813), .ZN(n11903) );
  OAI21_X1 U14391 ( .B1(n14813), .B2(n11904), .A(n11903), .ZN(P1_U3542) );
  XNOR2_X1 U14392 ( .A(n11905), .B(n12409), .ZN(n11906) );
  XNOR2_X1 U14393 ( .A(n6712), .B(n11906), .ZN(n11913) );
  NOR2_X1 U14394 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11908), .ZN(n14572) );
  AOI21_X1 U14395 ( .B1(n6439), .B2(n12990), .A(n14572), .ZN(n11910) );
  NAND2_X1 U14396 ( .A1(n12464), .A2(n12993), .ZN(n11909) );
  OAI211_X1 U14397 ( .C1(n7077), .C2(n12455), .A(n11910), .B(n11909), .ZN(
        n11911) );
  AOI21_X1 U14398 ( .B1(n13122), .B2(n12469), .A(n11911), .ZN(n11912) );
  OAI21_X1 U14399 ( .B1(n11913), .B2(n12471), .A(n11912), .ZN(P3_U3181) );
  NAND2_X1 U14400 ( .A1(n11915), .A2(n7120), .ZN(n11916) );
  INV_X1 U14401 ( .A(n11965), .ZN(n11917) );
  AOI21_X1 U14402 ( .B1(n11930), .B2(n11918), .A(n11917), .ZN(n14497) );
  AOI211_X1 U14403 ( .C1(n14654), .C2(n11919), .A(n14355), .B(n14372), .ZN(
        n14493) );
  OAI22_X1 U14404 ( .A1(n14350), .A2(n14474), .B1(n11920), .B2(n14400), .ZN(
        n14657) );
  AOI22_X1 U14405 ( .A1(n14657), .A2(n14377), .B1(n11921), .B2(n14323), .ZN(
        n11923) );
  NAND2_X1 U14406 ( .A1(n14325), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11922) );
  OAI211_X1 U14407 ( .C1(n11924), .C2(n14364), .A(n11923), .B(n11922), .ZN(
        n11925) );
  AOI21_X1 U14408 ( .B1(n14493), .B2(n14357), .A(n11925), .ZN(n11933) );
  OR2_X1 U14409 ( .A1(n14663), .A2(n14029), .ZN(n11928) );
  NAND2_X1 U14410 ( .A1(n11929), .A2(n11928), .ZN(n11931) );
  NAND2_X1 U14411 ( .A1(n11931), .A2(n11930), .ZN(n11986) );
  OAI21_X1 U14412 ( .B1(n11931), .B2(n11930), .A(n11986), .ZN(n14494) );
  NAND2_X1 U14413 ( .A1(n14494), .A2(n14337), .ZN(n11932) );
  OAI211_X1 U14414 ( .C1(n14497), .C2(n14346), .A(n11933), .B(n11932), .ZN(
        P1_U3277) );
  XNOR2_X1 U14415 ( .A(n11934), .B(n12507), .ZN(n11961) );
  NAND2_X1 U14416 ( .A1(n11935), .A2(n12507), .ZN(n11936) );
  NAND3_X1 U14417 ( .A1(n11937), .A2(n14991), .A3(n11936), .ZN(n11939) );
  AOI22_X1 U14418 ( .A1(n14987), .A2(n14577), .B1(n12980), .B2(n14988), .ZN(
        n11938) );
  NAND2_X1 U14419 ( .A1(n11939), .A2(n11938), .ZN(n11956) );
  INV_X1 U14420 ( .A(n11956), .ZN(n11940) );
  MUX2_X1 U14421 ( .A(n11941), .B(n11940), .S(n15051), .Z(n11943) );
  NAND2_X1 U14422 ( .A1(n12602), .A2(n8048), .ZN(n11942) );
  OAI211_X1 U14423 ( .C1(n13043), .C2(n11961), .A(n11943), .B(n11942), .ZN(
        P3_U3473) );
  XNOR2_X1 U14424 ( .A(n11945), .B(n11944), .ZN(n11953) );
  NAND2_X1 U14425 ( .A1(n11946), .A2(n14704), .ZN(n11948) );
  OAI211_X1 U14426 ( .C1(n14707), .C2(n11949), .A(n11948), .B(n11947), .ZN(
        n11950) );
  AOI21_X1 U14427 ( .B1(n11951), .B2(n14653), .A(n11950), .ZN(n11952) );
  OAI21_X1 U14428 ( .B1(n11953), .B2(n14699), .A(n11952), .ZN(P1_U3234) );
  MUX2_X1 U14429 ( .A(n11956), .B(P3_REG0_REG_14__SCAN_IN), .S(n15037), .Z(
        n11955) );
  OAI22_X1 U14430 ( .A1(n11961), .A2(n13125), .B1(n12601), .B2(n13097), .ZN(
        n11954) );
  OR2_X1 U14431 ( .A1(n11955), .A2(n11954), .ZN(P3_U3432) );
  MUX2_X1 U14432 ( .A(n11956), .B(P3_REG2_REG_14__SCAN_IN), .S(n15004), .Z(
        n11957) );
  INV_X1 U14433 ( .A(n11957), .ZN(n11960) );
  AOI22_X1 U14434 ( .A1(n12602), .A2(n12994), .B1(n14998), .B2(n11958), .ZN(
        n11959) );
  OAI211_X1 U14435 ( .C1(n11961), .C2(n12997), .A(n11960), .B(n11959), .ZN(
        P3_U3219) );
  INV_X1 U14436 ( .A(n12232), .ZN(n13789) );
  OAI222_X1 U14437 ( .A1(n14534), .A2(n13789), .B1(n11962), .B2(P1_U3086), 
        .C1(n12032), .C2(n14528), .ZN(P1_U3326) );
  INV_X1 U14438 ( .A(n12250), .ZN(n13793) );
  OAI222_X1 U14439 ( .A1(P1_U3086), .A2(n14055), .B1(n14534), .B2(n13793), 
        .C1(n11963), .C2(n14528), .ZN(P1_U3327) );
  NAND2_X1 U14440 ( .A1(n14654), .A2(n14382), .ZN(n11964) );
  INV_X1 U14441 ( .A(n11966), .ZN(n11968) );
  NAND2_X1 U14442 ( .A1(n14349), .A2(n14348), .ZN(n11970) );
  NAND2_X1 U14443 ( .A1(n14476), .A2(n14484), .ZN(n11969) );
  INV_X1 U14444 ( .A(n14326), .ZN(n14294) );
  NOR2_X1 U14445 ( .A1(n14455), .A2(n14294), .ZN(n11971) );
  NAND2_X1 U14446 ( .A1(n14285), .A2(n11994), .ZN(n11973) );
  NAND2_X1 U14447 ( .A1(n14449), .A2(n14278), .ZN(n11972) );
  NAND2_X1 U14448 ( .A1(n11973), .A2(n11972), .ZN(n14265) );
  NAND2_X1 U14449 ( .A1(n14280), .A2(n13996), .ZN(n11975) );
  INV_X1 U14450 ( .A(n14255), .ZN(n14006) );
  NOR2_X1 U14451 ( .A1(n14418), .A2(n14025), .ZN(n12040) );
  INV_X1 U14452 ( .A(n12002), .ZN(n11978) );
  NAND2_X1 U14453 ( .A1(n11979), .A2(n11978), .ZN(n12012) );
  NAND2_X1 U14454 ( .A1(n14022), .A2(n14739), .ZN(n11982) );
  NAND2_X1 U14455 ( .A1(n14024), .A2(n14483), .ZN(n11981) );
  AOI21_X2 U14456 ( .B1(n11984), .B2(n14489), .A(n11983), .ZN(n14409) );
  INV_X1 U14457 ( .A(n14412), .ZN(n13895) );
  OR2_X1 U14458 ( .A1(n14654), .A2(n14482), .ZN(n11985) );
  OR2_X1 U14459 ( .A1(n14322), .A2(n13939), .ZN(n11991) );
  OR2_X1 U14460 ( .A1(n14455), .A2(n14326), .ZN(n11992) );
  NAND2_X1 U14461 ( .A1(n11993), .A2(n11992), .ZN(n14288) );
  INV_X1 U14462 ( .A(n11994), .ZN(n14287) );
  OR2_X1 U14463 ( .A1(n14449), .A2(n14026), .ZN(n11995) );
  NAND2_X1 U14464 ( .A1(n14280), .A2(n14297), .ZN(n11996) );
  NAND2_X1 U14465 ( .A1(n14267), .A2(n11996), .ZN(n14243) );
  INV_X1 U14466 ( .A(n14243), .ZN(n11998) );
  INV_X1 U14467 ( .A(n14025), .ZN(n13952) );
  OAI21_X1 U14468 ( .B1(n12003), .B2(n12002), .A(n12015), .ZN(n14410) );
  OAI22_X1 U14469 ( .A1(n14377), .A2(n12004), .B1(n13930), .B2(n14374), .ZN(
        n12005) );
  AOI21_X1 U14470 ( .B1(n14407), .B2(n14384), .A(n12005), .ZN(n12008) );
  INV_X1 U14471 ( .A(n14280), .ZN(n14272) );
  INV_X1 U14472 ( .A(n14385), .ZN(n14487) );
  AND2_X1 U14473 ( .A1(n14372), .A2(n14487), .ZN(n14352) );
  NAND2_X1 U14474 ( .A1(n14272), .A2(n14291), .ZN(n14271) );
  NAND2_X1 U14475 ( .A1(n13925), .A2(n12045), .ZN(n12018) );
  OR2_X1 U14476 ( .A1(n13925), .A2(n12045), .ZN(n12006) );
  NAND2_X1 U14477 ( .A1(n14406), .A2(n14357), .ZN(n12007) );
  OAI211_X1 U14478 ( .C1(n14410), .C2(n14391), .A(n12008), .B(n12007), .ZN(
        n12009) );
  INV_X1 U14479 ( .A(n12009), .ZN(n12010) );
  OAI21_X1 U14480 ( .B1(n14409), .B2(n14325), .A(n12010), .ZN(P1_U3265) );
  NAND2_X1 U14481 ( .A1(n14398), .A2(n14337), .ZN(n12028) );
  AOI211_X1 U14482 ( .C1(n14404), .C2(n12018), .A(n14355), .B(n14208), .ZN(
        n14402) );
  NAND2_X1 U14483 ( .A1(n14404), .A2(n14384), .ZN(n12025) );
  INV_X1 U14484 ( .A(P1_B_REG_SCAN_IN), .ZN(n12019) );
  OR2_X1 U14485 ( .A1(n14524), .A2(n12019), .ZN(n12020) );
  AND2_X1 U14486 ( .A1(n14739), .A2(n12020), .ZN(n14203) );
  NAND2_X1 U14487 ( .A1(n14203), .A2(n14021), .ZN(n14399) );
  OAI22_X1 U14488 ( .A1(n12022), .A2(n14399), .B1(n12021), .B2(n14374), .ZN(
        n12023) );
  AOI21_X1 U14489 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14325), .A(n12023), 
        .ZN(n12024) );
  OAI211_X1 U14490 ( .C1(n14401), .C2(n14381), .A(n12025), .B(n12024), .ZN(
        n12026) );
  AOI21_X1 U14491 ( .B1(n14402), .B2(n14357), .A(n12026), .ZN(n12027) );
  OAI211_X1 U14492 ( .C1(n14405), .C2(n14346), .A(n12028), .B(n12027), .ZN(
        P1_U3356) );
  INV_X1 U14493 ( .A(n12029), .ZN(n12030) );
  NAND2_X1 U14494 ( .A1(n12032), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12033) );
  INV_X1 U14495 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12054) );
  NAND2_X1 U14496 ( .A1(n12054), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12481) );
  NAND2_X1 U14497 ( .A1(n12055), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12035) );
  NAND2_X1 U14498 ( .A1(n12481), .A2(n12035), .ZN(n12482) );
  XNOR2_X1 U14499 ( .A(n12483), .B(n12482), .ZN(n12478) );
  INV_X1 U14500 ( .A(n12478), .ZN(n12036) );
  OAI222_X1 U14501 ( .A1(n12037), .A2(P3_U3151), .B1(n13140), .B2(n12036), 
        .C1(n15053), .C2(n13142), .ZN(P3_U3265) );
  INV_X1 U14502 ( .A(n14415), .ZN(n12050) );
  OR3_X1 U14503 ( .A1(n14215), .A2(n12041), .A3(n12040), .ZN(n12042) );
  OAI22_X1 U14504 ( .A1(n13952), .A2(n14400), .B1(n14401), .B2(n14474), .ZN(
        n12044) );
  AOI211_X1 U14505 ( .C1(n14412), .C2(n14219), .A(n14355), .B(n12045), .ZN(
        n14411) );
  NOR2_X1 U14506 ( .A1(n13895), .A2(n14364), .ZN(n12048) );
  OAI22_X1 U14507 ( .A1(n14377), .A2(n12046), .B1(n13890), .B2(n14374), .ZN(
        n12047) );
  AOI211_X1 U14508 ( .C1(n14411), .C2(n14357), .A(n12048), .B(n12047), .ZN(
        n12052) );
  NAND2_X1 U14509 ( .A1(n12050), .A2(n12049), .ZN(n12051) );
  OAI211_X1 U14510 ( .C1(n14414), .C2(n14325), .A(n12052), .B(n12051), .ZN(
        P1_U3266) );
  INV_X1 U14511 ( .A(n12217), .ZN(n12057) );
  OAI222_X1 U14512 ( .A1(n13800), .A2(n12057), .B1(P2_U3088), .B2(n6687), .C1(
        n12054), .C2(n13803), .ZN(P2_U3297) );
  OAI222_X1 U14513 ( .A1(n14534), .A2(n12057), .B1(n12056), .B2(P1_U3086), 
        .C1(n12055), .C2(n14528), .ZN(P1_U3325) );
  OAI22_X1 U14514 ( .A1(n14631), .A2(n12276), .B1(n12150), .B2(n12277), .ZN(
        n12156) );
  NAND2_X1 U14515 ( .A1(n12064), .A2(n12072), .ZN(n12061) );
  NAND2_X1 U14516 ( .A1(n12103), .A2(n12059), .ZN(n12060) );
  NAND2_X1 U14517 ( .A1(n12064), .A2(n12063), .ZN(n12069) );
  INV_X1 U14518 ( .A(n12286), .ZN(n12067) );
  INV_X1 U14519 ( .A(n12065), .ZN(n12066) );
  NAND2_X1 U14520 ( .A1(n12069), .A2(n12068), .ZN(n12070) );
  AND2_X1 U14521 ( .A1(n12071), .A2(n12070), .ZN(n12080) );
  NAND2_X1 U14522 ( .A1(n13295), .A2(n12228), .ZN(n12075) );
  NAND2_X1 U14523 ( .A1(n12073), .A2(n6459), .ZN(n12074) );
  NAND2_X1 U14524 ( .A1(n12075), .A2(n12074), .ZN(n12084) );
  AOI22_X1 U14525 ( .A1(n6734), .A2(n12228), .B1(n6459), .B2(n12076), .ZN(
        n12077) );
  INV_X1 U14526 ( .A(n12077), .ZN(n12078) );
  OAI21_X1 U14527 ( .B1(n12080), .B2(n12079), .A(n12078), .ZN(n12081) );
  NAND2_X1 U14528 ( .A1(n12082), .A2(n12081), .ZN(n12086) );
  NAND2_X1 U14529 ( .A1(n12086), .A2(n12085), .ZN(n12089) );
  NAND2_X1 U14530 ( .A1(n12089), .A2(n12090), .ZN(n12094) );
  OAI22_X1 U14531 ( .A1(n12088), .A2(n12276), .B1(n12087), .B2(n12228), .ZN(
        n12093) );
  INV_X1 U14532 ( .A(n12089), .ZN(n12092) );
  INV_X1 U14533 ( .A(n12090), .ZN(n12091) );
  AOI22_X1 U14534 ( .A1(n12095), .A2(n12254), .B1(n13293), .B2(n12228), .ZN(
        n12100) );
  OAI22_X1 U14535 ( .A1(n12097), .A2(n12276), .B1(n12096), .B2(n12277), .ZN(
        n12098) );
  AOI22_X1 U14536 ( .A1(n12102), .A2(n12228), .B1(n6459), .B2(n13292), .ZN(
        n12107) );
  OAI22_X1 U14537 ( .A1(n12109), .A2(n12277), .B1(n12108), .B2(n12276), .ZN(
        n12110) );
  NAND2_X1 U14538 ( .A1(n12111), .A2(n12110), .ZN(n12114) );
  OAI22_X1 U14539 ( .A1(n12109), .A2(n12276), .B1(n12108), .B2(n12277), .ZN(
        n12113) );
  AOI22_X1 U14540 ( .A1(n12115), .A2(n12277), .B1(n12103), .B2(n13290), .ZN(
        n12119) );
  OAI22_X1 U14541 ( .A1(n12117), .A2(n12277), .B1(n12116), .B2(n12276), .ZN(
        n12118) );
  OAI21_X1 U14542 ( .B1(n12120), .B2(n12119), .A(n12118), .ZN(n12122) );
  NAND2_X1 U14543 ( .A1(n12120), .A2(n12119), .ZN(n12121) );
  NAND2_X1 U14544 ( .A1(n12122), .A2(n12121), .ZN(n12124) );
  NAND2_X1 U14545 ( .A1(n12124), .A2(n12125), .ZN(n12129) );
  OAI22_X1 U14546 ( .A1(n14897), .A2(n12276), .B1(n12123), .B2(n12277), .ZN(
        n12128) );
  INV_X1 U14547 ( .A(n12124), .ZN(n12127) );
  INV_X1 U14548 ( .A(n12125), .ZN(n12126) );
  AOI22_X1 U14549 ( .A1(n12130), .A2(n12277), .B1(n6459), .B2(n13288), .ZN(
        n12134) );
  OAI22_X1 U14550 ( .A1(n12132), .A2(n12277), .B1(n12131), .B2(n12276), .ZN(
        n12133) );
  AOI22_X1 U14551 ( .A1(n13655), .A2(n12276), .B1(n13287), .B2(n12277), .ZN(
        n12140) );
  INV_X1 U14552 ( .A(n12140), .ZN(n12139) );
  OAI22_X1 U14553 ( .A1(n14908), .A2(n12276), .B1(n12141), .B2(n12277), .ZN(
        n12145) );
  NAND2_X1 U14554 ( .A1(n12144), .A2(n12145), .ZN(n12143) );
  OAI22_X1 U14555 ( .A1(n14908), .A2(n12277), .B1(n12141), .B2(n12276), .ZN(
        n12142) );
  NAND2_X1 U14556 ( .A1(n12143), .A2(n12142), .ZN(n12149) );
  INV_X1 U14557 ( .A(n12144), .ZN(n12147) );
  INV_X1 U14558 ( .A(n12145), .ZN(n12146) );
  NAND2_X1 U14559 ( .A1(n12147), .A2(n12146), .ZN(n12148) );
  OAI22_X1 U14560 ( .A1(n14631), .A2(n12277), .B1(n12150), .B2(n12276), .ZN(
        n12153) );
  INV_X1 U14561 ( .A(n12153), .ZN(n12151) );
  NAND2_X1 U14562 ( .A1(n12152), .A2(n12153), .ZN(n12155) );
  INV_X1 U14563 ( .A(n12152), .ZN(n12154) );
  AOI22_X1 U14564 ( .A1(n12157), .A2(n12277), .B1(n12276), .B2(n13284), .ZN(
        n12161) );
  OAI22_X1 U14565 ( .A1(n12159), .A2(n12277), .B1(n12158), .B2(n12276), .ZN(
        n12160) );
  OAI21_X1 U14566 ( .B1(n12162), .B2(n12161), .A(n12160), .ZN(n12164) );
  AOI22_X1 U14567 ( .A1(n14620), .A2(n12254), .B1(n13388), .B2(n12277), .ZN(
        n12167) );
  INV_X1 U14568 ( .A(n12167), .ZN(n12166) );
  OAI22_X1 U14569 ( .A1(n13781), .A2(n12276), .B1(n13389), .B2(n12277), .ZN(
        n12169) );
  NOR2_X1 U14570 ( .A1(n12170), .A2(n12169), .ZN(n12172) );
  AOI22_X1 U14571 ( .A1(n13644), .A2(n12254), .B1(n13350), .B2(n12277), .ZN(
        n12168) );
  OAI22_X1 U14572 ( .A1(n13390), .A2(n12277), .B1(n13633), .B2(n12276), .ZN(
        n12174) );
  NOR2_X1 U14573 ( .A1(n12175), .A2(n12174), .ZN(n12177) );
  INV_X1 U14574 ( .A(n13633), .ZN(n13353) );
  AOI22_X1 U14575 ( .A1(n13775), .A2(n12277), .B1(n12254), .B2(n13353), .ZN(
        n12173) );
  OAI22_X1 U14576 ( .A1(n13604), .A2(n12276), .B1(n13393), .B2(n12277), .ZN(
        n12179) );
  INV_X1 U14577 ( .A(n13393), .ZN(n13355) );
  AOI22_X1 U14578 ( .A1(n13730), .A2(n12254), .B1(n13355), .B2(n12277), .ZN(
        n12178) );
  OAI22_X1 U14579 ( .A1(n13593), .A2(n12277), .B1(n13396), .B2(n12276), .ZN(
        n12180) );
  OAI22_X1 U14580 ( .A1(n13593), .A2(n12276), .B1(n13396), .B2(n12277), .ZN(
        n12182) );
  INV_X1 U14581 ( .A(n12180), .ZN(n12181) );
  INV_X1 U14582 ( .A(n12186), .ZN(n12183) );
  NAND2_X1 U14583 ( .A1(n12183), .A2(n12184), .ZN(n12188) );
  OAI22_X1 U14584 ( .A1(n13578), .A2(n12277), .B1(n13247), .B2(n12276), .ZN(
        n12187) );
  INV_X1 U14585 ( .A(n12184), .ZN(n12185) );
  AOI22_X1 U14586 ( .A1(n13715), .A2(n12254), .B1(n13543), .B2(n12277), .ZN(
        n12190) );
  INV_X1 U14587 ( .A(n13715), .ZN(n13564) );
  INV_X1 U14588 ( .A(n13543), .ZN(n13364) );
  OAI22_X1 U14589 ( .A1(n13564), .A2(n12276), .B1(n13364), .B2(n12277), .ZN(
        n12189) );
  OAI22_X1 U14590 ( .A1(n13552), .A2(n12276), .B1(n13403), .B2(n12277), .ZN(
        n12193) );
  INV_X1 U14591 ( .A(n12193), .ZN(n12192) );
  OAI22_X1 U14592 ( .A1(n13552), .A2(n12277), .B1(n13403), .B2(n12276), .ZN(
        n12191) );
  NAND2_X1 U14593 ( .A1(n12194), .A2(n12192), .ZN(n12195) );
  NAND2_X1 U14594 ( .A1(n12196), .A2(n12195), .ZN(n12199) );
  OAI22_X1 U14595 ( .A1(n13526), .A2(n12277), .B1(n13233), .B2(n12276), .ZN(
        n12198) );
  OAI22_X1 U14596 ( .A1(n13512), .A2(n12276), .B1(n13406), .B2(n12277), .ZN(
        n12200) );
  OAI22_X1 U14597 ( .A1(n13512), .A2(n12277), .B1(n13406), .B2(n12276), .ZN(
        n12201) );
  AOI22_X1 U14598 ( .A1(n13692), .A2(n12254), .B1(n13408), .B2(n12277), .ZN(
        n12203) );
  INV_X1 U14599 ( .A(n13692), .ZN(n13500) );
  INV_X1 U14600 ( .A(n13408), .ZN(n13474) );
  OAI22_X1 U14601 ( .A1(n13500), .A2(n12276), .B1(n13474), .B2(n12277), .ZN(
        n12202) );
  OAI21_X1 U14602 ( .B1(n12204), .B2(n12203), .A(n12202), .ZN(n12206) );
  NAND2_X1 U14603 ( .A1(n12204), .A2(n12203), .ZN(n12205) );
  AOI22_X1 U14604 ( .A1(n13763), .A2(n12277), .B1(n12254), .B2(n13455), .ZN(
        n12208) );
  AOI22_X1 U14605 ( .A1(n13763), .A2(n12254), .B1(n13455), .B2(n12277), .ZN(
        n12207) );
  INV_X1 U14606 ( .A(n12208), .ZN(n12209) );
  AND2_X1 U14607 ( .A1(n13456), .A2(n12277), .ZN(n12210) );
  AOI21_X1 U14608 ( .B1(n13446), .B2(n12254), .A(n12210), .ZN(n12261) );
  NAND2_X1 U14609 ( .A1(n13446), .A2(n12277), .ZN(n12212) );
  NAND2_X1 U14610 ( .A1(n13456), .A2(n12254), .ZN(n12211) );
  NAND2_X1 U14611 ( .A1(n12212), .A2(n12211), .ZN(n12259) );
  AND2_X1 U14612 ( .A1(n13472), .A2(n12277), .ZN(n12213) );
  AOI21_X1 U14613 ( .B1(n13681), .B2(n12254), .A(n12213), .ZN(n12256) );
  NAND2_X1 U14614 ( .A1(n13681), .A2(n12228), .ZN(n12215) );
  NAND2_X1 U14615 ( .A1(n13472), .A2(n12254), .ZN(n12214) );
  NAND2_X1 U14616 ( .A1(n12215), .A2(n12214), .ZN(n12255) );
  AOI22_X1 U14617 ( .A1(n12261), .A2(n12259), .B1(n12256), .B2(n12255), .ZN(
        n12216) );
  INV_X1 U14618 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13668) );
  OR2_X1 U14619 ( .A1(n12218), .A2(n13668), .ZN(n12223) );
  INV_X1 U14620 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n12219) );
  OR2_X1 U14621 ( .A1(n12239), .A2(n12219), .ZN(n12222) );
  INV_X1 U14622 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13753) );
  OR2_X1 U14623 ( .A1(n12220), .A2(n13753), .ZN(n12221) );
  AND3_X1 U14624 ( .A1(n12223), .A2(n12222), .A3(n12221), .ZN(n12224) );
  OAI22_X1 U14625 ( .A1(n13755), .A2(n12276), .B1(n12224), .B2(n12277), .ZN(
        n12274) );
  INV_X1 U14626 ( .A(n13755), .ZN(n12289) );
  INV_X1 U14627 ( .A(n12224), .ZN(n13377) );
  INV_X1 U14628 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n12227) );
  NAND2_X1 U14629 ( .A1(n6647), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U14630 ( .A1(n12236), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12225) );
  OAI211_X1 U14631 ( .C1(n12239), .C2(n12227), .A(n12226), .B(n12225), .ZN(
        n13340) );
  NAND2_X1 U14632 ( .A1(n13340), .A2(n12228), .ZN(n12278) );
  OR2_X1 U14633 ( .A1(n12229), .A2(n12295), .ZN(n12230) );
  NAND4_X1 U14634 ( .A1(n12278), .A2(n12283), .A3(n12285), .A4(n12230), .ZN(
        n12231) );
  AOI22_X1 U14635 ( .A1(n12289), .A2(n12254), .B1(n13377), .B2(n12231), .ZN(
        n12273) );
  NAND2_X1 U14636 ( .A1(n12232), .A2(n12249), .ZN(n12234) );
  NAND2_X1 U14637 ( .A1(n12251), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12233) );
  NAND2_X1 U14638 ( .A1(n13383), .A2(n9026), .ZN(n12243) );
  INV_X1 U14639 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U14640 ( .A1(n6647), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n12238) );
  NAND2_X1 U14641 ( .A1(n12236), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n12237) );
  OAI211_X1 U14642 ( .C1(n12240), .C2(n12239), .A(n12238), .B(n12237), .ZN(
        n12241) );
  INV_X1 U14643 ( .A(n12241), .ZN(n12242) );
  NAND2_X1 U14644 ( .A1(n12243), .A2(n12242), .ZN(n13420) );
  AND2_X1 U14645 ( .A1(n13420), .A2(n12228), .ZN(n12244) );
  AOI21_X1 U14646 ( .B1(n13335), .B2(n12254), .A(n12244), .ZN(n12266) );
  NAND2_X1 U14647 ( .A1(n13335), .A2(n12277), .ZN(n12246) );
  NAND2_X1 U14648 ( .A1(n13420), .A2(n12254), .ZN(n12245) );
  NAND2_X1 U14649 ( .A1(n12246), .A2(n12245), .ZN(n12265) );
  NAND2_X1 U14650 ( .A1(n13782), .A2(n12249), .ZN(n12248) );
  NAND2_X1 U14651 ( .A1(n12251), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12247) );
  XNOR2_X1 U14652 ( .A(n13336), .B(n13340), .ZN(n12324) );
  NAND2_X1 U14653 ( .A1(n12250), .A2(n12249), .ZN(n12253) );
  NAND2_X1 U14654 ( .A1(n12251), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U14655 ( .A1(n13674), .A2(n12228), .B1(n12254), .B2(n13379), .ZN(
        n12268) );
  OAI22_X1 U14656 ( .A1(n13428), .A2(n12277), .B1(n13436), .B2(n12276), .ZN(
        n12267) );
  INV_X1 U14657 ( .A(n12255), .ZN(n12258) );
  INV_X1 U14658 ( .A(n12256), .ZN(n12257) );
  NAND2_X1 U14659 ( .A1(n12258), .A2(n12257), .ZN(n12260) );
  NOR2_X1 U14660 ( .A1(n12261), .A2(n12260), .ZN(n12263) );
  AOI21_X1 U14661 ( .B1(n12261), .B2(n12260), .A(n12259), .ZN(n12262) );
  AOI211_X1 U14662 ( .C1(n12268), .C2(n12267), .A(n12263), .B(n12262), .ZN(
        n12264) );
  INV_X1 U14663 ( .A(n12265), .ZN(n12270) );
  INV_X1 U14664 ( .A(n12266), .ZN(n12269) );
  OAI22_X1 U14665 ( .A1(n12270), .A2(n12269), .B1(n12268), .B2(n12267), .ZN(
        n12271) );
  NAND2_X1 U14666 ( .A1(n13340), .A2(n12276), .ZN(n12280) );
  NAND2_X1 U14667 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  MUX2_X1 U14668 ( .A(n12280), .B(n12279), .S(n13336), .Z(n12281) );
  INV_X1 U14669 ( .A(n12337), .ZN(n12288) );
  NAND2_X1 U14670 ( .A1(n12283), .A2(n12334), .ZN(n12284) );
  OAI211_X1 U14671 ( .C1(n12286), .C2(n12343), .A(n12285), .B(n12284), .ZN(
        n12287) );
  XNOR2_X1 U14672 ( .A(n12289), .B(n13377), .ZN(n12325) );
  NAND2_X1 U14673 ( .A1(n13674), .A2(n13436), .ZN(n12290) );
  NAND2_X1 U14674 ( .A1(n13411), .A2(n13472), .ZN(n12291) );
  NAND2_X1 U14675 ( .A1(n13681), .A2(n13435), .ZN(n13372) );
  NAND2_X1 U14676 ( .A1(n12291), .A2(n13372), .ZN(n13347) );
  INV_X1 U14677 ( .A(n13455), .ZN(n12292) );
  NAND2_X1 U14678 ( .A1(n13763), .A2(n12292), .ZN(n13371) );
  OR2_X1 U14679 ( .A1(n13763), .A2(n12292), .ZN(n12293) );
  NAND2_X1 U14680 ( .A1(n13371), .A2(n12293), .ZN(n13478) );
  XNOR2_X1 U14681 ( .A(n13692), .B(n13408), .ZN(n13493) );
  NAND2_X1 U14682 ( .A1(n13698), .A2(n13406), .ZN(n13369) );
  OR2_X1 U14683 ( .A1(n13698), .A2(n13406), .ZN(n12294) );
  XNOR2_X1 U14684 ( .A(n13702), .B(n13233), .ZN(n13535) );
  XNOR2_X1 U14685 ( .A(n13710), .B(n13524), .ZN(n13553) );
  XNOR2_X1 U14686 ( .A(n13725), .B(n13359), .ZN(n13585) );
  NAND4_X1 U14687 ( .A1(n12296), .A2(n12297), .A3(n12295), .A4(n14882), .ZN(
        n12299) );
  NOR2_X1 U14688 ( .A1(n12299), .A2(n12298), .ZN(n12302) );
  NAND4_X1 U14689 ( .A1(n12303), .A2(n12302), .A3(n12301), .A4(n12300), .ZN(
        n12304) );
  NOR2_X1 U14690 ( .A1(n12305), .A2(n12304), .ZN(n12308) );
  NAND4_X1 U14691 ( .A1(n12309), .A2(n12308), .A3(n12307), .A4(n12306), .ZN(
        n12310) );
  NOR2_X1 U14692 ( .A1(n12311), .A2(n12310), .ZN(n12314) );
  NAND4_X1 U14693 ( .A1(n12315), .A2(n12314), .A3(n12313), .A4(n12312), .ZN(
        n12316) );
  XNOR2_X1 U14694 ( .A(n13775), .B(n13633), .ZN(n13612) );
  NOR2_X1 U14695 ( .A1(n12316), .A2(n13612), .ZN(n12317) );
  XNOR2_X1 U14696 ( .A(n13730), .B(n13355), .ZN(n13606) );
  AND4_X1 U14697 ( .A1(n13585), .A2(n12317), .A3(n13606), .A4(n13645), .ZN(
        n12318) );
  XNOR2_X1 U14698 ( .A(n13715), .B(n13543), .ZN(n13565) );
  INV_X1 U14699 ( .A(n13247), .ZN(n13362) );
  NAND2_X1 U14700 ( .A1(n13720), .A2(n13362), .ZN(n13397) );
  NAND2_X1 U14701 ( .A1(n13398), .A2(n13397), .ZN(n13579) );
  NAND4_X1 U14702 ( .A1(n13553), .A2(n12318), .A3(n13565), .A4(n13579), .ZN(
        n12319) );
  NOR2_X1 U14703 ( .A1(n13535), .A2(n12319), .ZN(n12320) );
  NAND3_X1 U14704 ( .A1(n13493), .A2(n13516), .A3(n12320), .ZN(n12321) );
  NOR3_X1 U14705 ( .A1(n13347), .A2(n13478), .A3(n12321), .ZN(n12322) );
  XNOR2_X1 U14706 ( .A(n13446), .B(n13456), .ZN(n13447) );
  AND3_X1 U14707 ( .A1(n13417), .A2(n12322), .A3(n13447), .ZN(n12323) );
  XNOR2_X1 U14708 ( .A(n13335), .B(n13420), .ZN(n13414) );
  NAND4_X1 U14709 ( .A1(n12325), .A2(n12324), .A3(n12323), .A4(n13414), .ZN(
        n12327) );
  OAI21_X1 U14710 ( .B1(n12334), .B2(n12331), .A(n12327), .ZN(n12328) );
  NAND2_X1 U14711 ( .A1(n12333), .A2(n12328), .ZN(n12338) );
  AOI21_X1 U14712 ( .B1(n12331), .B2(n6756), .A(n12329), .ZN(n12332) );
  NOR2_X1 U14713 ( .A1(n12335), .A2(n12334), .ZN(n12336) );
  NAND4_X1 U14714 ( .A1(n14881), .A2(n12341), .A3(n12340), .A4(n13542), .ZN(
        n12342) );
  OAI211_X1 U14715 ( .C1(n12343), .C2(n7433), .A(n12342), .B(P2_B_REG_SCAN_IN), 
        .ZN(n12344) );
  XNOR2_X1 U14716 ( .A(n12346), .B(n12345), .ZN(n12347) );
  NAND2_X1 U14717 ( .A1(n12347), .A2(n12449), .ZN(n12352) );
  AOI22_X1 U14718 ( .A1(n6439), .A2(n12871), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12348) );
  OAI21_X1 U14719 ( .B1(n12349), .B2(n12455), .A(n12348), .ZN(n12350) );
  AOI21_X1 U14720 ( .B1(n12845), .B2(n12464), .A(n12350), .ZN(n12351) );
  OAI211_X1 U14721 ( .C1(n12848), .C2(n12459), .A(n12352), .B(n12351), .ZN(
        P3_U3154) );
  XNOR2_X1 U14722 ( .A(n12423), .B(n12422), .ZN(n12424) );
  XNOR2_X1 U14723 ( .A(n12424), .B(n12903), .ZN(n12357) );
  AOI22_X1 U14724 ( .A1(n12463), .A2(n12892), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12354) );
  NAND2_X1 U14725 ( .A1(n12464), .A2(n12896), .ZN(n12353) );
  OAI211_X1 U14726 ( .C1(n12467), .C2(n12914), .A(n12354), .B(n12353), .ZN(
        n12355) );
  AOI21_X1 U14727 ( .B1(n13077), .B2(n12469), .A(n12355), .ZN(n12356) );
  OAI21_X1 U14728 ( .B1(n12357), .B2(n12471), .A(n12356), .ZN(P3_U3156) );
  OAI211_X1 U14729 ( .C1(n12360), .C2(n12359), .A(n12358), .B(n12449), .ZN(
        n12369) );
  NAND2_X1 U14730 ( .A1(n6439), .A2(n12699), .ZN(n12361) );
  NAND2_X1 U14731 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n14945)
         );
  OAI211_X1 U14732 ( .C1(n12362), .C2(n12455), .A(n12361), .B(n14945), .ZN(
        n12363) );
  INV_X1 U14733 ( .A(n12363), .ZN(n12368) );
  NAND2_X1 U14734 ( .A1(n12464), .A2(n12364), .ZN(n12367) );
  OR2_X1 U14735 ( .A1(n12459), .A2(n12365), .ZN(n12366) );
  NAND4_X1 U14736 ( .A1(n12369), .A2(n12368), .A3(n12367), .A4(n12366), .ZN(
        P3_U3157) );
  OAI211_X1 U14737 ( .C1(n12372), .C2(n12371), .A(n12370), .B(n12449), .ZN(
        n12376) );
  NAND2_X1 U14738 ( .A1(n6439), .A2(n12969), .ZN(n12373) );
  NAND2_X1 U14739 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12807)
         );
  OAI211_X1 U14740 ( .C1(n12940), .C2(n12455), .A(n12373), .B(n12807), .ZN(
        n12374) );
  AOI21_X1 U14741 ( .B1(n12946), .B2(n12464), .A(n12374), .ZN(n12375) );
  OAI211_X1 U14742 ( .C1(n12459), .C2(n13098), .A(n12376), .B(n12375), .ZN(
        P3_U3159) );
  OAI211_X1 U14743 ( .C1(n12379), .C2(n12378), .A(n12377), .B(n12449), .ZN(
        n12386) );
  AOI21_X1 U14744 ( .B1(n12469), .B2(n12381), .A(n12380), .ZN(n12385) );
  AOI22_X1 U14745 ( .A1(n6439), .A2(n12701), .B1(n12463), .B2(n12699), .ZN(
        n12384) );
  NAND2_X1 U14746 ( .A1(n12464), .A2(n12382), .ZN(n12383) );
  NAND4_X1 U14747 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        P3_U3161) );
  OAI211_X1 U14748 ( .C1(n12389), .C2(n12388), .A(n12387), .B(n12449), .ZN(
        n12394) );
  AOI22_X1 U14749 ( .A1(n6439), .A2(n12698), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12391) );
  NAND2_X1 U14750 ( .A1(n12464), .A2(n12917), .ZN(n12390) );
  OAI211_X1 U14751 ( .C1(n12914), .C2(n12455), .A(n12391), .B(n12390), .ZN(
        n12392) );
  AOI21_X1 U14752 ( .B1(n13021), .B2(n12469), .A(n12392), .ZN(n12393) );
  NAND2_X1 U14753 ( .A1(n12394), .A2(n12393), .ZN(P3_U3163) );
  XOR2_X1 U14754 ( .A(n12396), .B(n12395), .Z(n12402) );
  AOI22_X1 U14755 ( .A1(n12463), .A2(n12871), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12398) );
  NAND2_X1 U14756 ( .A1(n12464), .A2(n12875), .ZN(n12397) );
  OAI211_X1 U14757 ( .C1(n12467), .C2(n12399), .A(n12398), .B(n12397), .ZN(
        n12400) );
  AOI21_X1 U14758 ( .B1(n13008), .B2(n12469), .A(n12400), .ZN(n12401) );
  OAI21_X1 U14759 ( .B1(n12402), .B2(n12471), .A(n12401), .ZN(P3_U3165) );
  NAND2_X1 U14760 ( .A1(n12404), .A2(n12403), .ZN(n12406) );
  XOR2_X1 U14761 ( .A(n12406), .B(n12405), .Z(n12412) );
  AND2_X1 U14762 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12731) );
  AOI21_X1 U14763 ( .B1(n12463), .B2(n12981), .A(n12731), .ZN(n12408) );
  NAND2_X1 U14764 ( .A1(n12464), .A2(n12984), .ZN(n12407) );
  OAI211_X1 U14765 ( .C1(n12467), .C2(n12409), .A(n12408), .B(n12407), .ZN(
        n12410) );
  AOI21_X1 U14766 ( .B1(n13115), .B2(n12469), .A(n12410), .ZN(n12411) );
  OAI21_X1 U14767 ( .B1(n12412), .B2(n12471), .A(n12411), .ZN(P3_U3166) );
  INV_X1 U14768 ( .A(n13109), .ZN(n12421) );
  OAI211_X1 U14769 ( .C1(n12415), .C2(n12414), .A(n12413), .B(n12449), .ZN(
        n12420) );
  NOR2_X1 U14770 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12416), .ZN(n12757) );
  AOI21_X1 U14771 ( .B1(n12463), .B2(n12969), .A(n12757), .ZN(n12417) );
  OAI21_X1 U14772 ( .B1(n12467), .B2(n7077), .A(n12417), .ZN(n12418) );
  AOI21_X1 U14773 ( .B1(n12972), .B2(n12464), .A(n12418), .ZN(n12419) );
  OAI211_X1 U14774 ( .C1(n12421), .C2(n12459), .A(n12420), .B(n12419), .ZN(
        P3_U3168) );
  OAI22_X1 U14775 ( .A1(n12424), .A2(n12697), .B1(n12423), .B2(n12422), .ZN(
        n12427) );
  XNOR2_X1 U14776 ( .A(n12425), .B(n12892), .ZN(n12426) );
  XNOR2_X1 U14777 ( .A(n12427), .B(n12426), .ZN(n12432) );
  AOI22_X1 U14778 ( .A1(n12463), .A2(n12881), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12429) );
  NAND2_X1 U14779 ( .A1(n12464), .A2(n12886), .ZN(n12428) );
  OAI211_X1 U14780 ( .C1(n12467), .C2(n12903), .A(n12429), .B(n12428), .ZN(
        n12430) );
  AOI21_X1 U14781 ( .B1(n13071), .B2(n12469), .A(n12430), .ZN(n12431) );
  OAI21_X1 U14782 ( .B1(n12432), .B2(n12471), .A(n12431), .ZN(P3_U3169) );
  INV_X1 U14783 ( .A(n12932), .ZN(n13091) );
  OAI211_X1 U14784 ( .C1(n12435), .C2(n12434), .A(n12433), .B(n12449), .ZN(
        n12442) );
  OAI22_X1 U14785 ( .A1(n12455), .A2(n12902), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12436), .ZN(n12440) );
  INV_X1 U14786 ( .A(n12931), .ZN(n12437) );
  NOR2_X1 U14787 ( .A1(n12438), .A2(n12437), .ZN(n12439) );
  AOI211_X1 U14788 ( .C1(n6439), .C2(n12926), .A(n12440), .B(n12439), .ZN(
        n12441) );
  OAI211_X1 U14789 ( .C1(n13091), .C2(n12459), .A(n12442), .B(n12441), .ZN(
        P3_U3173) );
  XNOR2_X1 U14790 ( .A(n12443), .B(n12893), .ZN(n12448) );
  AOI22_X1 U14791 ( .A1(n6439), .A2(n12927), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12445) );
  NAND2_X1 U14792 ( .A1(n12464), .A2(n12907), .ZN(n12444) );
  OAI211_X1 U14793 ( .C1(n12903), .C2(n12455), .A(n12445), .B(n12444), .ZN(
        n12446) );
  AOI21_X1 U14794 ( .B1(n13082), .B2(n12469), .A(n12446), .ZN(n12447) );
  OAI21_X1 U14795 ( .B1(n12448), .B2(n12471), .A(n12447), .ZN(P3_U3175) );
  INV_X1 U14796 ( .A(n13032), .ZN(n12460) );
  OAI211_X1 U14797 ( .C1(n12452), .C2(n12451), .A(n12450), .B(n12449), .ZN(
        n12458) );
  NAND2_X1 U14798 ( .A1(n6439), .A2(n12981), .ZN(n12454) );
  NAND2_X1 U14799 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12774)
         );
  OAI211_X1 U14800 ( .C1(n12957), .C2(n12455), .A(n12454), .B(n12774), .ZN(
        n12456) );
  AOI21_X1 U14801 ( .B1(n12959), .B2(n12464), .A(n12456), .ZN(n12457) );
  OAI211_X1 U14802 ( .C1(n12460), .C2(n12459), .A(n12458), .B(n12457), .ZN(
        P3_U3178) );
  XOR2_X1 U14803 ( .A(n12462), .B(n12461), .Z(n12472) );
  AOI22_X1 U14804 ( .A1(n12463), .A2(n12696), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12466) );
  NAND2_X1 U14805 ( .A1(n12464), .A2(n12861), .ZN(n12465) );
  OAI211_X1 U14806 ( .C1(n12467), .C2(n12651), .A(n12466), .B(n12465), .ZN(
        n12468) );
  AOI21_X1 U14807 ( .B1(n13060), .B2(n12469), .A(n12468), .ZN(n12470) );
  OAI21_X1 U14808 ( .B1(n12472), .B2(n12471), .A(n12470), .ZN(P3_U3180) );
  NAND2_X1 U14809 ( .A1(n6449), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U14810 ( .A1(n6447), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12475) );
  NAND2_X1 U14811 ( .A1(n8931), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12474) );
  INV_X1 U14812 ( .A(n12817), .ZN(n12694) );
  NAND2_X1 U14813 ( .A1(n12478), .A2(n12486), .ZN(n12480) );
  OR2_X1 U14814 ( .A1(n12487), .A2(n15053), .ZN(n12479) );
  INV_X1 U14815 ( .A(n12493), .ZN(n12695) );
  NAND2_X1 U14816 ( .A1(n13001), .A2(n12695), .ZN(n12490) );
  OAI21_X1 U14817 ( .B1(n12483), .B2(n12482), .A(n12481), .ZN(n12485) );
  XNOR2_X1 U14818 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12484) );
  XNOR2_X1 U14819 ( .A(n12485), .B(n12484), .ZN(n13135) );
  NAND2_X1 U14820 ( .A1(n13135), .A2(n12486), .ZN(n12489) );
  OR2_X1 U14821 ( .A1(n12487), .A2(n13130), .ZN(n12488) );
  NAND2_X1 U14822 ( .A1(n12489), .A2(n12488), .ZN(n12492) );
  AOI21_X1 U14823 ( .B1(n12694), .B2(n12490), .A(n13046), .ZN(n12678) );
  INV_X1 U14824 ( .A(n12678), .ZN(n12491) );
  INV_X1 U14825 ( .A(n12671), .ZN(n12518) );
  OR2_X1 U14826 ( .A1(n12492), .A2(n12817), .ZN(n12672) );
  NAND2_X1 U14827 ( .A1(n13047), .A2(n12493), .ZN(n12494) );
  NAND2_X1 U14828 ( .A1(n12672), .A2(n12494), .ZN(n12670) );
  INV_X1 U14829 ( .A(n12670), .ZN(n12517) );
  NAND2_X1 U14830 ( .A1(n12639), .A2(n12640), .ZN(n12900) );
  INV_X1 U14831 ( .A(n6779), .ZN(n12496) );
  NAND4_X1 U14832 ( .A1(n12497), .A2(n12496), .A3(n12534), .A4(n12495), .ZN(
        n12500) );
  NAND3_X1 U14833 ( .A1(n12547), .A2(n12498), .A3(n12552), .ZN(n12499) );
  NOR2_X1 U14834 ( .A1(n12500), .A2(n12499), .ZN(n12503) );
  AND4_X1 U14835 ( .A1(n12503), .A2(n12502), .A3(n12501), .A4(n12567), .ZN(
        n12504) );
  NAND4_X1 U14836 ( .A1(n14583), .A2(n12504), .A3(n12572), .A4(n14595), .ZN(
        n12505) );
  NOR2_X1 U14837 ( .A1(n12506), .A2(n12505), .ZN(n12508) );
  NAND4_X1 U14838 ( .A1(n12979), .A2(n12988), .A3(n12508), .A4(n12507), .ZN(
        n12509) );
  OR4_X1 U14839 ( .A1(n12938), .A2(n12626), .A3(n12966), .A4(n12509), .ZN(
        n12510) );
  OR4_X1 U14840 ( .A1(n12900), .A2(n12925), .A3(n7970), .A4(n12510), .ZN(
        n12511) );
  NOR2_X1 U14841 ( .A1(n12512), .A2(n12511), .ZN(n12513) );
  NAND4_X1 U14842 ( .A1(n12854), .A2(n12879), .A3(n12513), .A4(n12868), .ZN(
        n12514) );
  NOR4_X1 U14843 ( .A1(n12515), .A2(n12663), .A3(n12659), .A4(n12514), .ZN(
        n12516) );
  NAND3_X1 U14844 ( .A1(n12518), .A2(n12517), .A3(n12516), .ZN(n12519) );
  XNOR2_X1 U14845 ( .A(n12519), .B(n12680), .ZN(n12685) );
  NOR2_X1 U14846 ( .A1(n12520), .A2(n12656), .ZN(n12523) );
  AOI21_X1 U14847 ( .B1(n12523), .B2(n12522), .A(n12521), .ZN(n12667) );
  INV_X1 U14848 ( .A(n12524), .ZN(n12527) );
  OAI21_X1 U14849 ( .B1(n6779), .B2(n12525), .A(n12532), .ZN(n12526) );
  NAND3_X1 U14850 ( .A1(n6657), .A2(n12529), .A3(n12528), .ZN(n12530) );
  OAI21_X1 U14851 ( .B1(n14985), .B2(n12531), .A(n12530), .ZN(n12533) );
  NAND2_X1 U14852 ( .A1(n12533), .A2(n12532), .ZN(n12535) );
  NAND2_X1 U14853 ( .A1(n12535), .A2(n12534), .ZN(n12542) );
  NAND2_X1 U14854 ( .A1(n12545), .A2(n12536), .ZN(n12539) );
  NAND2_X1 U14855 ( .A1(n12544), .A2(n12537), .ZN(n12538) );
  INV_X1 U14856 ( .A(n12540), .ZN(n12541) );
  MUX2_X1 U14857 ( .A(n12545), .B(n12544), .S(n6458), .Z(n12546) );
  MUX2_X1 U14858 ( .A(n12550), .B(n12549), .S(n6458), .Z(n12551) );
  NAND2_X1 U14859 ( .A1(n12560), .A2(n12553), .ZN(n12554) );
  NAND2_X1 U14860 ( .A1(n12554), .A2(n6458), .ZN(n12555) );
  AOI21_X1 U14861 ( .B1(n12558), .B2(n12556), .A(n6458), .ZN(n12557) );
  AOI21_X1 U14862 ( .B1(n12559), .B2(n12558), .A(n12557), .ZN(n12563) );
  NOR2_X1 U14863 ( .A1(n12560), .A2(n6458), .ZN(n12562) );
  MUX2_X1 U14864 ( .A(n12565), .B(n12564), .S(n6458), .Z(n12566) );
  NAND3_X1 U14865 ( .A1(n12568), .A2(n12567), .A3(n12566), .ZN(n12573) );
  MUX2_X1 U14866 ( .A(n12570), .B(n12569), .S(n6458), .Z(n12571) );
  NAND3_X1 U14867 ( .A1(n12573), .A2(n12572), .A3(n12571), .ZN(n12579) );
  NAND2_X1 U14868 ( .A1(n12574), .A2(n6458), .ZN(n12576) );
  OR2_X1 U14869 ( .A1(n12574), .A2(n6458), .ZN(n12575) );
  MUX2_X1 U14870 ( .A(n12576), .B(n12575), .S(n12699), .Z(n12578) );
  INV_X1 U14871 ( .A(n12585), .ZN(n12581) );
  NAND3_X1 U14872 ( .A1(n12581), .A2(n14595), .A3(n12580), .ZN(n12588) );
  NAND2_X1 U14873 ( .A1(n14595), .A2(n12582), .ZN(n12584) );
  OAI211_X1 U14874 ( .C1(n12585), .C2(n12584), .A(n12589), .B(n12583), .ZN(
        n12586) );
  INV_X1 U14875 ( .A(n12586), .ZN(n12587) );
  MUX2_X1 U14876 ( .A(n12588), .B(n12587), .S(n6458), .Z(n12598) );
  MUX2_X1 U14877 ( .A(n12593), .B(n12589), .S(n12656), .Z(n12590) );
  NAND2_X1 U14878 ( .A1(n12591), .A2(n12590), .ZN(n12597) );
  AOI21_X1 U14879 ( .B1(n12593), .B2(n12592), .A(n12597), .ZN(n12595) );
  OAI21_X1 U14880 ( .B1(n12595), .B2(n12594), .A(n12656), .ZN(n12596) );
  INV_X1 U14881 ( .A(n12599), .ZN(n12600) );
  OAI33_X1 U14882 ( .A1(n12990), .A2(n12601), .A3(n12656), .B1(n12604), .B2(
        n7959), .B3(n12600), .ZN(n12609) );
  OAI22_X1 U14883 ( .A1(n12604), .A2(n7959), .B1(n12603), .B2(n12602), .ZN(
        n12605) );
  NAND2_X1 U14884 ( .A1(n12605), .A2(n12988), .ZN(n12607) );
  OAI211_X1 U14885 ( .C1(n7077), .C2(n13115), .A(n12607), .B(n12606), .ZN(
        n12608) );
  AOI21_X1 U14886 ( .B1(n12611), .B2(n12610), .A(n12656), .ZN(n12613) );
  NAND2_X1 U14887 ( .A1(n12991), .A2(n6458), .ZN(n12612) );
  OAI22_X1 U14888 ( .A1(n12614), .A2(n12613), .B1(n13115), .B2(n12612), .ZN(
        n12619) );
  INV_X1 U14889 ( .A(n12615), .ZN(n12617) );
  NAND3_X1 U14890 ( .A1(n12629), .A2(n6458), .A3(n12616), .ZN(n12621) );
  AOI22_X1 U14891 ( .A1(n12619), .A2(n12618), .B1(n12617), .B2(n12621), .ZN(
        n12627) );
  AND3_X1 U14892 ( .A1(n12628), .A2(n12656), .A3(n12622), .ZN(n12625) );
  INV_X1 U14893 ( .A(n12620), .ZN(n12623) );
  AOI21_X1 U14894 ( .B1(n12623), .B2(n12622), .A(n12621), .ZN(n12624) );
  OAI22_X1 U14895 ( .A1(n12627), .A2(n12626), .B1(n12625), .B2(n12624), .ZN(
        n12631) );
  MUX2_X1 U14896 ( .A(n12629), .B(n12628), .S(n6458), .Z(n12630) );
  NAND2_X1 U14897 ( .A1(n12932), .A2(n12940), .ZN(n12633) );
  MUX2_X1 U14898 ( .A(n12633), .B(n12632), .S(n6458), .Z(n12634) );
  MUX2_X1 U14899 ( .A(n12636), .B(n12635), .S(n12656), .Z(n12637) );
  MUX2_X1 U14900 ( .A(n12640), .B(n12639), .S(n6458), .Z(n12641) );
  OAI21_X1 U14901 ( .B1(n12642), .B2(n12644), .A(n12868), .ZN(n12655) );
  NAND2_X1 U14902 ( .A1(n13077), .A2(n12903), .ZN(n12643) );
  OAI21_X1 U14903 ( .B1(n12644), .B2(n12643), .A(n12645), .ZN(n12650) );
  INV_X1 U14904 ( .A(n12645), .ZN(n12646) );
  AOI21_X1 U14905 ( .B1(n12648), .B2(n12647), .A(n12646), .ZN(n12649) );
  MUX2_X1 U14906 ( .A(n12650), .B(n12649), .S(n12656), .Z(n12654) );
  MUX2_X1 U14907 ( .A(n6458), .B(n12651), .S(n13008), .Z(n12652) );
  OAI21_X1 U14908 ( .B1(n12656), .B2(n12881), .A(n12652), .ZN(n12653) );
  OAI211_X1 U14909 ( .C1(n12655), .C2(n12654), .A(n12854), .B(n12653), .ZN(
        n12661) );
  MUX2_X1 U14910 ( .A(n12658), .B(n12657), .S(n12656), .Z(n12660) );
  AOI21_X1 U14911 ( .B1(n12661), .B2(n12660), .A(n12659), .ZN(n12665) );
  NOR3_X1 U14912 ( .A1(n12662), .A2(n12857), .A3(n6458), .ZN(n12664) );
  INV_X1 U14913 ( .A(n12668), .ZN(n12669) );
  NOR2_X1 U14914 ( .A1(n12670), .A2(n12669), .ZN(n12679) );
  XNOR2_X1 U14915 ( .A(n12681), .B(n12680), .ZN(n12683) );
  NOR2_X1 U14916 ( .A1(n12683), .A2(n12682), .ZN(n12684) );
  NOR3_X1 U14917 ( .A1(n12689), .A2(n12688), .A3(n6710), .ZN(n12692) );
  OAI21_X1 U14918 ( .B1(n12693), .B2(n12690), .A(P3_B_REG_SCAN_IN), .ZN(n12691) );
  MUX2_X1 U14919 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12694), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14920 ( .A(n12695), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12706), .Z(
        P3_U3521) );
  MUX2_X1 U14921 ( .A(n12696), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12706), .Z(
        P3_U3518) );
  MUX2_X1 U14922 ( .A(n12871), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12706), .Z(
        P3_U3517) );
  MUX2_X1 U14923 ( .A(n12881), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12706), .Z(
        P3_U3516) );
  MUX2_X1 U14924 ( .A(n12892), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12706), .Z(
        P3_U3515) );
  MUX2_X1 U14925 ( .A(n12697), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12706), .Z(
        P3_U3514) );
  MUX2_X1 U14926 ( .A(n12893), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12706), .Z(
        P3_U3513) );
  MUX2_X1 U14927 ( .A(n12927), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12706), .Z(
        P3_U3512) );
  MUX2_X1 U14928 ( .A(n12698), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12706), .Z(
        P3_U3511) );
  MUX2_X1 U14929 ( .A(n12926), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12706), .Z(
        P3_U3510) );
  MUX2_X1 U14930 ( .A(n12969), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12706), .Z(
        P3_U3509) );
  MUX2_X1 U14931 ( .A(n12981), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12706), .Z(
        P3_U3508) );
  MUX2_X1 U14932 ( .A(n12980), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12706), .Z(
        P3_U3506) );
  MUX2_X1 U14933 ( .A(n12990), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12706), .Z(
        P3_U3505) );
  MUX2_X1 U14934 ( .A(n14577), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12706), .Z(
        P3_U3504) );
  MUX2_X1 U14935 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n14591), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14936 ( .A(n14576), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12706), .Z(
        P3_U3502) );
  MUX2_X1 U14937 ( .A(n14590), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12706), .Z(
        P3_U3501) );
  MUX2_X1 U14938 ( .A(n12699), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12706), .Z(
        P3_U3500) );
  MUX2_X1 U14939 ( .A(n12700), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12706), .Z(
        P3_U3499) );
  MUX2_X1 U14940 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12701), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14941 ( .A(n12702), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12706), .Z(
        P3_U3497) );
  MUX2_X1 U14942 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12703), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14943 ( .A(n12704), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12706), .Z(
        P3_U3495) );
  MUX2_X1 U14944 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n14989), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14945 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12705), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14946 ( .A(n6657), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12706), .Z(
        P3_U3491) );
  NAND2_X1 U14947 ( .A1(n14954), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U14948 ( .A1(n14923), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n12715) );
  NOR2_X1 U14949 ( .A1(n12707), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n12708) );
  OAI22_X1 U14950 ( .A1(n12709), .A2(n14936), .B1(n12712), .B2(n12708), .ZN(
        n12714) );
  OAI21_X1 U14951 ( .B1(n12712), .B2(n12711), .A(n12710), .ZN(n12713) );
  NAND4_X1 U14952 ( .A1(n12716), .A2(n12715), .A3(n12714), .A4(n12713), .ZN(
        P3_U3182) );
  INV_X1 U14953 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14563) );
  INV_X1 U14954 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13038) );
  OR2_X1 U14955 ( .A1(n12740), .A2(n13038), .ZN(n12750) );
  NAND2_X1 U14956 ( .A1(n12740), .A2(n13038), .ZN(n12719) );
  NAND2_X1 U14957 ( .A1(n12750), .A2(n12719), .ZN(n12721) );
  INV_X1 U14958 ( .A(n12751), .ZN(n12720) );
  AOI21_X1 U14959 ( .B1(n12722), .B2(n12721), .A(n12720), .ZN(n12749) );
  MUX2_X1 U14960 ( .A(n12736), .B(n12723), .S(n11411), .Z(n12724) );
  NAND2_X1 U14961 ( .A1(n12725), .A2(n12724), .ZN(n12726) );
  INV_X1 U14962 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14558) );
  MUX2_X1 U14963 ( .A(n14558), .B(n14563), .S(n11411), .Z(n14564) );
  NOR2_X1 U14964 ( .A1(n12727), .A2(n14567), .ZN(n12761) );
  INV_X1 U14965 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12983) );
  MUX2_X1 U14966 ( .A(n12983), .B(n13038), .S(n11411), .Z(n12728) );
  NAND2_X1 U14967 ( .A1(n12740), .A2(n12728), .ZN(n12760) );
  NOR2_X1 U14968 ( .A1(n12740), .A2(n12728), .ZN(n12762) );
  INV_X1 U14969 ( .A(n12762), .ZN(n12729) );
  NAND2_X1 U14970 ( .A1(n12760), .A2(n12729), .ZN(n12730) );
  XNOR2_X1 U14971 ( .A(n12761), .B(n12730), .ZN(n12747) );
  AOI21_X1 U14972 ( .B1(n14923), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12731), 
        .ZN(n12732) );
  OAI21_X1 U14973 ( .B1(n14966), .B2(n12733), .A(n12732), .ZN(n12746) );
  NOR2_X1 U14974 ( .A1(n12737), .A2(n12738), .ZN(n12739) );
  OR2_X1 U14975 ( .A1(n12740), .A2(n12983), .ZN(n12753) );
  NAND2_X1 U14976 ( .A1(n12740), .A2(n12983), .ZN(n12741) );
  NAND2_X1 U14977 ( .A1(n12753), .A2(n12741), .ZN(n12742) );
  NAND2_X1 U14978 ( .A1(n12743), .A2(n12742), .ZN(n12744) );
  AOI21_X1 U14979 ( .B1(n12754), .B2(n12744), .A(n14983), .ZN(n12745) );
  AOI211_X1 U14980 ( .C1(n14936), .C2(n12747), .A(n12746), .B(n12745), .ZN(
        n12748) );
  OAI21_X1 U14981 ( .B1(n12749), .B2(n14977), .A(n12748), .ZN(P3_U3198) );
  INV_X1 U14982 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13035) );
  AOI21_X1 U14983 ( .B1(n13035), .B2(n12752), .A(n12770), .ZN(n12768) );
  INV_X1 U14984 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12755) );
  AOI21_X1 U14985 ( .B1(n12756), .B2(n12755), .A(n12786), .ZN(n12759) );
  AOI21_X1 U14986 ( .B1(n14923), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12757), 
        .ZN(n12758) );
  OAI21_X1 U14987 ( .B1(n12759), .B2(n14983), .A(n12758), .ZN(n12766) );
  MUX2_X1 U14988 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n11411), .Z(n12777) );
  XNOR2_X1 U14989 ( .A(n12778), .B(n12777), .ZN(n12763) );
  NOR2_X1 U14990 ( .A1(n12764), .A2(n12763), .ZN(n12776) );
  AOI211_X1 U14991 ( .C1(n12764), .C2(n12763), .A(n12776), .B(n14975), .ZN(
        n12765) );
  AOI211_X1 U14992 ( .C1(n14954), .C2(n12785), .A(n12766), .B(n12765), .ZN(
        n12767) );
  OAI21_X1 U14993 ( .B1(n12768), .B2(n14977), .A(n12767), .ZN(P3_U3199) );
  NOR2_X1 U14994 ( .A1(n12785), .A2(n12769), .ZN(n12771) );
  NAND2_X1 U14995 ( .A1(n12788), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12795) );
  OAI21_X1 U14996 ( .B1(n12788), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12795), 
        .ZN(n12772) );
  NOR2_X1 U14997 ( .A1(n12773), .A2(n12772), .ZN(n12797) );
  AOI21_X1 U14998 ( .B1(n12773), .B2(n12772), .A(n12797), .ZN(n12794) );
  OAI21_X1 U14999 ( .B1(n14967), .B2(n12775), .A(n12774), .ZN(n12783) );
  MUX2_X1 U15000 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n11411), .Z(n12780) );
  XNOR2_X1 U15001 ( .A(n12803), .B(n12802), .ZN(n12779) );
  NOR2_X1 U15002 ( .A1(n12779), .A2(n12780), .ZN(n12801) );
  AOI21_X1 U15003 ( .B1(n12780), .B2(n12779), .A(n12801), .ZN(n12781) );
  NOR2_X1 U15004 ( .A1(n12781), .A2(n14975), .ZN(n12782) );
  AOI211_X1 U15005 ( .C1(n14954), .C2(n12802), .A(n12783), .B(n12782), .ZN(
        n12793) );
  NOR2_X1 U15006 ( .A1(n12785), .A2(n12784), .ZN(n12787) );
  NAND2_X1 U15007 ( .A1(n12788), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12809) );
  OAI21_X1 U15008 ( .B1(n12788), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12809), 
        .ZN(n12789) );
  AOI21_X1 U15009 ( .B1(n12790), .B2(n12789), .A(n12810), .ZN(n12791) );
  OR2_X1 U15010 ( .A1(n12791), .A2(n14983), .ZN(n12792) );
  OAI211_X1 U15011 ( .C1(n12794), .C2(n14977), .A(n12793), .B(n12792), .ZN(
        P3_U3200) );
  INV_X1 U15012 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13025) );
  XNOR2_X1 U15013 ( .A(n12808), .B(n13025), .ZN(n12800) );
  INV_X1 U15014 ( .A(n12795), .ZN(n12796) );
  INV_X1 U15015 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12798) );
  MUX2_X1 U15016 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n12798), .S(n12808), .Z(
        n12811) );
  MUX2_X1 U15017 ( .A(n12811), .B(n12800), .S(n11411), .Z(n12805) );
  AOI21_X1 U15018 ( .B1(n12803), .B2(n12802), .A(n12801), .ZN(n12804) );
  NAND2_X1 U15019 ( .A1(n14923), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12806) );
  OAI211_X1 U15020 ( .C1(n14966), .C2(n12808), .A(n12807), .B(n12806), .ZN(
        n12812) );
  OAI21_X1 U15021 ( .B1(n12815), .B2(n14977), .A(n12814), .ZN(P3_U3201) );
  NAND2_X1 U15022 ( .A1(n14998), .A2(n12818), .ZN(n12823) );
  OAI21_X1 U15023 ( .B1(n15004), .B2(n13044), .A(n12823), .ZN(n12820) );
  AOI21_X1 U15024 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15004), .A(n12820), 
        .ZN(n12819) );
  OAI21_X1 U15025 ( .B1(n13046), .B2(n12847), .A(n12819), .ZN(P3_U3202) );
  AOI21_X1 U15026 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n15004), .A(n12820), 
        .ZN(n12821) );
  OAI21_X1 U15027 ( .B1(n13001), .B2(n12847), .A(n12821), .ZN(P3_U3203) );
  NAND2_X1 U15028 ( .A1(n12822), .A2(n15002), .ZN(n12828) );
  INV_X1 U15029 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12824) );
  OAI21_X1 U15030 ( .B1(n15002), .B2(n12824), .A(n12823), .ZN(n12825) );
  AOI21_X1 U15031 ( .B1(n12826), .B2(n14598), .A(n12825), .ZN(n12827) );
  OAI211_X1 U15032 ( .C1(n12829), .C2(n12997), .A(n12828), .B(n12827), .ZN(
        P3_U3204) );
  XNOR2_X1 U15033 ( .A(n12830), .B(n12833), .ZN(n13057) );
  NAND2_X1 U15034 ( .A1(n12832), .A2(n12831), .ZN(n12834) );
  NAND2_X1 U15035 ( .A1(n12834), .A2(n12833), .ZN(n12836) );
  OAI22_X1 U15036 ( .A1(n12837), .A2(n12958), .B1(n12857), .B2(n12956), .ZN(
        n12838) );
  INV_X1 U15037 ( .A(n12838), .ZN(n12839) );
  AND2_X2 U15038 ( .A1(n12840), .A2(n12839), .ZN(n13052) );
  AOI22_X1 U15039 ( .A1(n13054), .A2(n12994), .B1(n14998), .B2(n12841), .ZN(
        n12842) );
  OAI211_X1 U15040 ( .C1(n13057), .C2(n12997), .A(n12843), .B(n12842), .ZN(
        P3_U3205) );
  INV_X1 U15041 ( .A(n12844), .ZN(n12851) );
  AOI22_X1 U15042 ( .A1(n15004), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n14998), 
        .B2(n12845), .ZN(n12846) );
  OAI21_X1 U15043 ( .B1(n12848), .B2(n12847), .A(n12846), .ZN(n12849) );
  AOI21_X1 U15044 ( .B1(n6763), .B2(n14999), .A(n12849), .ZN(n12850) );
  OAI21_X1 U15045 ( .B1(n12851), .B2(n15004), .A(n12850), .ZN(P3_U3206) );
  INV_X1 U15046 ( .A(n12854), .ZN(n12852) );
  XNOR2_X1 U15047 ( .A(n12853), .B(n12852), .ZN(n13063) );
  XNOR2_X1 U15048 ( .A(n12855), .B(n12854), .ZN(n12859) );
  NAND2_X1 U15049 ( .A1(n12881), .A2(n14987), .ZN(n12856) );
  OAI21_X1 U15050 ( .B1(n12857), .B2(n12958), .A(n12856), .ZN(n12858) );
  AOI21_X1 U15051 ( .B1(n12859), .B2(n14991), .A(n12858), .ZN(n13059) );
  INV_X1 U15052 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12860) );
  MUX2_X1 U15053 ( .A(n13059), .B(n12860), .S(n15004), .Z(n12863) );
  AOI22_X1 U15054 ( .A1(n13060), .A2(n12994), .B1(n14998), .B2(n12861), .ZN(
        n12862) );
  OAI211_X1 U15055 ( .C1(n13063), .C2(n12997), .A(n12863), .B(n12862), .ZN(
        P3_U3207) );
  OR2_X1 U15056 ( .A1(n12864), .A2(n12868), .ZN(n12865) );
  AND2_X1 U15057 ( .A1(n12866), .A2(n12865), .ZN(n13066) );
  NAND2_X1 U15058 ( .A1(n12869), .A2(n12868), .ZN(n12870) );
  NAND3_X1 U15059 ( .A1(n12867), .A2(n14991), .A3(n12870), .ZN(n12873) );
  AOI22_X1 U15060 ( .A1(n14988), .A2(n12871), .B1(n12892), .B2(n14987), .ZN(
        n12872) );
  NAND2_X1 U15061 ( .A1(n12873), .A2(n12872), .ZN(n13064) );
  MUX2_X1 U15062 ( .A(n13064), .B(P3_REG2_REG_25__SCAN_IN), .S(n15004), .Z(
        n12874) );
  INV_X1 U15063 ( .A(n12874), .ZN(n12877) );
  AOI22_X1 U15064 ( .A1(n13008), .A2(n12994), .B1(n14998), .B2(n12875), .ZN(
        n12876) );
  OAI211_X1 U15065 ( .C1(n13066), .C2(n12997), .A(n12877), .B(n12876), .ZN(
        P3_U3208) );
  XNOR2_X1 U15066 ( .A(n12878), .B(n12879), .ZN(n13074) );
  INV_X1 U15067 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12885) );
  XNOR2_X1 U15068 ( .A(n12880), .B(n12879), .ZN(n12884) );
  NAND2_X1 U15069 ( .A1(n12881), .A2(n14988), .ZN(n12882) );
  OAI21_X1 U15070 ( .B1(n12903), .B2(n12956), .A(n12882), .ZN(n12883) );
  AOI21_X1 U15071 ( .B1(n12884), .B2(n14991), .A(n12883), .ZN(n13069) );
  MUX2_X1 U15072 ( .A(n12885), .B(n13069), .S(n15002), .Z(n12888) );
  AOI22_X1 U15073 ( .A1(n13071), .A2(n12994), .B1(n14998), .B2(n12886), .ZN(
        n12887) );
  OAI211_X1 U15074 ( .C1(n13074), .C2(n12997), .A(n12888), .B(n12887), .ZN(
        P3_U3209) );
  XNOR2_X1 U15075 ( .A(n12889), .B(n12891), .ZN(n13080) );
  INV_X1 U15076 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12895) );
  XNOR2_X1 U15077 ( .A(n12890), .B(n12891), .ZN(n12894) );
  AOI222_X1 U15078 ( .A1(n14991), .A2(n12894), .B1(n12893), .B2(n14987), .C1(
        n12892), .C2(n14988), .ZN(n13075) );
  MUX2_X1 U15079 ( .A(n12895), .B(n13075), .S(n15002), .Z(n12898) );
  AOI22_X1 U15080 ( .A1(n13077), .A2(n12994), .B1(n14998), .B2(n12896), .ZN(
        n12897) );
  OAI211_X1 U15081 ( .C1(n13080), .C2(n12997), .A(n12898), .B(n12897), .ZN(
        P3_U3210) );
  XOR2_X1 U15082 ( .A(n12899), .B(n12900), .Z(n13085) );
  XNOR2_X1 U15083 ( .A(n12901), .B(n12900), .ZN(n12905) );
  OAI22_X1 U15084 ( .A1(n12903), .A2(n12958), .B1(n12902), .B2(n12956), .ZN(
        n12904) );
  AOI21_X1 U15085 ( .B1(n12905), .B2(n14991), .A(n12904), .ZN(n13081) );
  INV_X1 U15086 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12906) );
  MUX2_X1 U15087 ( .A(n13081), .B(n12906), .S(n15004), .Z(n12909) );
  AOI22_X1 U15088 ( .A1(n13082), .A2(n12994), .B1(n14998), .B2(n12907), .ZN(
        n12908) );
  OAI211_X1 U15089 ( .C1(n13085), .C2(n12997), .A(n12909), .B(n12908), .ZN(
        P3_U3211) );
  INV_X1 U15090 ( .A(n12910), .ZN(n12911) );
  AOI21_X1 U15091 ( .B1(n12915), .B2(n12912), .A(n12911), .ZN(n12913) );
  OAI222_X1 U15092 ( .A1(n12958), .A2(n12914), .B1(n12956), .B2(n12940), .C1(
        n12954), .C2(n12913), .ZN(n13020) );
  XNOR2_X1 U15093 ( .A(n12916), .B(n12915), .ZN(n13089) );
  AOI22_X1 U15094 ( .A1(n15004), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n14998), 
        .B2(n12917), .ZN(n12919) );
  NAND2_X1 U15095 ( .A1(n13021), .A2(n12994), .ZN(n12918) );
  OAI211_X1 U15096 ( .C1(n13089), .C2(n12997), .A(n12919), .B(n12918), .ZN(
        n12920) );
  AOI21_X1 U15097 ( .B1(n13020), .B2(n15002), .A(n12920), .ZN(n12921) );
  INV_X1 U15098 ( .A(n12921), .ZN(P3_U3212) );
  XNOR2_X1 U15099 ( .A(n12922), .B(n12925), .ZN(n13092) );
  OAI211_X1 U15100 ( .C1(n12925), .C2(n12924), .A(n12923), .B(n14991), .ZN(
        n12929) );
  AOI22_X1 U15101 ( .A1(n12927), .A2(n14988), .B1(n14987), .B2(n12926), .ZN(
        n12928) );
  NAND2_X1 U15102 ( .A1(n12929), .A2(n12928), .ZN(n13090) );
  MUX2_X1 U15103 ( .A(n13090), .B(P3_REG2_REG_20__SCAN_IN), .S(n15004), .Z(
        n12930) );
  INV_X1 U15104 ( .A(n12930), .ZN(n12934) );
  AOI22_X1 U15105 ( .A1(n12932), .A2(n12994), .B1(n14998), .B2(n12931), .ZN(
        n12933) );
  OAI211_X1 U15106 ( .C1(n13092), .C2(n12997), .A(n12934), .B(n12933), .ZN(
        P3_U3213) );
  INV_X1 U15107 ( .A(n12938), .ZN(n12935) );
  XNOR2_X1 U15108 ( .A(n12936), .B(n12935), .ZN(n13099) );
  OAI211_X1 U15109 ( .C1(n12939), .C2(n12938), .A(n12937), .B(n14991), .ZN(
        n12944) );
  OAI22_X1 U15110 ( .A1(n12941), .A2(n12956), .B1(n12940), .B2(n12958), .ZN(
        n12942) );
  INV_X1 U15111 ( .A(n12942), .ZN(n12943) );
  NAND2_X1 U15112 ( .A1(n12944), .A2(n12943), .ZN(n13095) );
  MUX2_X1 U15113 ( .A(n13095), .B(P3_REG2_REG_19__SCAN_IN), .S(n15004), .Z(
        n12945) );
  INV_X1 U15114 ( .A(n12945), .ZN(n12949) );
  INV_X1 U15115 ( .A(n13098), .ZN(n12947) );
  AOI22_X1 U15116 ( .A1(n12947), .A2(n12994), .B1(n14998), .B2(n12946), .ZN(
        n12948) );
  OAI211_X1 U15117 ( .C1(n13099), .C2(n12997), .A(n12949), .B(n12948), .ZN(
        P3_U3214) );
  OAI21_X1 U15118 ( .B1(n6592), .B2(n12952), .A(n12950), .ZN(n13106) );
  AOI21_X1 U15119 ( .B1(n12952), .B2(n12951), .A(n6541), .ZN(n12953) );
  OAI222_X1 U15120 ( .A1(n12958), .A2(n12957), .B1(n12956), .B2(n12955), .C1(
        n12954), .C2(n12953), .ZN(n13031) );
  NAND2_X1 U15121 ( .A1(n13031), .A2(n15002), .ZN(n12964) );
  INV_X1 U15122 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12961) );
  INV_X1 U15123 ( .A(n12959), .ZN(n12960) );
  OAI22_X1 U15124 ( .A1(n15002), .A2(n12961), .B1(n12960), .B2(n14580), .ZN(
        n12962) );
  AOI21_X1 U15125 ( .B1(n13032), .B2(n12994), .A(n12962), .ZN(n12963) );
  OAI211_X1 U15126 ( .C1(n13106), .C2(n12997), .A(n12964), .B(n12963), .ZN(
        P3_U3215) );
  XNOR2_X1 U15127 ( .A(n12965), .B(n12966), .ZN(n13112) );
  XNOR2_X1 U15128 ( .A(n12967), .B(n12966), .ZN(n12968) );
  NAND2_X1 U15129 ( .A1(n12968), .A2(n14991), .ZN(n12971) );
  AOI22_X1 U15130 ( .A1(n12969), .A2(n14988), .B1(n14987), .B2(n12991), .ZN(
        n12970) );
  MUX2_X1 U15131 ( .A(n12755), .B(n13107), .S(n15002), .Z(n12974) );
  AOI22_X1 U15132 ( .A1(n13109), .A2(n12994), .B1(n14998), .B2(n12972), .ZN(
        n12973) );
  OAI211_X1 U15133 ( .C1(n13112), .C2(n12997), .A(n12974), .B(n12973), .ZN(
        P3_U3216) );
  OAI21_X1 U15134 ( .B1(n12976), .B2(n12979), .A(n12975), .ZN(n12977) );
  INV_X1 U15135 ( .A(n12977), .ZN(n13118) );
  XNOR2_X1 U15136 ( .A(n6766), .B(n12979), .ZN(n12982) );
  AOI222_X1 U15137 ( .A1(n14991), .A2(n12982), .B1(n12981), .B2(n14988), .C1(
        n12980), .C2(n14987), .ZN(n13113) );
  MUX2_X1 U15138 ( .A(n12983), .B(n13113), .S(n15002), .Z(n12986) );
  AOI22_X1 U15139 ( .A1(n13115), .A2(n12994), .B1(n14998), .B2(n12984), .ZN(
        n12985) );
  OAI211_X1 U15140 ( .C1(n13118), .C2(n12997), .A(n12986), .B(n12985), .ZN(
        P3_U3217) );
  XOR2_X1 U15141 ( .A(n12987), .B(n12988), .Z(n13126) );
  XNOR2_X1 U15142 ( .A(n12989), .B(n12988), .ZN(n12992) );
  AOI222_X1 U15143 ( .A1(n14991), .A2(n12992), .B1(n12991), .B2(n14988), .C1(
        n12990), .C2(n14987), .ZN(n13119) );
  MUX2_X1 U15144 ( .A(n14558), .B(n13119), .S(n15002), .Z(n12996) );
  AOI22_X1 U15145 ( .A1(n13122), .A2(n12994), .B1(n14998), .B2(n12993), .ZN(
        n12995) );
  OAI211_X1 U15146 ( .C1(n13126), .C2(n12997), .A(n12996), .B(n12995), .ZN(
        P3_U3218) );
  NOR2_X1 U15147 ( .A1(n15049), .A2(n13044), .ZN(n12999) );
  AOI21_X1 U15148 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15049), .A(n12999), 
        .ZN(n12998) );
  OAI21_X1 U15149 ( .B1(n13046), .B2(n13027), .A(n12998), .ZN(P3_U3490) );
  AOI21_X1 U15150 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15049), .A(n12999), 
        .ZN(n13000) );
  OAI21_X1 U15151 ( .B1(n13001), .B2(n13027), .A(n13000), .ZN(P3_U3489) );
  INV_X1 U15152 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13002) );
  MUX2_X1 U15153 ( .A(n13002), .B(n13052), .S(n15051), .Z(n13004) );
  NAND2_X1 U15154 ( .A1(n13054), .A2(n8048), .ZN(n13003) );
  INV_X1 U15155 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13005) );
  MUX2_X1 U15156 ( .A(n13059), .B(n13005), .S(n15049), .Z(n13007) );
  NAND2_X1 U15157 ( .A1(n13060), .A2(n8048), .ZN(n13006) );
  OAI211_X1 U15158 ( .C1(n13043), .C2(n13063), .A(n13007), .B(n13006), .ZN(
        P3_U3485) );
  MUX2_X1 U15159 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13064), .S(n15051), .Z(
        n13010) );
  INV_X1 U15160 ( .A(n13008), .ZN(n13065) );
  OAI22_X1 U15161 ( .A1(n13066), .A2(n13043), .B1(n13065), .B2(n13027), .ZN(
        n13009) );
  OR2_X1 U15162 ( .A1(n13010), .A2(n13009), .ZN(P3_U3484) );
  INV_X1 U15163 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13011) );
  MUX2_X1 U15164 ( .A(n13011), .B(n13069), .S(n15051), .Z(n13013) );
  NAND2_X1 U15165 ( .A1(n13071), .A2(n8048), .ZN(n13012) );
  OAI211_X1 U15166 ( .C1(n13074), .C2(n13043), .A(n13013), .B(n13012), .ZN(
        P3_U3483) );
  INV_X1 U15167 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13014) );
  MUX2_X1 U15168 ( .A(n13014), .B(n13075), .S(n15051), .Z(n13016) );
  NAND2_X1 U15169 ( .A1(n13077), .A2(n8048), .ZN(n13015) );
  OAI211_X1 U15170 ( .C1(n13043), .C2(n13080), .A(n13016), .B(n13015), .ZN(
        P3_U3482) );
  INV_X1 U15171 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13017) );
  MUX2_X1 U15172 ( .A(n13017), .B(n13081), .S(n15051), .Z(n13019) );
  NAND2_X1 U15173 ( .A1(n13082), .A2(n8048), .ZN(n13018) );
  OAI211_X1 U15174 ( .C1(n13085), .C2(n13043), .A(n13019), .B(n13018), .ZN(
        P3_U3481) );
  INV_X1 U15175 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n15123) );
  AOI21_X1 U15176 ( .B1(n15015), .B2(n13021), .A(n13020), .ZN(n13086) );
  MUX2_X1 U15177 ( .A(n15123), .B(n13086), .S(n15051), .Z(n13022) );
  OAI21_X1 U15178 ( .B1(n13089), .B2(n13043), .A(n13022), .ZN(P3_U3480) );
  MUX2_X1 U15179 ( .A(n13090), .B(P3_REG1_REG_20__SCAN_IN), .S(n15049), .Z(
        n13024) );
  OAI22_X1 U15180 ( .A1(n13092), .A2(n13043), .B1(n13091), .B2(n13027), .ZN(
        n13023) );
  OR2_X1 U15181 ( .A1(n13024), .A2(n13023), .ZN(P3_U3479) );
  INV_X1 U15182 ( .A(n13095), .ZN(n13026) );
  MUX2_X1 U15183 ( .A(n13026), .B(n13025), .S(n15049), .Z(n13030) );
  OAI22_X1 U15184 ( .A1(n13099), .A2(n13043), .B1(n13098), .B2(n13027), .ZN(
        n13028) );
  INV_X1 U15185 ( .A(n13028), .ZN(n13029) );
  NAND2_X1 U15186 ( .A1(n13030), .A2(n13029), .ZN(P3_U3478) );
  INV_X1 U15187 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13033) );
  AOI21_X1 U15188 ( .B1(n15015), .B2(n13032), .A(n13031), .ZN(n13103) );
  MUX2_X1 U15189 ( .A(n13033), .B(n13103), .S(n15051), .Z(n13034) );
  OAI21_X1 U15190 ( .B1(n13043), .B2(n13106), .A(n13034), .ZN(P3_U3477) );
  MUX2_X1 U15191 ( .A(n13035), .B(n13107), .S(n15051), .Z(n13037) );
  NAND2_X1 U15192 ( .A1(n13109), .A2(n8048), .ZN(n13036) );
  OAI211_X1 U15193 ( .C1(n13043), .C2(n13112), .A(n13037), .B(n13036), .ZN(
        P3_U3476) );
  MUX2_X1 U15194 ( .A(n13038), .B(n13113), .S(n15051), .Z(n13040) );
  NAND2_X1 U15195 ( .A1(n13115), .A2(n8048), .ZN(n13039) );
  OAI211_X1 U15196 ( .C1(n13118), .C2(n13043), .A(n13040), .B(n13039), .ZN(
        P3_U3475) );
  MUX2_X1 U15197 ( .A(n14563), .B(n13119), .S(n15051), .Z(n13042) );
  NAND2_X1 U15198 ( .A1(n13122), .A2(n8048), .ZN(n13041) );
  OAI211_X1 U15199 ( .C1(n13043), .C2(n13126), .A(n13042), .B(n13041), .ZN(
        P3_U3474) );
  NOR2_X1 U15200 ( .A1(n15037), .A2(n13044), .ZN(n13048) );
  AOI21_X1 U15201 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15037), .A(n13048), 
        .ZN(n13045) );
  OAI21_X1 U15202 ( .B1(n13046), .B2(n13097), .A(n13045), .ZN(P3_U3458) );
  INV_X1 U15203 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13051) );
  NAND2_X1 U15204 ( .A1(n13047), .A2(n13121), .ZN(n13050) );
  INV_X1 U15205 ( .A(n13048), .ZN(n13049) );
  OAI211_X1 U15206 ( .C1(n13051), .C2(n15039), .A(n13050), .B(n13049), .ZN(
        P3_U3457) );
  INV_X1 U15207 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13053) );
  MUX2_X1 U15208 ( .A(n13053), .B(n13052), .S(n15039), .Z(n13056) );
  NAND2_X1 U15209 ( .A1(n13054), .A2(n13121), .ZN(n13055) );
  INV_X1 U15210 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13058) );
  MUX2_X1 U15211 ( .A(n13059), .B(n13058), .S(n15037), .Z(n13062) );
  NAND2_X1 U15212 ( .A1(n13060), .A2(n13121), .ZN(n13061) );
  OAI211_X1 U15213 ( .C1(n13063), .C2(n13125), .A(n13062), .B(n13061), .ZN(
        P3_U3453) );
  MUX2_X1 U15214 ( .A(n13064), .B(P3_REG0_REG_25__SCAN_IN), .S(n15037), .Z(
        n13068) );
  OAI22_X1 U15215 ( .A1(n13066), .A2(n13125), .B1(n13065), .B2(n13097), .ZN(
        n13067) );
  OR2_X1 U15216 ( .A1(n13068), .A2(n13067), .ZN(P3_U3452) );
  INV_X1 U15217 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13070) );
  MUX2_X1 U15218 ( .A(n13070), .B(n13069), .S(n15039), .Z(n13073) );
  NAND2_X1 U15219 ( .A1(n13071), .A2(n13121), .ZN(n13072) );
  OAI211_X1 U15220 ( .C1(n13074), .C2(n13125), .A(n13073), .B(n13072), .ZN(
        P3_U3451) );
  INV_X1 U15221 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13076) );
  MUX2_X1 U15222 ( .A(n13076), .B(n13075), .S(n15039), .Z(n13079) );
  NAND2_X1 U15223 ( .A1(n13077), .A2(n13121), .ZN(n13078) );
  OAI211_X1 U15224 ( .C1(n13080), .C2(n13125), .A(n13079), .B(n13078), .ZN(
        P3_U3450) );
  INV_X1 U15225 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n15095) );
  MUX2_X1 U15226 ( .A(n13081), .B(n15095), .S(n15037), .Z(n13084) );
  NAND2_X1 U15227 ( .A1(n13082), .A2(n13121), .ZN(n13083) );
  OAI211_X1 U15228 ( .C1(n13085), .C2(n13125), .A(n13084), .B(n13083), .ZN(
        P3_U3449) );
  INV_X1 U15229 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13087) );
  MUX2_X1 U15230 ( .A(n13087), .B(n13086), .S(n15039), .Z(n13088) );
  OAI21_X1 U15231 ( .B1(n13089), .B2(n13125), .A(n13088), .ZN(P3_U3448) );
  MUX2_X1 U15232 ( .A(n13090), .B(P3_REG0_REG_20__SCAN_IN), .S(n15037), .Z(
        n13094) );
  OAI22_X1 U15233 ( .A1(n13092), .A2(n13125), .B1(n13091), .B2(n13097), .ZN(
        n13093) );
  OR2_X1 U15234 ( .A1(n13094), .A2(n13093), .ZN(P3_U3447) );
  MUX2_X1 U15235 ( .A(n13095), .B(P3_REG0_REG_19__SCAN_IN), .S(n15037), .Z(
        n13096) );
  INV_X1 U15236 ( .A(n13096), .ZN(n13102) );
  OAI22_X1 U15237 ( .A1(n13099), .A2(n13125), .B1(n13098), .B2(n13097), .ZN(
        n13100) );
  INV_X1 U15238 ( .A(n13100), .ZN(n13101) );
  NAND2_X1 U15239 ( .A1(n13102), .A2(n13101), .ZN(P3_U3446) );
  INV_X1 U15240 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13104) );
  MUX2_X1 U15241 ( .A(n13104), .B(n13103), .S(n15039), .Z(n13105) );
  OAI21_X1 U15242 ( .B1(n13106), .B2(n13125), .A(n13105), .ZN(P3_U3444) );
  INV_X1 U15243 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13108) );
  MUX2_X1 U15244 ( .A(n13108), .B(n13107), .S(n15039), .Z(n13111) );
  NAND2_X1 U15245 ( .A1(n13109), .A2(n13121), .ZN(n13110) );
  OAI211_X1 U15246 ( .C1(n13112), .C2(n13125), .A(n13111), .B(n13110), .ZN(
        P3_U3441) );
  INV_X1 U15247 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13114) );
  MUX2_X1 U15248 ( .A(n13114), .B(n13113), .S(n15039), .Z(n13117) );
  NAND2_X1 U15249 ( .A1(n13115), .A2(n13121), .ZN(n13116) );
  OAI211_X1 U15250 ( .C1(n13118), .C2(n13125), .A(n13117), .B(n13116), .ZN(
        P3_U3438) );
  INV_X1 U15251 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13120) );
  MUX2_X1 U15252 ( .A(n13120), .B(n13119), .S(n15039), .Z(n13124) );
  NAND2_X1 U15253 ( .A1(n13122), .A2(n13121), .ZN(n13123) );
  OAI211_X1 U15254 ( .C1(n13126), .C2(n13125), .A(n13124), .B(n13123), .ZN(
        P3_U3435) );
  MUX2_X1 U15255 ( .A(n13128), .B(P3_D_REG_0__SCAN_IN), .S(n13127), .Z(
        P3_U3376) );
  NAND3_X1 U15256 ( .A1(n13129), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13131) );
  OAI22_X1 U15257 ( .A1(n13132), .A2(n13131), .B1(n13130), .B2(n13142), .ZN(
        n13133) );
  AOI21_X1 U15258 ( .B1(n13135), .B2(n13134), .A(n13133), .ZN(n13136) );
  INV_X1 U15259 ( .A(n13136), .ZN(P3_U3264) );
  INV_X1 U15260 ( .A(n13137), .ZN(n13139) );
  OAI222_X1 U15261 ( .A1(n13142), .A2(n13141), .B1(n13140), .B2(n13139), .C1(
        P3_U3151), .C2(n13138), .ZN(P3_U3266) );
  INV_X1 U15262 ( .A(n13406), .ZN(n13523) );
  AOI22_X1 U15263 ( .A1(n13143), .A2(n9485), .B1(n13270), .B2(n13523), .ZN(
        n13149) );
  NOR2_X1 U15264 ( .A1(n13233), .A2(n13630), .ZN(n13144) );
  AOI21_X1 U15265 ( .B1(n13408), .B2(n13544), .A(n13144), .ZN(n13518) );
  INV_X1 U15266 ( .A(n13145), .ZN(n13510) );
  AOI22_X1 U15267 ( .A1(n13510), .A2(n13240), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13146) );
  OAI21_X1 U15268 ( .B1(n13518), .B2(n13199), .A(n13146), .ZN(n13147) );
  AOI21_X1 U15269 ( .B1(n13698), .B2(n13281), .A(n13147), .ZN(n13148) );
  OAI21_X1 U15270 ( .B1(n13150), .B2(n13149), .A(n13148), .ZN(P2_U3188) );
  XNOR2_X1 U15271 ( .A(n6803), .B(n13152), .ZN(n13153) );
  XNOR2_X1 U15272 ( .A(n13222), .B(n13153), .ZN(n13160) );
  INV_X1 U15273 ( .A(n13576), .ZN(n13157) );
  NAND2_X1 U15274 ( .A1(n13543), .A2(n13544), .ZN(n13155) );
  NAND2_X1 U15275 ( .A1(n13359), .A2(n13542), .ZN(n13154) );
  NAND2_X1 U15276 ( .A1(n13155), .A2(n13154), .ZN(n13571) );
  NAND2_X1 U15277 ( .A1(n13571), .A2(n13251), .ZN(n13156) );
  NAND2_X1 U15278 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13333)
         );
  OAI211_X1 U15279 ( .C1(n13276), .C2(n13157), .A(n13156), .B(n13333), .ZN(
        n13158) );
  AOI21_X1 U15280 ( .B1(n13720), .B2(n13281), .A(n13158), .ZN(n13159) );
  OAI21_X1 U15281 ( .B1(n13160), .B2(n13272), .A(n13159), .ZN(P2_U3191) );
  INV_X1 U15282 ( .A(n13161), .ZN(n13162) );
  NAND2_X1 U15283 ( .A1(n13379), .A2(n9321), .ZN(n13165) );
  XNOR2_X1 U15284 ( .A(n13165), .B(n13164), .ZN(n13166) );
  XNOR2_X1 U15285 ( .A(n13428), .B(n13166), .ZN(n13167) );
  XNOR2_X1 U15286 ( .A(n13168), .B(n13167), .ZN(n13174) );
  OAI22_X1 U15287 ( .A1(n13423), .A2(n13276), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13169), .ZN(n13171) );
  INV_X1 U15288 ( .A(n13456), .ZN(n13373) );
  NOR2_X1 U15289 ( .A1(n13373), .A2(n13277), .ZN(n13170) );
  AOI211_X1 U15290 ( .C1(n13261), .C2(n13420), .A(n13171), .B(n13170), .ZN(
        n13173) );
  NAND2_X1 U15291 ( .A1(n13674), .A2(n13281), .ZN(n13172) );
  OAI211_X1 U15292 ( .C1(n13174), .C2(n13272), .A(n13173), .B(n13172), .ZN(
        P2_U3192) );
  AOI21_X1 U15293 ( .B1(n13176), .B2(n13175), .A(n13272), .ZN(n13178) );
  NAND2_X1 U15294 ( .A1(n13178), .A2(n13177), .ZN(n13182) );
  NOR2_X1 U15295 ( .A1(n13549), .A2(n13276), .ZN(n13180) );
  OAI22_X1 U15296 ( .A1(n13233), .A2(n13278), .B1(n13364), .B2(n13277), .ZN(
        n13179) );
  AOI211_X1 U15297 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(P2_U3088), .A(n13180), 
        .B(n13179), .ZN(n13181) );
  OAI211_X1 U15298 ( .C1(n13552), .C2(n13258), .A(n13182), .B(n13181), .ZN(
        P2_U3195) );
  INV_X1 U15299 ( .A(n13763), .ZN(n13486) );
  OAI21_X1 U15300 ( .B1(n13213), .B2(n13183), .A(n9485), .ZN(n13186) );
  NAND3_X1 U15301 ( .A1(n13184), .A2(n13270), .A3(n13408), .ZN(n13185) );
  INV_X1 U15302 ( .A(n13187), .ZN(n13483) );
  AOI22_X1 U15303 ( .A1(n13483), .A2(n13240), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13188) );
  OAI21_X1 U15304 ( .B1(n13474), .B2(n13277), .A(n13188), .ZN(n13189) );
  AOI21_X1 U15305 ( .B1(n13261), .B2(n13472), .A(n13189), .ZN(n13190) );
  OAI211_X1 U15306 ( .C1(n13486), .C2(n13258), .A(n13191), .B(n13190), .ZN(
        P2_U3197) );
  OAI21_X1 U15307 ( .B1(n13194), .B2(n13193), .A(n13192), .ZN(n13195) );
  NAND2_X1 U15308 ( .A1(n13195), .A2(n9485), .ZN(n13203) );
  INV_X1 U15309 ( .A(n13618), .ZN(n13201) );
  OR2_X1 U15310 ( .A1(n13393), .A2(n13632), .ZN(n13197) );
  NAND2_X1 U15311 ( .A1(n13350), .A2(n13542), .ZN(n13196) );
  NAND2_X1 U15312 ( .A1(n13197), .A2(n13196), .ZN(n13616) );
  INV_X1 U15313 ( .A(n13616), .ZN(n13736) );
  OAI22_X1 U15314 ( .A1(n13736), .A2(n13199), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13198), .ZN(n13200) );
  AOI21_X1 U15315 ( .B1(n13201), .B2(n13240), .A(n13200), .ZN(n13202) );
  OAI211_X1 U15316 ( .C1(n13390), .C2(n13258), .A(n13203), .B(n13202), .ZN(
        P2_U3198) );
  OAI21_X1 U15317 ( .B1(n13206), .B2(n13205), .A(n13204), .ZN(n13207) );
  NAND2_X1 U15318 ( .A1(n13207), .A2(n9485), .ZN(n13212) );
  OAI22_X1 U15319 ( .A1(n13396), .A2(n13632), .B1(n13633), .B2(n13630), .ZN(
        n13598) );
  INV_X1 U15320 ( .A(n13601), .ZN(n13208) );
  NOR2_X1 U15321 ( .A1(n13276), .A2(n13208), .ZN(n13209) );
  AOI211_X1 U15322 ( .C1(n13598), .C2(n13251), .A(n13210), .B(n13209), .ZN(
        n13211) );
  OAI211_X1 U15323 ( .C1(n13604), .C2(n13258), .A(n13212), .B(n13211), .ZN(
        P2_U3200) );
  NAND2_X1 U15324 ( .A1(n13455), .A2(n13544), .ZN(n13217) );
  NAND2_X1 U15325 ( .A1(n13523), .A2(n13542), .ZN(n13216) );
  NAND2_X1 U15326 ( .A1(n13217), .A2(n13216), .ZN(n13491) );
  INV_X1 U15327 ( .A(n13497), .ZN(n13219) );
  OAI22_X1 U15328 ( .A1(n13219), .A2(n13276), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13218), .ZN(n13220) );
  AOI21_X1 U15329 ( .B1(n13491), .B2(n13251), .A(n13220), .ZN(n13221) );
  INV_X1 U15330 ( .A(n13222), .ZN(n13225) );
  INV_X1 U15331 ( .A(n13223), .ZN(n13224) );
  OAI33_X1 U15332 ( .A1(n13272), .A2(n13225), .A3(n6803), .B1(n13262), .B2(
        n13224), .B3(n13247), .ZN(n13230) );
  AOI22_X1 U15333 ( .A1(n13240), .A2(n13562), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13227) );
  OAI22_X1 U15334 ( .A1(n13403), .A2(n13632), .B1(n13247), .B2(n13630), .ZN(
        n13559) );
  NAND2_X1 U15335 ( .A1(n13559), .A2(n13251), .ZN(n13226) );
  OAI211_X1 U15336 ( .C1(n13564), .C2(n13258), .A(n13227), .B(n13226), .ZN(
        n13228) );
  AOI21_X1 U15337 ( .B1(n13230), .B2(n13229), .A(n13228), .ZN(n13231) );
  OAI21_X1 U15338 ( .B1(n13232), .B2(n13272), .A(n13231), .ZN(P2_U3205) );
  INV_X1 U15339 ( .A(n13233), .ZN(n13545) );
  NAND2_X1 U15340 ( .A1(n13545), .A2(n13270), .ZN(n13237) );
  NAND2_X1 U15341 ( .A1(n13234), .A2(n9485), .ZN(n13236) );
  MUX2_X1 U15342 ( .A(n13237), .B(n13236), .S(n13235), .Z(n13244) );
  NOR2_X1 U15343 ( .A1(n13238), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13239) );
  AOI21_X1 U15344 ( .B1(n13530), .B2(n13240), .A(n13239), .ZN(n13241) );
  OAI21_X1 U15345 ( .B1(n13403), .B2(n13277), .A(n13241), .ZN(n13242) );
  AOI21_X1 U15346 ( .B1(n13523), .B2(n13261), .A(n13242), .ZN(n13243) );
  OAI211_X1 U15347 ( .C1(n13526), .C2(n13258), .A(n13244), .B(n13243), .ZN(
        P2_U3207) );
  XNOR2_X1 U15348 ( .A(n13246), .B(n13245), .ZN(n13253) );
  OAI22_X1 U15349 ( .A1(n13247), .A2(n13632), .B1(n13393), .B2(n13630), .ZN(
        n13587) );
  OAI22_X1 U15350 ( .A1(n13276), .A2(n13589), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13248), .ZN(n13250) );
  NOR2_X1 U15351 ( .A1(n13593), .A2(n13258), .ZN(n13249) );
  AOI211_X1 U15352 ( .C1(n13251), .C2(n13587), .A(n13250), .B(n13249), .ZN(
        n13252) );
  OAI21_X1 U15353 ( .B1(n13253), .B2(n13272), .A(n13252), .ZN(P2_U3210) );
  OAI21_X1 U15354 ( .B1(n13264), .B2(n13255), .A(n13254), .ZN(n13256) );
  INV_X1 U15355 ( .A(n13256), .ZN(n13269) );
  OAI22_X1 U15356 ( .A1(n13459), .A2(n13276), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13257), .ZN(n13260) );
  NOR2_X1 U15357 ( .A1(n13411), .A2(n13258), .ZN(n13259) );
  AOI211_X1 U15358 ( .C1(n13261), .C2(n13456), .A(n13260), .B(n13259), .ZN(
        n13268) );
  NOR3_X1 U15359 ( .A1(n13264), .A2(n13263), .A3(n13262), .ZN(n13266) );
  OAI21_X1 U15360 ( .B1(n13266), .B2(n13265), .A(n13455), .ZN(n13267) );
  OAI211_X1 U15361 ( .C1(n13269), .C2(n13272), .A(n13268), .B(n13267), .ZN(
        P2_U3212) );
  NAND2_X1 U15362 ( .A1(n13270), .A2(n13350), .ZN(n13275) );
  OR2_X1 U15363 ( .A1(n13272), .A2(n13271), .ZN(n13274) );
  MUX2_X1 U15364 ( .A(n13275), .B(n13274), .S(n13273), .Z(n13283) );
  OAI22_X1 U15365 ( .A1(n13276), .A2(n13637), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9270), .ZN(n13280) );
  OAI22_X1 U15366 ( .A1(n13278), .A2(n13633), .B1(n13631), .B2(n13277), .ZN(
        n13279) );
  AOI211_X1 U15367 ( .C1(n13644), .C2(n13281), .A(n13280), .B(n13279), .ZN(
        n13282) );
  NAND2_X1 U15368 ( .A1(n13283), .A2(n13282), .ZN(P2_U3213) );
  MUX2_X1 U15369 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13340), .S(n6457), .Z(
        P2_U3562) );
  MUX2_X1 U15370 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13377), .S(n6457), .Z(
        P2_U3561) );
  MUX2_X1 U15371 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13420), .S(n6457), .Z(
        P2_U3560) );
  MUX2_X1 U15372 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13379), .S(n6457), .Z(
        P2_U3559) );
  MUX2_X1 U15373 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13456), .S(n6457), .Z(
        P2_U3558) );
  MUX2_X1 U15374 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13472), .S(n6457), .Z(
        P2_U3557) );
  MUX2_X1 U15375 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13455), .S(n6457), .Z(
        P2_U3556) );
  MUX2_X1 U15376 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13408), .S(n6457), .Z(
        P2_U3555) );
  MUX2_X1 U15377 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13523), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15378 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13545), .S(n6457), .Z(
        P2_U3553) );
  MUX2_X1 U15379 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13524), .S(n6457), .Z(
        P2_U3552) );
  MUX2_X1 U15380 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13543), .S(n6457), .Z(
        P2_U3551) );
  MUX2_X1 U15381 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13362), .S(n6457), .Z(
        P2_U3550) );
  MUX2_X1 U15382 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13359), .S(n6457), .Z(
        P2_U3549) );
  MUX2_X1 U15383 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13355), .S(n6457), .Z(
        P2_U3548) );
  MUX2_X1 U15384 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13353), .S(n6457), .Z(
        P2_U3547) );
  MUX2_X1 U15385 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13350), .S(n6457), .Z(
        P2_U3546) );
  MUX2_X1 U15386 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13388), .S(n6457), .Z(
        P2_U3545) );
  MUX2_X1 U15387 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13284), .S(n6457), .Z(
        P2_U3544) );
  MUX2_X1 U15388 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13285), .S(n6457), .Z(
        P2_U3543) );
  MUX2_X1 U15389 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13286), .S(n6457), .Z(
        P2_U3542) );
  MUX2_X1 U15390 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13287), .S(n6457), .Z(
        P2_U3541) );
  MUX2_X1 U15391 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13288), .S(n6457), .Z(
        P2_U3540) );
  MUX2_X1 U15392 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13289), .S(n6457), .Z(
        P2_U3539) );
  MUX2_X1 U15393 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13290), .S(n6457), .Z(
        P2_U3538) );
  MUX2_X1 U15394 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13291), .S(n6457), .Z(
        P2_U3537) );
  MUX2_X1 U15395 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13292), .S(n6457), .Z(
        P2_U3536) );
  MUX2_X1 U15396 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13293), .S(n6457), .Z(
        P2_U3535) );
  MUX2_X1 U15397 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13294), .S(n6457), .Z(
        P2_U3534) );
  MUX2_X1 U15398 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13295), .S(n6457), .Z(
        P2_U3533) );
  MUX2_X1 U15399 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6734), .S(n6457), .Z(
        P2_U3532) );
  MUX2_X1 U15400 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n12064), .S(n6457), .Z(
        P2_U3531) );
  INV_X1 U15401 ( .A(n13297), .ZN(n13300) );
  NOR2_X1 U15402 ( .A1(n14820), .A2(n13298), .ZN(n13299) );
  AOI211_X1 U15403 ( .C1(n14859), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n13300), .B(
        n13299), .ZN(n13311) );
  OAI211_X1 U15404 ( .C1(n13303), .C2(n13302), .A(n13301), .B(n14865), .ZN(
        n13310) );
  OR3_X1 U15405 ( .A1(n13306), .A2(n13305), .A3(n13304), .ZN(n13307) );
  NAND3_X1 U15406 ( .A1(n13308), .A2(n14868), .A3(n13307), .ZN(n13309) );
  NAND3_X1 U15407 ( .A1(n13311), .A2(n13310), .A3(n13309), .ZN(P2_U3220) );
  XNOR2_X1 U15408 ( .A(n14864), .B(n13314), .ZN(n14862) );
  NAND2_X1 U15409 ( .A1(n13314), .A2(n13321), .ZN(n13315) );
  NAND2_X1 U15410 ( .A1(n14860), .A2(n13315), .ZN(n13316) );
  XNOR2_X1 U15411 ( .A(n13316), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13326) );
  INV_X1 U15412 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13317) );
  OAI22_X1 U15413 ( .A1(n13320), .A2(n13319), .B1(n13318), .B2(n13317), .ZN(
        n13322) );
  XNOR2_X1 U15414 ( .A(n13322), .B(n13321), .ZN(n14869) );
  NAND2_X1 U15415 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14869), .ZN(n14867) );
  NAND2_X1 U15416 ( .A1(n14864), .A2(n13322), .ZN(n13323) );
  NAND2_X1 U15417 ( .A1(n14867), .A2(n13323), .ZN(n13325) );
  XNOR2_X1 U15418 ( .A(n13325), .B(n13324), .ZN(n13329) );
  AOI22_X1 U15419 ( .A1(n13326), .A2(n14865), .B1(n14868), .B2(n13329), .ZN(
        n13332) );
  INV_X1 U15420 ( .A(n13326), .ZN(n13327) );
  MUX2_X1 U15421 ( .A(n13332), .B(n13331), .S(n13330), .Z(n13334) );
  OAI211_X1 U15422 ( .C1(n7495), .C2(n14857), .A(n13334), .B(n13333), .ZN(
        P2_U3233) );
  NAND2_X1 U15423 ( .A1(n13411), .A2(n13482), .ZN(n13462) );
  NAND2_X1 U15424 ( .A1(n13755), .A2(n13382), .ZN(n13343) );
  XNOR2_X1 U15425 ( .A(n13343), .B(n13751), .ZN(n13337) );
  NAND2_X1 U15426 ( .A1(n13337), .A2(n13639), .ZN(n13664) );
  INV_X1 U15427 ( .A(P2_B_REG_SCAN_IN), .ZN(n13338) );
  NOR2_X1 U15428 ( .A1(n13795), .A2(n13338), .ZN(n13339) );
  NOR2_X1 U15429 ( .A1(n13632), .A2(n13339), .ZN(n13378) );
  NAND2_X1 U15430 ( .A1(n13340), .A2(n13378), .ZN(n13666) );
  NOR2_X1 U15431 ( .A1(n13649), .A2(n13666), .ZN(n13345) );
  NOR2_X1 U15432 ( .A1(n13751), .A2(n13603), .ZN(n13341) );
  AOI211_X1 U15433 ( .C1(n13649), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13345), 
        .B(n13341), .ZN(n13342) );
  OAI21_X1 U15434 ( .B1(n13664), .B2(n13641), .A(n13342), .ZN(P2_U3234) );
  OAI211_X1 U15435 ( .C1(n13755), .C2(n13382), .A(n13639), .B(n13343), .ZN(
        n13667) );
  NOR2_X1 U15436 ( .A1(n13755), .A2(n13603), .ZN(n13344) );
  AOI211_X1 U15437 ( .C1(n13649), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13345), 
        .B(n13344), .ZN(n13346) );
  OAI21_X1 U15438 ( .B1(n13641), .B2(n13667), .A(n13346), .ZN(P2_U3235) );
  OR2_X1 U15439 ( .A1(n13781), .A2(n13350), .ZN(n13351) );
  NAND2_X1 U15440 ( .A1(n13390), .A2(n13353), .ZN(n13352) );
  OR2_X1 U15441 ( .A1(n13390), .A2(n13353), .ZN(n13354) );
  NAND2_X1 U15442 ( .A1(n13597), .A2(n13606), .ZN(n13357) );
  OR2_X1 U15443 ( .A1(n13604), .A2(n13355), .ZN(n13356) );
  NOR2_X1 U15444 ( .A1(n13593), .A2(n13359), .ZN(n13358) );
  NAND2_X1 U15445 ( .A1(n13593), .A2(n13359), .ZN(n13360) );
  AND2_X1 U15446 ( .A1(n13578), .A2(n13362), .ZN(n13361) );
  OR2_X1 U15447 ( .A1(n13578), .A2(n13362), .ZN(n13363) );
  AND2_X1 U15448 ( .A1(n13715), .A2(n13364), .ZN(n13365) );
  NAND2_X1 U15449 ( .A1(n13710), .A2(n13403), .ZN(n13367) );
  AND2_X1 U15450 ( .A1(n13552), .A2(n13524), .ZN(n13366) );
  NAND2_X1 U15451 ( .A1(n13526), .A2(n13545), .ZN(n13368) );
  NAND2_X1 U15452 ( .A1(n13692), .A2(n13474), .ZN(n13370) );
  NAND2_X1 U15453 ( .A1(n13489), .A2(n13370), .ZN(n13468) );
  INV_X1 U15454 ( .A(n13478), .ZN(n13469) );
  NAND2_X1 U15455 ( .A1(n13468), .A2(n13469), .ZN(n13471) );
  NAND2_X1 U15456 ( .A1(n13454), .A2(n13453), .ZN(n13452) );
  NAND2_X1 U15457 ( .A1(n13446), .A2(n13373), .ZN(n13418) );
  NAND2_X1 U15458 ( .A1(n13419), .A2(n13374), .ZN(n13376) );
  INV_X1 U15459 ( .A(n13335), .ZN(n13385) );
  AOI22_X1 U15460 ( .A1(n13383), .A2(n15200), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13649), .ZN(n13384) );
  OAI21_X1 U15461 ( .B1(n13385), .B2(n13603), .A(n13384), .ZN(n13415) );
  INV_X1 U15462 ( .A(n13447), .ZN(n13413) );
  NOR2_X1 U15463 ( .A1(n14620), .A2(n13388), .ZN(n13386) );
  NAND2_X1 U15464 ( .A1(n13611), .A2(n13612), .ZN(n13610) );
  OR2_X1 U15465 ( .A1(n13390), .A2(n13633), .ZN(n13391) );
  NOR2_X1 U15466 ( .A1(n13604), .A2(n13393), .ZN(n13392) );
  NAND2_X1 U15467 ( .A1(n13604), .A2(n13393), .ZN(n13394) );
  INV_X1 U15468 ( .A(n13585), .ZN(n13395) );
  NAND2_X1 U15469 ( .A1(n13580), .A2(n13397), .ZN(n13399) );
  NAND2_X1 U15470 ( .A1(n13399), .A2(n13398), .ZN(n13566) );
  NAND2_X1 U15471 ( .A1(n13715), .A2(n13543), .ZN(n13400) );
  NAND2_X1 U15472 ( .A1(n13566), .A2(n13400), .ZN(n13402) );
  OR2_X1 U15473 ( .A1(n13715), .A2(n13543), .ZN(n13401) );
  INV_X1 U15474 ( .A(n13553), .ZN(n13540) );
  AND2_X1 U15475 ( .A1(n13552), .A2(n13403), .ZN(n13404) );
  NAND2_X1 U15476 ( .A1(n13702), .A2(n13545), .ZN(n13405) );
  NAND2_X1 U15477 ( .A1(n13512), .A2(n13406), .ZN(n13407) );
  NAND2_X1 U15478 ( .A1(n13692), .A2(n13408), .ZN(n13409) );
  OR2_X1 U15479 ( .A1(n13763), .A2(n13455), .ZN(n13410) );
  NOR2_X1 U15480 ( .A1(n13681), .A2(n13472), .ZN(n13412) );
  XNOR2_X1 U15481 ( .A(n13416), .B(n13417), .ZN(n13675) );
  NAND2_X1 U15482 ( .A1(n13419), .A2(n13635), .ZN(n13422) );
  AOI22_X1 U15483 ( .A1(n13456), .A2(n13542), .B1(n13544), .B2(n13420), .ZN(
        n13421) );
  NOR2_X1 U15484 ( .A1(n13423), .A2(n13651), .ZN(n13424) );
  OAI21_X1 U15485 ( .B1(n13672), .B2(n13424), .A(n15210), .ZN(n13431) );
  OR2_X1 U15486 ( .A1(n13428), .A2(n13443), .ZN(n13425) );
  AND3_X1 U15487 ( .A1(n13426), .A2(n13639), .A3(n13425), .ZN(n13673) );
  OAI22_X1 U15488 ( .A1(n13428), .A2(n13603), .B1(n15210), .B2(n13427), .ZN(
        n13429) );
  AOI21_X1 U15489 ( .B1(n13673), .B2(n13658), .A(n13429), .ZN(n13430) );
  OAI211_X1 U15490 ( .C1(n13627), .C2(n13675), .A(n13431), .B(n13430), .ZN(
        P2_U3237) );
  OR2_X1 U15491 ( .A1(n13433), .A2(n13447), .ZN(n13434) );
  NAND2_X1 U15492 ( .A1(n13432), .A2(n13434), .ZN(n13438) );
  OAI22_X1 U15493 ( .A1(n13436), .A2(n13632), .B1(n13435), .B2(n13630), .ZN(
        n13437) );
  OAI22_X1 U15494 ( .A1(n13440), .A2(n13651), .B1(n13439), .B2(n15210), .ZN(
        n13445) );
  NAND2_X1 U15495 ( .A1(n13446), .A2(n13462), .ZN(n13441) );
  NAND2_X1 U15496 ( .A1(n13441), .A2(n13639), .ZN(n13442) );
  OR2_X1 U15497 ( .A1(n13443), .A2(n13442), .ZN(n13677) );
  NOR2_X1 U15498 ( .A1(n13677), .A2(n13641), .ZN(n13444) );
  AOI211_X1 U15499 ( .C1(n13654), .C2(n13446), .A(n13445), .B(n13444), .ZN(
        n13450) );
  XNOR2_X1 U15500 ( .A(n13448), .B(n13447), .ZN(n13676) );
  NAND2_X1 U15501 ( .A1(n13676), .A2(n13656), .ZN(n13449) );
  OAI211_X1 U15502 ( .C1(n13679), .C2(n13649), .A(n13450), .B(n13449), .ZN(
        P2_U3238) );
  XNOR2_X1 U15503 ( .A(n13454), .B(n13451), .ZN(n13684) );
  OAI21_X1 U15504 ( .B1(n13454), .B2(n13453), .A(n13452), .ZN(n13457) );
  AOI222_X1 U15505 ( .A1(n13635), .A2(n13457), .B1(n13456), .B2(n13544), .C1(
        n13455), .C2(n13542), .ZN(n13683) );
  OAI22_X1 U15506 ( .A1(n13459), .A2(n13651), .B1(n13458), .B2(n15210), .ZN(
        n13460) );
  AOI21_X1 U15507 ( .B1(n13681), .B2(n13654), .A(n13460), .ZN(n13465) );
  INV_X1 U15508 ( .A(n13482), .ZN(n13461) );
  AOI21_X1 U15509 ( .B1(n13461), .B2(n13681), .A(n13620), .ZN(n13463) );
  AND2_X1 U15510 ( .A1(n13463), .A2(n13462), .ZN(n13680) );
  NAND2_X1 U15511 ( .A1(n13680), .A2(n13658), .ZN(n13464) );
  OAI211_X1 U15512 ( .C1(n13683), .C2(n13649), .A(n13465), .B(n13464), .ZN(
        n13466) );
  INV_X1 U15513 ( .A(n13466), .ZN(n13467) );
  OAI21_X1 U15514 ( .B1(n13684), .B2(n13627), .A(n13467), .ZN(P2_U3239) );
  OR2_X1 U15515 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  NAND2_X1 U15516 ( .A1(n13471), .A2(n13470), .ZN(n13476) );
  NAND2_X1 U15517 ( .A1(n13472), .A2(n13544), .ZN(n13473) );
  OAI21_X1 U15518 ( .B1(n13474), .B2(n13630), .A(n13473), .ZN(n13475) );
  AOI21_X1 U15519 ( .B1(n13476), .B2(n13635), .A(n13475), .ZN(n13687) );
  OAI21_X1 U15520 ( .B1(n13479), .B2(n13478), .A(n13477), .ZN(n13686) );
  NAND2_X1 U15521 ( .A1(n13763), .A2(n13496), .ZN(n13480) );
  NAND2_X1 U15522 ( .A1(n13480), .A2(n13639), .ZN(n13481) );
  NOR2_X1 U15523 ( .A1(n13482), .A2(n13481), .ZN(n13685) );
  NAND2_X1 U15524 ( .A1(n13685), .A2(n13658), .ZN(n13485) );
  AOI22_X1 U15525 ( .A1(n13483), .A2(n15200), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13649), .ZN(n13484) );
  OAI211_X1 U15526 ( .C1(n13486), .C2(n13603), .A(n13485), .B(n13484), .ZN(
        n13487) );
  AOI21_X1 U15527 ( .B1(n13656), .B2(n13686), .A(n13487), .ZN(n13488) );
  OAI21_X1 U15528 ( .B1(n13649), .B2(n13687), .A(n13488), .ZN(P2_U3240) );
  OAI21_X1 U15529 ( .B1(n13490), .B2(n13493), .A(n13489), .ZN(n13492) );
  AOI21_X1 U15530 ( .B1(n13492), .B2(n13635), .A(n13491), .ZN(n13694) );
  OAI21_X1 U15531 ( .B1(n6631), .B2(n6445), .A(n13494), .ZN(n13695) );
  INV_X1 U15532 ( .A(n13695), .ZN(n13502) );
  AOI21_X1 U15533 ( .B1(n13692), .B2(n13508), .A(n13620), .ZN(n13495) );
  AND2_X1 U15534 ( .A1(n13496), .A2(n13495), .ZN(n13691) );
  NAND2_X1 U15535 ( .A1(n13691), .A2(n13658), .ZN(n13499) );
  AOI22_X1 U15536 ( .A1(n13497), .A2(n15200), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13649), .ZN(n13498) );
  OAI211_X1 U15537 ( .C1(n13500), .C2(n13603), .A(n13499), .B(n13498), .ZN(
        n13501) );
  AOI21_X1 U15538 ( .B1(n13502), .B2(n13656), .A(n13501), .ZN(n13503) );
  OAI21_X1 U15539 ( .B1(n13649), .B2(n13694), .A(n13503), .ZN(P2_U3241) );
  INV_X1 U15540 ( .A(n13504), .ZN(n13505) );
  AOI21_X1 U15541 ( .B1(n13516), .B2(n13506), .A(n13505), .ZN(n13701) );
  INV_X1 U15542 ( .A(n13507), .ZN(n13529) );
  INV_X1 U15543 ( .A(n13508), .ZN(n13509) );
  AOI211_X1 U15544 ( .C1(n13698), .C2(n13529), .A(n13620), .B(n13509), .ZN(
        n13696) );
  AOI22_X1 U15545 ( .A1(n13510), .A2(n15200), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n13649), .ZN(n13511) );
  OAI21_X1 U15546 ( .B1(n13512), .B2(n13603), .A(n13511), .ZN(n13513) );
  AOI21_X1 U15547 ( .B1(n13696), .B2(n13658), .A(n13513), .ZN(n13521) );
  OAI21_X1 U15548 ( .B1(n13516), .B2(n13515), .A(n13514), .ZN(n13517) );
  NAND2_X1 U15549 ( .A1(n13517), .A2(n13635), .ZN(n13699) );
  INV_X1 U15550 ( .A(n13699), .ZN(n13519) );
  INV_X1 U15551 ( .A(n13518), .ZN(n13697) );
  OAI21_X1 U15552 ( .B1(n13519), .B2(n13697), .A(n15210), .ZN(n13520) );
  OAI211_X1 U15553 ( .C1(n13701), .C2(n13627), .A(n13521), .B(n13520), .ZN(
        P2_U3242) );
  XOR2_X1 U15554 ( .A(n13522), .B(n13535), .Z(n13525) );
  AOI222_X1 U15555 ( .A1(n13635), .A2(n13525), .B1(n13524), .B2(n13542), .C1(
        n13523), .C2(n13544), .ZN(n13708) );
  OAI21_X1 U15556 ( .B1(n13526), .B2(n13547), .A(n13639), .ZN(n13527) );
  INV_X1 U15557 ( .A(n13527), .ZN(n13528) );
  NAND2_X1 U15558 ( .A1(n13529), .A2(n13528), .ZN(n13705) );
  NAND2_X1 U15559 ( .A1(n13530), .A2(n15200), .ZN(n13531) );
  OAI21_X1 U15560 ( .B1(n15210), .B2(n13532), .A(n13531), .ZN(n13533) );
  AOI21_X1 U15561 ( .B1(n13702), .B2(n13654), .A(n13533), .ZN(n13537) );
  OR2_X1 U15562 ( .A1(n13535), .A2(n13534), .ZN(n13704) );
  NAND3_X1 U15563 ( .A1(n13704), .A2(n13656), .A3(n6755), .ZN(n13536) );
  OAI211_X1 U15564 ( .C1(n13705), .C2(n13641), .A(n13537), .B(n13536), .ZN(
        n13538) );
  INV_X1 U15565 ( .A(n13538), .ZN(n13539) );
  OAI21_X1 U15566 ( .B1(n13708), .B2(n13649), .A(n13539), .ZN(P2_U3243) );
  XNOR2_X1 U15567 ( .A(n6614), .B(n13540), .ZN(n13546) );
  AOI222_X1 U15568 ( .A1(n13635), .A2(n13546), .B1(n13545), .B2(n13544), .C1(
        n13543), .C2(n13542), .ZN(n13712) );
  INV_X1 U15569 ( .A(n13561), .ZN(n13548) );
  AOI211_X1 U15570 ( .C1(n13710), .C2(n13548), .A(n13620), .B(n13547), .ZN(
        n13709) );
  INV_X1 U15571 ( .A(n13549), .ZN(n13550) );
  AOI22_X1 U15572 ( .A1(n13550), .A2(n15200), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n13649), .ZN(n13551) );
  OAI21_X1 U15573 ( .B1(n13552), .B2(n13603), .A(n13551), .ZN(n13556) );
  XNOR2_X1 U15574 ( .A(n13554), .B(n13553), .ZN(n13713) );
  NOR2_X1 U15575 ( .A1(n13713), .A2(n13627), .ZN(n13555) );
  AOI211_X1 U15576 ( .C1(n13709), .C2(n13658), .A(n13556), .B(n13555), .ZN(
        n13557) );
  OAI21_X1 U15577 ( .B1(n13712), .B2(n13649), .A(n13557), .ZN(P2_U3244) );
  XNOR2_X1 U15578 ( .A(n13558), .B(n13565), .ZN(n13560) );
  AOI21_X1 U15579 ( .B1(n13560), .B2(n13635), .A(n13559), .ZN(n13717) );
  AOI211_X1 U15580 ( .C1(n13715), .C2(n13573), .A(n13620), .B(n13561), .ZN(
        n13714) );
  AOI22_X1 U15581 ( .A1(n13562), .A2(n15200), .B1(n13649), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n13563) );
  OAI21_X1 U15582 ( .B1(n13564), .B2(n13603), .A(n13563), .ZN(n13568) );
  XNOR2_X1 U15583 ( .A(n13566), .B(n13565), .ZN(n13718) );
  NOR2_X1 U15584 ( .A1(n13718), .A2(n13627), .ZN(n13567) );
  AOI211_X1 U15585 ( .C1(n13714), .C2(n13658), .A(n13568), .B(n13567), .ZN(
        n13569) );
  OAI21_X1 U15586 ( .B1(n13649), .B2(n13717), .A(n13569), .ZN(P2_U3245) );
  XOR2_X1 U15587 ( .A(n13570), .B(n13579), .Z(n13572) );
  AOI21_X1 U15588 ( .B1(n13572), .B2(n13635), .A(n13571), .ZN(n13722) );
  INV_X1 U15589 ( .A(n13591), .ZN(n13575) );
  INV_X1 U15590 ( .A(n13573), .ZN(n13574) );
  AOI211_X1 U15591 ( .C1(n13720), .C2(n13575), .A(n13620), .B(n13574), .ZN(
        n13719) );
  AOI22_X1 U15592 ( .A1(n13649), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13576), 
        .B2(n15200), .ZN(n13577) );
  OAI21_X1 U15593 ( .B1(n13578), .B2(n13603), .A(n13577), .ZN(n13582) );
  XNOR2_X1 U15594 ( .A(n13580), .B(n13579), .ZN(n13723) );
  NOR2_X1 U15595 ( .A1(n13723), .A2(n13627), .ZN(n13581) );
  AOI211_X1 U15596 ( .C1(n13719), .C2(n13658), .A(n13582), .B(n13581), .ZN(
        n13583) );
  OAI21_X1 U15597 ( .B1(n13649), .B2(n13722), .A(n13583), .ZN(P2_U3246) );
  XNOR2_X1 U15598 ( .A(n13584), .B(n13585), .ZN(n13728) );
  XNOR2_X1 U15599 ( .A(n13586), .B(n13585), .ZN(n13588) );
  AOI21_X1 U15600 ( .B1(n13588), .B2(n13635), .A(n13587), .ZN(n13727) );
  OAI21_X1 U15601 ( .B1(n13589), .B2(n13651), .A(n13727), .ZN(n13590) );
  NAND2_X1 U15602 ( .A1(n13590), .A2(n15210), .ZN(n13596) );
  INV_X1 U15603 ( .A(n13600), .ZN(n13592) );
  AOI211_X1 U15604 ( .C1(n13725), .C2(n13592), .A(n13620), .B(n13591), .ZN(
        n13724) );
  OAI22_X1 U15605 ( .A1(n13593), .A2(n13603), .B1(n15210), .B2(n14861), .ZN(
        n13594) );
  AOI21_X1 U15606 ( .B1(n13724), .B2(n13658), .A(n13594), .ZN(n13595) );
  OAI211_X1 U15607 ( .C1(n13728), .C2(n13627), .A(n13596), .B(n13595), .ZN(
        P2_U3247) );
  XNOR2_X1 U15608 ( .A(n13597), .B(n13606), .ZN(n13599) );
  AOI21_X1 U15609 ( .B1(n13599), .B2(n13635), .A(n13598), .ZN(n13732) );
  AOI211_X1 U15610 ( .C1(n13730), .C2(n13621), .A(n13620), .B(n13600), .ZN(
        n13729) );
  AOI22_X1 U15611 ( .A1(n13649), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13601), 
        .B2(n15200), .ZN(n13602) );
  OAI21_X1 U15612 ( .B1(n13604), .B2(n13603), .A(n13602), .ZN(n13608) );
  XOR2_X1 U15613 ( .A(n13605), .B(n13606), .Z(n13733) );
  NOR2_X1 U15614 ( .A1(n13733), .A2(n13627), .ZN(n13607) );
  AOI211_X1 U15615 ( .C1(n13729), .C2(n13658), .A(n13608), .B(n13607), .ZN(
        n13609) );
  OAI21_X1 U15616 ( .B1(n13649), .B2(n13732), .A(n13609), .ZN(P2_U3248) );
  OAI21_X1 U15617 ( .B1(n13611), .B2(n13612), .A(n13610), .ZN(n13735) );
  INV_X1 U15618 ( .A(n13612), .ZN(n13613) );
  XNOR2_X1 U15619 ( .A(n13614), .B(n13613), .ZN(n13615) );
  NAND2_X1 U15620 ( .A1(n13615), .A2(n13635), .ZN(n13738) );
  INV_X1 U15621 ( .A(n13738), .ZN(n13617) );
  OAI21_X1 U15622 ( .B1(n13617), .B2(n13616), .A(n15210), .ZN(n13626) );
  INV_X1 U15623 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13619) );
  OAI22_X1 U15624 ( .A1(n15210), .A2(n13619), .B1(n13618), .B2(n13651), .ZN(
        n13624) );
  AOI21_X1 U15625 ( .B1(n13638), .B2(n13775), .A(n13620), .ZN(n13622) );
  NAND2_X1 U15626 ( .A1(n13622), .A2(n13621), .ZN(n13737) );
  NOR2_X1 U15627 ( .A1(n13737), .A2(n13641), .ZN(n13623) );
  AOI211_X1 U15628 ( .C1(n13654), .C2(n13775), .A(n13624), .B(n13623), .ZN(
        n13625) );
  OAI211_X1 U15629 ( .C1(n13735), .C2(n13627), .A(n13626), .B(n13625), .ZN(
        P2_U3249) );
  OAI21_X1 U15630 ( .B1(n13629), .B2(n13645), .A(n13628), .ZN(n13636) );
  OAI22_X1 U15631 ( .A1(n13633), .A2(n13632), .B1(n13631), .B2(n13630), .ZN(
        n13634) );
  AOI21_X1 U15632 ( .B1(n13636), .B2(n13635), .A(n13634), .ZN(n13747) );
  OAI22_X1 U15633 ( .A1(n15210), .A2(n11529), .B1(n13637), .B2(n13651), .ZN(
        n13643) );
  OAI211_X1 U15634 ( .C1(n13781), .C2(n13640), .A(n13639), .B(n13638), .ZN(
        n13745) );
  NOR2_X1 U15635 ( .A1(n13745), .A2(n13641), .ZN(n13642) );
  AOI211_X1 U15636 ( .C1(n13654), .C2(n13644), .A(n13643), .B(n13642), .ZN(
        n13648) );
  XNOR2_X1 U15637 ( .A(n13646), .B(n13645), .ZN(n13744) );
  NAND2_X1 U15638 ( .A1(n13744), .A2(n13656), .ZN(n13647) );
  OAI211_X1 U15639 ( .C1(n13747), .C2(n13649), .A(n13648), .B(n13647), .ZN(
        P2_U3250) );
  NAND2_X1 U15640 ( .A1(n13650), .A2(n15210), .ZN(n13663) );
  OAI22_X1 U15641 ( .A1(n15210), .A2(n10061), .B1(n13652), .B2(n13651), .ZN(
        n13653) );
  AOI21_X1 U15642 ( .B1(n13655), .B2(n13654), .A(n13653), .ZN(n13662) );
  NAND2_X1 U15643 ( .A1(n13657), .A2(n13656), .ZN(n13661) );
  NAND2_X1 U15644 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  NAND4_X1 U15645 ( .A1(n13663), .A2(n13662), .A3(n13661), .A4(n13660), .ZN(
        P2_U3255) );
  OAI21_X1 U15646 ( .B1(n13751), .B2(n13749), .A(n13665), .ZN(P2_U3530) );
  AND2_X1 U15647 ( .A1(n13667), .A2(n13666), .ZN(n13752) );
  MUX2_X1 U15648 ( .A(n13668), .B(n13752), .S(n14922), .Z(n13669) );
  OAI21_X1 U15649 ( .B1(n13755), .B2(n13749), .A(n13669), .ZN(P2_U3529) );
  MUX2_X1 U15650 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13757), .S(n14922), .Z(
        P2_U3527) );
  NAND2_X1 U15651 ( .A1(n13676), .A2(n14623), .ZN(n13678) );
  NAND3_X1 U15652 ( .A1(n13679), .A2(n13678), .A3(n13677), .ZN(n13758) );
  AOI21_X1 U15653 ( .B1(n14889), .B2(n13681), .A(n13680), .ZN(n13682) );
  OAI211_X1 U15654 ( .C1(n13734), .C2(n13684), .A(n13683), .B(n13682), .ZN(
        n13760) );
  MUX2_X1 U15655 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13760), .S(n14922), .Z(
        P2_U3525) );
  AOI21_X1 U15656 ( .B1(n13686), .B2(n14623), .A(n13685), .ZN(n13688) );
  NAND2_X1 U15657 ( .A1(n13688), .A2(n13687), .ZN(n13761) );
  MUX2_X1 U15658 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13761), .S(n14922), .Z(
        n13689) );
  AOI21_X1 U15659 ( .B1(n13742), .B2(n13763), .A(n13689), .ZN(n13690) );
  INV_X1 U15660 ( .A(n13690), .ZN(P2_U3524) );
  AOI21_X1 U15661 ( .B1(n14889), .B2(n13692), .A(n13691), .ZN(n13693) );
  OAI211_X1 U15662 ( .C1(n13695), .C2(n13734), .A(n13694), .B(n13693), .ZN(
        n13765) );
  MUX2_X1 U15663 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13765), .S(n14922), .Z(
        P2_U3523) );
  AOI211_X1 U15664 ( .C1(n14889), .C2(n13698), .A(n13697), .B(n13696), .ZN(
        n13700) );
  OAI211_X1 U15665 ( .C1(n13734), .C2(n13701), .A(n13700), .B(n13699), .ZN(
        n13766) );
  MUX2_X1 U15666 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13766), .S(n14922), .Z(
        P2_U3522) );
  NAND2_X1 U15667 ( .A1(n13702), .A2(n14889), .ZN(n13707) );
  NAND3_X1 U15668 ( .A1(n13704), .A2(n14623), .A3(n6755), .ZN(n13706) );
  NAND4_X1 U15669 ( .A1(n13708), .A2(n13707), .A3(n13706), .A4(n13705), .ZN(
        n13767) );
  MUX2_X1 U15670 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13767), .S(n14922), .Z(
        P2_U3521) );
  AOI21_X1 U15671 ( .B1(n14889), .B2(n13710), .A(n13709), .ZN(n13711) );
  OAI211_X1 U15672 ( .C1(n13734), .C2(n13713), .A(n13712), .B(n13711), .ZN(
        n13768) );
  MUX2_X1 U15673 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13768), .S(n14922), .Z(
        P2_U3520) );
  AOI21_X1 U15674 ( .B1(n14889), .B2(n13715), .A(n13714), .ZN(n13716) );
  OAI211_X1 U15675 ( .C1(n13734), .C2(n13718), .A(n13717), .B(n13716), .ZN(
        n13769) );
  MUX2_X1 U15676 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13769), .S(n14922), .Z(
        P2_U3519) );
  AOI21_X1 U15677 ( .B1(n14889), .B2(n13720), .A(n13719), .ZN(n13721) );
  OAI211_X1 U15678 ( .C1(n13734), .C2(n13723), .A(n13722), .B(n13721), .ZN(
        n13770) );
  MUX2_X1 U15679 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13770), .S(n14922), .Z(
        P2_U3518) );
  AOI21_X1 U15680 ( .B1(n14889), .B2(n13725), .A(n13724), .ZN(n13726) );
  OAI211_X1 U15681 ( .C1(n13728), .C2(n13734), .A(n13727), .B(n13726), .ZN(
        n13771) );
  MUX2_X1 U15682 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13771), .S(n14922), .Z(
        P2_U3517) );
  AOI21_X1 U15683 ( .B1(n14889), .B2(n13730), .A(n13729), .ZN(n13731) );
  OAI211_X1 U15684 ( .C1(n13733), .C2(n13734), .A(n13732), .B(n13731), .ZN(
        n13772) );
  MUX2_X1 U15685 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13772), .S(n14922), .Z(
        P2_U3516) );
  OR2_X1 U15686 ( .A1(n13735), .A2(n13734), .ZN(n13740) );
  AND2_X1 U15687 ( .A1(n13737), .A2(n13736), .ZN(n13739) );
  NAND3_X1 U15688 ( .A1(n13740), .A2(n13739), .A3(n13738), .ZN(n13773) );
  MUX2_X1 U15689 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13773), .S(n14922), .Z(
        n13741) );
  AOI21_X1 U15690 ( .B1(n13742), .B2(n13775), .A(n13741), .ZN(n13743) );
  INV_X1 U15691 ( .A(n13743), .ZN(P2_U3515) );
  NAND2_X1 U15692 ( .A1(n13744), .A2(n14623), .ZN(n13746) );
  AND3_X1 U15693 ( .A1(n13747), .A2(n13746), .A3(n13745), .ZN(n13777) );
  MUX2_X1 U15694 ( .A(n11600), .B(n13777), .S(n14922), .Z(n13748) );
  OAI21_X1 U15695 ( .B1(n13781), .B2(n13749), .A(n13748), .ZN(P2_U3514) );
  OAI21_X1 U15696 ( .B1(n13751), .B2(n13780), .A(n13750), .ZN(P2_U3498) );
  MUX2_X1 U15697 ( .A(n13753), .B(n13752), .S(n14915), .Z(n13754) );
  OAI21_X1 U15698 ( .B1(n13755), .B2(n13780), .A(n13754), .ZN(P2_U3497) );
  MUX2_X1 U15699 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13757), .S(n14915), .Z(
        P2_U3495) );
  MUX2_X1 U15700 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13760), .S(n14915), .Z(
        P2_U3493) );
  MUX2_X1 U15701 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13761), .S(n14915), .Z(
        n13762) );
  AOI21_X1 U15702 ( .B1(n6641), .B2(n13763), .A(n13762), .ZN(n13764) );
  INV_X1 U15703 ( .A(n13764), .ZN(P2_U3492) );
  MUX2_X1 U15704 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13765), .S(n14915), .Z(
        P2_U3491) );
  MUX2_X1 U15705 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13766), .S(n14915), .Z(
        P2_U3490) );
  MUX2_X1 U15706 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13767), .S(n14915), .Z(
        P2_U3489) );
  MUX2_X1 U15707 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13768), .S(n14915), .Z(
        P2_U3488) );
  MUX2_X1 U15708 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13769), .S(n14915), .Z(
        P2_U3487) );
  MUX2_X1 U15709 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13770), .S(n14915), .Z(
        P2_U3486) );
  MUX2_X1 U15710 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13771), .S(n14915), .Z(
        P2_U3484) );
  MUX2_X1 U15711 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13772), .S(n14915), .Z(
        P2_U3481) );
  MUX2_X1 U15712 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13773), .S(n14915), .Z(
        n13774) );
  AOI21_X1 U15713 ( .B1(n6641), .B2(n13775), .A(n13774), .ZN(n13776) );
  INV_X1 U15714 ( .A(n13776), .ZN(P2_U3478) );
  INV_X1 U15715 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13778) );
  MUX2_X1 U15716 ( .A(n13778), .B(n13777), .S(n14915), .Z(n13779) );
  OAI21_X1 U15717 ( .B1(n13781), .B2(n13780), .A(n13779), .ZN(P2_U3475) );
  INV_X1 U15718 ( .A(n13782), .ZN(n14521) );
  NOR4_X1 U15719 ( .A1(n13783), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13784), .A4(
        P2_U3088), .ZN(n13785) );
  AOI21_X1 U15720 ( .B1(n13790), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13785), 
        .ZN(n13786) );
  OAI21_X1 U15721 ( .B1(n14521), .B2(n13800), .A(n13786), .ZN(P2_U3296) );
  OAI222_X1 U15722 ( .A1(n13800), .A2(n13789), .B1(P2_U3088), .B2(n13788), 
        .C1(n13787), .C2(n13803), .ZN(P2_U3298) );
  NAND2_X1 U15723 ( .A1(n13790), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13791) );
  OAI211_X1 U15724 ( .C1(n13793), .C2(n13800), .A(n13792), .B(n13791), .ZN(
        P2_U3299) );
  INV_X1 U15725 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13796) );
  INV_X1 U15726 ( .A(n13794), .ZN(n14523) );
  OAI222_X1 U15727 ( .A1(n13803), .A2(n13796), .B1(n13800), .B2(n14523), .C1(
        P2_U3088), .C2(n13795), .ZN(P2_U3300) );
  OAI222_X1 U15728 ( .A1(n13798), .A2(P2_U3088), .B1(n13800), .B2(n14526), 
        .C1(n13797), .C2(n13803), .ZN(P2_U3301) );
  INV_X1 U15729 ( .A(n9411), .ZN(n14530) );
  OAI222_X1 U15730 ( .A1(n13803), .A2(n13801), .B1(n13800), .B2(n14530), .C1(
        n13799), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15731 ( .A(n13802), .ZN(n14533) );
  OAI222_X1 U15732 ( .A1(n13805), .A2(P2_U3088), .B1(n13800), .B2(n14533), 
        .C1(n13804), .C2(n13803), .ZN(P2_U3303) );
  MUX2_X1 U15733 ( .A(n13806), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15734 ( .A1(n14412), .A2(n6456), .ZN(n13808) );
  NAND2_X1 U15735 ( .A1(n14024), .A2(n13868), .ZN(n13807) );
  NAND2_X1 U15736 ( .A1(n13808), .A2(n13807), .ZN(n13809) );
  XNOR2_X1 U15737 ( .A(n13809), .B(n13921), .ZN(n13813) );
  NAND2_X1 U15738 ( .A1(n14412), .A2(n9675), .ZN(n13811) );
  NAND2_X1 U15739 ( .A1(n9680), .A2(n14024), .ZN(n13810) );
  NAND2_X1 U15740 ( .A1(n13811), .A2(n13810), .ZN(n13812) );
  NOR2_X1 U15741 ( .A1(n13813), .A2(n13812), .ZN(n13918) );
  NAND2_X1 U15742 ( .A1(n14470), .A2(n6456), .ZN(n13815) );
  NAND2_X1 U15743 ( .A1(n14361), .A2(n13880), .ZN(n13814) );
  NAND2_X1 U15744 ( .A1(n13815), .A2(n13814), .ZN(n13816) );
  XNOR2_X1 U15745 ( .A(n13816), .B(n13865), .ZN(n13822) );
  AND2_X1 U15746 ( .A1(n14361), .A2(n9680), .ZN(n13817) );
  AOI21_X1 U15747 ( .B1(n14470), .B2(n13829), .A(n13817), .ZN(n13821) );
  XNOR2_X1 U15748 ( .A(n13822), .B(n13821), .ZN(n13910) );
  NOR2_X1 U15749 ( .A1(n13819), .A2(n13818), .ZN(n13911) );
  NOR2_X1 U15750 ( .A1(n13910), .A2(n13911), .ZN(n13820) );
  OR2_X1 U15751 ( .A1(n13822), .A2(n13821), .ZN(n13823) );
  OAI22_X1 U15752 ( .A1(n14322), .A2(n13923), .B1(n13939), .B2(n13920), .ZN(
        n13825) );
  OAI22_X1 U15753 ( .A1(n14322), .A2(n13924), .B1(n13939), .B2(n13923), .ZN(
        n13824) );
  XNOR2_X1 U15754 ( .A(n13824), .B(n13921), .ZN(n13826) );
  XOR2_X1 U15755 ( .A(n13825), .B(n13826), .Z(n13980) );
  NAND2_X1 U15756 ( .A1(n13826), .A2(n13825), .ZN(n13827) );
  AOI22_X1 U15757 ( .A1(n14455), .A2(n6456), .B1(n13829), .B2(n14326), .ZN(
        n13830) );
  XNOR2_X1 U15758 ( .A(n13830), .B(n13921), .ZN(n13832) );
  AOI22_X1 U15759 ( .A1(n14455), .A2(n13868), .B1(n9680), .B2(n14326), .ZN(
        n13831) );
  NAND2_X1 U15760 ( .A1(n13832), .A2(n13831), .ZN(n13990) );
  OAI21_X1 U15761 ( .B1(n13832), .B2(n13831), .A(n13990), .ZN(n13938) );
  NAND2_X1 U15762 ( .A1(n14449), .A2(n6456), .ZN(n13834) );
  NAND2_X1 U15763 ( .A1(n14026), .A2(n13880), .ZN(n13833) );
  NAND2_X1 U15764 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  XNOR2_X1 U15765 ( .A(n13835), .B(n13865), .ZN(n13837) );
  AND2_X1 U15766 ( .A1(n9680), .A2(n14026), .ZN(n13836) );
  AOI21_X1 U15767 ( .B1(n14449), .B2(n13868), .A(n13836), .ZN(n13838) );
  NAND2_X1 U15768 ( .A1(n13837), .A2(n13838), .ZN(n13897) );
  INV_X1 U15769 ( .A(n13837), .ZN(n13840) );
  INV_X1 U15770 ( .A(n13838), .ZN(n13839) );
  NAND2_X1 U15771 ( .A1(n13840), .A2(n13839), .ZN(n13841) );
  AND2_X1 U15772 ( .A1(n13897), .A2(n13841), .ZN(n13991) );
  NAND2_X1 U15773 ( .A1(n13842), .A2(n13991), .ZN(n13896) );
  NAND2_X1 U15774 ( .A1(n13896), .A2(n13897), .ZN(n13852) );
  NAND2_X1 U15775 ( .A1(n14280), .A2(n6456), .ZN(n13844) );
  NAND2_X1 U15776 ( .A1(n14297), .A2(n13829), .ZN(n13843) );
  NAND2_X1 U15777 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  XNOR2_X1 U15778 ( .A(n13845), .B(n13865), .ZN(n13847) );
  AND2_X1 U15779 ( .A1(n9680), .A2(n14297), .ZN(n13846) );
  AOI21_X1 U15780 ( .B1(n14280), .B2(n9675), .A(n13846), .ZN(n13848) );
  NAND2_X1 U15781 ( .A1(n13847), .A2(n13848), .ZN(n13968) );
  INV_X1 U15782 ( .A(n13847), .ZN(n13850) );
  INV_X1 U15783 ( .A(n13848), .ZN(n13849) );
  NAND2_X1 U15784 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  NAND2_X1 U15785 ( .A1(n13852), .A2(n13898), .ZN(n13900) );
  NAND2_X1 U15786 ( .A1(n13900), .A2(n13968), .ZN(n13862) );
  NAND2_X1 U15787 ( .A1(n14251), .A2(n6456), .ZN(n13854) );
  NAND2_X1 U15788 ( .A1(n14276), .A2(n13868), .ZN(n13853) );
  NAND2_X1 U15789 ( .A1(n13854), .A2(n13853), .ZN(n13855) );
  XNOR2_X1 U15790 ( .A(n13855), .B(n13865), .ZN(n13857) );
  AND2_X1 U15791 ( .A1(n9680), .A2(n14276), .ZN(n13856) );
  AOI21_X1 U15792 ( .B1(n14251), .B2(n13868), .A(n13856), .ZN(n13858) );
  NAND2_X1 U15793 ( .A1(n13857), .A2(n13858), .ZN(n13946) );
  INV_X1 U15794 ( .A(n13857), .ZN(n13860) );
  INV_X1 U15795 ( .A(n13858), .ZN(n13859) );
  NAND2_X1 U15796 ( .A1(n13860), .A2(n13859), .ZN(n13861) );
  NAND2_X1 U15797 ( .A1(n13862), .A2(n13969), .ZN(n13945) );
  NAND2_X1 U15798 ( .A1(n13945), .A2(n13946), .ZN(n13874) );
  NAND2_X1 U15799 ( .A1(n14425), .A2(n6456), .ZN(n13864) );
  NAND2_X1 U15800 ( .A1(n14255), .A2(n13880), .ZN(n13863) );
  NAND2_X1 U15801 ( .A1(n13864), .A2(n13863), .ZN(n13866) );
  XNOR2_X1 U15802 ( .A(n13866), .B(n13865), .ZN(n13869) );
  AND2_X1 U15803 ( .A1(n9680), .A2(n14255), .ZN(n13867) );
  AOI21_X1 U15804 ( .B1(n14425), .B2(n13868), .A(n13867), .ZN(n13870) );
  NAND2_X1 U15805 ( .A1(n13869), .A2(n13870), .ZN(n13875) );
  INV_X1 U15806 ( .A(n13869), .ZN(n13872) );
  INV_X1 U15807 ( .A(n13870), .ZN(n13871) );
  NAND2_X1 U15808 ( .A1(n13872), .A2(n13871), .ZN(n13873) );
  NAND2_X1 U15809 ( .A1(n13874), .A2(n13947), .ZN(n13949) );
  NAND2_X1 U15810 ( .A1(n14225), .A2(n6456), .ZN(n13878) );
  NAND2_X1 U15811 ( .A1(n14025), .A2(n13880), .ZN(n13877) );
  NAND2_X1 U15812 ( .A1(n13878), .A2(n13877), .ZN(n13879) );
  XNOR2_X1 U15813 ( .A(n13879), .B(n13921), .ZN(n13884) );
  NAND2_X1 U15814 ( .A1(n14225), .A2(n13829), .ZN(n13882) );
  NAND2_X1 U15815 ( .A1(n9680), .A2(n14025), .ZN(n13881) );
  NAND2_X1 U15816 ( .A1(n13882), .A2(n13881), .ZN(n13883) );
  NOR2_X1 U15817 ( .A1(n13884), .A2(n13883), .ZN(n13885) );
  AOI21_X1 U15818 ( .B1(n13884), .B2(n13883), .A(n13885), .ZN(n14003) );
  INV_X1 U15819 ( .A(n13885), .ZN(n13886) );
  OAI21_X1 U15820 ( .B1(n13888), .B2(n13887), .A(n13919), .ZN(n13889) );
  NAND2_X1 U15821 ( .A1(n13889), .A2(n14655), .ZN(n13894) );
  NOR2_X1 U15822 ( .A1(n14707), .A2(n13890), .ZN(n13892) );
  OAI22_X1 U15823 ( .A1(n14401), .A2(n13975), .B1(n13974), .B2(n13952), .ZN(
        n13891) );
  AOI211_X1 U15824 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n13892), 
        .B(n13891), .ZN(n13893) );
  OAI211_X1 U15825 ( .C1(n13895), .C2(n14015), .A(n13894), .B(n13893), .ZN(
        P1_U3214) );
  NAND2_X1 U15826 ( .A1(n14280), .A2(n14793), .ZN(n14439) );
  INV_X1 U15827 ( .A(n13896), .ZN(n13994) );
  INV_X1 U15828 ( .A(n13897), .ZN(n13899) );
  NOR3_X1 U15829 ( .A1(n13994), .A2(n13899), .A3(n13898), .ZN(n13901) );
  INV_X1 U15830 ( .A(n13900), .ZN(n13971) );
  OAI21_X1 U15831 ( .B1(n13901), .B2(n13971), .A(n14655), .ZN(n13907) );
  NAND2_X1 U15832 ( .A1(n14026), .A2(n14483), .ZN(n13903) );
  NAND2_X1 U15833 ( .A1(n14276), .A2(n14739), .ZN(n13902) );
  NAND2_X1 U15834 ( .A1(n13903), .A2(n13902), .ZN(n14438) );
  INV_X1 U15835 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13904) );
  OAI22_X1 U15836 ( .A1(n14707), .A2(n14273), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13904), .ZN(n13905) );
  AOI21_X1 U15837 ( .B1(n14704), .B2(n14438), .A(n13905), .ZN(n13906) );
  OAI211_X1 U15838 ( .C1(n13908), .C2(n14439), .A(n13907), .B(n13906), .ZN(
        P1_U3216) );
  INV_X1 U15839 ( .A(n14470), .ZN(n14342) );
  INV_X1 U15840 ( .A(n13909), .ZN(n13912) );
  OAI21_X1 U15841 ( .B1(n13912), .B2(n13911), .A(n13910), .ZN(n13914) );
  NAND3_X1 U15842 ( .A1(n13914), .A2(n14655), .A3(n13913), .ZN(n13917) );
  OAI22_X1 U15843 ( .A1(n13939), .A2(n14474), .B1(n13964), .B2(n14400), .ZN(
        n14469) );
  NAND2_X1 U15844 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14198)
         );
  OAI21_X1 U15845 ( .B1(n14707), .B2(n14338), .A(n14198), .ZN(n13915) );
  AOI21_X1 U15846 ( .B1(n14469), .B2(n14704), .A(n13915), .ZN(n13916) );
  OAI211_X1 U15847 ( .C1(n14342), .C2(n14015), .A(n13917), .B(n13916), .ZN(
        P1_U3219) );
  OAI22_X1 U15848 ( .A1(n13925), .A2(n13923), .B1(n14401), .B2(n13920), .ZN(
        n13922) );
  XNOR2_X1 U15849 ( .A(n13922), .B(n13921), .ZN(n13927) );
  OAI22_X1 U15850 ( .A1(n13925), .A2(n13924), .B1(n14401), .B2(n13923), .ZN(
        n13926) );
  XNOR2_X1 U15851 ( .A(n13927), .B(n13926), .ZN(n13928) );
  OAI22_X1 U15852 ( .A1(n14707), .A2(n13930), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13929), .ZN(n13933) );
  INV_X1 U15853 ( .A(n14022), .ZN(n13931) );
  OAI22_X1 U15854 ( .A1(n13931), .A2(n13975), .B1(n13974), .B2(n14005), .ZN(
        n13932) );
  AOI211_X1 U15855 ( .C1(n14407), .C2(n14653), .A(n13933), .B(n13932), .ZN(
        n13934) );
  OAI21_X1 U15856 ( .B1(n13935), .B2(n14699), .A(n13934), .ZN(P1_U3220) );
  INV_X1 U15857 ( .A(n13937), .ZN(n13993) );
  AOI21_X1 U15858 ( .B1(n13936), .B2(n13938), .A(n13993), .ZN(n13944) );
  OAI22_X1 U15859 ( .A1(n13939), .A2(n14400), .B1(n14278), .B2(n14474), .ZN(
        n14454) );
  INV_X1 U15860 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13940) );
  OAI22_X1 U15861 ( .A1(n14707), .A2(n14308), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13940), .ZN(n13941) );
  AOI21_X1 U15862 ( .B1(n14454), .B2(n14704), .A(n13941), .ZN(n13943) );
  NAND2_X1 U15863 ( .A1(n14455), .A2(n14653), .ZN(n13942) );
  OAI211_X1 U15864 ( .C1(n13944), .C2(n14699), .A(n13943), .B(n13942), .ZN(
        P1_U3223) );
  INV_X1 U15865 ( .A(n14425), .ZN(n14240) );
  INV_X1 U15866 ( .A(n13945), .ZN(n13972) );
  INV_X1 U15867 ( .A(n13946), .ZN(n13948) );
  NOR3_X1 U15868 ( .A1(n13972), .A2(n13948), .A3(n13947), .ZN(n13951) );
  INV_X1 U15869 ( .A(n13949), .ZN(n13950) );
  OAI21_X1 U15870 ( .B1(n13951), .B2(n13950), .A(n14655), .ZN(n13956) );
  OAI22_X1 U15871 ( .A1(n11999), .A2(n14400), .B1(n13952), .B2(n14474), .ZN(
        n14424) );
  OAI22_X1 U15872 ( .A1(n14707), .A2(n14235), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13953), .ZN(n13954) );
  AOI21_X1 U15873 ( .B1(n14424), .B2(n14704), .A(n13954), .ZN(n13955) );
  OAI211_X1 U15874 ( .C1(n14240), .C2(n14015), .A(n13956), .B(n13955), .ZN(
        P1_U3225) );
  INV_X1 U15875 ( .A(n13957), .ZN(n14649) );
  INV_X1 U15876 ( .A(n13958), .ZN(n13960) );
  NOR3_X1 U15877 ( .A1(n14649), .A2(n13960), .A3(n13959), .ZN(n13963) );
  INV_X1 U15878 ( .A(n13961), .ZN(n13962) );
  OAI21_X1 U15879 ( .B1(n13963), .B2(n13962), .A(n14655), .ZN(n13967) );
  AND2_X1 U15880 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14732) );
  OAI22_X1 U15881 ( .A1(n14382), .A2(n13974), .B1(n13975), .B2(n13964), .ZN(
        n13965) );
  AOI211_X1 U15882 ( .C1(n13982), .C2(n14373), .A(n14732), .B(n13965), .ZN(
        n13966) );
  OAI211_X1 U15883 ( .C1(n14487), .C2(n14015), .A(n13967), .B(n13966), .ZN(
        P1_U3228) );
  INV_X1 U15884 ( .A(n13968), .ZN(n13970) );
  NOR3_X1 U15885 ( .A1(n13971), .A2(n13970), .A3(n13969), .ZN(n13973) );
  OAI21_X1 U15886 ( .B1(n13973), .B2(n13972), .A(n14655), .ZN(n13979) );
  NOR2_X1 U15887 ( .A1(n14707), .A2(n14246), .ZN(n13977) );
  OAI22_X1 U15888 ( .A1(n14006), .A2(n13975), .B1(n13974), .B2(n13996), .ZN(
        n13976) );
  AOI211_X1 U15889 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n13977), 
        .B(n13976), .ZN(n13978) );
  OAI211_X1 U15890 ( .C1(n12000), .C2(n14015), .A(n13979), .B(n13978), .ZN(
        P1_U3229) );
  XOR2_X1 U15891 ( .A(n13981), .B(n13980), .Z(n13988) );
  AOI22_X1 U15892 ( .A1(n13982), .A2(n14324), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13986) );
  NAND2_X1 U15893 ( .A1(n14361), .A2(n14483), .ZN(n13984) );
  NAND2_X1 U15894 ( .A1(n14326), .A2(n14739), .ZN(n13983) );
  NAND2_X1 U15895 ( .A1(n13984), .A2(n13983), .ZN(n14461) );
  NAND2_X1 U15896 ( .A1(n14461), .A2(n14704), .ZN(n13985) );
  OAI211_X1 U15897 ( .C1(n14322), .C2(n14015), .A(n13986), .B(n13985), .ZN(
        n13987) );
  AOI21_X1 U15898 ( .B1(n13988), .B2(n14655), .A(n13987), .ZN(n13989) );
  INV_X1 U15899 ( .A(n13989), .ZN(P1_U3233) );
  INV_X1 U15900 ( .A(n13990), .ZN(n13992) );
  NOR3_X1 U15901 ( .A1(n13993), .A2(n13992), .A3(n13991), .ZN(n13995) );
  OAI21_X1 U15902 ( .B1(n13995), .B2(n13994), .A(n14655), .ZN(n14000) );
  OAI22_X1 U15903 ( .A1(n14294), .A2(n14400), .B1(n13996), .B2(n14474), .ZN(
        n14448) );
  INV_X1 U15904 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13997) );
  OAI22_X1 U15905 ( .A1(n14707), .A2(n14292), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13997), .ZN(n13998) );
  AOI21_X1 U15906 ( .B1(n14448), .B2(n14704), .A(n13998), .ZN(n13999) );
  OAI211_X1 U15907 ( .C1(n14015), .C2(n14300), .A(n14000), .B(n13999), .ZN(
        P1_U3235) );
  OAI21_X1 U15908 ( .B1(n14003), .B2(n14002), .A(n14001), .ZN(n14004) );
  NAND2_X1 U15909 ( .A1(n14004), .A2(n14655), .ZN(n14010) );
  OAI22_X1 U15910 ( .A1(n14006), .A2(n14400), .B1(n14005), .B2(n14474), .ZN(
        n14221) );
  OAI22_X1 U15911 ( .A1(n14707), .A2(n14222), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14007), .ZN(n14008) );
  AOI21_X1 U15912 ( .B1(n14221), .B2(n14704), .A(n14008), .ZN(n14009) );
  OAI211_X1 U15913 ( .C1(n14418), .C2(n14015), .A(n14010), .B(n14009), .ZN(
        P1_U3240) );
  XNOR2_X1 U15914 ( .A(n14012), .B(n14011), .ZN(n14020) );
  OAI22_X1 U15915 ( .A1(n14707), .A2(n14014), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14013), .ZN(n14018) );
  NOR2_X1 U15916 ( .A1(n14016), .A2(n14015), .ZN(n14017) );
  AOI211_X1 U15917 ( .C1(n14704), .C2(n14662), .A(n14018), .B(n14017), .ZN(
        n14019) );
  OAI21_X1 U15918 ( .B1(n14020), .B2(n14699), .A(n14019), .ZN(P1_U3241) );
  MUX2_X1 U15919 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14204), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15920 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14021), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15921 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14022), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15922 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14023), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15923 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14024), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15924 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14025), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15925 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14255), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15926 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14276), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15927 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14297), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15928 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14026), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15929 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14326), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15930 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14027), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15931 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14361), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15932 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14484), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15933 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14028), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15934 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14482), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15935 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14029), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15936 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14030), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15937 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14031), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15938 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14032), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15939 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14033), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15940 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14034), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15941 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14035), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15942 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14036), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15943 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14037), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15944 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14038), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15945 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14740), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15946 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6450), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15947 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6651), .S(P1_U4016), .Z(
        P1_U3560) );
  AOI211_X1 U15948 ( .C1(n14042), .C2(n14041), .A(n14040), .B(n14729), .ZN(
        n14043) );
  INV_X1 U15949 ( .A(n14043), .ZN(n14051) );
  AOI22_X1 U15950 ( .A1(n14733), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14050) );
  NAND2_X1 U15951 ( .A1(n14722), .A2(n14044), .ZN(n14049) );
  NAND2_X1 U15952 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14053) );
  INV_X1 U15953 ( .A(n14053), .ZN(n14047) );
  OAI211_X1 U15954 ( .C1(n14047), .C2(n14046), .A(n14724), .B(n14045), .ZN(
        n14048) );
  NAND4_X1 U15955 ( .A1(n14051), .A2(n14050), .A3(n14049), .A4(n14048), .ZN(
        P1_U3244) );
  MUX2_X1 U15956 ( .A(n14053), .B(n14052), .S(n14524), .Z(n14056) );
  NOR2_X1 U15957 ( .A1(n14524), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14054) );
  OR2_X1 U15958 ( .A1(n14055), .A2(n14054), .ZN(n14709) );
  NAND2_X1 U15959 ( .A1(n14709), .A2(n14711), .ZN(n14714) );
  OAI211_X1 U15960 ( .C1(n14056), .C2(n14055), .A(P1_U4016), .B(n14714), .ZN(
        n14101) );
  INV_X1 U15961 ( .A(n14057), .ZN(n14060) );
  OAI22_X1 U15962 ( .A1(n14199), .A2(n14058), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10796), .ZN(n14059) );
  AOI21_X1 U15963 ( .B1(n14060), .B2(n14722), .A(n14059), .ZN(n14068) );
  OAI211_X1 U15964 ( .C1(n14062), .C2(n14061), .A(n14724), .B(n14070), .ZN(
        n14067) );
  AOI211_X1 U15965 ( .C1(n14064), .C2(n14063), .A(n14079), .B(n14729), .ZN(
        n14065) );
  INV_X1 U15966 ( .A(n14065), .ZN(n14066) );
  NAND4_X1 U15967 ( .A1(n14101), .A2(n14068), .A3(n14067), .A4(n14066), .ZN(
        P1_U3245) );
  MUX2_X1 U15968 ( .A(n10038), .B(P1_REG2_REG_3__SCAN_IN), .S(n14074), .Z(
        n14071) );
  NAND3_X1 U15969 ( .A1(n14071), .A2(n14070), .A3(n14069), .ZN(n14072) );
  NAND3_X1 U15970 ( .A1(n14724), .A2(n14095), .A3(n14072), .ZN(n14083) );
  NOR2_X1 U15971 ( .A1(n14073), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14695) );
  AOI21_X1 U15972 ( .B1(n14733), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14695), .ZN(
        n14082) );
  NAND2_X1 U15973 ( .A1(n14722), .A2(n14074), .ZN(n14081) );
  MUX2_X1 U15974 ( .A(n10024), .B(P1_REG1_REG_3__SCAN_IN), .S(n14074), .Z(
        n14077) );
  INV_X1 U15975 ( .A(n14075), .ZN(n14076) );
  NAND2_X1 U15976 ( .A1(n14077), .A2(n14076), .ZN(n14078) );
  OAI211_X1 U15977 ( .C1(n14079), .C2(n14078), .A(n14194), .B(n14090), .ZN(
        n14080) );
  NAND4_X1 U15978 ( .A1(n14083), .A2(n14082), .A3(n14081), .A4(n14080), .ZN(
        P1_U3246) );
  INV_X1 U15979 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14085) );
  OAI21_X1 U15980 ( .B1(n14199), .B2(n14085), .A(n14084), .ZN(n14086) );
  AOI21_X1 U15981 ( .B1(n14093), .B2(n14722), .A(n14086), .ZN(n14100) );
  INV_X1 U15982 ( .A(n14087), .ZN(n14092) );
  NAND3_X1 U15983 ( .A1(n14090), .A2(n14089), .A3(n14088), .ZN(n14091) );
  NAND3_X1 U15984 ( .A1(n14194), .A2(n14092), .A3(n14091), .ZN(n14099) );
  MUX2_X1 U15985 ( .A(n11097), .B(P1_REG2_REG_4__SCAN_IN), .S(n14093), .Z(
        n14096) );
  NAND3_X1 U15986 ( .A1(n14096), .A2(n14095), .A3(n14094), .ZN(n14097) );
  NAND3_X1 U15987 ( .A1(n14724), .A2(n14112), .A3(n14097), .ZN(n14098) );
  NAND4_X1 U15988 ( .A1(n14101), .A2(n14100), .A3(n14099), .A4(n14098), .ZN(
        P1_U3247) );
  INV_X1 U15989 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14103) );
  OAI21_X1 U15990 ( .B1(n14199), .B2(n14103), .A(n14102), .ZN(n14104) );
  AOI21_X1 U15991 ( .B1(n14109), .B2(n14722), .A(n14104), .ZN(n14116) );
  OAI21_X1 U15992 ( .B1(n14107), .B2(n14106), .A(n14105), .ZN(n14108) );
  NAND2_X1 U15993 ( .A1(n14108), .A2(n14194), .ZN(n14115) );
  MUX2_X1 U15994 ( .A(n10047), .B(P1_REG2_REG_5__SCAN_IN), .S(n14109), .Z(
        n14110) );
  NAND3_X1 U15995 ( .A1(n14112), .A2(n14111), .A3(n14110), .ZN(n14113) );
  NAND3_X1 U15996 ( .A1(n14724), .A2(n14128), .A3(n14113), .ZN(n14114) );
  NAND3_X1 U15997 ( .A1(n14116), .A2(n14115), .A3(n14114), .ZN(P1_U3248) );
  INV_X1 U15998 ( .A(n14117), .ZN(n14121) );
  MUX2_X1 U15999 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n14118), .S(n14125), .Z(
        n14120) );
  OAI211_X1 U16000 ( .C1(n14121), .C2(n14120), .A(n14194), .B(n14119), .ZN(
        n14133) );
  OAI21_X1 U16001 ( .B1(n14199), .B2(n14123), .A(n14122), .ZN(n14124) );
  AOI21_X1 U16002 ( .B1(n14125), .B2(n14722), .A(n14124), .ZN(n14132) );
  MUX2_X1 U16003 ( .A(n11172), .B(P1_REG2_REG_6__SCAN_IN), .S(n14125), .Z(
        n14127) );
  NAND3_X1 U16004 ( .A1(n14128), .A2(n14127), .A3(n14126), .ZN(n14129) );
  NAND3_X1 U16005 ( .A1(n14724), .A2(n14130), .A3(n14129), .ZN(n14131) );
  NAND3_X1 U16006 ( .A1(n14133), .A2(n14132), .A3(n14131), .ZN(P1_U3249) );
  OAI21_X1 U16007 ( .B1(n14135), .B2(n14134), .A(n14150), .ZN(n14136) );
  NAND2_X1 U16008 ( .A1(n14136), .A2(n14194), .ZN(n14147) );
  OAI21_X1 U16009 ( .B1(n14199), .B2(n14138), .A(n14137), .ZN(n14139) );
  AOI21_X1 U16010 ( .B1(n14140), .B2(n14722), .A(n14139), .ZN(n14146) );
  MUX2_X1 U16011 ( .A(n10294), .B(P1_REG2_REG_8__SCAN_IN), .S(n14140), .Z(
        n14141) );
  NAND3_X1 U16012 ( .A1(n14143), .A2(n14142), .A3(n14141), .ZN(n14144) );
  NAND3_X1 U16013 ( .A1(n14724), .A2(n14156), .A3(n14144), .ZN(n14145) );
  NAND3_X1 U16014 ( .A1(n14147), .A2(n14146), .A3(n14145), .ZN(P1_U3251) );
  AND3_X1 U16015 ( .A1(n14150), .A2(n14149), .A3(n14148), .ZN(n14151) );
  OAI21_X1 U16016 ( .B1(n14152), .B2(n14151), .A(n14194), .ZN(n14163) );
  AOI21_X1 U16017 ( .B1(n14733), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n14153), .ZN(
        n14162) );
  MUX2_X1 U16018 ( .A(n11483), .B(P1_REG2_REG_9__SCAN_IN), .S(n14159), .Z(
        n14154) );
  NAND3_X1 U16019 ( .A1(n14156), .A2(n14155), .A3(n14154), .ZN(n14157) );
  NAND3_X1 U16020 ( .A1(n14724), .A2(n14158), .A3(n14157), .ZN(n14161) );
  NAND2_X1 U16021 ( .A1(n14722), .A2(n14159), .ZN(n14160) );
  NAND4_X1 U16022 ( .A1(n14163), .A2(n14162), .A3(n14161), .A4(n14160), .ZN(
        P1_U3252) );
  NAND2_X1 U16023 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14658)
         );
  XNOR2_X1 U16024 ( .A(n14165), .B(n14164), .ZN(n14166) );
  NAND2_X1 U16025 ( .A1(n14166), .A2(n14194), .ZN(n14167) );
  AND2_X1 U16026 ( .A1(n14658), .A2(n14167), .ZN(n14175) );
  AOI22_X1 U16027 ( .A1(n14722), .A2(n14168), .B1(n14733), .B2(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n14174) );
  MUX2_X1 U16028 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n14169), .S(n14168), .Z(
        n14171) );
  OAI211_X1 U16029 ( .C1(n14172), .C2(n14171), .A(n14170), .B(n14724), .ZN(
        n14173) );
  NAND3_X1 U16030 ( .A1(n14175), .A2(n14174), .A3(n14173), .ZN(P1_U3259) );
  INV_X1 U16031 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14181) );
  INV_X1 U16032 ( .A(n14176), .ZN(n14177) );
  NAND2_X1 U16033 ( .A1(n14177), .A2(n14184), .ZN(n14179) );
  NAND2_X1 U16034 ( .A1(n14179), .A2(n14178), .ZN(n14180) );
  INV_X1 U16035 ( .A(n14182), .ZN(n14183) );
  NAND2_X1 U16036 ( .A1(n14183), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14187) );
  NAND2_X1 U16037 ( .A1(n14185), .A2(n14184), .ZN(n14186) );
  NAND2_X1 U16038 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  XOR2_X1 U16039 ( .A(n14188), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14191) );
  AOI22_X1 U16040 ( .A1(n14189), .A2(n14194), .B1(n14191), .B2(n14724), .ZN(
        n14197) );
  INV_X1 U16041 ( .A(n14189), .ZN(n14193) );
  NOR2_X1 U16042 ( .A1(n14191), .A2(n14190), .ZN(n14192) );
  AOI211_X1 U16043 ( .C1(n14194), .C2(n14193), .A(n14722), .B(n14192), .ZN(
        n14196) );
  NAND2_X1 U16044 ( .A1(n14397), .A2(n14208), .ZN(n14207) );
  XOR2_X1 U16045 ( .A(n14392), .B(n14207), .Z(n14201) );
  NAND2_X1 U16046 ( .A1(n14201), .A2(n14370), .ZN(n14393) );
  NOR2_X1 U16047 ( .A1(n14377), .A2(n14202), .ZN(n14205) );
  NAND2_X1 U16048 ( .A1(n14204), .A2(n14203), .ZN(n14395) );
  NOR2_X1 U16049 ( .A1(n14325), .A2(n14395), .ZN(n14209) );
  AOI211_X1 U16050 ( .C1(n14392), .C2(n14384), .A(n14205), .B(n14209), .ZN(
        n14206) );
  OAI21_X1 U16051 ( .B1(n14393), .B2(n14387), .A(n14206), .ZN(P1_U3263) );
  OAI211_X1 U16052 ( .C1(n14397), .C2(n14208), .A(n14370), .B(n14207), .ZN(
        n14396) );
  AOI21_X1 U16053 ( .B1(n14325), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14209), 
        .ZN(n14212) );
  NAND2_X1 U16054 ( .A1(n14210), .A2(n14384), .ZN(n14211) );
  OAI211_X1 U16055 ( .C1(n14396), .C2(n14387), .A(n14212), .B(n14211), .ZN(
        P1_U3264) );
  XNOR2_X1 U16056 ( .A(n14213), .B(n14217), .ZN(n14422) );
  INV_X1 U16057 ( .A(n14214), .ZN(n14218) );
  INV_X1 U16058 ( .A(n14215), .ZN(n14216) );
  OAI21_X1 U16059 ( .B1(n14218), .B2(n14217), .A(n14216), .ZN(n14420) );
  OAI211_X1 U16060 ( .C1(n14418), .C2(n14234), .A(n14370), .B(n14219), .ZN(
        n14417) );
  NOR2_X1 U16061 ( .A1(n14377), .A2(n14220), .ZN(n14224) );
  INV_X1 U16062 ( .A(n14221), .ZN(n14416) );
  OAI22_X1 U16063 ( .A1(n14416), .A2(n14325), .B1(n14222), .B2(n14374), .ZN(
        n14223) );
  AOI211_X1 U16064 ( .C1(n14225), .C2(n14384), .A(n14224), .B(n14223), .ZN(
        n14226) );
  OAI21_X1 U16065 ( .B1(n14417), .B2(n14387), .A(n14226), .ZN(n14227) );
  AOI21_X1 U16066 ( .B1(n14420), .B2(n14389), .A(n14227), .ZN(n14228) );
  OAI21_X1 U16067 ( .B1(n14391), .B2(n14422), .A(n14228), .ZN(P1_U3267) );
  XOR2_X1 U16068 ( .A(n14231), .B(n6499), .Z(n14429) );
  AOI21_X1 U16069 ( .B1(n14231), .B2(n14230), .A(n14229), .ZN(n14426) );
  NAND2_X1 U16070 ( .A1(n14425), .A2(n6483), .ZN(n14232) );
  NAND2_X1 U16071 ( .A1(n14232), .A2(n14370), .ZN(n14233) );
  NOR2_X1 U16072 ( .A1(n14234), .A2(n14233), .ZN(n14423) );
  NAND2_X1 U16073 ( .A1(n14423), .A2(n14357), .ZN(n14239) );
  INV_X1 U16074 ( .A(n14424), .ZN(n14236) );
  OAI22_X1 U16075 ( .A1(n14236), .A2(n14325), .B1(n14235), .B2(n14374), .ZN(
        n14237) );
  AOI21_X1 U16076 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n14325), .A(n14237), 
        .ZN(n14238) );
  OAI211_X1 U16077 ( .C1(n14240), .C2(n14364), .A(n14239), .B(n14238), .ZN(
        n14241) );
  AOI21_X1 U16078 ( .B1(n14426), .B2(n14337), .A(n14241), .ZN(n14242) );
  OAI21_X1 U16079 ( .B1(n14346), .B2(n14429), .A(n14242), .ZN(P1_U3268) );
  NAND2_X1 U16080 ( .A1(n14243), .A2(n14253), .ZN(n14244) );
  NAND2_X1 U16081 ( .A1(n14245), .A2(n14244), .ZN(n14431) );
  INV_X1 U16082 ( .A(n14431), .ZN(n14263) );
  OAI22_X1 U16083 ( .A1(n14377), .A2(n14247), .B1(n14246), .B2(n14374), .ZN(
        n14250) );
  AOI21_X1 U16084 ( .B1(n14251), .B2(n14271), .A(n14355), .ZN(n14248) );
  NAND2_X1 U16085 ( .A1(n14248), .A2(n6483), .ZN(n14432) );
  NOR2_X1 U16086 ( .A1(n14432), .A2(n14387), .ZN(n14249) );
  AOI211_X1 U16087 ( .C1(n14384), .C2(n14251), .A(n14250), .B(n14249), .ZN(
        n14261) );
  OAI21_X1 U16088 ( .B1(n14253), .B2(n14252), .A(n14489), .ZN(n14258) );
  NAND2_X1 U16089 ( .A1(n14431), .A2(n14254), .ZN(n14257) );
  AOI22_X1 U16090 ( .A1(n14483), .A2(n14297), .B1(n14255), .B2(n14739), .ZN(
        n14256) );
  OAI211_X1 U16091 ( .C1(n14259), .C2(n14258), .A(n14257), .B(n14256), .ZN(
        n14435) );
  NAND2_X1 U16092 ( .A1(n14435), .A2(n14377), .ZN(n14260) );
  OAI211_X1 U16093 ( .C1(n14263), .C2(n14262), .A(n14261), .B(n14260), .ZN(
        P1_U3269) );
  OAI21_X1 U16094 ( .B1(n14265), .B2(n14270), .A(n14264), .ZN(n14266) );
  AND2_X1 U16095 ( .A1(n14266), .A2(n14489), .ZN(n14443) );
  INV_X1 U16096 ( .A(n14443), .ZN(n14284) );
  INV_X1 U16097 ( .A(n14267), .ZN(n14268) );
  AOI21_X1 U16098 ( .B1(n14270), .B2(n14269), .A(n14268), .ZN(n14444) );
  OAI211_X1 U16099 ( .C1(n14272), .C2(n14291), .A(n14370), .B(n14271), .ZN(
        n14441) );
  OAI22_X1 U16100 ( .A1(n14377), .A2(n14274), .B1(n14273), .B2(n14374), .ZN(
        n14275) );
  AOI21_X1 U16101 ( .B1(n14379), .B2(n14276), .A(n14275), .ZN(n14277) );
  OAI21_X1 U16102 ( .B1(n14278), .B2(n14381), .A(n14277), .ZN(n14279) );
  AOI21_X1 U16103 ( .B1(n14280), .B2(n14384), .A(n14279), .ZN(n14281) );
  OAI21_X1 U16104 ( .B1(n14441), .B2(n14387), .A(n14281), .ZN(n14282) );
  AOI21_X1 U16105 ( .B1(n14444), .B2(n14337), .A(n14282), .ZN(n14283) );
  OAI21_X1 U16106 ( .B1(n14325), .B2(n14284), .A(n14283), .ZN(P1_U3270) );
  XNOR2_X1 U16107 ( .A(n14285), .B(n14287), .ZN(n14452) );
  OAI21_X1 U16108 ( .B1(n14288), .B2(n14287), .A(n14286), .ZN(n14446) );
  NAND2_X1 U16109 ( .A1(n14449), .A2(n14306), .ZN(n14289) );
  NAND2_X1 U16110 ( .A1(n14289), .A2(n14370), .ZN(n14290) );
  NOR2_X1 U16111 ( .A1(n14291), .A2(n14290), .ZN(n14447) );
  NAND2_X1 U16112 ( .A1(n14447), .A2(n14357), .ZN(n14299) );
  OAI22_X1 U16113 ( .A1(n14377), .A2(n14293), .B1(n14292), .B2(n14374), .ZN(
        n14296) );
  NOR2_X1 U16114 ( .A1(n14381), .A2(n14294), .ZN(n14295) );
  AOI211_X1 U16115 ( .C1(n14379), .C2(n14297), .A(n14296), .B(n14295), .ZN(
        n14298) );
  OAI211_X1 U16116 ( .C1(n14364), .C2(n14300), .A(n14299), .B(n14298), .ZN(
        n14301) );
  AOI21_X1 U16117 ( .B1(n14446), .B2(n14337), .A(n14301), .ZN(n14302) );
  OAI21_X1 U16118 ( .B1(n14452), .B2(n14346), .A(n14302), .ZN(P1_U3271) );
  XNOR2_X1 U16119 ( .A(n14303), .B(n14304), .ZN(n14459) );
  XNOR2_X1 U16120 ( .A(n14305), .B(n14304), .ZN(n14456) );
  NAND2_X1 U16121 ( .A1(n14456), .A2(n14337), .ZN(n14314) );
  INV_X1 U16122 ( .A(n14306), .ZN(n14307) );
  AOI211_X1 U16123 ( .C1(n14455), .C2(n14321), .A(n14355), .B(n14307), .ZN(
        n14453) );
  OAI22_X1 U16124 ( .A1(n14377), .A2(n14309), .B1(n14308), .B2(n14374), .ZN(
        n14310) );
  AOI21_X1 U16125 ( .B1(n14454), .B2(n14377), .A(n14310), .ZN(n14311) );
  OAI21_X1 U16126 ( .B1(n6865), .B2(n14364), .A(n14311), .ZN(n14312) );
  AOI21_X1 U16127 ( .B1(n14453), .B2(n14357), .A(n14312), .ZN(n14313) );
  OAI211_X1 U16128 ( .C1(n14459), .C2(n14346), .A(n14314), .B(n14313), .ZN(
        P1_U3272) );
  OAI211_X1 U16129 ( .C1(n14316), .C2(n14320), .A(n14489), .B(n14315), .ZN(
        n14464) );
  INV_X1 U16130 ( .A(n14317), .ZN(n14318) );
  AOI21_X1 U16131 ( .B1(n14320), .B2(n14319), .A(n14318), .ZN(n14460) );
  OAI211_X1 U16132 ( .C1(n14322), .C2(n6586), .A(n14370), .B(n14321), .ZN(
        n14463) );
  AOI22_X1 U16133 ( .A1(n14325), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14324), 
        .B2(n14323), .ZN(n14328) );
  NAND2_X1 U16134 ( .A1(n14379), .A2(n14326), .ZN(n14327) );
  OAI211_X1 U16135 ( .C1(n14475), .C2(n14381), .A(n14328), .B(n14327), .ZN(
        n14329) );
  AOI21_X1 U16136 ( .B1(n14462), .B2(n14384), .A(n14329), .ZN(n14330) );
  OAI21_X1 U16137 ( .B1(n14463), .B2(n14387), .A(n14330), .ZN(n14331) );
  AOI21_X1 U16138 ( .B1(n14460), .B2(n14337), .A(n14331), .ZN(n14332) );
  OAI21_X1 U16139 ( .B1(n14325), .B2(n14464), .A(n14332), .ZN(P1_U3273) );
  XNOR2_X1 U16140 ( .A(n14334), .B(n14333), .ZN(n14473) );
  XNOR2_X1 U16141 ( .A(n14336), .B(n14335), .ZN(n14467) );
  NAND2_X1 U16142 ( .A1(n14467), .A2(n14337), .ZN(n14345) );
  AOI211_X1 U16143 ( .C1(n14470), .C2(n14353), .A(n14355), .B(n6586), .ZN(
        n14468) );
  INV_X1 U16144 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14339) );
  OAI22_X1 U16145 ( .A1(n14377), .A2(n14339), .B1(n14338), .B2(n14374), .ZN(
        n14340) );
  AOI21_X1 U16146 ( .B1(n14469), .B2(n14377), .A(n14340), .ZN(n14341) );
  OAI21_X1 U16147 ( .B1(n14342), .B2(n14364), .A(n14341), .ZN(n14343) );
  AOI21_X1 U16148 ( .B1(n14468), .B2(n14357), .A(n14343), .ZN(n14344) );
  OAI211_X1 U16149 ( .C1(n14473), .C2(n14346), .A(n14345), .B(n14344), .ZN(
        P1_U3274) );
  XOR2_X1 U16150 ( .A(n14347), .B(n14348), .Z(n14481) );
  XNOR2_X1 U16151 ( .A(n14349), .B(n14348), .ZN(n14351) );
  OAI22_X1 U16152 ( .A1(n14351), .A2(n14795), .B1(n14350), .B2(n14400), .ZN(
        n14479) );
  INV_X1 U16153 ( .A(n14352), .ZN(n14371) );
  INV_X1 U16154 ( .A(n14353), .ZN(n14354) );
  AOI211_X1 U16155 ( .C1(n14356), .C2(n14371), .A(n14355), .B(n14354), .ZN(
        n14478) );
  NAND2_X1 U16156 ( .A1(n14478), .A2(n14357), .ZN(n14363) );
  OAI22_X1 U16157 ( .A1(n14377), .A2(n14359), .B1(n14358), .B2(n14374), .ZN(
        n14360) );
  AOI21_X1 U16158 ( .B1(n14379), .B2(n14361), .A(n14360), .ZN(n14362) );
  OAI211_X1 U16159 ( .C1(n14476), .C2(n14364), .A(n14363), .B(n14362), .ZN(
        n14365) );
  AOI21_X1 U16160 ( .B1(n14479), .B2(n14377), .A(n14365), .ZN(n14366) );
  OAI21_X1 U16161 ( .B1(n14481), .B2(n14391), .A(n14366), .ZN(P1_U3275) );
  XNOR2_X1 U16162 ( .A(n14367), .B(n14368), .ZN(n14492) );
  XNOR2_X1 U16163 ( .A(n14369), .B(n14368), .ZN(n14490) );
  OAI211_X1 U16164 ( .C1(n14487), .C2(n14372), .A(n14371), .B(n14370), .ZN(
        n14486) );
  INV_X1 U16165 ( .A(n14373), .ZN(n14375) );
  OAI22_X1 U16166 ( .A1(n14377), .A2(n14376), .B1(n14375), .B2(n14374), .ZN(
        n14378) );
  AOI21_X1 U16167 ( .B1(n14379), .B2(n14484), .A(n14378), .ZN(n14380) );
  OAI21_X1 U16168 ( .B1(n14382), .B2(n14381), .A(n14380), .ZN(n14383) );
  AOI21_X1 U16169 ( .B1(n14385), .B2(n14384), .A(n14383), .ZN(n14386) );
  OAI21_X1 U16170 ( .B1(n14486), .B2(n14387), .A(n14386), .ZN(n14388) );
  AOI21_X1 U16171 ( .B1(n14490), .B2(n14389), .A(n14388), .ZN(n14390) );
  OAI21_X1 U16172 ( .B1(n14492), .B2(n14391), .A(n14390), .ZN(P1_U3276) );
  INV_X1 U16173 ( .A(n14392), .ZN(n14394) );
  OAI211_X1 U16174 ( .C1(n14394), .C2(n14775), .A(n14393), .B(n14395), .ZN(
        n14498) );
  MUX2_X1 U16175 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14498), .S(n14813), .Z(
        P1_U3559) );
  OAI211_X1 U16176 ( .C1(n14397), .C2(n14775), .A(n14396), .B(n14395), .ZN(
        n14499) );
  MUX2_X1 U16177 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14499), .S(n14813), .Z(
        P1_U3558) );
  OAI21_X1 U16178 ( .B1(n14401), .B2(n14400), .A(n14399), .ZN(n14403) );
  AOI21_X1 U16179 ( .B1(n14793), .B2(n14407), .A(n14406), .ZN(n14408) );
  OAI211_X1 U16180 ( .C1(n14753), .C2(n14410), .A(n14409), .B(n14408), .ZN(
        n14500) );
  MUX2_X1 U16181 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14500), .S(n14813), .Z(
        P1_U3556) );
  AOI21_X1 U16182 ( .B1(n14793), .B2(n14412), .A(n14411), .ZN(n14413) );
  OAI211_X1 U16183 ( .C1(n14415), .C2(n14430), .A(n14414), .B(n14413), .ZN(
        n14501) );
  MUX2_X1 U16184 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14501), .S(n14813), .Z(
        P1_U3555) );
  OAI211_X1 U16185 ( .C1(n14418), .C2(n14775), .A(n14417), .B(n14416), .ZN(
        n14419) );
  AOI21_X1 U16186 ( .B1(n14420), .B2(n14489), .A(n14419), .ZN(n14421) );
  OAI21_X1 U16187 ( .B1(n14753), .B2(n14422), .A(n14421), .ZN(n14502) );
  MUX2_X1 U16188 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14502), .S(n14813), .Z(
        P1_U3554) );
  AOI211_X1 U16189 ( .C1(n14793), .C2(n14425), .A(n14424), .B(n14423), .ZN(
        n14428) );
  NAND2_X1 U16190 ( .A1(n14426), .A2(n14799), .ZN(n14427) );
  OAI211_X1 U16191 ( .C1(n14429), .C2(n14795), .A(n14428), .B(n14427), .ZN(
        n14503) );
  MUX2_X1 U16192 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14503), .S(n14813), .Z(
        P1_U3553) );
  INV_X1 U16193 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14436) );
  INV_X1 U16194 ( .A(n14430), .ZN(n14785) );
  NAND2_X1 U16195 ( .A1(n14431), .A2(n14785), .ZN(n14433) );
  OAI211_X1 U16196 ( .C1(n12000), .C2(n14775), .A(n14433), .B(n14432), .ZN(
        n14434) );
  NOR2_X1 U16197 ( .A1(n14435), .A2(n14434), .ZN(n14504) );
  MUX2_X1 U16198 ( .A(n14436), .B(n14504), .S(n14813), .Z(n14437) );
  INV_X1 U16199 ( .A(n14437), .ZN(P1_U3552) );
  INV_X1 U16200 ( .A(n14438), .ZN(n14440) );
  NAND3_X1 U16201 ( .A1(n14441), .A2(n14440), .A3(n14439), .ZN(n14442) );
  AOI211_X1 U16202 ( .C1(n14444), .C2(n14799), .A(n14443), .B(n14442), .ZN(
        n14445) );
  INV_X1 U16203 ( .A(n14445), .ZN(n14507) );
  MUX2_X1 U16204 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14507), .S(n14813), .Z(
        P1_U3551) );
  NAND2_X1 U16205 ( .A1(n14446), .A2(n14799), .ZN(n14451) );
  AOI211_X1 U16206 ( .C1(n14793), .C2(n14449), .A(n14448), .B(n14447), .ZN(
        n14450) );
  OAI211_X1 U16207 ( .C1(n14795), .C2(n14452), .A(n14451), .B(n14450), .ZN(
        n14508) );
  MUX2_X1 U16208 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14508), .S(n14813), .Z(
        P1_U3550) );
  AOI211_X1 U16209 ( .C1(n14793), .C2(n14455), .A(n14454), .B(n14453), .ZN(
        n14458) );
  NAND2_X1 U16210 ( .A1(n14456), .A2(n14799), .ZN(n14457) );
  OAI211_X1 U16211 ( .C1(n14795), .C2(n14459), .A(n14458), .B(n14457), .ZN(
        n14509) );
  MUX2_X1 U16212 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14509), .S(n14813), .Z(
        P1_U3549) );
  NAND2_X1 U16213 ( .A1(n14460), .A2(n14799), .ZN(n14466) );
  AOI21_X1 U16214 ( .B1(n14462), .B2(n14793), .A(n14461), .ZN(n14465) );
  NAND4_X1 U16215 ( .A1(n14466), .A2(n14465), .A3(n14464), .A4(n14463), .ZN(
        n14510) );
  MUX2_X1 U16216 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14510), .S(n14813), .Z(
        P1_U3548) );
  NAND2_X1 U16217 ( .A1(n14467), .A2(n14799), .ZN(n14472) );
  AOI211_X1 U16218 ( .C1(n14793), .C2(n14470), .A(n14469), .B(n14468), .ZN(
        n14471) );
  OAI211_X1 U16219 ( .C1(n14795), .C2(n14473), .A(n14472), .B(n14471), .ZN(
        n14511) );
  MUX2_X1 U16220 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14511), .S(n14813), .Z(
        P1_U3547) );
  OAI22_X1 U16221 ( .A1(n14476), .A2(n14775), .B1(n14475), .B2(n14474), .ZN(
        n14477) );
  NOR3_X1 U16222 ( .A1(n14479), .A2(n14478), .A3(n14477), .ZN(n14480) );
  OAI21_X1 U16223 ( .B1(n14481), .B2(n14753), .A(n14480), .ZN(n14512) );
  MUX2_X1 U16224 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14512), .S(n14813), .Z(
        P1_U3546) );
  AOI22_X1 U16225 ( .A1(n14484), .A2(n14739), .B1(n14483), .B2(n14482), .ZN(
        n14485) );
  OAI211_X1 U16226 ( .C1(n14487), .C2(n14775), .A(n14486), .B(n14485), .ZN(
        n14488) );
  AOI21_X1 U16227 ( .B1(n14490), .B2(n14489), .A(n14488), .ZN(n14491) );
  OAI21_X1 U16228 ( .B1(n14492), .B2(n14753), .A(n14491), .ZN(n14513) );
  MUX2_X1 U16229 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14513), .S(n14813), .Z(
        P1_U3545) );
  AOI211_X1 U16230 ( .C1(n14793), .C2(n14654), .A(n14657), .B(n14493), .ZN(
        n14496) );
  NAND2_X1 U16231 ( .A1(n14494), .A2(n14799), .ZN(n14495) );
  OAI211_X1 U16232 ( .C1(n14497), .C2(n14795), .A(n14496), .B(n14495), .ZN(
        n14514) );
  MUX2_X1 U16233 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14514), .S(n14813), .Z(
        P1_U3544) );
  MUX2_X1 U16234 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14498), .S(n14802), .Z(
        P1_U3527) );
  MUX2_X1 U16235 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14499), .S(n14802), .Z(
        P1_U3526) );
  MUX2_X1 U16236 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14500), .S(n14802), .Z(
        P1_U3524) );
  MUX2_X1 U16237 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14501), .S(n14802), .Z(
        P1_U3523) );
  MUX2_X1 U16238 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14502), .S(n14802), .Z(
        P1_U3522) );
  MUX2_X1 U16239 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14503), .S(n14802), .Z(
        P1_U3521) );
  MUX2_X1 U16240 ( .A(n14505), .B(n14504), .S(n14802), .Z(n14506) );
  INV_X1 U16241 ( .A(n14506), .ZN(P1_U3520) );
  MUX2_X1 U16242 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14507), .S(n14802), .Z(
        P1_U3519) );
  MUX2_X1 U16243 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14508), .S(n14802), .Z(
        P1_U3518) );
  MUX2_X1 U16244 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14509), .S(n14802), .Z(
        P1_U3517) );
  MUX2_X1 U16245 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14510), .S(n14802), .Z(
        P1_U3516) );
  MUX2_X1 U16246 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14511), .S(n14802), .Z(
        P1_U3515) );
  MUX2_X1 U16247 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14512), .S(n14802), .Z(
        P1_U3513) );
  MUX2_X1 U16248 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14513), .S(n14802), .Z(
        P1_U3510) );
  MUX2_X1 U16249 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14514), .S(n14802), .Z(
        P1_U3507) );
  INV_X1 U16250 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14515) );
  NAND3_X1 U16251 ( .A1(n14515), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n14517) );
  OAI22_X1 U16252 ( .A1(n14518), .A2(n14517), .B1(n14516), .B2(n14528), .ZN(
        n14519) );
  INV_X1 U16253 ( .A(n14519), .ZN(n14520) );
  OAI21_X1 U16254 ( .B1(n14521), .B2(n14534), .A(n14520), .ZN(P1_U3324) );
  OAI222_X1 U16255 ( .A1(P1_U3086), .A2(n14524), .B1(n14534), .B2(n14523), 
        .C1(n14522), .C2(n14528), .ZN(P1_U3328) );
  OAI222_X1 U16256 ( .A1(n14527), .A2(P1_U3086), .B1(n14534), .B2(n14526), 
        .C1(n14525), .C2(n14528), .ZN(P1_U3329) );
  OAI222_X1 U16257 ( .A1(P1_U3086), .A2(n14531), .B1(n14534), .B2(n14530), 
        .C1(n14529), .C2(n14528), .ZN(P1_U3330) );
  OAI222_X1 U16258 ( .A1(n14535), .A2(P1_U3086), .B1(n14534), .B2(n14533), 
        .C1(n14532), .C2(n14528), .ZN(P1_U3331) );
  MUX2_X1 U16259 ( .A(n14537), .B(n14536), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16260 ( .A(n14538), .ZN(n14539) );
  MUX2_X1 U16261 ( .A(n14539), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U16262 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14540), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16263 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14541) );
  OAI21_X1 U16264 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14541), 
        .ZN(U28) );
  AOI21_X1 U16265 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14542) );
  OAI21_X1 U16266 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14542), 
        .ZN(U29) );
  OAI21_X1 U16267 ( .B1(n14545), .B2(n14544), .A(n14543), .ZN(n14546) );
  XNOR2_X1 U16268 ( .A(n14546), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  XOR2_X1 U16269 ( .A(n14548), .B(n14547), .Z(SUB_1596_U57) );
  XNOR2_X1 U16270 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14549), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16271 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14550), .Z(SUB_1596_U54) );
  XOR2_X1 U16272 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14551), .Z(SUB_1596_U70)
         );
  OAI21_X1 U16273 ( .B1(n14554), .B2(n14553), .A(n14552), .ZN(n14555) );
  XNOR2_X1 U16274 ( .A(n14555), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  AOI21_X1 U16275 ( .B1(n14558), .B2(n14557), .A(n14556), .ZN(n14574) );
  OAI22_X1 U16276 ( .A1(n14560), .A2(n14967), .B1(n14966), .B2(n14559), .ZN(
        n14571) );
  AOI21_X1 U16277 ( .B1(n14563), .B2(n14562), .A(n14561), .ZN(n14569) );
  NOR2_X1 U16278 ( .A1(n14565), .A2(n14564), .ZN(n14566) );
  OAI21_X1 U16279 ( .B1(n14567), .B2(n14566), .A(n14936), .ZN(n14568) );
  OAI21_X1 U16280 ( .B1(n14569), .B2(n14977), .A(n14568), .ZN(n14570) );
  NOR3_X1 U16281 ( .A1(n14572), .A2(n14571), .A3(n14570), .ZN(n14573) );
  OAI21_X1 U16282 ( .B1(n14574), .B2(n14983), .A(n14573), .ZN(P3_U3197) );
  XNOR2_X1 U16283 ( .A(n14575), .B(n14583), .ZN(n14578) );
  AOI222_X1 U16284 ( .A1(n14991), .A2(n14578), .B1(n14577), .B2(n14988), .C1(
        n14576), .C2(n14987), .ZN(n14607) );
  OAI22_X1 U16285 ( .A1(n15002), .A2(n11417), .B1(n14580), .B2(n14579), .ZN(
        n14581) );
  INV_X1 U16286 ( .A(n14581), .ZN(n14588) );
  OAI21_X1 U16287 ( .B1(n14584), .B2(n14583), .A(n14582), .ZN(n14610) );
  INV_X1 U16288 ( .A(n14585), .ZN(n14586) );
  NOR2_X1 U16289 ( .A1(n14586), .A2(n15026), .ZN(n14609) );
  AOI22_X1 U16290 ( .A1(n14610), .A2(n14599), .B1(n14598), .B2(n14609), .ZN(
        n14587) );
  OAI211_X1 U16291 ( .C1(n15004), .C2(n14607), .A(n14588), .B(n14587), .ZN(
        P3_U3221) );
  XNOR2_X1 U16292 ( .A(n14589), .B(n14595), .ZN(n14592) );
  AOI222_X1 U16293 ( .A1(n14991), .A2(n14592), .B1(n14591), .B2(n14988), .C1(
        n14590), .C2(n14987), .ZN(n14611) );
  AOI22_X1 U16294 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n15004), .B1(n14998), 
        .B2(n14593), .ZN(n14601) );
  OAI21_X1 U16295 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(n14614) );
  NOR2_X1 U16296 ( .A1(n14597), .A2(n15026), .ZN(n14613) );
  AOI22_X1 U16297 ( .A1(n14614), .A2(n14599), .B1(n14598), .B2(n14613), .ZN(
        n14600) );
  OAI211_X1 U16298 ( .C1(n15004), .C2(n14611), .A(n14601), .B(n14600), .ZN(
        P3_U3222) );
  OAI22_X1 U16299 ( .A1(n14604), .A2(n14603), .B1(n14602), .B2(n15026), .ZN(
        n14605) );
  NOR2_X1 U16300 ( .A1(n14606), .A2(n14605), .ZN(n14615) );
  AOI22_X1 U16301 ( .A1(n15051), .A2(n14615), .B1(n14971), .B2(n15049), .ZN(
        P3_U3472) );
  INV_X1 U16302 ( .A(n14607), .ZN(n14608) );
  AOI211_X1 U16303 ( .C1(n15032), .C2(n14610), .A(n14609), .B(n14608), .ZN(
        n14617) );
  AOI22_X1 U16304 ( .A1(n15051), .A2(n14617), .B1(n11405), .B2(n15049), .ZN(
        P3_U3471) );
  INV_X1 U16305 ( .A(n14611), .ZN(n14612) );
  AOI211_X1 U16306 ( .C1(n15032), .C2(n14614), .A(n14613), .B(n14612), .ZN(
        n14619) );
  AOI22_X1 U16307 ( .A1(n15051), .A2(n14619), .B1(n11312), .B2(n15049), .ZN(
        P3_U3470) );
  INV_X1 U16308 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15073) );
  AOI22_X1 U16309 ( .A1(n15039), .A2(n14615), .B1(n15073), .B2(n15037), .ZN(
        P3_U3429) );
  INV_X1 U16310 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14616) );
  AOI22_X1 U16311 ( .A1(n15039), .A2(n14617), .B1(n14616), .B2(n15037), .ZN(
        P3_U3426) );
  INV_X1 U16312 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14618) );
  AOI22_X1 U16313 ( .A1(n15039), .A2(n14619), .B1(n14618), .B2(n15037), .ZN(
        P3_U3423) );
  NAND2_X1 U16314 ( .A1(n14620), .A2(n14889), .ZN(n14621) );
  AND2_X1 U16315 ( .A1(n14622), .A2(n14621), .ZN(n14626) );
  NAND2_X1 U16316 ( .A1(n14624), .A2(n14623), .ZN(n14625) );
  AND3_X1 U16317 ( .A1(n14627), .A2(n14626), .A3(n14625), .ZN(n14636) );
  AOI22_X1 U16318 ( .A1(n14922), .A2(n14636), .B1(n14628), .B2(n14920), .ZN(
        P2_U3513) );
  INV_X1 U16319 ( .A(n14629), .ZN(n14634) );
  INV_X1 U16320 ( .A(n14889), .ZN(n14907) );
  OAI21_X1 U16321 ( .B1(n14631), .B2(n14907), .A(n14630), .ZN(n14633) );
  AOI211_X1 U16322 ( .C1(n14901), .C2(n14634), .A(n14633), .B(n14632), .ZN(
        n14638) );
  AOI22_X1 U16323 ( .A1(n14922), .A2(n14638), .B1(n9213), .B2(n14920), .ZN(
        P2_U3511) );
  INV_X1 U16324 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14635) );
  AOI22_X1 U16325 ( .A1(n14915), .A2(n14636), .B1(n14635), .B2(n14913), .ZN(
        P2_U3472) );
  INV_X1 U16326 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14637) );
  AOI22_X1 U16327 ( .A1(n14915), .A2(n14638), .B1(n14637), .B2(n14913), .ZN(
        P2_U3466) );
  NAND2_X1 U16328 ( .A1(n14641), .A2(n14640), .ZN(n14642) );
  NAND2_X1 U16329 ( .A1(n14639), .A2(n14642), .ZN(n14644) );
  AOI222_X1 U16330 ( .A1(n14645), .A2(n14704), .B1(n14644), .B2(n14655), .C1(
        n14643), .C2(n14653), .ZN(n14647) );
  OAI211_X1 U16331 ( .C1(n14707), .C2(n14648), .A(n14647), .B(n14646), .ZN(
        P1_U3215) );
  AOI21_X1 U16332 ( .B1(n14651), .B2(n14650), .A(n14649), .ZN(n14652) );
  INV_X1 U16333 ( .A(n14652), .ZN(n14656) );
  AOI222_X1 U16334 ( .A1(n14657), .A2(n14704), .B1(n14656), .B2(n14655), .C1(
        n14654), .C2(n14653), .ZN(n14659) );
  OAI211_X1 U16335 ( .C1(n14707), .C2(n14660), .A(n14659), .B(n14658), .ZN(
        P1_U3226) );
  AOI211_X1 U16336 ( .C1(n14793), .C2(n14663), .A(n14662), .B(n14661), .ZN(
        n14664) );
  OAI21_X1 U16337 ( .B1(n14795), .B2(n14665), .A(n14664), .ZN(n14666) );
  AOI21_X1 U16338 ( .B1(n14667), .B2(n14799), .A(n14666), .ZN(n14674) );
  AOI22_X1 U16339 ( .A1(n14813), .A2(n14674), .B1(n8434), .B2(n14811), .ZN(
        P1_U3543) );
  OAI21_X1 U16340 ( .B1(n14669), .B2(n14775), .A(n14668), .ZN(n14671) );
  AOI211_X1 U16341 ( .C1(n14799), .C2(n14672), .A(n14671), .B(n14670), .ZN(
        n14676) );
  AOI22_X1 U16342 ( .A1(n14813), .A2(n14676), .B1(n10317), .B2(n14811), .ZN(
        P1_U3539) );
  INV_X1 U16343 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14673) );
  AOI22_X1 U16344 ( .A1(n14802), .A2(n14674), .B1(n14673), .B2(n14800), .ZN(
        P1_U3504) );
  INV_X1 U16345 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14675) );
  AOI22_X1 U16346 ( .A1(n14802), .A2(n14676), .B1(n14675), .B2(n14800), .ZN(
        P1_U3492) );
  XOR2_X1 U16347 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14677), .Z(SUB_1596_U69)
         );
  XNOR2_X1 U16348 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14678), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16349 ( .B1(n6463), .B2(n14680), .A(n14679), .ZN(n14682) );
  XNOR2_X1 U16350 ( .A(n14682), .B(n14681), .ZN(SUB_1596_U67) );
  AOI21_X1 U16351 ( .B1(n14685), .B2(n14684), .A(n14683), .ZN(n14686) );
  XOR2_X1 U16352 ( .A(n14686), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16353 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  XOR2_X1 U16354 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14689), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16355 ( .B1(n14691), .B2(n14690), .A(n6579), .ZN(n14693) );
  XNOR2_X1 U16356 ( .A(n14693), .B(n14692), .ZN(SUB_1596_U64) );
  NAND2_X1 U16357 ( .A1(n14793), .A2(n14694), .ZN(n14747) );
  INV_X1 U16358 ( .A(n14747), .ZN(n14696) );
  AOI21_X1 U16359 ( .B1(n14697), .B2(n14696), .A(n14695), .ZN(n14706) );
  AOI211_X1 U16360 ( .C1(n14701), .C2(n14700), .A(n14699), .B(n14698), .ZN(
        n14702) );
  AOI21_X1 U16361 ( .B1(n14704), .B2(n14703), .A(n14702), .ZN(n14705) );
  OAI211_X1 U16362 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14707), .A(n14706), .B(
        n14705), .ZN(P1_U3218) );
  NOR2_X1 U16363 ( .A1(n14708), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n14710) );
  OR2_X1 U16364 ( .A1(n14709), .A2(n14710), .ZN(n14713) );
  INV_X1 U16365 ( .A(n14710), .ZN(n14712) );
  MUX2_X1 U16366 ( .A(n14713), .B(n14712), .S(n14711), .Z(n14715) );
  NAND2_X1 U16367 ( .A1(n14715), .A2(n14714), .ZN(n14717) );
  AOI22_X1 U16368 ( .A1(n14733), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14716) );
  OAI21_X1 U16369 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(P1_U3243) );
  XNOR2_X1 U16370 ( .A(n14720), .B(n14719), .ZN(n14730) );
  NAND2_X1 U16371 ( .A1(n14722), .A2(n14721), .ZN(n14728) );
  OAI211_X1 U16372 ( .C1(n14726), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        n14727) );
  OAI211_X1 U16373 ( .C1(n14730), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        n14731) );
  AOI211_X1 U16374 ( .C1(P1_ADDR_REG_17__SCAN_IN), .C2(n14733), .A(n14732), 
        .B(n14731), .ZN(n14734) );
  INV_X1 U16375 ( .A(n14734), .ZN(P1_U3260) );
  AND2_X1 U16376 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14736), .ZN(P1_U3294) );
  AND2_X1 U16377 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14736), .ZN(P1_U3295) );
  AND2_X1 U16378 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14736), .ZN(P1_U3296) );
  AND2_X1 U16379 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14736), .ZN(P1_U3297) );
  AND2_X1 U16380 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14736), .ZN(P1_U3298) );
  AND2_X1 U16381 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14736), .ZN(P1_U3299) );
  AND2_X1 U16382 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14736), .ZN(P1_U3300) );
  AND2_X1 U16383 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14736), .ZN(P1_U3301) );
  AND2_X1 U16384 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14736), .ZN(P1_U3302) );
  AND2_X1 U16385 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14736), .ZN(P1_U3303) );
  AND2_X1 U16386 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14736), .ZN(P1_U3304) );
  AND2_X1 U16387 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14736), .ZN(P1_U3305) );
  AND2_X1 U16388 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14736), .ZN(P1_U3306) );
  AND2_X1 U16389 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14736), .ZN(P1_U3307) );
  AND2_X1 U16390 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14736), .ZN(P1_U3308) );
  AND2_X1 U16391 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14736), .ZN(P1_U3309) );
  AND2_X1 U16392 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14736), .ZN(P1_U3310) );
  INV_X1 U16393 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15126) );
  NOR2_X1 U16394 ( .A1(n14735), .A2(n15126), .ZN(P1_U3311) );
  INV_X1 U16395 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15181) );
  NOR2_X1 U16396 ( .A1(n14735), .A2(n15181), .ZN(P1_U3312) );
  AND2_X1 U16397 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14736), .ZN(P1_U3313) );
  AND2_X1 U16398 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14736), .ZN(P1_U3314) );
  AND2_X1 U16399 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14736), .ZN(P1_U3315) );
  AND2_X1 U16400 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14736), .ZN(P1_U3316) );
  AND2_X1 U16401 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14736), .ZN(P1_U3317) );
  AND2_X1 U16402 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14736), .ZN(P1_U3318) );
  AND2_X1 U16403 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14736), .ZN(P1_U3319) );
  AND2_X1 U16404 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14736), .ZN(P1_U3320) );
  AND2_X1 U16405 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14736), .ZN(P1_U3321) );
  AND2_X1 U16406 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14736), .ZN(P1_U3322) );
  AND2_X1 U16407 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14736), .ZN(P1_U3323) );
  AOI22_X1 U16408 ( .A1(n14802), .A2(n14737), .B1(n8073), .B2(n14800), .ZN(
        P1_U3459) );
  AOI22_X1 U16409 ( .A1(n14740), .A2(n14739), .B1(n14738), .B2(n14793), .ZN(
        n14742) );
  NAND2_X1 U16410 ( .A1(n14742), .A2(n14741), .ZN(n14743) );
  AOI21_X1 U16411 ( .B1(n14744), .B2(n14785), .A(n14743), .ZN(n14745) );
  AND2_X1 U16412 ( .A1(n14746), .A2(n14745), .ZN(n14804) );
  AOI22_X1 U16413 ( .A1(n14802), .A2(n14804), .B1(n8094), .B2(n14800), .ZN(
        P1_U3462) );
  NAND2_X1 U16414 ( .A1(n14748), .A2(n14747), .ZN(n14750) );
  AOI211_X1 U16415 ( .C1(n14785), .C2(n14751), .A(n14750), .B(n14749), .ZN(
        n14805) );
  AOI22_X1 U16416 ( .A1(n14802), .A2(n14805), .B1(n8152), .B2(n14800), .ZN(
        P1_U3468) );
  INV_X1 U16417 ( .A(n14752), .ZN(n14758) );
  NOR2_X1 U16418 ( .A1(n14754), .A2(n14753), .ZN(n14757) );
  NOR4_X1 U16419 ( .A1(n14758), .A2(n14757), .A3(n14756), .A4(n14755), .ZN(
        n14806) );
  INV_X1 U16420 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14759) );
  AOI22_X1 U16421 ( .A1(n14802), .A2(n14806), .B1(n14759), .B2(n14800), .ZN(
        P1_U3471) );
  OAI21_X1 U16422 ( .B1(n14761), .B2(n14775), .A(n14760), .ZN(n14763) );
  AOI211_X1 U16423 ( .C1(n14785), .C2(n14764), .A(n14763), .B(n14762), .ZN(
        n14807) );
  AOI22_X1 U16424 ( .A1(n14802), .A2(n14807), .B1(n8212), .B2(n14800), .ZN(
        P1_U3474) );
  AND2_X1 U16425 ( .A1(n14765), .A2(n14793), .ZN(n14766) );
  OR2_X1 U16426 ( .A1(n14767), .A2(n14766), .ZN(n14768) );
  AOI21_X1 U16427 ( .B1(n14769), .B2(n14785), .A(n14768), .ZN(n14770) );
  INV_X1 U16428 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14772) );
  AOI22_X1 U16429 ( .A1(n14802), .A2(n14808), .B1(n14772), .B2(n14800), .ZN(
        P1_U3477) );
  INV_X1 U16430 ( .A(n14773), .ZN(n14774) );
  OAI21_X1 U16431 ( .B1(n14776), .B2(n14775), .A(n14774), .ZN(n14777) );
  AOI21_X1 U16432 ( .B1(n14778), .B2(n14785), .A(n14777), .ZN(n14779) );
  INV_X1 U16433 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14781) );
  AOI22_X1 U16434 ( .A1(n14802), .A2(n14809), .B1(n14781), .B2(n14800), .ZN(
        P1_U3480) );
  INV_X1 U16435 ( .A(n14782), .ZN(n14784) );
  AOI211_X1 U16436 ( .C1(n14786), .C2(n14785), .A(n14784), .B(n14783), .ZN(
        n14787) );
  AND2_X1 U16437 ( .A1(n14788), .A2(n14787), .ZN(n14810) );
  INV_X1 U16438 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14789) );
  AOI22_X1 U16439 ( .A1(n14802), .A2(n14810), .B1(n14789), .B2(n14800), .ZN(
        P1_U3486) );
  AOI211_X1 U16440 ( .C1(n14793), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14794) );
  OAI21_X1 U16441 ( .B1(n14796), .B2(n14795), .A(n14794), .ZN(n14797) );
  AOI21_X1 U16442 ( .B1(n14799), .B2(n14798), .A(n14797), .ZN(n14812) );
  INV_X1 U16443 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U16444 ( .A1(n14802), .A2(n14812), .B1(n14801), .B2(n14800), .ZN(
        P1_U3489) );
  AOI22_X1 U16445 ( .A1(n14813), .A2(n14804), .B1(n14803), .B2(n14811), .ZN(
        P1_U3529) );
  AOI22_X1 U16446 ( .A1(n14813), .A2(n14805), .B1(n10024), .B2(n14811), .ZN(
        P1_U3531) );
  AOI22_X1 U16447 ( .A1(n14813), .A2(n14806), .B1(n8181), .B2(n14811), .ZN(
        P1_U3532) );
  AOI22_X1 U16448 ( .A1(n14813), .A2(n14807), .B1(n8211), .B2(n14811), .ZN(
        P1_U3533) );
  AOI22_X1 U16449 ( .A1(n14813), .A2(n14808), .B1(n14118), .B2(n14811), .ZN(
        P1_U3534) );
  AOI22_X1 U16450 ( .A1(n14813), .A2(n14809), .B1(n8248), .B2(n14811), .ZN(
        P1_U3535) );
  AOI22_X1 U16451 ( .A1(n14813), .A2(n14810), .B1(n10308), .B2(n14811), .ZN(
        P1_U3537) );
  AOI22_X1 U16452 ( .A1(n14813), .A2(n14812), .B1(n10310), .B2(n14811), .ZN(
        P1_U3538) );
  NOR2_X1 U16453 ( .A1(n14859), .A2(P2_U3947), .ZN(P2_U3087) );
  NAND2_X1 U16454 ( .A1(P2_U3088), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n14818) );
  OAI211_X1 U16455 ( .C1(n14816), .C2(n14815), .A(n14865), .B(n14814), .ZN(
        n14817) );
  OAI211_X1 U16456 ( .C1(n14820), .C2(n14819), .A(n14818), .B(n14817), .ZN(
        n14821) );
  INV_X1 U16457 ( .A(n14821), .ZN(n14826) );
  OAI211_X1 U16458 ( .C1(n14824), .C2(n14823), .A(n14868), .B(n14822), .ZN(
        n14825) );
  OAI211_X1 U16459 ( .C1(n14857), .C2(n14827), .A(n14826), .B(n14825), .ZN(
        P2_U3216) );
  INV_X1 U16460 ( .A(n14828), .ZN(n14829) );
  OAI211_X1 U16461 ( .C1(n14831), .C2(n14830), .A(n14829), .B(n14865), .ZN(
        n14834) );
  INV_X1 U16462 ( .A(n14832), .ZN(n14833) );
  OAI211_X1 U16463 ( .C1(n14836), .C2(n14835), .A(n14834), .B(n14833), .ZN(
        n14837) );
  INV_X1 U16464 ( .A(n14837), .ZN(n14842) );
  OAI211_X1 U16465 ( .C1(n14840), .C2(n14839), .A(n14838), .B(n14868), .ZN(
        n14841) );
  OAI211_X1 U16466 ( .C1(n14857), .C2(n7130), .A(n14842), .B(n14841), .ZN(
        P2_U3221) );
  INV_X1 U16467 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14858) );
  OAI21_X1 U16468 ( .B1(n14845), .B2(n14844), .A(n14843), .ZN(n14854) );
  INV_X1 U16469 ( .A(n14846), .ZN(n14851) );
  OAI21_X1 U16470 ( .B1(n14849), .B2(n14848), .A(n14847), .ZN(n14850) );
  NAND2_X1 U16471 ( .A1(n14851), .A2(n14850), .ZN(n14852) );
  AOI222_X1 U16472 ( .A1(n14854), .A2(n14868), .B1(n14853), .B2(n14863), .C1(
        n14852), .C2(n14865), .ZN(n14856) );
  OAI211_X1 U16473 ( .C1(n14858), .C2(n14857), .A(n14856), .B(n14855), .ZN(
        P2_U3223) );
  AOI22_X1 U16474 ( .A1(n14859), .A2(P2_ADDR_REG_18__SCAN_IN), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(P2_U3088), .ZN(n14872) );
  OAI21_X1 U16475 ( .B1(n14862), .B2(n14861), .A(n14860), .ZN(n14866) );
  AOI22_X1 U16476 ( .A1(n14866), .A2(n14865), .B1(n14864), .B2(n14863), .ZN(
        n14871) );
  OAI211_X1 U16477 ( .C1(n14869), .C2(P2_REG1_REG_18__SCAN_IN), .A(n14868), 
        .B(n14867), .ZN(n14870) );
  NAND3_X1 U16478 ( .A1(n14872), .A2(n14871), .A3(n14870), .ZN(P2_U3232) );
  AND2_X1 U16479 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14875), .ZN(P2_U3266) );
  AND2_X1 U16480 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14875), .ZN(P2_U3267) );
  AND2_X1 U16481 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14875), .ZN(P2_U3268) );
  AND2_X1 U16482 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14875), .ZN(P2_U3269) );
  AND2_X1 U16483 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14875), .ZN(P2_U3270) );
  AND2_X1 U16484 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14875), .ZN(P2_U3271) );
  AND2_X1 U16485 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14875), .ZN(P2_U3272) );
  AND2_X1 U16486 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14875), .ZN(P2_U3273) );
  AND2_X1 U16487 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14875), .ZN(P2_U3274) );
  INV_X1 U16488 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15071) );
  NOR2_X1 U16489 ( .A1(n14874), .A2(n15071), .ZN(P2_U3275) );
  AND2_X1 U16490 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14875), .ZN(P2_U3276) );
  AND2_X1 U16491 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14875), .ZN(P2_U3277) );
  AND2_X1 U16492 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14875), .ZN(P2_U3278) );
  AND2_X1 U16493 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14875), .ZN(P2_U3279) );
  AND2_X1 U16494 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14875), .ZN(P2_U3280) );
  AND2_X1 U16495 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14875), .ZN(P2_U3281) );
  AND2_X1 U16496 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14875), .ZN(P2_U3282) );
  INV_X1 U16497 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15058) );
  NOR2_X1 U16498 ( .A1(n14874), .A2(n15058), .ZN(P2_U3283) );
  AND2_X1 U16499 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14875), .ZN(P2_U3284) );
  AND2_X1 U16500 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14875), .ZN(P2_U3285) );
  INV_X1 U16501 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15102) );
  NOR2_X1 U16502 ( .A1(n14874), .A2(n15102), .ZN(P2_U3286) );
  AND2_X1 U16503 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14875), .ZN(P2_U3287) );
  AND2_X1 U16504 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14875), .ZN(P2_U3288) );
  AND2_X1 U16505 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14875), .ZN(P2_U3289) );
  AND2_X1 U16506 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14875), .ZN(P2_U3290) );
  AND2_X1 U16507 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14875), .ZN(P2_U3291) );
  AND2_X1 U16508 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14875), .ZN(P2_U3292) );
  AND2_X1 U16509 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14875), .ZN(P2_U3293) );
  AND2_X1 U16510 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14875), .ZN(P2_U3294) );
  AND2_X1 U16511 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14875), .ZN(P2_U3295) );
  AOI22_X1 U16512 ( .A1(n14881), .A2(n14877), .B1(n14876), .B2(n14878), .ZN(
        P2_U3416) );
  AOI22_X1 U16513 ( .A1(n14881), .A2(n14880), .B1(n14879), .B2(n14878), .ZN(
        P2_U3417) );
  INV_X1 U16514 ( .A(n14882), .ZN(n14885) );
  AOI211_X1 U16515 ( .C1(n14885), .C2(n14901), .A(n14884), .B(n14883), .ZN(
        n14917) );
  INV_X1 U16516 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14886) );
  AOI22_X1 U16517 ( .A1(n14915), .A2(n14917), .B1(n14886), .B2(n14913), .ZN(
        P2_U3430) );
  AOI21_X1 U16518 ( .B1(n14889), .B2(n14888), .A(n14887), .ZN(n14890) );
  OAI211_X1 U16519 ( .C1(n14892), .C2(n14903), .A(n14891), .B(n14890), .ZN(
        n14893) );
  INV_X1 U16520 ( .A(n14893), .ZN(n14918) );
  INV_X1 U16521 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14894) );
  AOI22_X1 U16522 ( .A1(n14915), .A2(n14918), .B1(n14894), .B2(n14913), .ZN(
        P2_U3448) );
  INV_X1 U16523 ( .A(n14895), .ZN(n14900) );
  OAI21_X1 U16524 ( .B1(n14897), .B2(n14907), .A(n14896), .ZN(n14899) );
  AOI211_X1 U16525 ( .C1(n14901), .C2(n14900), .A(n14899), .B(n14898), .ZN(
        n14919) );
  INV_X1 U16526 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14902) );
  AOI22_X1 U16527 ( .A1(n14915), .A2(n14919), .B1(n14902), .B2(n14913), .ZN(
        P2_U3454) );
  NOR2_X1 U16528 ( .A1(n14904), .A2(n14903), .ZN(n14910) );
  OAI211_X1 U16529 ( .C1(n14908), .C2(n14907), .A(n14906), .B(n14905), .ZN(
        n14909) );
  AOI211_X1 U16530 ( .C1(n14912), .C2(n14911), .A(n14910), .B(n14909), .ZN(
        n14921) );
  INV_X1 U16531 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14914) );
  AOI22_X1 U16532 ( .A1(n14915), .A2(n14921), .B1(n14914), .B2(n14913), .ZN(
        P2_U3463) );
  AOI22_X1 U16533 ( .A1(n14922), .A2(n14917), .B1(n14916), .B2(n14920), .ZN(
        P2_U3499) );
  AOI22_X1 U16534 ( .A1(n14922), .A2(n14918), .B1(n10000), .B2(n14920), .ZN(
        P2_U3505) );
  AOI22_X1 U16535 ( .A1(n14922), .A2(n14919), .B1(n9142), .B2(n14920), .ZN(
        P2_U3507) );
  AOI22_X1 U16536 ( .A1(n14922), .A2(n14921), .B1(n9193), .B2(n14920), .ZN(
        P2_U3510) );
  NOR2_X1 U16537 ( .A1(P3_U3897), .A2(n14923), .ZN(P3_U3150) );
  INV_X1 U16538 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14940) );
  OAI21_X1 U16539 ( .B1(n14926), .B2(n14925), .A(n14924), .ZN(n14937) );
  AOI21_X1 U16540 ( .B1(n14929), .B2(n14928), .A(n14927), .ZN(n14930) );
  NOR2_X1 U16541 ( .A1(n14930), .A2(n14983), .ZN(n14935) );
  AOI21_X1 U16542 ( .B1(n14931), .B2(n15044), .A(n6602), .ZN(n14933) );
  OAI22_X1 U16543 ( .A1(n14933), .A2(n14977), .B1(n14932), .B2(n14966), .ZN(
        n14934) );
  AOI211_X1 U16544 ( .C1(n14937), .C2(n14936), .A(n14935), .B(n14934), .ZN(
        n14939) );
  OAI211_X1 U16545 ( .C1(n14940), .C2(n14967), .A(n14939), .B(n14938), .ZN(
        P3_U3189) );
  AOI21_X1 U16546 ( .B1(n14943), .B2(n14942), .A(n14941), .ZN(n14961) );
  INV_X1 U16547 ( .A(n14944), .ZN(n14953) );
  OAI21_X1 U16548 ( .B1(n14967), .B2(n14946), .A(n14945), .ZN(n14952) );
  NAND2_X1 U16549 ( .A1(n14948), .A2(n14947), .ZN(n14949) );
  AOI21_X1 U16550 ( .B1(n14950), .B2(n14949), .A(n14977), .ZN(n14951) );
  AOI211_X1 U16551 ( .C1(n14954), .C2(n14953), .A(n14952), .B(n14951), .ZN(
        n14960) );
  AOI21_X1 U16552 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n14958) );
  OR2_X1 U16553 ( .A1(n14958), .A2(n14975), .ZN(n14959) );
  OAI211_X1 U16554 ( .C1(n14961), .C2(n14983), .A(n14960), .B(n14959), .ZN(
        P3_U3192) );
  AOI21_X1 U16555 ( .B1(n14964), .B2(n14963), .A(n14962), .ZN(n14984) );
  OAI22_X1 U16556 ( .A1(n14968), .A2(n14967), .B1(n14966), .B2(n14965), .ZN(
        n14980) );
  AOI21_X1 U16557 ( .B1(n14971), .B2(n14970), .A(n14969), .ZN(n14978) );
  AOI21_X1 U16558 ( .B1(n14974), .B2(n14973), .A(n14972), .ZN(n14976) );
  OAI22_X1 U16559 ( .A1(n14978), .A2(n14977), .B1(n14976), .B2(n14975), .ZN(
        n14979) );
  NOR3_X1 U16560 ( .A1(n14981), .A2(n14980), .A3(n14979), .ZN(n14982) );
  OAI21_X1 U16561 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(P3_U3195) );
  NOR2_X1 U16562 ( .A1(n7939), .A2(n15026), .ZN(n15006) );
  XNOR2_X1 U16563 ( .A(n14985), .B(n6779), .ZN(n14997) );
  AOI22_X1 U16564 ( .A1(n14989), .A2(n14988), .B1(n14987), .B2(n6657), .ZN(
        n14994) );
  XNOR2_X1 U16565 ( .A(n14990), .B(n6779), .ZN(n14992) );
  NAND2_X1 U16566 ( .A1(n14992), .A2(n14991), .ZN(n14993) );
  OAI211_X1 U16567 ( .C1(n14997), .C2(n14995), .A(n14994), .B(n14993), .ZN(
        n15005) );
  AOI21_X1 U16568 ( .B1(n15006), .B2(n14996), .A(n15005), .ZN(n15003) );
  INV_X1 U16569 ( .A(n14997), .ZN(n15007) );
  AOI22_X1 U16570 ( .A1(n15007), .A2(n14999), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n14998), .ZN(n15000) );
  OAI221_X1 U16571 ( .B1(n15004), .B2(n15003), .C1(n15002), .C2(n15001), .A(
        n15000), .ZN(P3_U3232) );
  AOI211_X1 U16572 ( .C1(n15023), .C2(n15007), .A(n15006), .B(n15005), .ZN(
        n15041) );
  INV_X1 U16573 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U16574 ( .A1(n15039), .A2(n15041), .B1(n15008), .B2(n15037), .ZN(
        P3_U3393) );
  INV_X1 U16575 ( .A(n15009), .ZN(n15011) );
  AOI211_X1 U16576 ( .C1(n15023), .C2(n15012), .A(n15011), .B(n15010), .ZN(
        n15043) );
  INV_X1 U16577 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U16578 ( .A1(n15039), .A2(n15043), .B1(n15013), .B2(n15037), .ZN(
        P3_U3396) );
  AOI22_X1 U16579 ( .A1(n15016), .A2(n15032), .B1(n15015), .B2(n15014), .ZN(
        n15017) );
  AND2_X1 U16580 ( .A1(n15018), .A2(n15017), .ZN(n15045) );
  INV_X1 U16581 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U16582 ( .A1(n15039), .A2(n15045), .B1(n15115), .B2(n15037), .ZN(
        P3_U3411) );
  INV_X1 U16583 ( .A(n15019), .ZN(n15022) );
  AOI211_X1 U16584 ( .C1(n15022), .C2(n15023), .A(n15021), .B(n15020), .ZN(
        n15046) );
  INV_X1 U16585 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15182) );
  AOI22_X1 U16586 ( .A1(n15039), .A2(n15046), .B1(n15182), .B2(n15037), .ZN(
        P3_U3414) );
  NAND2_X1 U16587 ( .A1(n15030), .A2(n15023), .ZN(n15024) );
  OAI211_X1 U16588 ( .C1(n15027), .C2(n15026), .A(n15025), .B(n15024), .ZN(
        n15028) );
  AOI21_X1 U16589 ( .B1(n15030), .B2(n15029), .A(n15028), .ZN(n15048) );
  INV_X1 U16590 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15031) );
  AOI22_X1 U16591 ( .A1(n15039), .A2(n15048), .B1(n15031), .B2(n15037), .ZN(
        P3_U3417) );
  NAND2_X1 U16592 ( .A1(n15033), .A2(n15032), .ZN(n15034) );
  INV_X1 U16593 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15038) );
  AOI22_X1 U16594 ( .A1(n15039), .A2(n15050), .B1(n15038), .B2(n15037), .ZN(
        P3_U3420) );
  AOI22_X1 U16595 ( .A1(n15051), .A2(n15041), .B1(n15040), .B2(n15049), .ZN(
        P3_U3460) );
  AOI22_X1 U16596 ( .A1(n15051), .A2(n15043), .B1(n15042), .B2(n15049), .ZN(
        P3_U3461) );
  AOI22_X1 U16597 ( .A1(n15051), .A2(n15045), .B1(n15044), .B2(n15049), .ZN(
        P3_U3466) );
  AOI22_X1 U16598 ( .A1(n15051), .A2(n15046), .B1(n10532), .B2(n15049), .ZN(
        P3_U3467) );
  AOI22_X1 U16599 ( .A1(n15051), .A2(n15048), .B1(n15047), .B2(n15049), .ZN(
        P3_U3468) );
  AOI22_X1 U16600 ( .A1(n15051), .A2(n15050), .B1(n11333), .B2(n15049), .ZN(
        P3_U3469) );
  OAI22_X1 U16601 ( .A1(n15054), .A2(keyinput37), .B1(n15053), .B2(keyinput11), 
        .ZN(n15052) );
  AOI221_X1 U16602 ( .B1(n15054), .B2(keyinput37), .C1(keyinput11), .C2(n15053), .A(n15052), .ZN(n15065) );
  OAI22_X1 U16603 ( .A1(n7559), .A2(keyinput29), .B1(n15056), .B2(keyinput60), 
        .ZN(n15055) );
  AOI221_X1 U16604 ( .B1(n7559), .B2(keyinput29), .C1(keyinput60), .C2(n15056), 
        .A(n15055), .ZN(n15064) );
  OAI22_X1 U16605 ( .A1(n15058), .A2(keyinput27), .B1(n10047), .B2(keyinput47), 
        .ZN(n15057) );
  AOI221_X1 U16606 ( .B1(n15058), .B2(keyinput27), .C1(keyinput47), .C2(n10047), .A(n15057), .ZN(n15063) );
  INV_X1 U16607 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n15061) );
  OAI22_X1 U16608 ( .A1(n15061), .A2(keyinput33), .B1(n15060), .B2(keyinput48), 
        .ZN(n15059) );
  AOI221_X1 U16609 ( .B1(n15061), .B2(keyinput33), .C1(keyinput48), .C2(n15060), .A(n15059), .ZN(n15062) );
  NAND4_X1 U16610 ( .A1(n15065), .A2(n15064), .A3(n15063), .A4(n15062), .ZN(
        n15198) );
  OAI22_X1 U16611 ( .A1(n15067), .A2(keyinput56), .B1(n12895), .B2(keyinput23), 
        .ZN(n15066) );
  AOI221_X1 U16612 ( .B1(n15067), .B2(keyinput56), .C1(keyinput23), .C2(n12895), .A(n15066), .ZN(n15078) );
  OAI22_X1 U16613 ( .A1(n12885), .A2(keyinput10), .B1(n6955), .B2(keyinput40), 
        .ZN(n15068) );
  AOI221_X1 U16614 ( .B1(n12885), .B2(keyinput10), .C1(keyinput40), .C2(n6955), 
        .A(n15068), .ZN(n15077) );
  OAI22_X1 U16615 ( .A1(n15071), .A2(keyinput14), .B1(n15070), .B2(keyinput30), 
        .ZN(n15069) );
  AOI221_X1 U16616 ( .B1(n15071), .B2(keyinput14), .C1(keyinput30), .C2(n15070), .A(n15069), .ZN(n15076) );
  OAI22_X1 U16617 ( .A1(n15074), .A2(keyinput4), .B1(n15073), .B2(keyinput51), 
        .ZN(n15072) );
  AOI221_X1 U16618 ( .B1(n15074), .B2(keyinput4), .C1(keyinput51), .C2(n15073), 
        .A(n15072), .ZN(n15075) );
  NAND4_X1 U16619 ( .A1(n15078), .A2(n15077), .A3(n15076), .A4(n15075), .ZN(
        n15197) );
  INV_X1 U16620 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15081) );
  INV_X1 U16621 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n15080) );
  AOI22_X1 U16622 ( .A1(n15081), .A2(keyinput62), .B1(n15080), .B2(keyinput2), 
        .ZN(n15079) );
  OAI221_X1 U16623 ( .B1(n15081), .B2(keyinput62), .C1(n15080), .C2(keyinput2), 
        .A(n15079), .ZN(n15093) );
  INV_X1 U16624 ( .A(keyinput19), .ZN(n15083) );
  AOI22_X1 U16625 ( .A1(n15084), .A2(keyinput58), .B1(P3_DATAO_REG_3__SCAN_IN), 
        .B2(n15083), .ZN(n15082) );
  OAI221_X1 U16626 ( .B1(n15084), .B2(keyinput58), .C1(n15083), .C2(
        P3_DATAO_REG_3__SCAN_IN), .A(n15082), .ZN(n15092) );
  INV_X1 U16627 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15087) );
  INV_X1 U16628 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n15086) );
  AOI22_X1 U16629 ( .A1(n15087), .A2(keyinput43), .B1(n15086), .B2(keyinput15), 
        .ZN(n15085) );
  OAI221_X1 U16630 ( .B1(n15087), .B2(keyinput43), .C1(n15086), .C2(keyinput15), .A(n15085), .ZN(n15091) );
  XNOR2_X1 U16631 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput24), .ZN(n15089) );
  XNOR2_X1 U16632 ( .A(keyinput5), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U16633 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  NOR4_X1 U16634 ( .A1(n15093), .A2(n15092), .A3(n15091), .A4(n15090), .ZN(
        n15140) );
  AOI22_X1 U16635 ( .A1(n15095), .A2(keyinput0), .B1(keyinput31), .B2(n9884), 
        .ZN(n15094) );
  OAI221_X1 U16636 ( .B1(n15095), .B2(keyinput0), .C1(n9884), .C2(keyinput31), 
        .A(n15094), .ZN(n15106) );
  AOI22_X1 U16637 ( .A1(n15098), .A2(keyinput7), .B1(n15097), .B2(keyinput13), 
        .ZN(n15096) );
  OAI221_X1 U16638 ( .B1(n15098), .B2(keyinput7), .C1(n15097), .C2(keyinput13), 
        .A(n15096), .ZN(n15105) );
  XNOR2_X1 U16639 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput55), .ZN(n15101)
         );
  XNOR2_X1 U16640 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput49), .ZN(n15100) );
  XNOR2_X1 U16641 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput45), .ZN(n15099) );
  NAND3_X1 U16642 ( .A1(n15101), .A2(n15100), .A3(n15099), .ZN(n15104) );
  XNOR2_X1 U16643 ( .A(n15102), .B(keyinput35), .ZN(n15103) );
  NOR4_X1 U16644 ( .A1(n15106), .A2(n15105), .A3(n15104), .A4(n15103), .ZN(
        n15139) );
  INV_X1 U16645 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U16646 ( .A1(n15109), .A2(keyinput21), .B1(keyinput8), .B2(n15108), 
        .ZN(n15107) );
  OAI221_X1 U16647 ( .B1(n15109), .B2(keyinput21), .C1(n15108), .C2(keyinput8), 
        .A(n15107), .ZN(n15121) );
  AOI22_X1 U16648 ( .A1(n10992), .A2(keyinput12), .B1(n15111), .B2(keyinput28), 
        .ZN(n15110) );
  OAI221_X1 U16649 ( .B1(n10992), .B2(keyinput12), .C1(n15111), .C2(keyinput28), .A(n15110), .ZN(n15120) );
  INV_X1 U16650 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U16651 ( .A1(n15114), .A2(keyinput63), .B1(n15113), .B2(keyinput20), 
        .ZN(n15112) );
  OAI221_X1 U16652 ( .B1(n15114), .B2(keyinput63), .C1(n15113), .C2(keyinput20), .A(n15112), .ZN(n15119) );
  XOR2_X1 U16653 ( .A(n15115), .B(keyinput54), .Z(n15117) );
  XNOR2_X1 U16654 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput18), .ZN(n15116) );
  NAND2_X1 U16655 ( .A1(n15117), .A2(n15116), .ZN(n15118) );
  NOR4_X1 U16656 ( .A1(n15121), .A2(n15120), .A3(n15119), .A4(n15118), .ZN(
        n15138) );
  AOI22_X1 U16657 ( .A1(n15124), .A2(keyinput16), .B1(keyinput6), .B2(n15123), 
        .ZN(n15122) );
  OAI221_X1 U16658 ( .B1(n15124), .B2(keyinput16), .C1(n15123), .C2(keyinput6), 
        .A(n15122), .ZN(n15136) );
  AOI22_X1 U16659 ( .A1(n15127), .A2(keyinput1), .B1(n15126), .B2(keyinput36), 
        .ZN(n15125) );
  OAI221_X1 U16660 ( .B1(n15127), .B2(keyinput1), .C1(n15126), .C2(keyinput36), 
        .A(n15125), .ZN(n15135) );
  AOI22_X1 U16661 ( .A1(n15129), .A2(keyinput57), .B1(keyinput39), .B2(n12824), 
        .ZN(n15128) );
  OAI221_X1 U16662 ( .B1(n15129), .B2(keyinput57), .C1(n12824), .C2(keyinput39), .A(n15128), .ZN(n15134) );
  AOI22_X1 U16663 ( .A1(n15132), .A2(keyinput41), .B1(keyinput26), .B2(n15131), 
        .ZN(n15130) );
  OAI221_X1 U16664 ( .B1(n15132), .B2(keyinput41), .C1(n15131), .C2(keyinput26), .A(n15130), .ZN(n15133) );
  NOR4_X1 U16665 ( .A1(n15136), .A2(n15135), .A3(n15134), .A4(n15133), .ZN(
        n15137) );
  NAND4_X1 U16666 ( .A1(n15140), .A2(n15139), .A3(n15138), .A4(n15137), .ZN(
        n15196) );
  NOR4_X1 U16667 ( .A1(keyinput9), .A2(keyinput29), .A3(keyinput25), .A4(
        keyinput37), .ZN(n15144) );
  NOR4_X1 U16668 ( .A1(keyinput33), .A2(keyinput53), .A3(keyinput61), .A4(
        keyinput60), .ZN(n15143) );
  NOR4_X1 U16669 ( .A1(keyinput48), .A2(keyinput56), .A3(keyinput32), .A4(
        keyinput42), .ZN(n15142) );
  NOR4_X1 U16670 ( .A1(keyinput46), .A2(keyinput38), .A3(keyinput50), .A4(
        keyinput10), .ZN(n15141) );
  NAND4_X1 U16671 ( .A1(n15144), .A2(n15143), .A3(n15142), .A4(n15141), .ZN(
        n15194) );
  NAND3_X1 U16672 ( .A1(keyinput43), .A2(keyinput15), .A3(keyinput2), .ZN(
        n15146) );
  NAND3_X1 U16673 ( .A1(keyinput31), .A2(keyinput35), .A3(keyinput49), .ZN(
        n15145) );
  NOR4_X1 U16674 ( .A1(keyinput62), .A2(keyinput0), .A3(n15146), .A4(n15145), 
        .ZN(n15164) );
  NAND2_X1 U16675 ( .A1(keyinput19), .A2(keyinput24), .ZN(n15149) );
  NOR2_X1 U16676 ( .A1(keyinput13), .A2(keyinput45), .ZN(n15147) );
  NAND3_X1 U16677 ( .A1(keyinput7), .A2(keyinput55), .A3(n15147), .ZN(n15148)
         );
  NOR4_X1 U16678 ( .A1(keyinput58), .A2(keyinput5), .A3(n15149), .A4(n15148), 
        .ZN(n15163) );
  NAND3_X1 U16679 ( .A1(keyinput54), .A2(keyinput18), .A3(keyinput63), .ZN(
        n15155) );
  NOR2_X1 U16680 ( .A1(keyinput16), .A2(keyinput6), .ZN(n15150) );
  NAND3_X1 U16681 ( .A1(keyinput1), .A2(keyinput36), .A3(n15150), .ZN(n15154)
         );
  NOR3_X1 U16682 ( .A1(keyinput12), .A2(keyinput28), .A3(keyinput21), .ZN(
        n15152) );
  NOR3_X1 U16683 ( .A1(keyinput57), .A2(keyinput41), .A3(keyinput26), .ZN(
        n15151) );
  NAND4_X1 U16684 ( .A1(keyinput8), .A2(n15152), .A3(keyinput39), .A4(n15151), 
        .ZN(n15153) );
  NOR4_X1 U16685 ( .A1(keyinput20), .A2(n15155), .A3(n15154), .A4(n15153), 
        .ZN(n15162) );
  NOR2_X1 U16686 ( .A1(keyinput3), .A2(keyinput27), .ZN(n15156) );
  NAND3_X1 U16687 ( .A1(keyinput17), .A2(keyinput4), .A3(n15156), .ZN(n15160)
         );
  NAND4_X1 U16688 ( .A1(keyinput40), .A2(keyinput52), .A3(keyinput44), .A4(
        keyinput47), .ZN(n15159) );
  NAND4_X1 U16689 ( .A1(keyinput34), .A2(keyinput59), .A3(keyinput51), .A4(
        keyinput11), .ZN(n15158) );
  NAND4_X1 U16690 ( .A1(keyinput14), .A2(keyinput30), .A3(keyinput23), .A4(
        keyinput22), .ZN(n15157) );
  NOR4_X1 U16691 ( .A1(n15160), .A2(n15159), .A3(n15158), .A4(n15157), .ZN(
        n15161) );
  NAND4_X1 U16692 ( .A1(n15164), .A2(n15163), .A3(n15162), .A4(n15161), .ZN(
        n15193) );
  AOI22_X1 U16693 ( .A1(n11309), .A2(keyinput52), .B1(keyinput59), .B2(n13130), 
        .ZN(n15165) );
  OAI221_X1 U16694 ( .B1(n11309), .B2(keyinput52), .C1(n13130), .C2(keyinput59), .A(n15165), .ZN(n15176) );
  INV_X1 U16695 ( .A(keyinput53), .ZN(n15167) );
  AOI22_X1 U16696 ( .A1(n15168), .A2(keyinput25), .B1(P3_DATAO_REG_16__SCAN_IN), .B2(n15167), .ZN(n15166) );
  OAI221_X1 U16697 ( .B1(n15168), .B2(keyinput25), .C1(n15167), .C2(
        P3_DATAO_REG_16__SCAN_IN), .A(n15166), .ZN(n15175) );
  XOR2_X1 U16698 ( .A(n9391), .B(keyinput32), .Z(n15171) );
  XNOR2_X1 U16699 ( .A(P3_IR_REG_20__SCAN_IN), .B(keyinput22), .ZN(n15170) );
  XNOR2_X1 U16700 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput61), .ZN(n15169) );
  NAND3_X1 U16701 ( .A1(n15171), .A2(n15170), .A3(n15169), .ZN(n15174) );
  XNOR2_X1 U16702 ( .A(n15172), .B(keyinput3), .ZN(n15173) );
  NOR4_X1 U16703 ( .A1(n15176), .A2(n15175), .A3(n15174), .A4(n15173), .ZN(
        n15192) );
  AOI22_X1 U16704 ( .A1(P2_U3088), .A2(keyinput50), .B1(keyinput44), .B2(
        n15178), .ZN(n15177) );
  OAI221_X1 U16705 ( .B1(P2_U3088), .B2(keyinput50), .C1(n15178), .C2(
        keyinput44), .A(n15177), .ZN(n15190) );
  AOI22_X1 U16706 ( .A1(n15181), .A2(keyinput38), .B1(n15180), .B2(keyinput34), 
        .ZN(n15179) );
  OAI221_X1 U16707 ( .B1(n15181), .B2(keyinput38), .C1(n15180), .C2(keyinput34), .A(n15179), .ZN(n15189) );
  XOR2_X1 U16708 ( .A(n15182), .B(keyinput46), .Z(n15185) );
  XNOR2_X1 U16709 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput9), .ZN(n15184) );
  XNOR2_X1 U16710 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput42), .ZN(n15183) );
  NAND3_X1 U16711 ( .A1(n15185), .A2(n15184), .A3(n15183), .ZN(n15188) );
  XNOR2_X1 U16712 ( .A(n15186), .B(keyinput17), .ZN(n15187) );
  NOR4_X1 U16713 ( .A1(n15190), .A2(n15189), .A3(n15188), .A4(n15187), .ZN(
        n15191) );
  OAI211_X1 U16714 ( .C1(n15194), .C2(n15193), .A(n15192), .B(n15191), .ZN(
        n15195) );
  NOR4_X1 U16715 ( .A1(n15198), .A2(n15197), .A3(n15196), .A4(n15195), .ZN(
        n15213) );
  INV_X1 U16716 ( .A(n15199), .ZN(n15204) );
  AOI22_X1 U16717 ( .A1(n15202), .A2(n15201), .B1(n15200), .B2(n10377), .ZN(
        n15203) );
  OAI21_X1 U16718 ( .B1(n15204), .B2(n9321), .A(n15203), .ZN(n15207) );
  INV_X1 U16719 ( .A(n15205), .ZN(n15206) );
  AOI211_X1 U16720 ( .C1(n15209), .C2(n15208), .A(n15207), .B(n15206), .ZN(
        n15211) );
  AOI22_X1 U16721 ( .A1(n13649), .A2(n9884), .B1(n15211), .B2(n15210), .ZN(
        n15212) );
  XOR2_X1 U16722 ( .A(n15213), .B(n15212), .Z(P2_U3262) );
  XOR2_X1 U16723 ( .A(n15215), .B(n15214), .Z(SUB_1596_U59) );
  XNOR2_X1 U16724 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15216), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16725 ( .B1(n15218), .B2(n15217), .A(n15223), .ZN(SUB_1596_U53) );
  XOR2_X1 U16726 ( .A(n15219), .B(n15220), .Z(SUB_1596_U56) );
  XNOR2_X1 U16727 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15221), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16728 ( .A(n15223), .B(n15222), .Z(SUB_1596_U5) );
  CLKBUF_X2 U7196 ( .A(n8352), .Z(n8791) );
  CLKBUF_X2 U7198 ( .A(n13876), .Z(n6456) );
  NAND3_X1 U7211 ( .A1(n6929), .A2(n6503), .A3(n6688), .ZN(n10911) );
  CLKBUF_X1 U7241 ( .A(n7434), .Z(n6804) );
  CLKBUF_X3 U7248 ( .A(n7662), .Z(n8930) );
  CLKBUF_X1 U7253 ( .A(n12235), .Z(n6647) );
  MUX2_X1 U7314 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7476), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7478) );
  CLKBUF_X1 U7417 ( .A(n10089), .Z(n12331) );
  OR2_X1 U7468 ( .A1(n9797), .A2(n9905), .ZN(n15228) );
endmodule

