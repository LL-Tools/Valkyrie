

module b14_C_gen_AntiSAT_k_128_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755;

  OAI21_X1 U2286 ( .B1(n3391), .B2(n3390), .A(n3389), .ZN(n3392) );
  INV_X2 U2287 ( .A(n2047), .ZN(n2049) );
  OAI22_X1 U2288 ( .A1(n2905), .A2(n2904), .B1(n4562), .B2(n2903), .ZN(n3953)
         );
  NAND2_X1 U2289 ( .A1(n2874), .A2(n2873), .ZN(n2875) );
  NAND2_X1 U2290 ( .A1(n3808), .A2(n3811), .ZN(n3768) );
  CLKBUF_X2 U2291 ( .A(n2364), .Z(n2596) );
  AND2_X1 U2292 ( .A1(n2638), .A2(n2667), .ZN(n2934) );
  NAND2_X1 U2293 ( .A1(n2692), .A2(IR_REG_31__SCAN_IN), .ZN(n2693) );
  AND2_X1 U2294 ( .A1(n2105), .A2(n2103), .ZN(n4388) );
  NAND2_X1 U2295 ( .A1(n2634), .A2(IR_REG_31__SCAN_IN), .ZN(n2636) );
  BUF_X1 U2296 ( .A(n2947), .Z(n2045) );
  NAND2_X1 U2298 ( .A1(n2836), .A2(n2934), .ZN(n3499) );
  XNOR2_X1 U2299 ( .A(n2857), .B(n3472), .ZN(n2870) );
  NAND2_X1 U2300 ( .A1(n3660), .A2(n3662), .ZN(n3659) );
  INV_X1 U2301 ( .A(n3896), .ZN(n3148) );
  INV_X1 U2302 ( .A(n2046), .ZN(n3742) );
  NAND2_X1 U2303 ( .A1(n4273), .A2(n2587), .ZN(n4085) );
  AOI21_X1 U2304 ( .B1(n2409), .B2(n2220), .A(n2070), .ZN(n2219) );
  AND2_X1 U2305 ( .A1(n2936), .A2(n3872), .ZN(n4537) );
  INV_X1 U2306 ( .A(IR_REG_31__SCAN_IN), .ZN(n2760) );
  XNOR2_X1 U2307 ( .A(n2636), .B(n2635), .ZN(n3798) );
  AOI211_X1 U2308 ( .C1(n2273), .C2(n3904), .A(n3885), .B(n2888), .ZN(n2921)
         );
  INV_X1 U2309 ( .A(n2074), .ZN(n3472) );
  INV_X1 U2311 ( .A(n3499), .ZN(n3542) );
  CLKBUF_X3 U2312 ( .A(n2363), .Z(n3738) );
  NOR2_X2 U2314 ( .A1(n2561), .A2(IR_REG_18__SCAN_IN), .ZN(n2633) );
  NOR2_X1 U2315 ( .A1(n2325), .A2(n2326), .ZN(n2354) );
  XNOR2_X2 U2316 ( .A(n2320), .B(IR_REG_30__SCAN_IN), .ZN(n2325) );
  NOR2_X1 U2317 ( .A1(n3553), .A2(n4537), .ZN(n2044) );
  AND2_X1 U2319 ( .A1(n3818), .A2(n3821), .ZN(n3772) );
  INV_X1 U2320 ( .A(n3897), .ZN(n2982) );
  NAND4_X1 U2321 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), .ZN(n3896)
         );
  INV_X1 U2322 ( .A(n3894), .ZN(n3215) );
  AND4_X1 U2323 ( .A1(n2368), .A2(n2367), .A3(n2366), .A4(n2365), .ZN(n2867)
         );
  INV_X2 U2324 ( .A(n2046), .ZN(n2487) );
  CLKBUF_X3 U2325 ( .A(n2354), .Z(n3737) );
  CLKBUF_X1 U2326 ( .A(n2638), .Z(n3872) );
  INV_X2 U2327 ( .A(IR_REG_0__SCAN_IN), .ZN(n2273) );
  NAND2_X1 U2328 ( .A1(n3536), .A2(n3530), .ZN(n3649) );
  NOR2_X1 U2329 ( .A1(n4054), .A2(n2599), .ZN(n2600) );
  NAND2_X1 U2330 ( .A1(n4118), .A2(n4117), .ZN(n4273) );
  NOR2_X1 U2331 ( .A1(n4468), .A2(n3971), .ZN(n4477) );
  NOR2_X1 U2332 ( .A1(n4467), .A2(REG1_REG_16__SCAN_IN), .ZN(n4468) );
  XNOR2_X1 U2333 ( .A(n3970), .B(n3969), .ZN(n4467) );
  AND2_X1 U2334 ( .A1(n4152), .A2(n4133), .ZN(n4128) );
  AOI21_X1 U2335 ( .B1(n2166), .B2(n2168), .A(n2076), .ZN(n2165) );
  NAND2_X1 U2336 ( .A1(n2255), .A2(n2256), .ZN(n2254) );
  AOI21_X1 U2337 ( .B1(n2284), .B2(n2287), .A(n2282), .ZN(n2281) );
  INV_X1 U2338 ( .A(n2284), .ZN(n2283) );
  AND2_X1 U2339 ( .A1(n2285), .A2(n2286), .ZN(n2284) );
  NAND2_X2 U2340 ( .A1(n2933), .A2(n4494), .ZN(n4200) );
  BUF_X4 U2341 ( .A(n3472), .Z(n2050) );
  INV_X1 U2342 ( .A(n3898), .ZN(n3036) );
  OR2_X1 U2343 ( .A1(n2596), .A2(n3137), .ZN(n2399) );
  NAND4_X1 U2344 ( .A1(n2389), .A2(n2388), .A3(n2387), .A4(n2386), .ZN(n3897)
         );
  AND2_X1 U2345 ( .A1(n2191), .A2(n2190), .ZN(n2799) );
  NAND4_X1 U2346 ( .A1(n2375), .A2(n2374), .A3(n2373), .A4(n2372), .ZN(n3898)
         );
  NAND4_X1 U2347 ( .A1(n2360), .A2(n2359), .A3(n2358), .A4(n2357), .ZN(n3901)
         );
  CLKBUF_X3 U2348 ( .A(n2355), .Z(n2558) );
  OR2_X1 U2349 ( .A1(n2823), .A2(n4380), .ZN(n2856) );
  INV_X1 U2350 ( .A(n3798), .ZN(n2667) );
  INV_X1 U2351 ( .A(n2326), .ZN(n2758) );
  INV_X2 U2352 ( .A(n2370), .ZN(n2046) );
  NAND2_X1 U2353 ( .A1(n2321), .A2(n2324), .ZN(n2326) );
  INV_X1 U2354 ( .A(n2673), .ZN(n2100) );
  OAI21_X1 U2355 ( .B1(n2691), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2698) );
  NAND2_X1 U2356 ( .A1(n2129), .A2(n2323), .ZN(n2324) );
  XNOR2_X1 U2357 ( .A(n2629), .B(IR_REG_19__SCAN_IN), .ZN(n4380) );
  AND2_X1 U2358 ( .A1(n2687), .A2(n2316), .ZN(n2673) );
  OAI211_X1 U2359 ( .C1(IR_REG_31__SCAN_IN), .C2(IR_REG_26__SCAN_IN), .A(n2687), .B(n2186), .ZN(n2769) );
  NAND2_X1 U2360 ( .A1(n2321), .A2(IR_REG_31__SCAN_IN), .ZN(n2320) );
  AND2_X1 U2361 ( .A1(n2315), .A2(n2060), .ZN(n2677) );
  OR2_X1 U2362 ( .A1(n2675), .A2(n2297), .ZN(n2674) );
  AND2_X1 U2363 ( .A1(n2313), .A2(n2251), .ZN(n2315) );
  INV_X1 U2364 ( .A(IR_REG_7__SCAN_IN), .ZN(n2430) );
  INV_X1 U2365 ( .A(IR_REG_3__SCAN_IN), .ZN(n2377) );
  NOR2_X1 U2366 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2495)
         );
  INV_X1 U2367 ( .A(IR_REG_5__SCAN_IN), .ZN(n2406) );
  INV_X1 U2368 ( .A(IR_REG_6__SCAN_IN), .ZN(n2417) );
  AND2_X1 U2369 ( .A1(n2860), .A2(n2837), .ZN(n2839) );
  OR2_X2 U2370 ( .A1(n3052), .A2(n3046), .ZN(n3053) );
  AOI21_X1 U2371 ( .B1(n2730), .B2(n3806), .A(n2299), .ZN(n3992) );
  XNOR2_X1 U2372 ( .A(n2730), .B(n2729), .ZN(n4004) );
  NAND2_X1 U2373 ( .A1(n2843), .A2(n2842), .ZN(n2861) );
  NAND2_X2 U2374 ( .A1(n2697), .A2(n2696), .ZN(n2836) );
  OAI21_X2 U2375 ( .B1(n3333), .B2(n2228), .A(n2226), .ZN(n3299) );
  NAND2_X2 U2376 ( .A1(n3322), .A2(n3321), .ZN(n3391) );
  MUX2_X2 U2377 ( .A(n2208), .B(n2207), .S(n2370), .Z(n3078) );
  OAI22_X1 U2378 ( .A1(n2867), .A2(n2951), .B1(n3499), .B2(n2869), .ZN(n2942)
         );
  INV_X1 U2379 ( .A(n3553), .ZN(n2947) );
  NOR2_X2 U2380 ( .A1(n3142), .A2(n3141), .ZN(n3166) );
  AOI21_X2 U2381 ( .B1(n2058), .B2(n2254), .A(n3130), .ZN(n3142) );
  AOI21_X1 U2382 ( .B1(n2859), .B2(n2044), .A(n2858), .ZN(n2871) );
  XNOR2_X2 U2383 ( .A(n2693), .B(IR_REG_24__SCAN_IN), .ZN(n2696) );
  NOR3_X2 U2384 ( .A1(n4045), .A2(n4236), .A3(n2737), .ZN(n2739) );
  XNOR2_X1 U2385 ( .A(n2806), .B(n2187), .ZN(n2801) );
  INV_X1 U2386 ( .A(n4383), .ZN(n2187) );
  INV_X1 U2387 ( .A(n2212), .ZN(n2211) );
  AOI21_X1 U2388 ( .B1(n2212), .B2(n2210), .A(n2081), .ZN(n2209) );
  NOR2_X1 U2389 ( .A1(n2597), .A2(n2082), .ZN(n2212) );
  NOR2_X1 U2390 ( .A1(n2588), .A2(n4603), .ZN(n2589) );
  AOI21_X1 U2391 ( .B1(n3774), .B2(n2478), .A(n2061), .ZN(n2229) );
  AND2_X1 U2392 ( .A1(n2064), .A2(n2219), .ZN(n2218) );
  NAND2_X1 U2393 ( .A1(n2854), .A2(n3070), .ZN(n3811) );
  AND2_X1 U2394 ( .A1(n2251), .A2(n2314), .ZN(n2250) );
  NAND2_X1 U2395 ( .A1(n2633), .A2(n2625), .ZN(n2691) );
  NAND2_X1 U2396 ( .A1(n2161), .A2(n2160), .ZN(n2403) );
  AND2_X1 U2397 ( .A1(n2377), .A2(n2302), .ZN(n2160) );
  INV_X1 U2398 ( .A(n3600), .ZN(n3503) );
  INV_X1 U2399 ( .A(n4386), .ZN(n2787) );
  NOR2_X1 U2400 ( .A1(n2796), .A2(n2189), .ZN(n2188) );
  INV_X1 U2401 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2189) );
  NAND2_X1 U2402 ( .A1(n4458), .A2(n3968), .ZN(n3970) );
  NOR2_X1 U2403 ( .A1(n2078), .A2(n2233), .ZN(n2232) );
  NOR2_X1 U2404 ( .A1(n2234), .A2(n3761), .ZN(n2233) );
  NAND2_X1 U2405 ( .A1(n3884), .A2(n2586), .ZN(n2587) );
  OR2_X1 U2406 ( .A1(n2766), .A2(D_REG_1__SCAN_IN), .ZN(n2929) );
  INV_X1 U2407 ( .A(n3893), .ZN(n3182) );
  NAND2_X1 U2408 ( .A1(n4471), .A2(n4473), .ZN(n4472) );
  NOR2_X1 U2409 ( .A1(n3800), .A2(n2093), .ZN(n2092) );
  NAND2_X1 U2410 ( .A1(n3799), .A2(n2077), .ZN(n2093) );
  NAND2_X1 U2411 ( .A1(n2177), .A2(n2181), .ZN(n2176) );
  INV_X1 U2412 ( .A(n2178), .ZN(n2177) );
  AND2_X1 U2413 ( .A1(n3462), .A2(n3448), .ZN(n2178) );
  NOR2_X1 U2414 ( .A1(n3673), .A2(n2170), .ZN(n2169) );
  INV_X1 U2415 ( .A(n3608), .ZN(n2170) );
  AND2_X1 U2416 ( .A1(n3588), .A2(n3586), .ZN(n3534) );
  NOR2_X1 U2417 ( .A1(n2340), .A2(n4690), .ZN(n2099) );
  NOR2_X1 U2418 ( .A1(n3553), .A2(n4537), .ZN(n3023) );
  OR2_X1 U2419 ( .A1(n2788), .A2(n2787), .ZN(n2115) );
  NAND2_X1 U2420 ( .A1(n4415), .A2(n3936), .ZN(n3937) );
  INV_X1 U2421 ( .A(n4433), .ZN(n2106) );
  NAND2_X1 U2422 ( .A1(n2235), .A2(n2236), .ZN(n2234) );
  OR2_X1 U2423 ( .A1(n4012), .A2(n4236), .ZN(n2235) );
  NAND2_X1 U2424 ( .A1(n3752), .A2(n2139), .ZN(n2138) );
  INV_X1 U2425 ( .A(n3780), .ZN(n2139) );
  NAND2_X1 U2426 ( .A1(n2589), .A2(REG3_REG_24__SCAN_IN), .ZN(n2340) );
  AND2_X1 U2427 ( .A1(n4139), .A2(n2658), .ZN(n3849) );
  AND2_X1 U2428 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2316)
         );
  NOR2_X1 U2429 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2632)
         );
  INV_X1 U2430 ( .A(IR_REG_17__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U2431 ( .A1(n2288), .A2(n3167), .ZN(n2286) );
  NOR2_X1 U2432 ( .A1(n2288), .A2(n3167), .ZN(n2287) );
  AND2_X1 U2433 ( .A1(n3534), .A2(n2167), .ZN(n2166) );
  NAND2_X1 U2434 ( .A1(n2169), .A2(n2293), .ZN(n2167) );
  INV_X1 U2435 ( .A(n2169), .ZN(n2168) );
  AOI21_X1 U2436 ( .B1(n3681), .B2(n3683), .A(n3682), .ZN(n3495) );
  INV_X1 U2437 ( .A(n3558), .ZN(n2263) );
  AOI21_X1 U2438 ( .B1(n2267), .B2(n2266), .A(n2054), .ZN(n2265) );
  INV_X1 U2439 ( .A(n2269), .ZN(n2266) );
  NOR2_X1 U2440 ( .A1(n2603), .A2(n4580), .ZN(n2610) );
  INV_X1 U2441 ( .A(DATAI_1_), .ZN(n2208) );
  INV_X1 U2442 ( .A(n4388), .ZN(n2207) );
  INV_X1 U2443 ( .A(DATAI_0_), .ZN(n2101) );
  NOR2_X1 U2444 ( .A1(n2080), .A2(n2291), .ZN(n2290) );
  AND2_X1 U2445 ( .A1(n2294), .A2(n2292), .ZN(n2291) );
  INV_X1 U2446 ( .A(n2099), .ZN(n2601) );
  NAND2_X1 U2447 ( .A1(n2099), .A2(REG3_REG_26__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U2448 ( .A1(n2891), .A2(n2777), .ZN(n2778) );
  AOI21_X1 U2449 ( .B1(n2197), .B2(n2383), .A(n2790), .ZN(n2116) );
  NAND2_X1 U2450 ( .A1(n2122), .A2(n2121), .ZN(n2120) );
  NAND2_X1 U2451 ( .A1(n4382), .A2(REG2_REG_7__SCAN_IN), .ZN(n2121) );
  INV_X1 U2452 ( .A(n2907), .ZN(n2122) );
  NAND2_X1 U2453 ( .A1(n4408), .A2(n3959), .ZN(n4413) );
  NAND2_X1 U2454 ( .A1(n4413), .A2(n4414), .ZN(n4412) );
  NAND2_X1 U2455 ( .A1(n4425), .A2(REG2_REG_12__SCAN_IN), .ZN(n4424) );
  OR2_X1 U2456 ( .A1(n4446), .A2(n3940), .ZN(n2127) );
  OAI21_X1 U2457 ( .B1(n4446), .B2(n2125), .A(n2124), .ZN(n3942) );
  NAND2_X1 U2458 ( .A1(n4454), .A2(n2128), .ZN(n2124) );
  OR2_X1 U2459 ( .A1(n3940), .A2(n2193), .ZN(n2125) );
  INV_X1 U2460 ( .A(n3864), .ZN(n2140) );
  OR2_X1 U2461 ( .A1(n4070), .A2(n2138), .ZN(n2137) );
  AND2_X1 U2462 ( .A1(n2140), .A2(n4022), .ZN(n2136) );
  AND2_X1 U2463 ( .A1(n4262), .A2(n4062), .ZN(n2599) );
  AOI21_X1 U2464 ( .B1(n2241), .B2(n2239), .A(n2079), .ZN(n2238) );
  NOR2_X1 U2465 ( .A1(n2244), .A2(n3781), .ZN(n2243) );
  NOR2_X1 U2466 ( .A1(n2056), .A2(n2562), .ZN(n2244) );
  AOI21_X1 U2467 ( .B1(n2243), .B2(n2056), .A(n2242), .ZN(n2241) );
  INV_X1 U2468 ( .A(n3782), .ZN(n2242) );
  NAND2_X1 U2469 ( .A1(n2563), .A2(REG3_REG_20__SCAN_IN), .ZN(n2578) );
  OAI21_X1 U2470 ( .B1(n2652), .B2(n2132), .A(n2130), .ZN(n3443) );
  INV_X1 U2471 ( .A(n2131), .ZN(n2130) );
  OAI21_X1 U2472 ( .B1(n2053), .B2(n2132), .A(n3793), .ZN(n2131) );
  INV_X1 U2473 ( .A(n3725), .ZN(n2132) );
  NAND2_X1 U2474 ( .A1(n2652), .A2(n2053), .ZN(n3412) );
  AOI21_X1 U2475 ( .B1(n2229), .B2(n2227), .A(n2069), .ZN(n2226) );
  INV_X1 U2476 ( .A(n2229), .ZN(n2228) );
  NAND2_X1 U2477 ( .A1(n2231), .A2(n2230), .ZN(n3331) );
  INV_X1 U2478 ( .A(n3774), .ZN(n2230) );
  INV_X1 U2479 ( .A(n3333), .ZN(n2231) );
  OAI21_X1 U2480 ( .B1(n3157), .B2(n2154), .A(n2150), .ZN(n3335) );
  AOI21_X1 U2481 ( .B1(n2153), .B2(n2152), .A(n2151), .ZN(n2150) );
  INV_X1 U2482 ( .A(n3834), .ZN(n2152) );
  INV_X1 U2483 ( .A(n3842), .ZN(n2151) );
  OAI21_X1 U2484 ( .B1(n3110), .B2(n2644), .A(n3830), .ZN(n3221) );
  INV_X1 U2485 ( .A(n2394), .ZN(n2220) );
  INV_X1 U2486 ( .A(n2409), .ZN(n2221) );
  OAI21_X1 U2487 ( .B1(n3045), .B2(n2642), .A(n3821), .ZN(n2979) );
  AND2_X1 U2488 ( .A1(n2821), .A2(n2820), .ZN(n2931) );
  AND2_X1 U2489 ( .A1(n2668), .A2(n3755), .ZN(n4172) );
  INV_X1 U2490 ( .A(n3213), .ZN(n3228) );
  NAND2_X1 U2491 ( .A1(n2751), .A2(n2695), .ZN(n2766) );
  NAND2_X1 U2492 ( .A1(n2322), .A2(IR_REG_31__SCAN_IN), .ZN(n2323) );
  OAI21_X1 U2493 ( .B1(n2677), .B2(n2760), .A(IR_REG_29__SCAN_IN), .ZN(n2129)
         );
  NOR2_X1 U2494 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2310)
         );
  NOR2_X1 U2495 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2309)
         );
  INV_X1 U2496 ( .A(IR_REG_23__SCAN_IN), .ZN(n2699) );
  XNOR2_X1 U2497 ( .A(n2627), .B(n2626), .ZN(n2823) );
  OR2_X1 U2498 ( .A1(n2633), .A2(n2760), .ZN(n2629) );
  AND2_X1 U2499 ( .A1(n2532), .A2(n2523), .ZN(n3948) );
  INV_X1 U2500 ( .A(IR_REG_9__SCAN_IN), .ZN(n2455) );
  INV_X1 U2501 ( .A(n3890), .ZN(n3405) );
  INV_X1 U2502 ( .A(n4095), .ZN(n4058) );
  INV_X1 U2503 ( .A(n3700), .ZN(n3707) );
  INV_X1 U2504 ( .A(n4317), .ZN(n3711) );
  OAI21_X1 U2505 ( .B1(n3874), .B2(n3872), .A(n2097), .ZN(n2096) );
  INV_X1 U2506 ( .A(n2098), .ZN(n2097) );
  OAI21_X1 U2507 ( .B1(n3873), .B2(n2754), .A(n3875), .ZN(n2098) );
  INV_X1 U2508 ( .A(n4262), .ZN(n4246) );
  OAI21_X1 U2509 ( .B1(n3591), .B2(n2596), .A(n2595), .ZN(n4259) );
  OR2_X1 U2510 ( .A1(n2517), .A2(n2516), .ZN(n3886) );
  NAND4_X1 U2511 ( .A1(n2439), .A2(n2438), .A3(n2437), .A4(n2436), .ZN(n3893)
         );
  INV_X1 U2512 ( .A(n2783), .ZN(n2190) );
  NAND2_X1 U2513 ( .A1(n4396), .A2(n4397), .ZN(n4395) );
  XNOR2_X1 U2514 ( .A(n3942), .B(n3969), .ZN(n4464) );
  NAND2_X1 U2515 ( .A1(n4464), .A2(n2525), .ZN(n4463) );
  NAND2_X1 U2516 ( .A1(n2202), .A2(n4435), .ZN(n2201) );
  NAND2_X1 U2517 ( .A1(n2203), .A2(n4484), .ZN(n2202) );
  NAND2_X1 U2518 ( .A1(n4472), .A2(n2204), .ZN(n2203) );
  AOI21_X1 U2519 ( .B1(n4486), .B2(ADDR_REG_18__SCAN_IN), .A(n4485), .ZN(n2200) );
  AND2_X1 U2520 ( .A1(n4472), .A2(n2088), .ZN(n4483) );
  INV_X1 U2521 ( .A(n2204), .ZN(n2123) );
  AND2_X1 U2522 ( .A1(n3906), .A2(n3902), .ZN(n4488) );
  NOR2_X1 U2523 ( .A1(n4016), .A2(n2158), .ZN(n2744) );
  NAND2_X1 U2524 ( .A1(n2159), .A2(n2735), .ZN(n2158) );
  NAND2_X1 U2525 ( .A1(n4004), .A2(n4546), .ZN(n2159) );
  NAND2_X1 U2526 ( .A1(n2744), .A2(n4554), .ZN(n2157) );
  INV_X1 U2527 ( .A(n2823), .ZN(n3879) );
  INV_X1 U2528 ( .A(n3946), .ZN(n4516) );
  AND2_X1 U2529 ( .A1(n2390), .A2(n2379), .ZN(n4386) );
  INV_X1 U2530 ( .A(n3202), .ZN(n2285) );
  NOR2_X1 U2531 ( .A1(n3200), .A2(n3201), .ZN(n2282) );
  INV_X1 U2532 ( .A(n3673), .ZN(n2296) );
  INV_X1 U2533 ( .A(n3662), .ZN(n2292) );
  NOR2_X1 U2534 ( .A1(n3801), .A2(n2091), .ZN(n2090) );
  NAND2_X1 U2535 ( .A1(n2094), .A2(n2092), .ZN(n2091) );
  OR2_X1 U2536 ( .A1(n2578), .A2(n2318), .ZN(n2588) );
  NOR2_X1 U2537 ( .A1(n2513), .A2(n2512), .ZN(n2526) );
  NAND2_X1 U2538 ( .A1(n2115), .A2(n2110), .ZN(n2109) );
  NAND2_X1 U2539 ( .A1(n3921), .A2(n2779), .ZN(n2780) );
  INV_X1 U2540 ( .A(n2598), .ZN(n2210) );
  AOI21_X1 U2541 ( .B1(n2148), .B2(n2144), .A(n2143), .ZN(n2142) );
  INV_X1 U2542 ( .A(n3856), .ZN(n2143) );
  INV_X1 U2543 ( .A(n3849), .ZN(n2144) );
  INV_X1 U2544 ( .A(n2148), .ZN(n2145) );
  INV_X1 U2545 ( .A(n2241), .ZN(n2240) );
  INV_X1 U2546 ( .A(n2243), .ZN(n2239) );
  AOI21_X1 U2547 ( .B1(n3849), .B2(n3727), .A(n2149), .ZN(n2148) );
  INV_X1 U2548 ( .A(n3729), .ZN(n2149) );
  NAND2_X1 U2549 ( .A1(n2526), .A2(REG3_REG_16__SCAN_IN), .ZN(n2537) );
  INV_X1 U2550 ( .A(n2478), .ZN(n2227) );
  NAND2_X1 U2551 ( .A1(n3834), .A2(n3156), .ZN(n2155) );
  NAND2_X1 U2552 ( .A1(n2224), .A2(n2371), .ZN(n2222) );
  INV_X1 U2553 ( .A(n3665), .ZN(n4153) );
  NAND2_X1 U2554 ( .A1(n2102), .A2(n3634), .ZN(n3437) );
  NOR2_X1 U2555 ( .A1(n3415), .A2(n4317), .ZN(n2102) );
  AND2_X1 U2556 ( .A1(n2312), .A2(n2252), .ZN(n2251) );
  INV_X1 U2557 ( .A(IR_REG_26__SCAN_IN), .ZN(n2252) );
  NOR2_X1 U2558 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2304)
         );
  NOR2_X1 U2559 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2305)
         );
  NOR2_X1 U2560 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2306)
         );
  NOR2_X1 U2561 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2307)
         );
  NOR2_X1 U2562 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2308)
         );
  XNOR2_X1 U2563 ( .A(n2631), .B(n2630), .ZN(n2638) );
  INV_X1 U2564 ( .A(IR_REG_20__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U2565 ( .A1(n2253), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U2566 ( .A1(n2629), .A2(n2628), .ZN(n2253) );
  OR3_X1 U2567 ( .A1(n2497), .A2(IR_REG_12__SCAN_IN), .A3(n2496), .ZN(n2507)
         );
  INV_X1 U2568 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2422) );
  OR2_X1 U2569 ( .A1(n2489), .A2(n2488), .ZN(n2501) );
  OR2_X1 U2570 ( .A1(n2501), .A2(n4693), .ZN(n2513) );
  AOI22_X1 U2571 ( .A1(n2178), .A2(n3449), .B1(n2180), .B2(n2182), .ZN(n2174)
         );
  NAND2_X1 U2572 ( .A1(n2184), .A2(n2183), .ZN(n2182) );
  INV_X1 U2573 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U2574 ( .A1(n2947), .A2(n3071), .ZN(n2860) );
  NAND2_X1 U2575 ( .A1(n2479), .A2(REG3_REG_12__SCAN_IN), .ZN(n2489) );
  NOR2_X1 U2576 ( .A1(n2076), .A2(n3530), .ZN(n3531) );
  NAND2_X1 U2577 ( .A1(n2173), .A2(n2172), .ZN(n2255) );
  INV_X1 U2578 ( .A(n3031), .ZN(n2173) );
  OAI22_X1 U2579 ( .A1(n3579), .A2(n2048), .B1(n2049), .B2(n3456), .ZN(n3461)
         );
  XNOR2_X1 U2580 ( .A(n2868), .B(n2050), .ZN(n2943) );
  OAI22_X1 U2581 ( .A1(n2869), .A2(n3553), .B1(n2867), .B2(n3499), .ZN(n2868)
         );
  NAND2_X1 U2582 ( .A1(n2674), .A2(n2206), .ZN(n2205) );
  AND2_X1 U2583 ( .A1(n2277), .A2(n3640), .ZN(n2275) );
  NAND2_X1 U2584 ( .A1(n3482), .A2(n3641), .ZN(n2277) );
  NOR2_X1 U2585 ( .A1(n2396), .A2(n2089), .ZN(n2410) );
  NAND2_X1 U2586 ( .A1(n2410), .A2(REG3_REG_6__SCAN_IN), .ZN(n2423) );
  AND2_X1 U2587 ( .A1(n2916), .A2(REG1_REG_4__SCAN_IN), .ZN(n2914) );
  CLKBUF_X1 U2588 ( .A(n2403), .Z(n2404) );
  NAND2_X1 U2589 ( .A1(n2114), .A2(n2113), .ZN(n2197) );
  AOI21_X1 U2590 ( .B1(n2115), .B2(n2789), .A(n2920), .ZN(n2113) );
  OR2_X1 U2591 ( .A1(n2914), .A2(n2192), .ZN(n2191) );
  AND2_X1 U2592 ( .A1(n2780), .A2(n4385), .ZN(n2192) );
  AND2_X1 U2593 ( .A1(n2196), .A2(n2195), .ZN(n2811) );
  NAND2_X1 U2594 ( .A1(n4384), .A2(REG2_REG_5__SCAN_IN), .ZN(n2195) );
  XNOR2_X1 U2595 ( .A(n2120), .B(n4381), .ZN(n3932) );
  INV_X1 U2596 ( .A(n4526), .ZN(n3951) );
  NAND2_X1 U2597 ( .A1(n4412), .A2(n3960), .ZN(n3962) );
  NAND2_X1 U2598 ( .A1(n2107), .A2(n2198), .ZN(n3939) );
  OR2_X1 U2599 ( .A1(n3949), .A2(REG2_REG_13__SCAN_IN), .ZN(n2198) );
  NAND2_X1 U2600 ( .A1(n4424), .A2(n2065), .ZN(n2107) );
  NAND2_X1 U2601 ( .A1(n4517), .A2(n2541), .ZN(n2204) );
  NAND2_X1 U2602 ( .A1(n2739), .A2(n3995), .ZN(n4231) );
  AND2_X1 U2603 ( .A1(n4240), .A2(n2737), .ZN(n3736) );
  NAND2_X1 U2604 ( .A1(n2135), .A2(n2134), .ZN(n2731) );
  AOI21_X1 U2605 ( .B1(n2136), .B2(n2138), .A(n3735), .ZN(n2134) );
  NAND2_X1 U2606 ( .A1(n4070), .A2(n2136), .ZN(n2135) );
  NAND2_X1 U2607 ( .A1(n2141), .A2(n2148), .ZN(n4124) );
  NAND2_X1 U2608 ( .A1(n4205), .A2(n3849), .ZN(n2141) );
  AND2_X1 U2609 ( .A1(n2570), .A2(n2569), .ZN(n4132) );
  AND2_X1 U2610 ( .A1(n2556), .A2(REG3_REG_19__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U2611 ( .A1(n2147), .A2(n2146), .ZN(n4140) );
  INV_X1 U2612 ( .A(n3727), .ZN(n2146) );
  INV_X1 U2613 ( .A(n4205), .ZN(n2147) );
  NOR2_X1 U2614 ( .A1(n2055), .A2(n2547), .ZN(n2556) );
  NOR2_X1 U2615 ( .A1(n2460), .A2(n2459), .ZN(n2468) );
  AND2_X1 U2616 ( .A1(n2468), .A2(REG3_REG_11__SCAN_IN), .ZN(n2479) );
  AOI21_X1 U2617 ( .B1(n2246), .B2(n2247), .A(n2063), .ZN(n2245) );
  INV_X1 U2618 ( .A(n2444), .ZN(n2246) );
  OR2_X1 U2619 ( .A1(n2447), .A2(n2446), .ZN(n2460) );
  NAND2_X1 U2620 ( .A1(n3221), .A2(n3833), .ZN(n2645) );
  INV_X1 U2621 ( .A(n3248), .ZN(n3255) );
  NOR2_X1 U2622 ( .A1(n2423), .A2(n2422), .ZN(n2434) );
  NAND2_X1 U2623 ( .A1(n2217), .A2(n2215), .ZN(n3121) );
  AND2_X1 U2624 ( .A1(n2216), .A2(n2420), .ZN(n2215) );
  OR2_X1 U2625 ( .A1(n3895), .A2(n3145), .ZN(n2420) );
  NAND2_X1 U2626 ( .A1(n2643), .A2(n3827), .ZN(n3110) );
  AND2_X1 U2627 ( .A1(n3828), .A2(n3830), .ZN(n3773) );
  AOI21_X1 U2628 ( .B1(n2979), .B2(n3825), .A(n2977), .ZN(n2992) );
  NAND2_X1 U2629 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2396) );
  NAND2_X1 U2630 ( .A1(n2641), .A2(n3817), .ZN(n3045) );
  NAND2_X1 U2631 ( .A1(n2225), .A2(n2640), .ZN(n3003) );
  INV_X1 U2632 ( .A(n3005), .ZN(n2225) );
  AND2_X1 U2633 ( .A1(n3901), .A2(n3071), .ZN(n3072) );
  NAND2_X1 U2634 ( .A1(n3768), .A2(n3072), .ZN(n3074) );
  NAND2_X1 U2635 ( .A1(n4064), .A2(n4048), .ZN(n4045) );
  INV_X1 U2636 ( .A(n4012), .ZN(n4249) );
  AND2_X1 U2637 ( .A1(n4074), .A2(n4062), .ZN(n4064) );
  NOR2_X1 U2638 ( .A1(n4100), .A2(n4258), .ZN(n4074) );
  INV_X1 U2639 ( .A(n4079), .ZN(n4258) );
  OR2_X1 U2640 ( .A1(n4114), .A2(n4098), .ZN(n4100) );
  NAND2_X1 U2641 ( .A1(n4128), .A2(n4112), .ZN(n4114) );
  NOR2_X2 U2642 ( .A1(n4176), .A2(n4153), .ZN(n4152) );
  NAND2_X1 U2643 ( .A1(n4211), .A2(n4195), .ZN(n4194) );
  INV_X1 U2644 ( .A(n2102), .ZN(n3438) );
  NAND2_X1 U2645 ( .A1(n3380), .A2(n3577), .ZN(n3415) );
  INV_X1 U2646 ( .A(n3464), .ZN(n3577) );
  AND2_X1 U2647 ( .A1(n3311), .A2(n3456), .ZN(n3380) );
  NOR2_X1 U2648 ( .A1(n3341), .A2(n3395), .ZN(n3311) );
  NAND2_X1 U2649 ( .A1(n2085), .A2(n3342), .ZN(n3341) );
  INV_X1 U2650 ( .A(n3284), .ZN(n3292) );
  INV_X1 U2651 ( .A(n4323), .ZN(n4278) );
  AND2_X1 U2652 ( .A1(n3226), .A2(n3255), .ZN(n3191) );
  NOR2_X2 U2653 ( .A1(n3227), .A2(n3228), .ZN(n3226) );
  INV_X1 U2654 ( .A(n3145), .ZN(n3149) );
  INV_X1 U2655 ( .A(n3132), .ZN(n2984) );
  AND2_X1 U2656 ( .A1(n2886), .A2(n2774), .ZN(n4319) );
  INV_X1 U2657 ( .A(n2963), .ZN(n2968) );
  NAND2_X1 U2658 ( .A1(n3012), .A2(n2968), .ZN(n3052) );
  NOR2_X1 U2659 ( .A1(n3068), .A2(n3013), .ZN(n3012) );
  AND3_X1 U2660 ( .A1(n2713), .A2(n2712), .A3(n2821), .ZN(n2723) );
  INV_X1 U2661 ( .A(IR_REG_21__SCAN_IN), .ZN(n2635) );
  NAND4_X1 U2662 ( .A1(n2441), .A2(n2430), .A3(n2417), .A4(n2406), .ZN(n2303)
         );
  AOI21_X1 U2663 ( .B1(n3166), .B2(n2280), .A(n2279), .ZN(n2278) );
  INV_X1 U2664 ( .A(n2286), .ZN(n2279) );
  INV_X1 U2665 ( .A(n2287), .ZN(n2280) );
  OR2_X1 U2666 ( .A1(n2319), .A2(n2610), .ZN(n4025) );
  NAND2_X1 U2667 ( .A1(n2185), .A2(n3694), .ZN(n3565) );
  NAND2_X1 U2668 ( .A1(n3541), .A2(n2269), .ZN(n2185) );
  INV_X1 U2669 ( .A(n4093), .ZN(n4098) );
  AND2_X1 U2670 ( .A1(n3585), .A2(n3586), .ZN(n3589) );
  OR2_X1 U2671 ( .A1(n3659), .A2(n2168), .ZN(n2164) );
  AND2_X1 U2672 ( .A1(n2265), .A2(n2263), .ZN(n2259) );
  OAI21_X1 U2673 ( .B1(n2265), .B2(n3558), .A(n2261), .ZN(n2260) );
  NAND2_X1 U2674 ( .A1(n2265), .A2(n2262), .ZN(n2261) );
  NAND2_X1 U2675 ( .A1(n2268), .A2(n2263), .ZN(n2262) );
  NAND2_X1 U2676 ( .A1(n2267), .A2(n3558), .ZN(n2264) );
  INV_X1 U2677 ( .A(n3078), .ZN(n3070) );
  NAND2_X1 U2678 ( .A1(n3659), .A2(n3661), .ZN(n3612) );
  INV_X1 U2679 ( .A(n2925), .ZN(n3071) );
  NAND2_X1 U2680 ( .A1(n2355), .A2(REG0_REG_1__SCAN_IN), .ZN(n2350) );
  OR2_X1 U2681 ( .A1(n3450), .A2(n3449), .ZN(n2179) );
  NAND2_X1 U2682 ( .A1(n2171), .A2(n3608), .ZN(n3672) );
  NAND2_X1 U2683 ( .A1(n3659), .A2(n2294), .ZN(n2171) );
  NAND2_X1 U2684 ( .A1(n2870), .A2(n2872), .ZN(n2873) );
  INV_X1 U2685 ( .A(n2871), .ZN(n2872) );
  XNOR2_X1 U2686 ( .A(n2943), .B(n2942), .ZN(n2876) );
  OR2_X1 U2687 ( .A1(n2851), .A2(n2846), .ZN(n3700) );
  INV_X1 U2688 ( .A(n3716), .ZN(n3685) );
  OR2_X1 U2689 ( .A1(n2851), .A2(n2850), .ZN(n3699) );
  NAND2_X1 U2690 ( .A1(n2956), .A2(n2955), .ZN(n3713) );
  NAND2_X1 U2691 ( .A1(n2346), .A2(n2345), .ZN(n4095) );
  OR2_X1 U2692 ( .A1(n3653), .A2(n2596), .ZN(n2346) );
  NAND2_X1 U2693 ( .A1(n2576), .A2(n2575), .ZN(n4109) );
  INV_X1 U2694 ( .A(n4132), .ZN(n4279) );
  OR2_X1 U2695 ( .A1(n2543), .A2(n2542), .ZN(n4308) );
  INV_X1 U2696 ( .A(n4303), .ZN(n4320) );
  OR2_X1 U2697 ( .A1(n2748), .A2(n2836), .ZN(n3885) );
  NAND4_X1 U2698 ( .A1(n2506), .A2(n2505), .A3(n2504), .A4(n2503), .ZN(n3887)
         );
  OR2_X1 U2699 ( .A1(n3738), .A2(n3262), .ZN(n2482) );
  INV_X1 U2700 ( .A(n2867), .ZN(n3899) );
  AOI21_X1 U2701 ( .B1(n2913), .B2(REG2_REG_4__SCAN_IN), .A(n2194), .ZN(n2791)
         );
  INV_X1 U2702 ( .A(n2197), .ZN(n2194) );
  INV_X1 U2703 ( .A(n2191), .ZN(n2784) );
  XNOR2_X1 U2704 ( .A(n2811), .B(n4383), .ZN(n2813) );
  XNOR2_X1 U2705 ( .A(n3953), .B(n3952), .ZN(n3954) );
  OAI22_X1 U2706 ( .A1(n3932), .A2(n4496), .B1(n3952), .B2(n2119), .ZN(n4396)
         );
  INV_X1 U2707 ( .A(n2120), .ZN(n2119) );
  XNOR2_X1 U2708 ( .A(n3958), .B(n4525), .ZN(n4409) );
  NAND2_X1 U2709 ( .A1(n4409), .A2(REG1_REG_10__SCAN_IN), .ZN(n4408) );
  NAND2_X1 U2710 ( .A1(n4403), .A2(n3935), .ZN(n4416) );
  NAND2_X1 U2711 ( .A1(n4416), .A2(n4417), .ZN(n4415) );
  NAND2_X1 U2712 ( .A1(n4424), .A2(n3938), .ZN(n4437) );
  XNOR2_X1 U2713 ( .A(n3939), .B(n4520), .ZN(n4447) );
  INV_X1 U2714 ( .A(n4454), .ZN(n2126) );
  INV_X1 U2715 ( .A(n2127), .ZN(n4455) );
  NAND2_X1 U2716 ( .A1(n4463), .A2(n3943), .ZN(n4471) );
  NOR2_X1 U2717 ( .A1(n4483), .A2(n2087), .ZN(n3944) );
  INV_X1 U2718 ( .A(n3806), .ZN(n2729) );
  NAND2_X1 U2719 ( .A1(n2137), .A2(n2136), .ZN(n4019) );
  AND2_X1 U2720 ( .A1(n2137), .A2(n2140), .ZN(n4020) );
  INV_X1 U2721 ( .A(n4240), .ZN(n4033) );
  AND2_X1 U2722 ( .A1(n2338), .A2(n2337), .ZN(n4262) );
  OR2_X1 U2723 ( .A1(n3622), .A2(n2596), .ZN(n2338) );
  AND2_X1 U2724 ( .A1(n2213), .A2(n2214), .ZN(n4072) );
  NAND2_X1 U2725 ( .A1(n4085), .A2(n2598), .ZN(n2213) );
  NAND2_X1 U2726 ( .A1(n2237), .A2(n2241), .ZN(n4126) );
  NAND2_X1 U2727 ( .A1(n4160), .A2(n2243), .ZN(n2237) );
  AOI21_X1 U2728 ( .B1(n4160), .B2(n2562), .A(n2056), .ZN(n4145) );
  NAND2_X1 U2729 ( .A1(n3412), .A2(n3725), .ZN(n3444) );
  INV_X1 U2730 ( .A(n3886), .ZN(n4310) );
  NAND2_X1 U2731 ( .A1(n2652), .A2(n3718), .ZN(n3411) );
  INV_X1 U2732 ( .A(n3887), .ZN(n4324) );
  NAND2_X1 U2733 ( .A1(n3331), .A2(n2478), .ZN(n3260) );
  NAND4_X1 U2734 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n3891)
         );
  NAND2_X1 U2735 ( .A1(n2249), .A2(n2445), .ZN(n3163) );
  NAND2_X1 U2736 ( .A1(n3220), .A2(n2444), .ZN(n2249) );
  OAI21_X1 U2737 ( .B1(n3042), .B2(n2221), .A(n2219), .ZN(n2989) );
  NAND2_X1 U2738 ( .A1(n3042), .A2(n2394), .ZN(n2978) );
  OR2_X1 U2739 ( .A1(n4196), .A2(n3114), .ZN(n4179) );
  OR2_X1 U2740 ( .A1(n2928), .A2(n2834), .ZN(n4494) );
  INV_X1 U2741 ( .A(n4179), .ZN(n4508) );
  NAND2_X1 U2742 ( .A1(n2686), .A2(n2067), .ZN(n2186) );
  NAND2_X1 U2743 ( .A1(n2766), .A2(n2765), .ZN(n4514) );
  AND2_X1 U2744 ( .A1(n2440), .A2(n2432), .ZN(n4382) );
  OR2_X1 U2745 ( .A1(n2353), .A2(n2760), .ZN(n2369) );
  NAND2_X1 U2746 ( .A1(n2057), .A2(IR_REG_1__SCAN_IN), .ZN(n2105) );
  NOR2_X1 U2747 ( .A1(n2353), .A2(n2104), .ZN(n2103) );
  INV_X1 U2748 ( .A(n2172), .ZN(n3032) );
  OAI21_X1 U2749 ( .B1(n2095), .B2(n3881), .A(n3880), .ZN(U3239) );
  XNOR2_X1 U2750 ( .A(n2096), .B(n4380), .ZN(n2095) );
  INV_X1 U2751 ( .A(n2199), .ZN(n4492) );
  OAI21_X1 U2752 ( .B1(n4483), .B2(n2201), .A(n2200), .ZN(n2199) );
  NOR2_X1 U2753 ( .A1(n4564), .A2(n2719), .ZN(n2720) );
  NAND2_X1 U2754 ( .A1(n2741), .A2(n2740), .ZN(n2742) );
  NOR2_X1 U2755 ( .A1(n4554), .A2(n2724), .ZN(n2725) );
  NAND2_X1 U2756 ( .A1(n2741), .A2(n2726), .ZN(n2746) );
  NAND2_X1 U2757 ( .A1(n2157), .A2(n2156), .ZN(n2747) );
  NAND2_X1 U2758 ( .A1(n4552), .A2(n2745), .ZN(n2156) );
  AND4_X1 U2759 ( .A1(n2304), .A2(n2305), .A3(n2306), .A4(n2495), .ZN(n2051)
         );
  OR2_X1 U2760 ( .A1(n2240), .A2(n2075), .ZN(n2052) );
  AND2_X1 U2761 ( .A1(n2133), .A2(n3718), .ZN(n2053) );
  NOR2_X1 U2762 ( .A1(n2295), .A2(n3607), .ZN(n2294) );
  INV_X1 U2763 ( .A(n2294), .ZN(n2293) );
  INV_X1 U2764 ( .A(n3334), .ZN(n3342) );
  AND2_X1 U2765 ( .A1(n3552), .A2(n3551), .ZN(n2054) );
  INV_X1 U2766 ( .A(n3462), .ZN(n2183) );
  OR2_X1 U2767 ( .A1(n2537), .A2(n2536), .ZN(n2055) );
  NOR2_X1 U2768 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2353)
         );
  AND4_X1 U2769 ( .A1(n2352), .A2(n2351), .A3(n2350), .A4(n2349), .ZN(n2854)
         );
  NOR2_X1 U2770 ( .A1(n4142), .A2(n4174), .ZN(n2056) );
  AND2_X1 U2771 ( .A1(n2327), .A2(n2326), .ZN(n2355) );
  AND2_X1 U2772 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2057)
         );
  NAND2_X1 U2773 ( .A1(n3126), .A2(n3125), .ZN(n2058) );
  OR2_X1 U2774 ( .A1(n4045), .A2(n4236), .ZN(n2059) );
  AND2_X1 U2775 ( .A1(n2206), .A2(n2314), .ZN(n2060) );
  AND2_X1 U2776 ( .A1(n3889), .A2(n3395), .ZN(n2061) );
  NOR2_X1 U2777 ( .A1(n4070), .A2(n3780), .ZN(n2062) );
  NAND2_X1 U2778 ( .A1(n2164), .A2(n2166), .ZN(n3587) );
  AND2_X1 U2779 ( .A1(n3293), .A2(n3255), .ZN(n2063) );
  NAND2_X1 U2780 ( .A1(n3895), .A2(n3145), .ZN(n2064) );
  OAI21_X1 U2781 ( .B1(n3660), .B2(n2293), .A(n2290), .ZN(n3585) );
  INV_X1 U2782 ( .A(n2313), .ZN(n2688) );
  AND2_X1 U2783 ( .A1(n3938), .A2(n2106), .ZN(n2065) );
  NAND2_X1 U2784 ( .A1(n3892), .A2(n3248), .ZN(n2066) );
  AND2_X1 U2785 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2067)
         );
  AND2_X1 U2786 ( .A1(n2127), .A2(n2126), .ZN(n2068) );
  AND2_X1 U2787 ( .A1(n2647), .A2(n3404), .ZN(n2069) );
  AND2_X1 U2788 ( .A1(n3896), .A2(n2984), .ZN(n2070) );
  INV_X1 U2789 ( .A(n2248), .ZN(n2247) );
  NAND2_X1 U2790 ( .A1(n2445), .A2(n2066), .ZN(n2248) );
  AND2_X1 U2791 ( .A1(n3290), .A2(n3282), .ZN(n2071) );
  AND2_X1 U2792 ( .A1(n2945), .A2(n2946), .ZN(n2072) );
  AND2_X1 U2793 ( .A1(n2060), .A2(n2322), .ZN(n2073) );
  INV_X1 U2794 ( .A(IR_REG_27__SCAN_IN), .ZN(n2314) );
  INV_X1 U2795 ( .A(IR_REG_29__SCAN_IN), .ZN(n2322) );
  INV_X1 U2796 ( .A(IR_REG_28__SCAN_IN), .ZN(n2206) );
  AND2_X2 U2797 ( .A1(n2856), .A2(n2855), .ZN(n2074) );
  INV_X1 U2798 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2089) );
  AND2_X1 U2799 ( .A1(n4144), .A2(n4133), .ZN(n2075) );
  OR2_X1 U2800 ( .A1(n3564), .A2(n3695), .ZN(n2268) );
  NAND2_X1 U2801 ( .A1(n2175), .A2(n2174), .ZN(n3571) );
  NAND2_X1 U2802 ( .A1(n2276), .A2(n3483), .ZN(n3639) );
  AND2_X1 U2803 ( .A1(n2179), .A2(n3448), .ZN(n3463) );
  AND2_X1 U2804 ( .A1(n3528), .A2(n3527), .ZN(n2076) );
  AND3_X1 U2805 ( .A1(n3797), .A2(n3869), .A3(n3798), .ZN(n2077) );
  XOR2_X1 U2806 ( .A(n2050), .B(n3452), .Z(n3462) );
  NOR2_X1 U2807 ( .A1(n4249), .A2(n4029), .ZN(n2078) );
  INV_X1 U2808 ( .A(n2181), .ZN(n2180) );
  OAI21_X1 U2809 ( .B1(n3462), .B2(n3448), .A(n3461), .ZN(n2181) );
  AND2_X1 U2810 ( .A1(n4109), .A2(n4277), .ZN(n2079) );
  NAND2_X1 U2811 ( .A1(n2296), .A2(n3608), .ZN(n2080) );
  NOR2_X1 U2812 ( .A1(n4095), .A2(n4258), .ZN(n2081) );
  NOR2_X1 U2813 ( .A1(n4058), .A2(n4079), .ZN(n2082) );
  INV_X1 U2814 ( .A(n2154), .ZN(n2153) );
  NAND2_X1 U2815 ( .A1(n2155), .A2(n3838), .ZN(n2154) );
  AND2_X1 U2816 ( .A1(n3631), .A2(n3641), .ZN(n2083) );
  INV_X1 U2817 ( .A(n2268), .ZN(n2267) );
  AND3_X1 U2818 ( .A1(n4090), .A2(n4166), .A3(n2090), .ZN(n2084) );
  INV_X1 U2819 ( .A(n3762), .ZN(n2236) );
  INV_X1 U2820 ( .A(n3449), .ZN(n2184) );
  INV_X1 U2821 ( .A(n3661), .ZN(n2295) );
  AND2_X1 U2822 ( .A1(n3191), .A2(n3292), .ZN(n2085) );
  OAI21_X1 U2823 ( .B1(n3245), .B2(n3246), .A(n3247), .ZN(n3277) );
  NAND2_X1 U2824 ( .A1(n3003), .A2(n2371), .ZN(n2961) );
  INV_X1 U2825 ( .A(n2278), .ZN(n3203) );
  INV_X1 U2826 ( .A(n4146), .ZN(n2094) );
  INV_X1 U2827 ( .A(n3769), .ZN(n2133) );
  NAND2_X1 U2828 ( .A1(n2289), .A2(n3282), .ZN(n3288) );
  AND2_X1 U2829 ( .A1(n2254), .A2(n2058), .ZN(n2086) );
  INV_X1 U2830 ( .A(n2597), .ZN(n2214) );
  AND2_X1 U2831 ( .A1(n3906), .A2(n3876), .ZN(n4435) );
  AND2_X1 U2832 ( .A1(n2313), .A2(n2250), .ZN(n2675) );
  NOR2_X1 U2833 ( .A1(n2876), .A2(n2875), .ZN(n2944) );
  INV_X1 U2834 ( .A(n2193), .ZN(n2128) );
  AND2_X1 U2835 ( .A1(n3948), .A2(REG2_REG_15__SCAN_IN), .ZN(n2193) );
  INV_X1 U2836 ( .A(n3973), .ZN(n4517) );
  AND2_X1 U2837 ( .A1(n3946), .A2(REG2_REG_18__SCAN_IN), .ZN(n2087) );
  NOR2_X1 U2838 ( .A1(n2123), .A2(n4484), .ZN(n2088) );
  NAND4_X1 U2839 ( .A1(n4022), .A2(n3993), .A3(n4073), .A4(n2084), .ZN(n3802)
         );
  NAND2_X1 U2840 ( .A1(n2434), .A2(REG3_REG_8__SCAN_IN), .ZN(n2447) );
  MUX2_X1 U2841 ( .A(n2101), .B(n2273), .S(n2370), .Z(n2925) );
  OAI21_X2 U2842 ( .B1(n2100), .B2(n2206), .A(n2205), .ZN(n2370) );
  NOR2_X2 U2843 ( .A1(n3053), .A2(n2984), .ZN(n2993) );
  NOR2_X2 U2844 ( .A1(n3437), .A2(n4299), .ZN(n4211) );
  AND3_X2 U2845 ( .A1(n2162), .A2(n2051), .A3(n2311), .ZN(n2313) );
  NOR2_X2 U2846 ( .A1(n2403), .A2(n2303), .ZN(n2162) );
  NAND2_X1 U2847 ( .A1(n4404), .A2(REG2_REG_10__SCAN_IN), .ZN(n4403) );
  MUX2_X1 U2848 ( .A(REG2_REG_1__SCAN_IN), .B(n2785), .S(n4388), .Z(n3912) );
  NOR2_X1 U2849 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2104)
         );
  OAI211_X1 U2850 ( .C1(n3923), .C2(n2112), .A(n2111), .B(n2108), .ZN(n2118)
         );
  OAI21_X1 U2851 ( .B1(n2115), .B2(n4385), .A(n2109), .ZN(n2108) );
  OR2_X1 U2852 ( .A1(n4385), .A2(REG2_REG_3__SCAN_IN), .ZN(n2110) );
  NAND3_X1 U2853 ( .A1(n3923), .A2(n2115), .A3(n2920), .ZN(n2111) );
  NAND2_X1 U2854 ( .A1(n4385), .A2(REG2_REG_3__SCAN_IN), .ZN(n2112) );
  NAND2_X1 U2855 ( .A1(n3923), .A2(n2115), .ZN(n2114) );
  INV_X1 U2856 ( .A(n2118), .ZN(n2913) );
  NAND2_X1 U2857 ( .A1(n2117), .A2(n2116), .ZN(n2196) );
  NAND2_X1 U2858 ( .A1(n2197), .A2(n2118), .ZN(n2117) );
  OAI21_X1 U2859 ( .B1(n4205), .B2(n2145), .A(n2142), .ZN(n2662) );
  OAI21_X1 U2860 ( .B1(n3157), .B2(n3156), .A(n3834), .ZN(n3189) );
  AND2_X1 U2861 ( .A1(n2162), .A2(n2051), .ZN(n2552) );
  INV_X1 U2862 ( .A(n2376), .ZN(n2161) );
  NAND2_X1 U2863 ( .A1(n2163), .A2(n2165), .ZN(n3536) );
  NAND2_X1 U2864 ( .A1(n3659), .A2(n2166), .ZN(n2163) );
  NAND2_X1 U2866 ( .A1(n3450), .A2(n2176), .ZN(n2175) );
  NAND2_X2 U2867 ( .A1(n3620), .A2(n3619), .ZN(n3541) );
  NAND2_X4 U2868 ( .A1(n2836), .A2(n2855), .ZN(n3553) );
  OAI21_X2 U2869 ( .B1(n3166), .B2(n2283), .A(n2281), .ZN(n3245) );
  INV_X1 U2870 ( .A(n2769), .ZN(n2751) );
  INV_X1 U2871 ( .A(n2315), .ZN(n2687) );
  NOR2_X2 U2872 ( .A1(n2799), .A2(n2188), .ZN(n2806) );
  NOR2_X1 U2873 ( .A1(n2801), .A2(n3094), .ZN(n2807) );
  AOI21_X1 U2874 ( .B1(n3983), .B2(n4488), .A(n3982), .ZN(n3984) );
  NOR2_X1 U2875 ( .A1(n3974), .A2(n4478), .ZN(n4489) );
  NOR2_X1 U2876 ( .A1(n4477), .A2(n4476), .ZN(n4478) );
  NAND2_X1 U2877 ( .A1(n3277), .A2(n3276), .ZN(n2289) );
  NAND2_X2 U2878 ( .A1(n3597), .A2(n3504), .ZN(n3660) );
  NAND2_X1 U2879 ( .A1(n2313), .A2(n2312), .ZN(n2686) );
  INV_X1 U2880 ( .A(n2196), .ZN(n2797) );
  OAI21_X2 U2881 ( .B1(n4085), .B2(n2211), .A(n2209), .ZN(n4054) );
  NAND2_X1 U2882 ( .A1(n2218), .A2(n3042), .ZN(n2217) );
  NAND3_X1 U2883 ( .A1(n2064), .A2(n2219), .A3(n2221), .ZN(n2216) );
  NAND2_X1 U2884 ( .A1(n3005), .A2(n2371), .ZN(n2223) );
  NAND3_X1 U2885 ( .A1(n2223), .A2(n2222), .A3(n2380), .ZN(n2382) );
  INV_X1 U2886 ( .A(n2640), .ZN(n2224) );
  OAI21_X1 U2887 ( .B1(n4042), .B2(n2234), .A(n2232), .ZN(n2730) );
  AOI21_X1 U2888 ( .B1(n4042), .B2(n3761), .A(n3762), .ZN(n4023) );
  OAI22_X2 U2889 ( .A1(n4160), .A2(n2052), .B1(n2238), .B2(n2075), .ZN(n4118)
         );
  OAI21_X2 U2890 ( .B1(n3220), .B2(n2248), .A(n2245), .ZN(n3190) );
  NAND2_X1 U2891 ( .A1(n2255), .A2(n3030), .ZN(n3033) );
  INV_X1 U2892 ( .A(n2254), .ZN(n3127) );
  NOR2_X1 U2893 ( .A1(n3034), .A2(n2257), .ZN(n2256) );
  INV_X1 U2894 ( .A(n3030), .ZN(n2257) );
  NAND2_X1 U2895 ( .A1(n3541), .A2(n2259), .ZN(n2258) );
  OAI211_X1 U2896 ( .C1(n3541), .C2(n2264), .A(n2260), .B(n2258), .ZN(n3563)
         );
  NAND2_X1 U2897 ( .A1(n3541), .A2(n3618), .ZN(n3693) );
  NOR2_X1 U2898 ( .A1(n3696), .A2(n2270), .ZN(n2269) );
  INV_X1 U2899 ( .A(n3618), .ZN(n2270) );
  INV_X1 U2900 ( .A(IR_REG_1__SCAN_IN), .ZN(n2272) );
  INV_X1 U2901 ( .A(IR_REG_2__SCAN_IN), .ZN(n2271) );
  NAND3_X1 U2902 ( .A1(n2273), .A2(n2272), .A3(n2271), .ZN(n2376) );
  NAND3_X1 U2903 ( .A1(n3628), .A2(n3481), .A3(n2083), .ZN(n2274) );
  NAND2_X1 U2904 ( .A1(n2274), .A2(n2275), .ZN(n3681) );
  NAND3_X1 U2905 ( .A1(n3628), .A2(n3481), .A3(n3631), .ZN(n2276) );
  INV_X1 U2906 ( .A(n3168), .ZN(n2288) );
  NAND2_X1 U2907 ( .A1(n2289), .A2(n2071), .ZN(n3322) );
  NAND2_X1 U2908 ( .A1(n2315), .A2(n2073), .ZN(n2321) );
  INV_X2 U2909 ( .A(n2934), .ZN(n2855) );
  NAND2_X1 U2910 ( .A1(n2552), .A2(n2551), .ZN(n2561) );
  AOI21_X1 U2911 ( .B1(n2685), .B2(n4546), .A(n2684), .ZN(n2728) );
  XNOR2_X1 U2912 ( .A(n3992), .B(n2623), .ZN(n2685) );
  OAI22_X1 U2913 ( .A1(n2854), .A2(n3499), .B1(n3553), .B2(n3078), .ZN(n2857)
         );
  OR2_X1 U2914 ( .A1(n2363), .A2(n2362), .ZN(n2367) );
  INV_X1 U2915 ( .A(n2363), .ZN(n2348) );
  NAND2_X1 U2916 ( .A1(n2325), .A2(n2326), .ZN(n2363) );
  NAND2_X1 U2917 ( .A1(n2325), .A2(n2758), .ZN(n2364) );
  NAND2_X2 U2918 ( .A1(n4183), .A2(n2555), .ZN(n4160) );
  AND2_X2 U2919 ( .A1(n2723), .A2(n2932), .ZN(n4554) );
  INV_X1 U2920 ( .A(n4378), .ZN(n2726) );
  AND2_X1 U2921 ( .A1(n2314), .A2(n2760), .ZN(n2297) );
  INV_X1 U2922 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2446) );
  AND2_X1 U2923 ( .A1(n4310), .A2(n3711), .ZN(n2298) );
  AND2_X1 U2924 ( .A1(n4033), .A2(n2737), .ZN(n2299) );
  NAND2_X1 U2925 ( .A1(n2393), .A2(n2392), .ZN(n3042) );
  AND2_X1 U2926 ( .A1(n3888), .A2(n3451), .ZN(n2300) );
  OR2_X1 U2927 ( .A1(n3888), .A2(n3451), .ZN(n2301) );
  INV_X1 U2928 ( .A(n3884), .ZN(n4283) );
  NAND2_X1 U2929 ( .A1(n2585), .A2(n2584), .ZN(n3884) );
  INV_X1 U2930 ( .A(n3998), .ZN(n2721) );
  AND2_X1 U2931 ( .A1(n3848), .A2(n3720), .ZN(n3793) );
  INV_X1 U2932 ( .A(n3793), .ZN(n2534) );
  INV_X1 U2933 ( .A(n4112), .ZN(n2586) );
  NOR2_X1 U2934 ( .A1(n3475), .A2(n3474), .ZN(n3473) );
  NAND2_X1 U2935 ( .A1(n3537), .A2(n3649), .ZN(n3620) );
  INV_X1 U2936 ( .A(n3535), .ZN(n3530) );
  INV_X1 U2937 ( .A(IR_REG_4__SCAN_IN), .ZN(n2302) );
  AND4_X1 U2938 ( .A1(n2310), .A2(n2309), .A3(n2308), .A4(n2307), .ZN(n2311)
         );
  INV_X1 U2939 ( .A(n3289), .ZN(n3290) );
  INV_X1 U2940 ( .A(n3023), .ZN(n2951) );
  INV_X1 U2941 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2512) );
  AND2_X1 U2942 ( .A1(n4259), .A2(n4098), .ZN(n2597) );
  INV_X1 U2943 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2488) );
  AND2_X1 U2944 ( .A1(n4279), .A2(n4153), .ZN(n3781) );
  NAND2_X1 U2945 ( .A1(n2382), .A2(n2381), .ZN(n3043) );
  NAND2_X1 U2946 ( .A1(n2867), .A2(n3013), .ZN(n3812) );
  INV_X1 U2947 ( .A(n4218), .ZN(n4299) );
  NAND2_X1 U2948 ( .A1(n2993), .A2(n3149), .ZN(n3116) );
  INV_X1 U2949 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4693) );
  AOI21_X1 U2950 ( .B1(n4209), .B2(n2546), .A(n2545), .ZN(n4185) );
  NAND2_X1 U2951 ( .A1(n3443), .A2(n3720), .ZN(n4205) );
  INV_X1 U2952 ( .A(n3891), .ZN(n3355) );
  INV_X1 U2953 ( .A(n3892), .ZN(n3293) );
  INV_X1 U2954 ( .A(n4319), .ZN(n4282) );
  OR2_X1 U2955 ( .A1(n2766), .A2(D_REG_0__SCAN_IN), .ZN(n2715) );
  INV_X1 U2956 ( .A(n2664), .ZN(n4062) );
  INV_X1 U2957 ( .A(n3451), .ZN(n3456) );
  OR2_X1 U2958 ( .A1(n2766), .A2(n2711), .ZN(n2821) );
  AND2_X1 U2959 ( .A1(n2611), .A2(n3997), .ZN(n4005) );
  INV_X1 U2960 ( .A(n3699), .ZN(n3708) );
  NAND2_X1 U2961 ( .A1(n2836), .A2(n4515), .ZN(n2928) );
  AND2_X1 U2962 ( .A1(n2603), .A2(n2602), .ZN(n4046) );
  AND2_X1 U2963 ( .A1(n2616), .A2(n2615), .ZN(n4240) );
  OR2_X1 U2964 ( .A1(n3674), .A2(n2596), .ZN(n2585) );
  AND4_X1 U2965 ( .A1(n2531), .A2(n2530), .A3(n2529), .A4(n2528), .ZN(n4303)
         );
  OR2_X1 U2966 ( .A1(n3738), .A2(n4496), .ZN(n2437) );
  INV_X1 U2967 ( .A(IR_REG_8__SCAN_IN), .ZN(n2441) );
  AND2_X1 U2968 ( .A1(n2782), .A2(n2781), .ZN(n3906) );
  INV_X1 U2969 ( .A(n4168), .ZN(n4318) );
  AND2_X1 U2970 ( .A1(n3268), .A2(n3270), .ZN(n3774) );
  INV_X1 U2971 ( .A(n4203), .ZN(n4210) );
  INV_X1 U2972 ( .A(n4172), .ZN(n4206) );
  INV_X1 U2973 ( .A(n4328), .ZN(n2740) );
  AND2_X1 U2974 ( .A1(n2715), .A2(n2714), .ZN(n2822) );
  INV_X1 U2975 ( .A(n4543), .ZN(n4532) );
  NAND2_X1 U2976 ( .A1(n4147), .A2(n4532), .ZN(n4546) );
  AND2_X1 U2977 ( .A1(n2938), .A2(n2823), .ZN(n4543) );
  INV_X1 U2978 ( .A(n2822), .ZN(n2932) );
  AND2_X1 U2979 ( .A1(n2477), .A2(n2485), .ZN(n4523) );
  AND2_X1 U2980 ( .A1(n2782), .A2(n2775), .ZN(n4486) );
  INV_X1 U2981 ( .A(n3713), .ZN(n3692) );
  OR2_X1 U2982 ( .A1(n2851), .A2(n2845), .ZN(n3716) );
  NAND2_X1 U2983 ( .A1(n2609), .A2(n2608), .ZN(n4237) );
  OAI211_X1 U2984 ( .C1(n3603), .C2(n2596), .A(n2560), .B(n2559), .ZN(n4142)
         );
  NAND4_X1 U2985 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n3889)
         );
  INV_X1 U2986 ( .A(n4435), .ZN(n4482) );
  AOI21_X1 U2987 ( .B1(n2721), .B2(n2740), .A(n2720), .ZN(n2722) );
  NAND2_X1 U2988 ( .A1(n4564), .A2(n4537), .ZN(n4328) );
  INV_X1 U2989 ( .A(n4564), .ZN(n4561) );
  AOI21_X1 U2990 ( .B1(n2721), .B2(n2726), .A(n2725), .ZN(n2727) );
  NAND2_X1 U2991 ( .A1(n4554), .A2(n4537), .ZN(n4378) );
  INV_X1 U2992 ( .A(n4554), .ZN(n4552) );
  INV_X1 U2993 ( .A(n2696), .ZN(n2770) );
  AND2_X1 U2994 ( .A1(n2773), .A2(STATE_REG_SCAN_IN), .ZN(n4515) );
  OR2_X1 U2995 ( .A1(n2457), .A2(n2456), .ZN(n4526) );
  AND2_X1 U2996 ( .A1(n2419), .A2(n2429), .ZN(n4383) );
  INV_X1 U2997 ( .A(IR_REG_25__SCAN_IN), .ZN(n2312) );
  INV_X1 U2998 ( .A(DATAI_27_), .ZN(n2317) );
  NOR2_X1 U2999 ( .A1(n2487), .A2(n2317), .ZN(n4236) );
  INV_X1 U3000 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2536) );
  INV_X1 U3001 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U3002 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2318) );
  INV_X1 U3003 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4603) );
  INV_X1 U3004 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4690) );
  INV_X1 U3005 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3698) );
  INV_X1 U3006 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4580) );
  AND2_X1 U3007 ( .A1(n2603), .A2(n4580), .ZN(n2319) );
  INV_X1 U3008 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4024) );
  NAND2_X1 U3009 ( .A1(n3737), .A2(REG1_REG_27__SCAN_IN), .ZN(n2329) );
  INV_X1 U3010 ( .A(n2325), .ZN(n2327) );
  NAND2_X1 U3011 ( .A1(n2558), .A2(REG0_REG_27__SCAN_IN), .ZN(n2328) );
  OAI211_X1 U3012 ( .C1(n4024), .C2(n3738), .A(n2329), .B(n2328), .ZN(n2330)
         );
  INV_X1 U3013 ( .A(n2330), .ZN(n2331) );
  OAI21_X1 U3014 ( .B1(n4025), .B2(n2596), .A(n2331), .ZN(n4012) );
  INV_X1 U3015 ( .A(DATAI_25_), .ZN(n4590) );
  NOR2_X1 U3016 ( .A1(n2487), .A2(n4590), .ZN(n2664) );
  NAND2_X1 U3017 ( .A1(n2340), .A2(n4690), .ZN(n2332) );
  NAND2_X1 U3018 ( .A1(n2601), .A2(n2332), .ZN(n3622) );
  INV_X1 U3019 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2335) );
  NAND2_X1 U3020 ( .A1(n3737), .A2(REG1_REG_25__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U3021 ( .A1(n2558), .A2(REG0_REG_25__SCAN_IN), .ZN(n2333) );
  OAI211_X1 U3022 ( .C1(n2335), .C2(n3738), .A(n2334), .B(n2333), .ZN(n2336)
         );
  INV_X1 U3023 ( .A(n2336), .ZN(n2337) );
  OR2_X1 U3024 ( .A1(n2589), .A2(REG3_REG_24__SCAN_IN), .ZN(n2339) );
  NAND2_X1 U3025 ( .A1(n2340), .A2(n2339), .ZN(n3653) );
  INV_X1 U3026 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2343) );
  NAND2_X1 U3027 ( .A1(n3737), .A2(REG1_REG_24__SCAN_IN), .ZN(n2342) );
  NAND2_X1 U3028 ( .A1(n2558), .A2(REG0_REG_24__SCAN_IN), .ZN(n2341) );
  OAI211_X1 U3029 ( .C1(n2343), .C2(n3738), .A(n2342), .B(n2341), .ZN(n2344)
         );
  INV_X1 U3030 ( .A(n2344), .ZN(n2345) );
  NAND2_X1 U3031 ( .A1(n2046), .A2(DATAI_24_), .ZN(n4079) );
  NAND2_X1 U3032 ( .A1(n2354), .A2(REG1_REG_1__SCAN_IN), .ZN(n2352) );
  INV_X1 U3033 ( .A(n2364), .ZN(n2347) );
  INV_X1 U3034 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U3035 ( .A1(n2347), .A2(REG3_REG_1__SCAN_IN), .ZN(n2351) );
  INV_X1 U3036 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2785) );
  NAND2_X1 U3037 ( .A1(n2348), .A2(REG2_REG_1__SCAN_IN), .ZN(n2349) );
  INV_X1 U3038 ( .A(n2854), .ZN(n2859) );
  INV_X1 U3039 ( .A(n2854), .ZN(n3900) );
  NAND2_X1 U3040 ( .A1(n3900), .A2(n3070), .ZN(n2361) );
  NAND2_X1 U3041 ( .A1(n2859), .A2(n3078), .ZN(n3808) );
  NAND2_X1 U3042 ( .A1(n2354), .A2(REG1_REG_0__SCAN_IN), .ZN(n2360) );
  NAND2_X1 U3043 ( .A1(n2355), .A2(REG0_REG_0__SCAN_IN), .ZN(n2359) );
  INV_X1 U3044 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2849) );
  OR2_X1 U3045 ( .A1(n2364), .A2(n2849), .ZN(n2358) );
  INV_X1 U3046 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2356) );
  OR2_X1 U3047 ( .A1(n2363), .A2(n2356), .ZN(n2357) );
  NAND2_X1 U3048 ( .A1(n2361), .A2(n3074), .ZN(n3005) );
  NAND2_X1 U3049 ( .A1(n2354), .A2(REG1_REG_2__SCAN_IN), .ZN(n2368) );
  INV_X1 U3050 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2362) );
  NAND2_X1 U3051 ( .A1(n2355), .A2(REG0_REG_2__SCAN_IN), .ZN(n2366) );
  INV_X1 U3052 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2877) );
  OR2_X1 U3053 ( .A1(n2364), .A2(n2877), .ZN(n2365) );
  XNOR2_X2 U3054 ( .A(n2369), .B(IR_REG_2__SCAN_IN), .ZN(n4387) );
  MUX2_X1 U3055 ( .A(DATAI_2_), .B(n4387), .S(n2370), .Z(n3013) );
  INV_X1 U3056 ( .A(n3013), .ZN(n2869) );
  NAND2_X1 U3057 ( .A1(n3899), .A2(n2869), .ZN(n3815) );
  NAND2_X1 U3058 ( .A1(n3815), .A2(n3812), .ZN(n2640) );
  NAND2_X1 U3059 ( .A1(n2867), .A2(n2869), .ZN(n2371) );
  NAND2_X1 U3060 ( .A1(n3737), .A2(REG1_REG_3__SCAN_IN), .ZN(n2375) );
  NAND2_X1 U3061 ( .A1(n2558), .A2(REG0_REG_3__SCAN_IN), .ZN(n2374) );
  OR2_X1 U3062 ( .A1(n2596), .A2(REG3_REG_3__SCAN_IN), .ZN(n2373) );
  INV_X1 U3063 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2789) );
  OR2_X1 U3064 ( .A1(n3738), .A2(n2789), .ZN(n2372) );
  NAND2_X1 U3065 ( .A1(n2376), .A2(IR_REG_31__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3066 ( .A1(n2378), .A2(n2377), .ZN(n2390) );
  OR2_X1 U3067 ( .A1(n2378), .A2(n2377), .ZN(n2379) );
  MUX2_X1 U3068 ( .A(DATAI_3_), .B(n4386), .S(n2370), .Z(n2963) );
  NAND2_X1 U3069 ( .A1(n3898), .A2(n2963), .ZN(n2380) );
  NAND2_X1 U3070 ( .A1(n3036), .A2(n2968), .ZN(n2381) );
  INV_X1 U3071 ( .A(n3043), .ZN(n2393) );
  NAND2_X1 U3072 ( .A1(n2354), .A2(REG1_REG_4__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U3073 ( .A1(n2558), .A2(REG0_REG_4__SCAN_IN), .ZN(n2388) );
  INV_X1 U3074 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2383) );
  OR2_X1 U3075 ( .A1(n2363), .A2(n2383), .ZN(n2387) );
  INV_X1 U3076 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3061) );
  INV_X1 U3077 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2384) );
  NAND2_X1 U3078 ( .A1(n3061), .A2(n2384), .ZN(n2385) );
  NAND2_X1 U3079 ( .A1(n2396), .A2(n2385), .ZN(n3056) );
  OR2_X1 U3080 ( .A1(n2596), .A2(n3056), .ZN(n2386) );
  NAND2_X1 U3081 ( .A1(n2390), .A2(IR_REG_31__SCAN_IN), .ZN(n2391) );
  XNOR2_X1 U3082 ( .A(n2391), .B(IR_REG_4__SCAN_IN), .ZN(n4385) );
  MUX2_X1 U3083 ( .A(DATAI_4_), .B(n4385), .S(n3742), .Z(n3046) );
  NAND2_X1 U3084 ( .A1(n2982), .A2(n3046), .ZN(n3818) );
  INV_X1 U3085 ( .A(n3046), .ZN(n3054) );
  NAND2_X1 U3086 ( .A1(n3897), .A2(n3054), .ZN(n3821) );
  INV_X1 U3087 ( .A(n3772), .ZN(n2392) );
  NAND2_X1 U3088 ( .A1(n3897), .A2(n3046), .ZN(n2394) );
  NAND2_X1 U3089 ( .A1(n3737), .A2(REG1_REG_5__SCAN_IN), .ZN(n2402) );
  NAND2_X1 U3090 ( .A1(n2558), .A2(REG0_REG_5__SCAN_IN), .ZN(n2401) );
  INV_X1 U3091 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2395) );
  OR2_X1 U3092 ( .A1(n3738), .A2(n2395), .ZN(n2400) );
  INV_X1 U3093 ( .A(n2410), .ZN(n2398) );
  NAND2_X1 U3094 ( .A1(n2396), .A2(n2089), .ZN(n2397) );
  NAND2_X1 U3095 ( .A1(n2398), .A2(n2397), .ZN(n3137) );
  INV_X1 U3096 ( .A(DATAI_5_), .ZN(n4633) );
  NAND2_X1 U3097 ( .A1(n2404), .A2(IR_REG_31__SCAN_IN), .ZN(n2405) );
  MUX2_X1 U3098 ( .A(n2405), .B(IR_REG_31__SCAN_IN), .S(n2406), .Z(n2408) );
  INV_X1 U3099 ( .A(n2404), .ZN(n2407) );
  NAND2_X1 U3100 ( .A1(n2407), .A2(n2406), .ZN(n2416) );
  NAND2_X1 U3101 ( .A1(n2408), .A2(n2416), .ZN(n2796) );
  MUX2_X1 U3102 ( .A(n4633), .B(n2796), .S(n2487), .Z(n3132) );
  NAND2_X1 U3103 ( .A1(n3148), .A2(n3132), .ZN(n2409) );
  NAND2_X1 U3104 ( .A1(n3737), .A2(REG1_REG_6__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U3105 ( .A1(n2558), .A2(REG0_REG_6__SCAN_IN), .ZN(n2413) );
  INV_X1 U3106 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2995) );
  OR2_X1 U3107 ( .A1(n3738), .A2(n2995), .ZN(n2412) );
  OAI21_X1 U3108 ( .B1(n2410), .B2(REG3_REG_6__SCAN_IN), .A(n2423), .ZN(n3155)
         );
  OR2_X1 U3109 ( .A1(n2596), .A2(n3155), .ZN(n2411) );
  NAND4_X1 U3110 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .ZN(n3895)
         );
  NAND2_X1 U3111 ( .A1(n2416), .A2(IR_REG_31__SCAN_IN), .ZN(n2415) );
  MUX2_X1 U3112 ( .A(n2415), .B(IR_REG_31__SCAN_IN), .S(n2417), .Z(n2419) );
  INV_X1 U3113 ( .A(n2416), .ZN(n2418) );
  NAND2_X1 U3114 ( .A1(n2418), .A2(n2417), .ZN(n2429) );
  MUX2_X1 U3115 ( .A(DATAI_6_), .B(n4383), .S(n2487), .Z(n3145) );
  NAND2_X1 U3116 ( .A1(n3737), .A2(REG1_REG_7__SCAN_IN), .ZN(n2428) );
  NAND2_X1 U3117 ( .A1(n2558), .A2(REG0_REG_7__SCAN_IN), .ZN(n2427) );
  INV_X1 U3118 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2421) );
  OR2_X1 U3119 ( .A1(n3738), .A2(n2421), .ZN(n2426) );
  AND2_X1 U3120 ( .A1(n2423), .A2(n2422), .ZN(n2424) );
  OR2_X1 U3121 ( .A1(n2424), .A2(n2434), .ZN(n3171) );
  OR2_X1 U3122 ( .A1(n2596), .A2(n3171), .ZN(n2425) );
  NAND4_X1 U3123 ( .A1(n2428), .A2(n2427), .A3(n2426), .A4(n2425), .ZN(n3894)
         );
  NAND2_X1 U3124 ( .A1(n2429), .A2(IR_REG_31__SCAN_IN), .ZN(n2431) );
  NAND2_X1 U3125 ( .A1(n2431), .A2(n2430), .ZN(n2440) );
  OR2_X1 U3126 ( .A1(n2431), .A2(n2430), .ZN(n2432) );
  MUX2_X1 U3127 ( .A(DATAI_7_), .B(n4382), .S(n2487), .Z(n3115) );
  NAND2_X1 U3128 ( .A1(n3215), .A2(n3115), .ZN(n3828) );
  INV_X1 U3129 ( .A(n3115), .ZN(n3175) );
  NAND2_X1 U3130 ( .A1(n3894), .A2(n3175), .ZN(n3830) );
  OR2_X2 U3131 ( .A1(n3121), .A2(n3773), .ZN(n4548) );
  NAND2_X1 U3132 ( .A1(n3894), .A2(n3115), .ZN(n2433) );
  NAND2_X2 U3133 ( .A1(n4548), .A2(n2433), .ZN(n3220) );
  NAND2_X1 U3134 ( .A1(n3737), .A2(REG1_REG_8__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U3135 ( .A1(n2558), .A2(REG0_REG_8__SCAN_IN), .ZN(n2438) );
  INV_X1 U3136 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4496) );
  OR2_X1 U3137 ( .A1(n2434), .A2(REG3_REG_8__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U3138 ( .A1(n2447), .A2(n2435), .ZN(n4495) );
  OR2_X1 U3139 ( .A1(n2596), .A2(n4495), .ZN(n2436) );
  INV_X1 U3140 ( .A(DATAI_8_), .ZN(n2443) );
  NAND2_X1 U3141 ( .A1(n2440), .A2(IR_REG_31__SCAN_IN), .ZN(n2442) );
  XNOR2_X1 U3142 ( .A(n2442), .B(n2441), .ZN(n3952) );
  MUX2_X1 U3143 ( .A(n2443), .B(n3952), .S(n2487), .Z(n3213) );
  NAND2_X1 U3144 ( .A1(n3182), .A2(n3213), .ZN(n2444) );
  NAND2_X1 U3145 ( .A1(n3893), .A2(n3228), .ZN(n2445) );
  NAND2_X1 U3146 ( .A1(n3737), .A2(REG1_REG_9__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U3147 ( .A1(n2558), .A2(REG0_REG_9__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U31480 ( .A1(n2447), .A2(n2446), .ZN(n2448) );
  NAND2_X1 U31490 ( .A1(n2460), .A2(n2448), .ZN(n3252) );
  OR2_X1 U3150 ( .A1(n2596), .A2(n3252), .ZN(n2451) );
  INV_X1 U3151 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2449) );
  OR2_X1 U3152 ( .A1(n3738), .A2(n2449), .ZN(n2450) );
  NAND4_X1 U3153 ( .A1(n2453), .A2(n2452), .A3(n2451), .A4(n2450), .ZN(n3892)
         );
  NOR2_X1 U3154 ( .A1(n2162), .A2(n2760), .ZN(n2454) );
  MUX2_X1 U3155 ( .A(n2760), .B(n2454), .S(IR_REG_9__SCAN_IN), .Z(n2457) );
  NAND2_X1 U3156 ( .A1(n2162), .A2(n2455), .ZN(n2497) );
  INV_X1 U3157 ( .A(n2497), .ZN(n2456) );
  MUX2_X1 U3158 ( .A(DATAI_9_), .B(n3951), .S(n2487), .Z(n3248) );
  NAND2_X1 U3159 ( .A1(n3737), .A2(REG1_REG_10__SCAN_IN), .ZN(n2465) );
  NAND2_X1 U3160 ( .A1(n2558), .A2(REG0_REG_10__SCAN_IN), .ZN(n2464) );
  INV_X1 U3161 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2458) );
  OR2_X1 U3162 ( .A1(n3738), .A2(n2458), .ZN(n2463) );
  AND2_X1 U3163 ( .A1(n2460), .A2(n2459), .ZN(n2461) );
  OR2_X1 U3164 ( .A1(n2461), .A2(n2468), .ZN(n3298) );
  OR2_X1 U3165 ( .A1(n2596), .A2(n3298), .ZN(n2462) );
  NAND2_X1 U3166 ( .A1(n2497), .A2(IR_REG_31__SCAN_IN), .ZN(n2466) );
  XNOR2_X1 U3167 ( .A(n2466), .B(IR_REG_10__SCAN_IN), .ZN(n3957) );
  MUX2_X1 U3168 ( .A(DATAI_10_), .B(n3957), .S(n2487), .Z(n3284) );
  NOR2_X1 U3169 ( .A1(n3891), .A2(n3284), .ZN(n2467) );
  OAI22_X1 U3170 ( .A1(n3190), .A2(n2467), .B1(n3355), .B2(n3292), .ZN(n3333)
         );
  NAND2_X1 U3171 ( .A1(n3737), .A2(REG1_REG_11__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3172 ( .A1(n2558), .A2(REG0_REG_11__SCAN_IN), .ZN(n2472) );
  INV_X1 U3173 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3340) );
  OR2_X1 U3174 ( .A1(n3738), .A2(n3340), .ZN(n2471) );
  NOR2_X1 U3175 ( .A1(n2468), .A2(REG3_REG_11__SCAN_IN), .ZN(n2469) );
  OR2_X1 U3176 ( .A1(n2479), .A2(n2469), .ZN(n3339) );
  OR2_X1 U3177 ( .A1(n2596), .A2(n3339), .ZN(n2470) );
  NAND4_X1 U3178 ( .A1(n2473), .A2(n2472), .A3(n2471), .A4(n2470), .ZN(n3890)
         );
  OR2_X1 U3179 ( .A1(n2497), .A2(IR_REG_10__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3180 ( .A1(n2474), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  INV_X1 U3181 ( .A(IR_REG_11__SCAN_IN), .ZN(n2475) );
  OR2_X1 U3182 ( .A1(n2476), .A2(n2475), .ZN(n2477) );
  NAND2_X1 U3183 ( .A1(n2476), .A2(n2475), .ZN(n2485) );
  MUX2_X1 U3184 ( .A(DATAI_11_), .B(n4523), .S(n2487), .Z(n3334) );
  NAND2_X1 U3185 ( .A1(n3405), .A2(n3334), .ZN(n3268) );
  NAND2_X1 U3186 ( .A1(n3890), .A2(n3342), .ZN(n3270) );
  NAND2_X1 U3187 ( .A1(n3405), .A2(n3342), .ZN(n2478) );
  NAND2_X1 U3188 ( .A1(n3737), .A2(REG1_REG_12__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3189 ( .A1(n2558), .A2(REG0_REG_12__SCAN_IN), .ZN(n2483) );
  INV_X1 U3190 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3262) );
  OR2_X1 U3191 ( .A1(n2479), .A2(REG3_REG_12__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3192 ( .A1(n2489), .A2(n2480), .ZN(n3410) );
  OR2_X1 U3193 ( .A1(n2596), .A2(n3410), .ZN(n2481) );
  NAND2_X1 U3194 ( .A1(n2485), .A2(IR_REG_31__SCAN_IN), .ZN(n2486) );
  XNOR2_X1 U3195 ( .A(n2486), .B(IR_REG_12__SCAN_IN), .ZN(n3961) );
  MUX2_X1 U3196 ( .A(DATAI_12_), .B(n3961), .S(n3742), .Z(n3395) );
  INV_X1 U3197 ( .A(n3889), .ZN(n2647) );
  INV_X1 U3198 ( .A(n3395), .ZN(n3404) );
  INV_X1 U3199 ( .A(n3299), .ZN(n2499) );
  NAND2_X1 U3200 ( .A1(n3737), .A2(REG1_REG_13__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U3201 ( .A1(n2558), .A2(REG0_REG_13__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3202 ( .A1(n2489), .A2(n2488), .ZN(n2490) );
  NAND2_X1 U3203 ( .A1(n2501), .A2(n2490), .ZN(n3313) );
  OR2_X1 U3204 ( .A1(n2596), .A2(n3313), .ZN(n2492) );
  INV_X1 U3205 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4434) );
  OR2_X1 U3206 ( .A1(n3738), .A2(n4434), .ZN(n2491) );
  NAND4_X1 U3207 ( .A1(n2494), .A2(n2493), .A3(n2492), .A4(n2491), .ZN(n3888)
         );
  INV_X1 U3208 ( .A(n2495), .ZN(n2496) );
  NAND2_X1 U3209 ( .A1(n2507), .A2(IR_REG_31__SCAN_IN), .ZN(n2498) );
  XNOR2_X1 U32100 ( .A(n2498), .B(IR_REG_13__SCAN_IN), .ZN(n3949) );
  MUX2_X1 U32110 ( .A(DATAI_13_), .B(n3949), .S(n2487), .Z(n3451) );
  AOI21_X2 U32120 ( .B1(n2499), .B2(n2301), .A(n2300), .ZN(n3379) );
  NAND2_X1 U32130 ( .A1(n3737), .A2(REG1_REG_14__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U32140 ( .A1(n2558), .A2(REG0_REG_14__SCAN_IN), .ZN(n2505) );
  INV_X1 U32150 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2500) );
  OR2_X1 U32160 ( .A1(n3738), .A2(n2500), .ZN(n2504) );
  NAND2_X1 U32170 ( .A1(n2501), .A2(n4693), .ZN(n2502) );
  NAND2_X1 U32180 ( .A1(n2513), .A2(n2502), .ZN(n3584) );
  OR2_X1 U32190 ( .A1(n2596), .A2(n3584), .ZN(n2503) );
  NOR2_X1 U32200 ( .A1(n2507), .A2(IR_REG_13__SCAN_IN), .ZN(n2519) );
  OR2_X1 U32210 ( .A1(n2519), .A2(n2760), .ZN(n2508) );
  XNOR2_X1 U32220 ( .A(n2508), .B(IR_REG_14__SCAN_IN), .ZN(n3965) );
  MUX2_X1 U32230 ( .A(DATAI_14_), .B(n3965), .S(n2487), .Z(n3464) );
  NAND2_X1 U32240 ( .A1(n4324), .A2(n3464), .ZN(n3718) );
  NAND2_X1 U32250 ( .A1(n3887), .A2(n3577), .ZN(n3726) );
  NAND2_X1 U32260 ( .A1(n3718), .A2(n3726), .ZN(n3378) );
  NAND2_X1 U32270 ( .A1(n3379), .A2(n3378), .ZN(n3377) );
  NAND2_X1 U32280 ( .A1(n4324), .A2(n3577), .ZN(n2509) );
  NAND2_X1 U32290 ( .A1(n3377), .A2(n2509), .ZN(n3414) );
  INV_X1 U32300 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U32310 ( .A1(n3737), .A2(REG1_REG_15__SCAN_IN), .ZN(n2510) );
  OAI21_X1 U32320 ( .B1(n2511), .B2(n3738), .A(n2510), .ZN(n2517) );
  AND2_X1 U32330 ( .A1(n2513), .A2(n2512), .ZN(n2514) );
  OR2_X1 U32340 ( .A1(n2514), .A2(n2526), .ZN(n3417) );
  NAND2_X1 U32350 ( .A1(n2558), .A2(REG0_REG_15__SCAN_IN), .ZN(n2515) );
  OAI21_X1 U32360 ( .B1(n3417), .B2(n2596), .A(n2515), .ZN(n2516) );
  INV_X1 U32370 ( .A(IR_REG_14__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U32380 ( .A1(n2519), .A2(n2518), .ZN(n2520) );
  NAND2_X1 U32390 ( .A1(n2520), .A2(IR_REG_31__SCAN_IN), .ZN(n2522) );
  INV_X1 U32400 ( .A(IR_REG_15__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U32410 ( .A1(n2522), .A2(n2521), .ZN(n2532) );
  OR2_X1 U32420 ( .A1(n2522), .A2(n2521), .ZN(n2523) );
  MUX2_X1 U32430 ( .A(DATAI_15_), .B(n3948), .S(n3742), .Z(n4317) );
  NAND2_X1 U32440 ( .A1(n3886), .A2(n4317), .ZN(n2524) );
  AOI21_X1 U32450 ( .B1(n3414), .B2(n2524), .A(n2298), .ZN(n3435) );
  NAND2_X1 U32460 ( .A1(n3737), .A2(REG1_REG_16__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32470 ( .A1(n2558), .A2(REG0_REG_16__SCAN_IN), .ZN(n2530) );
  INV_X1 U32480 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2525) );
  OR2_X1 U32490 ( .A1(n3738), .A2(n2525), .ZN(n2529) );
  OR2_X1 U32500 ( .A1(n2526), .A2(REG3_REG_16__SCAN_IN), .ZN(n2527) );
  NAND2_X1 U32510 ( .A1(n2537), .A2(n2527), .ZN(n3440) );
  OR2_X1 U32520 ( .A1(n3440), .A2(n2596), .ZN(n2528) );
  NAND2_X1 U32530 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  XNOR2_X1 U32540 ( .A(n2533), .B(IR_REG_16__SCAN_IN), .ZN(n3969) );
  MUX2_X1 U32550 ( .A(DATAI_16_), .B(n3969), .S(n2487), .Z(n4307) );
  NAND2_X1 U32560 ( .A1(n4303), .A2(n4307), .ZN(n3848) );
  INV_X1 U32570 ( .A(n4307), .ZN(n3634) );
  NAND2_X1 U32580 ( .A1(n4320), .A2(n3634), .ZN(n3720) );
  NAND2_X1 U32590 ( .A1(n3435), .A2(n2534), .ZN(n3436) );
  NAND2_X1 U32600 ( .A1(n4320), .A2(n4307), .ZN(n2535) );
  NAND2_X1 U32610 ( .A1(n3436), .A2(n2535), .ZN(n4209) );
  NAND2_X1 U32620 ( .A1(n2537), .A2(n2536), .ZN(n2538) );
  NAND2_X1 U32630 ( .A1(n2055), .A2(n2538), .ZN(n3643) );
  NAND2_X1 U32640 ( .A1(n2558), .A2(REG0_REG_17__SCAN_IN), .ZN(n2539) );
  OAI21_X1 U32650 ( .B1(n3643), .B2(n2596), .A(n2539), .ZN(n2543) );
  INV_X1 U32660 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32670 ( .A1(n3737), .A2(REG1_REG_17__SCAN_IN), .ZN(n2540) );
  OAI21_X1 U32680 ( .B1(n2541), .B2(n3738), .A(n2540), .ZN(n2542) );
  INV_X1 U32690 ( .A(n4308), .ZN(n3687) );
  INV_X1 U32700 ( .A(DATAI_17_), .ZN(n4734) );
  OR2_X1 U32710 ( .A1(n2552), .A2(n2760), .ZN(n2544) );
  XNOR2_X1 U32720 ( .A(n2544), .B(IR_REG_17__SCAN_IN), .ZN(n3973) );
  MUX2_X1 U32730 ( .A(n4734), .B(n4517), .S(n2487), .Z(n4218) );
  NAND2_X1 U32740 ( .A1(n3687), .A2(n4218), .ZN(n2546) );
  AND2_X1 U32750 ( .A1(n4308), .A2(n4299), .ZN(n2545) );
  AND2_X1 U32760 ( .A1(n2055), .A2(n2547), .ZN(n2548) );
  OR2_X1 U32770 ( .A1(n2548), .A2(n2556), .ZN(n4197) );
  AOI22_X1 U32780 ( .A1(n2348), .A2(REG2_REG_18__SCAN_IN), .B1(n3737), .B2(
        REG1_REG_18__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32790 ( .A1(n2558), .A2(REG0_REG_18__SCAN_IN), .ZN(n2549) );
  OAI211_X1 U32800 ( .C1(n4197), .C2(n2596), .A(n2550), .B(n2549), .ZN(n4300)
         );
  INV_X1 U32810 ( .A(DATAI_18_), .ZN(n2554) );
  NAND2_X1 U32820 ( .A1(n2561), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  XNOR2_X1 U32830 ( .A(n2553), .B(IR_REG_18__SCAN_IN), .ZN(n3946) );
  MUX2_X1 U32840 ( .A(n2554), .B(n4516), .S(n2487), .Z(n4195) );
  OR2_X1 U32850 ( .A1(n4300), .A2(n4195), .ZN(n4163) );
  NAND2_X1 U32860 ( .A1(n4300), .A2(n4195), .ZN(n4164) );
  NAND2_X1 U32870 ( .A1(n4163), .A2(n4164), .ZN(n4184) );
  NAND2_X1 U32880 ( .A1(n4185), .A2(n4184), .ZN(n4183) );
  INV_X1 U32890 ( .A(n4195), .ZN(n4189) );
  OR2_X1 U32900 ( .A1(n4300), .A2(n4189), .ZN(n2555) );
  NOR2_X1 U32910 ( .A1(n2556), .A2(REG3_REG_19__SCAN_IN), .ZN(n2557) );
  OR2_X1 U32920 ( .A1(n2563), .A2(n2557), .ZN(n3603) );
  AOI22_X1 U32930 ( .A1(n2348), .A2(REG2_REG_19__SCAN_IN), .B1(n3737), .B2(
        REG1_REG_19__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U32940 ( .A1(n2558), .A2(REG0_REG_19__SCAN_IN), .ZN(n2559) );
  MUX2_X1 U32950 ( .A(DATAI_19_), .B(n4380), .S(n2487), .Z(n4174) );
  NAND2_X1 U32960 ( .A1(n4142), .A2(n4174), .ZN(n2562) );
  OR2_X1 U32970 ( .A1(n2563), .A2(REG3_REG_20__SCAN_IN), .ZN(n2564) );
  AND2_X1 U32980 ( .A1(n2578), .A2(n2564), .ZN(n4151) );
  NAND2_X1 U32990 ( .A1(n4151), .A2(n2347), .ZN(n2570) );
  INV_X1 U33000 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U33010 ( .A1(n2558), .A2(REG0_REG_20__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U33020 ( .A1(n3737), .A2(REG1_REG_20__SCAN_IN), .ZN(n2565) );
  OAI211_X1 U33030 ( .C1(n3738), .C2(n2567), .A(n2566), .B(n2565), .ZN(n2568)
         );
  INV_X1 U33040 ( .A(n2568), .ZN(n2569) );
  NAND2_X1 U33050 ( .A1(n2046), .A2(DATAI_20_), .ZN(n3665) );
  NAND2_X1 U33060 ( .A1(n4132), .A2(n3665), .ZN(n3782) );
  XNOR2_X1 U33070 ( .A(n2578), .B(REG3_REG_21__SCAN_IN), .ZN(n4130) );
  NAND2_X1 U33080 ( .A1(n4130), .A2(n2347), .ZN(n2576) );
  INV_X1 U33090 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U33100 ( .A1(n2558), .A2(REG0_REG_21__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U33110 ( .A1(n3737), .A2(REG1_REG_21__SCAN_IN), .ZN(n2571) );
  OAI211_X1 U33120 ( .C1(n3738), .C2(n2573), .A(n2572), .B(n2571), .ZN(n2574)
         );
  INV_X1 U33130 ( .A(n2574), .ZN(n2575) );
  NAND2_X1 U33140 ( .A1(n2046), .A2(DATAI_21_), .ZN(n4133) );
  INV_X1 U33150 ( .A(n4133), .ZN(n4277) );
  INV_X1 U33160 ( .A(n4109), .ZN(n4144) );
  INV_X1 U33170 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2577) );
  INV_X1 U33180 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3676) );
  OAI21_X1 U33190 ( .B1(n2578), .B2(n2577), .A(n3676), .ZN(n2579) );
  NAND2_X1 U33200 ( .A1(n2579), .A2(n2588), .ZN(n3674) );
  INV_X1 U33210 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U33220 ( .A1(n2558), .A2(REG0_REG_22__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U33230 ( .A1(n3737), .A2(REG1_REG_22__SCAN_IN), .ZN(n2580) );
  OAI211_X1 U33240 ( .C1(n3738), .C2(n2582), .A(n2581), .B(n2580), .ZN(n2583)
         );
  INV_X1 U33250 ( .A(n2583), .ZN(n2584) );
  NAND2_X1 U33260 ( .A1(n2046), .A2(DATAI_22_), .ZN(n4112) );
  NAND2_X1 U33270 ( .A1(n4283), .A2(n2586), .ZN(n4088) );
  NAND2_X1 U33280 ( .A1(n3884), .A2(n4112), .ZN(n2659) );
  NAND2_X1 U33290 ( .A1(n4088), .A2(n2659), .ZN(n4117) );
  AND2_X1 U33300 ( .A1(n2588), .A2(n4603), .ZN(n2590) );
  OR2_X1 U33310 ( .A1(n2590), .A2(n2589), .ZN(n3591) );
  INV_X1 U33320 ( .A(REG2_REG_23__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U33330 ( .A1(n3737), .A2(REG1_REG_23__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U33340 ( .A1(n2558), .A2(REG0_REG_23__SCAN_IN), .ZN(n2591) );
  OAI211_X1 U33350 ( .C1(n2593), .C2(n3738), .A(n2592), .B(n2591), .ZN(n2594)
         );
  INV_X1 U33360 ( .A(n2594), .ZN(n2595) );
  INV_X1 U33370 ( .A(n4259), .ZN(n4107) );
  NAND2_X1 U33380 ( .A1(n2046), .A2(DATAI_23_), .ZN(n4093) );
  NAND2_X1 U33390 ( .A1(n4107), .A2(n4093), .ZN(n2598) );
  AOI21_X1 U33400 ( .B1(n2664), .B2(n4246), .A(n2600), .ZN(n4042) );
  NAND2_X1 U33410 ( .A1(n2601), .A2(n3698), .ZN(n2602) );
  NAND2_X1 U33420 ( .A1(n4046), .A2(n2347), .ZN(n2609) );
  INV_X1 U33430 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U33440 ( .A1(n3737), .A2(REG1_REG_26__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U33450 ( .A1(n2355), .A2(REG0_REG_26__SCAN_IN), .ZN(n2604) );
  OAI211_X1 U33460 ( .C1(n2606), .C2(n3738), .A(n2605), .B(n2604), .ZN(n2607)
         );
  INV_X1 U33470 ( .A(n2607), .ZN(n2608) );
  NAND2_X1 U33480 ( .A1(n2046), .A2(DATAI_26_), .ZN(n4048) );
  INV_X1 U33490 ( .A(n4048), .ZN(n4245) );
  NAND2_X1 U33500 ( .A1(n4237), .A2(n4245), .ZN(n3761) );
  NOR2_X1 U33510 ( .A1(n4237), .A2(n4245), .ZN(n3762) );
  INV_X1 U33520 ( .A(n4236), .ZN(n4029) );
  OR2_X1 U3353 ( .A1(n2610), .A2(REG3_REG_28__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U33540 ( .A1(n2610), .A2(REG3_REG_28__SCAN_IN), .ZN(n3997) );
  NAND2_X1 U3355 ( .A1(n4005), .A2(n2347), .ZN(n2616) );
  INV_X1 U3356 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4007) );
  NAND2_X1 U3357 ( .A1(n2355), .A2(REG0_REG_28__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U3358 ( .A1(n3737), .A2(REG1_REG_28__SCAN_IN), .ZN(n2612) );
  OAI211_X1 U3359 ( .C1(n3738), .C2(n4007), .A(n2613), .B(n2612), .ZN(n2614)
         );
  INV_X1 U3360 ( .A(n2614), .ZN(n2615) );
  NOR2_X1 U3361 ( .A1(n2487), .A2(n4717), .ZN(n2737) );
  INV_X1 U3362 ( .A(n3736), .ZN(n2617) );
  INV_X1 U3363 ( .A(n2737), .ZN(n4008) );
  NAND2_X1 U3364 ( .A1(n4033), .A2(n4008), .ZN(n3747) );
  NAND2_X1 U3365 ( .A1(n2617), .A2(n3747), .ZN(n3806) );
  NAND2_X1 U3366 ( .A1(n2046), .A2(DATAI_29_), .ZN(n3995) );
  OR2_X1 U3367 ( .A1(n3997), .A2(n2596), .ZN(n2622) );
  INV_X1 U3368 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3994) );
  NAND2_X1 U3369 ( .A1(n2558), .A2(REG0_REG_29__SCAN_IN), .ZN(n2619) );
  NAND2_X1 U3370 ( .A1(n3737), .A2(REG1_REG_29__SCAN_IN), .ZN(n2618) );
  OAI211_X1 U3371 ( .C1(n3738), .C2(n3994), .A(n2619), .B(n2618), .ZN(n2620)
         );
  INV_X1 U3372 ( .A(n2620), .ZN(n2621) );
  NAND2_X1 U3373 ( .A1(n2622), .A2(n2621), .ZN(n3883) );
  XOR2_X1 U3374 ( .A(n3995), .B(n3883), .Z(n3993) );
  INV_X1 U3375 ( .A(n3993), .ZN(n2623) );
  INV_X1 U3376 ( .A(n2632), .ZN(n2624) );
  NOR2_X1 U3377 ( .A1(IR_REG_21__SCAN_IN), .A2(n2624), .ZN(n2625) );
  NAND2_X1 U3378 ( .A1(n2691), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  INV_X1 U3379 ( .A(IR_REG_22__SCAN_IN), .ZN(n2626) );
  INV_X1 U3380 ( .A(IR_REG_19__SCAN_IN), .ZN(n2628) );
  NAND2_X1 U3381 ( .A1(n2633), .A2(n2632), .ZN(n2634) );
  XNOR2_X1 U3382 ( .A(n3879), .B(n2855), .ZN(n2637) );
  INV_X1 U3383 ( .A(n4380), .ZN(n3981) );
  NAND2_X1 U3384 ( .A1(n2637), .A2(n3981), .ZN(n4147) );
  AND2_X1 U3385 ( .A1(n3872), .A2(n4380), .ZN(n2938) );
  INV_X1 U3386 ( .A(n3901), .ZN(n2852) );
  NAND2_X1 U3387 ( .A1(n2852), .A2(n3071), .ZN(n3807) );
  OR2_X1 U3388 ( .A1(n3768), .A2(n3807), .ZN(n2639) );
  NAND2_X1 U3389 ( .A1(n2639), .A2(n3811), .ZN(n3007) );
  NAND2_X1 U3390 ( .A1(n3007), .A2(n2224), .ZN(n3006) );
  NAND2_X1 U3391 ( .A1(n3006), .A2(n3812), .ZN(n2962) );
  NAND2_X1 U3392 ( .A1(n3036), .A2(n2963), .ZN(n3817) );
  NAND2_X1 U3393 ( .A1(n3898), .A2(n2968), .ZN(n3814) );
  AND2_X1 U3394 ( .A1(n3817), .A2(n3814), .ZN(n3770) );
  NAND2_X1 U3395 ( .A1(n2962), .A2(n3770), .ZN(n2641) );
  INV_X1 U3396 ( .A(n3818), .ZN(n2642) );
  NAND2_X1 U3397 ( .A1(n3148), .A2(n2984), .ZN(n3825) );
  AND2_X1 U3398 ( .A1(n3896), .A2(n3132), .ZN(n2977) );
  NAND2_X1 U3399 ( .A1(n3895), .A2(n3149), .ZN(n3823) );
  NAND2_X1 U3400 ( .A1(n2992), .A2(n3823), .ZN(n2643) );
  INV_X1 U3401 ( .A(n3895), .ZN(n3143) );
  NAND2_X1 U3402 ( .A1(n3143), .A2(n3145), .ZN(n3827) );
  INV_X1 U3403 ( .A(n3828), .ZN(n2644) );
  NAND2_X1 U3404 ( .A1(n3182), .A2(n3228), .ZN(n3833) );
  NAND2_X1 U3405 ( .A1(n3893), .A2(n3213), .ZN(n3829) );
  NAND2_X1 U3406 ( .A1(n2645), .A2(n3829), .ZN(n3157) );
  AND2_X1 U3407 ( .A1(n3892), .A2(n3255), .ZN(n3156) );
  NAND2_X1 U3408 ( .A1(n3293), .A2(n3248), .ZN(n3834) );
  NAND2_X1 U3409 ( .A1(n3891), .A2(n3292), .ZN(n3838) );
  NAND2_X1 U3410 ( .A1(n3355), .A2(n3284), .ZN(n3842) );
  NAND2_X1 U3411 ( .A1(n3889), .A2(n3404), .ZN(n3303) );
  NAND2_X1 U3412 ( .A1(n3888), .A2(n3456), .ZN(n3300) );
  NAND2_X1 U3413 ( .A1(n3303), .A2(n3300), .ZN(n2648) );
  INV_X1 U3414 ( .A(n3270), .ZN(n2646) );
  NOR2_X1 U3415 ( .A1(n2648), .A2(n2646), .ZN(n3839) );
  NAND2_X1 U3416 ( .A1(n3335), .A2(n3839), .ZN(n2651) );
  NAND2_X1 U3417 ( .A1(n2647), .A2(n3395), .ZN(n3305) );
  NAND2_X1 U3418 ( .A1(n3268), .A2(n3305), .ZN(n2650) );
  INV_X1 U3419 ( .A(n2648), .ZN(n2649) );
  NOR2_X1 U3420 ( .A1(n3888), .A2(n3456), .ZN(n3301) );
  AOI21_X1 U3421 ( .B1(n2650), .B2(n2649), .A(n3301), .ZN(n3844) );
  NAND2_X1 U3422 ( .A1(n2651), .A2(n3844), .ZN(n3719) );
  INV_X1 U3423 ( .A(n3378), .ZN(n3791) );
  NAND2_X1 U3424 ( .A1(n3719), .A2(n3791), .ZN(n2652) );
  NAND2_X1 U3425 ( .A1(n4310), .A2(n4317), .ZN(n3722) );
  NAND2_X1 U3426 ( .A1(n3886), .A2(n3711), .ZN(n3725) );
  NAND2_X1 U3427 ( .A1(n3722), .A2(n3725), .ZN(n3769) );
  INV_X1 U3428 ( .A(n4174), .ZN(n4169) );
  NAND2_X1 U3429 ( .A1(n4142), .A2(n4169), .ZN(n2653) );
  NAND2_X1 U3430 ( .A1(n2653), .A2(n4164), .ZN(n2654) );
  AND2_X1 U3431 ( .A1(n4308), .A2(n4218), .ZN(n4162) );
  OR2_X1 U3432 ( .A1(n2654), .A2(n4162), .ZN(n3727) );
  INV_X1 U3433 ( .A(n2654), .ZN(n2657) );
  NAND2_X1 U3434 ( .A1(n3687), .A2(n4299), .ZN(n4161) );
  NAND2_X1 U3435 ( .A1(n4163), .A2(n4161), .ZN(n2656) );
  NOR2_X1 U3436 ( .A1(n4142), .A2(n4169), .ZN(n2655) );
  AOI21_X1 U3437 ( .B1(n2657), .B2(n2656), .A(n2655), .ZN(n4139) );
  NAND2_X1 U3438 ( .A1(n4132), .A2(n4153), .ZN(n2658) );
  NAND2_X1 U3439 ( .A1(n4279), .A2(n3665), .ZN(n3729) );
  OR2_X1 U3440 ( .A1(n4109), .A2(n4133), .ZN(n4086) );
  AND2_X1 U3441 ( .A1(n4088), .A2(n4086), .ZN(n3856) );
  NAND2_X1 U3442 ( .A1(n4259), .A2(n4093), .ZN(n3765) );
  AND2_X1 U3443 ( .A1(n3765), .A2(n2659), .ZN(n3861) );
  AND2_X1 U3444 ( .A1(n4109), .A2(n4133), .ZN(n4087) );
  NAND2_X1 U3445 ( .A1(n4088), .A2(n4087), .ZN(n2660) );
  NAND2_X1 U3446 ( .A1(n3861), .A2(n2660), .ZN(n3734) );
  INV_X1 U3447 ( .A(n3734), .ZN(n2661) );
  NAND2_X1 U3448 ( .A1(n2662), .A2(n2661), .ZN(n2663) );
  OR2_X1 U3449 ( .A1(n4259), .A2(n4093), .ZN(n3766) );
  NAND2_X1 U3450 ( .A1(n2663), .A2(n3766), .ZN(n4070) );
  NOR2_X1 U3451 ( .A1(n4095), .A2(n4079), .ZN(n3780) );
  NAND2_X1 U3452 ( .A1(n4262), .A2(n2664), .ZN(n4038) );
  OAI21_X1 U3453 ( .B1(n4237), .B2(n4048), .A(n4038), .ZN(n3859) );
  INV_X1 U3454 ( .A(n3859), .ZN(n3752) );
  NAND2_X1 U3455 ( .A1(n4246), .A2(n4062), .ZN(n3764) );
  NAND2_X1 U3456 ( .A1(n4095), .A2(n4079), .ZN(n3779) );
  AND2_X1 U3457 ( .A1(n3764), .A2(n3779), .ZN(n4037) );
  OR2_X1 U34580 ( .A1(n4037), .A2(n3859), .ZN(n2665) );
  NAND2_X1 U34590 ( .A1(n4237), .A2(n4048), .ZN(n3748) );
  NAND2_X1 U3460 ( .A1(n2665), .A2(n3748), .ZN(n3864) );
  XNOR2_X1 U3461 ( .A(n4012), .B(n4236), .ZN(n4022) );
  NOR2_X1 U3462 ( .A1(n4012), .A2(n4029), .ZN(n3735) );
  AOI21_X1 U3463 ( .B1(n2731), .B2(n3747), .A(n3736), .ZN(n2666) );
  XNOR2_X1 U3464 ( .A(n2666), .B(n3993), .ZN(n2680) );
  NAND2_X1 U3465 ( .A1(n3879), .A2(n4380), .ZN(n2668) );
  INV_X1 U3466 ( .A(n3872), .ZN(n2754) );
  NAND2_X1 U34670 ( .A1(n2667), .A2(n2754), .ZN(n3755) );
  NAND2_X1 U3468 ( .A1(n3737), .A2(REG1_REG_30__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U34690 ( .A1(n2558), .A2(REG0_REG_30__SCAN_IN), .ZN(n2671) );
  INV_X1 U3470 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2669) );
  OR2_X1 U34710 ( .A1(n3738), .A2(n2669), .ZN(n2670) );
  AND3_X1 U3472 ( .A1(n2672), .A2(n2671), .A3(n2670), .ZN(n3756) );
  INV_X1 U34730 ( .A(B_REG_SCAN_IN), .ZN(n2679) );
  OR2_X1 U3474 ( .A1(n2674), .A2(n2673), .ZN(n3902) );
  NOR2_X1 U34750 ( .A1(n2675), .A2(n2760), .ZN(n2676) );
  MUX2_X1 U3476 ( .A(n2760), .B(n2676), .S(IR_REG_28__SCAN_IN), .Z(n2678) );
  OR2_X1 U34770 ( .A1(n2678), .A2(n2677), .ZN(n2886) );
  NAND2_X1 U3478 ( .A1(n3879), .A2(n2667), .ZN(n2828) );
  INV_X1 U34790 ( .A(n2828), .ZN(n2774) );
  OAI21_X1 U3480 ( .B1(n2679), .B2(n3902), .A(n4319), .ZN(n3987) );
  OAI22_X1 U34810 ( .A1(n2680), .A2(n4172), .B1(n3756), .B2(n3987), .ZN(n4000)
         );
  INV_X1 U3482 ( .A(n4000), .ZN(n2683) );
  INV_X1 U34830 ( .A(n2886), .ZN(n2883) );
  NAND2_X1 U3484 ( .A1(n2883), .A2(n2774), .ZN(n4323) );
  NAND2_X1 U34850 ( .A1(n2823), .A2(n3798), .ZN(n2827) );
  OR2_X1 U3486 ( .A1(n2827), .A2(n3872), .ZN(n4168) );
  OAI22_X1 U34870 ( .A1(n4240), .A2(n4323), .B1(n3995), .B2(n4168), .ZN(n2681)
         );
  INV_X1 U3488 ( .A(n2681), .ZN(n2682) );
  NAND2_X1 U34890 ( .A1(n2683), .A2(n2682), .ZN(n2684) );
  NAND2_X1 U3490 ( .A1(n2688), .A2(IR_REG_31__SCAN_IN), .ZN(n2689) );
  MUX2_X1 U34910 ( .A(IR_REG_31__SCAN_IN), .B(n2689), .S(IR_REG_25__SCAN_IN), 
        .Z(n2690) );
  NAND2_X1 U3492 ( .A1(n2690), .A2(n2686), .ZN(n2750) );
  NAND2_X1 U34930 ( .A1(n2750), .A2(B_REG_SCAN_IN), .ZN(n2694) );
  NAND2_X1 U3494 ( .A1(n2698), .A2(n2699), .ZN(n2692) );
  MUX2_X1 U34950 ( .A(n2694), .B(B_REG_SCAN_IN), .S(n2696), .Z(n2695) );
  NAND2_X1 U3496 ( .A1(n2769), .A2(n2750), .ZN(n2820) );
  NAND2_X1 U34970 ( .A1(n2929), .A2(n2820), .ZN(n2713) );
  NOR2_X1 U3498 ( .A1(n2769), .A2(n2750), .ZN(n2697) );
  XNOR2_X1 U34990 ( .A(n2698), .B(n2699), .ZN(n2773) );
  NAND2_X1 U3500 ( .A1(n4543), .A2(n3798), .ZN(n2834) );
  AND2_X1 U35010 ( .A1(n3872), .A2(n3981), .ZN(n2826) );
  OR2_X1 U3502 ( .A1(n2828), .A2(n2826), .ZN(n2926) );
  NAND2_X1 U35030 ( .A1(n2834), .A2(n2926), .ZN(n2700) );
  NOR2_X1 U3504 ( .A1(n2928), .A2(n2700), .ZN(n2712) );
  NOR4_X1 U35050 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2704) );
  NOR4_X1 U35060 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2703) );
  NOR4_X1 U35070 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2702) );
  NOR4_X1 U35080 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2701) );
  NAND4_X1 U35090 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n2710)
         );
  NOR2_X1 U35100 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2708) );
  NOR4_X1 U35110 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2707) );
  NOR4_X1 U35120 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2706) );
  NOR4_X1 U35130 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2705) );
  NAND4_X1 U35140 ( .A1(n2708), .A2(n2707), .A3(n2706), .A4(n2705), .ZN(n2709)
         );
  NOR2_X1 U35150 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  NAND2_X1 U35160 ( .A1(n2770), .A2(n2769), .ZN(n2714) );
  AND2_X2 U35170 ( .A1(n2723), .A2(n2822), .ZN(n4564) );
  NAND2_X1 U35180 ( .A1(n3078), .A2(n2925), .ZN(n3068) );
  OR2_X2 U35190 ( .A1(n3116), .A2(n3115), .ZN(n3227) );
  OR2_X2 U35200 ( .A1(n4194), .A2(n4174), .ZN(n4176) );
  INV_X1 U35210 ( .A(n2739), .ZN(n2717) );
  INV_X1 U35220 ( .A(n3995), .ZN(n2716) );
  NAND2_X1 U35230 ( .A1(n2717), .A2(n2716), .ZN(n2718) );
  NAND2_X1 U35240 ( .A1(n4231), .A2(n2718), .ZN(n3998) );
  INV_X1 U35250 ( .A(n2827), .ZN(n2936) );
  INV_X1 U35260 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2719) );
  OAI21_X1 U35270 ( .B1(n2728), .B2(n4561), .A(n2722), .ZN(U3547) );
  INV_X1 U35280 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2724) );
  OAI21_X1 U35290 ( .B1(n2728), .B2(n4552), .A(n2727), .ZN(U3515) );
  INV_X1 U35300 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2736) );
  XNOR2_X1 U35310 ( .A(n2731), .B(n3806), .ZN(n2732) );
  NOR2_X1 U35320 ( .A1(n2732), .A2(n4172), .ZN(n4016) );
  AOI22_X1 U35330 ( .A1(n3883), .A2(n4319), .B1(n2737), .B2(n4318), .ZN(n2733)
         );
  OAI21_X1 U35340 ( .B1(n4249), .B2(n4323), .A(n2733), .ZN(n2734) );
  INV_X1 U35350 ( .A(n2734), .ZN(n2735) );
  MUX2_X1 U35360 ( .A(n2736), .B(n2744), .S(n4564), .Z(n2743) );
  AND2_X1 U35370 ( .A1(n2059), .A2(n2737), .ZN(n2738) );
  OR2_X1 U35380 ( .A1(n2739), .A2(n2738), .ZN(n4014) );
  INV_X1 U35390 ( .A(n4014), .ZN(n2741) );
  NAND2_X1 U35400 ( .A1(n2743), .A2(n2742), .ZN(U3546) );
  INV_X1 U35410 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2745) );
  NAND2_X1 U35420 ( .A1(n2747), .A2(n2746), .ZN(U3514) );
  INV_X2 U35430 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U35440 ( .A(n4515), .ZN(n2748) );
  INV_X2 U35450 ( .A(n3885), .ZN(U4043) );
  NAND2_X1 U35460 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2749) );
  OAI21_X1 U35470 ( .B1(n2750), .B2(U3149), .A(n2749), .ZN(U3327) );
  INV_X1 U35480 ( .A(DATAI_26_), .ZN(n4578) );
  NAND2_X1 U35490 ( .A1(n2751), .A2(STATE_REG_SCAN_IN), .ZN(n2752) );
  OAI21_X1 U35500 ( .B1(STATE_REG_SCAN_IN), .B2(n4578), .A(n2752), .ZN(U3326)
         );
  INV_X1 U35510 ( .A(DATAI_22_), .ZN(n4589) );
  NAND2_X1 U35520 ( .A1(n3879), .A2(STATE_REG_SCAN_IN), .ZN(n2753) );
  OAI21_X1 U35530 ( .B1(STATE_REG_SCAN_IN), .B2(n4589), .A(n2753), .ZN(U3330)
         );
  INV_X1 U35540 ( .A(DATAI_20_), .ZN(n4716) );
  NAND2_X1 U35550 ( .A1(n2754), .A2(STATE_REG_SCAN_IN), .ZN(n2755) );
  OAI21_X1 U35560 ( .B1(STATE_REG_SCAN_IN), .B2(n4716), .A(n2755), .ZN(U3332)
         );
  INV_X1 U35570 ( .A(DATAI_24_), .ZN(n4728) );
  NAND2_X1 U35580 ( .A1(n2696), .A2(STATE_REG_SCAN_IN), .ZN(n2756) );
  OAI21_X1 U35590 ( .B1(STATE_REG_SCAN_IN), .B2(n4728), .A(n2756), .ZN(U3328)
         );
  INV_X1 U35600 ( .A(n3902), .ZN(n2887) );
  NAND2_X1 U35610 ( .A1(n2887), .A2(STATE_REG_SCAN_IN), .ZN(n2757) );
  OAI21_X1 U35620 ( .B1(STATE_REG_SCAN_IN), .B2(n2317), .A(n2757), .ZN(U3325)
         );
  INV_X1 U35630 ( .A(DATAI_29_), .ZN(n4601) );
  NAND2_X1 U35640 ( .A1(n2758), .A2(STATE_REG_SCAN_IN), .ZN(n2759) );
  OAI21_X1 U35650 ( .B1(STATE_REG_SCAN_IN), .B2(n4601), .A(n2759), .ZN(U3323)
         );
  INV_X1 U35660 ( .A(DATAI_31_), .ZN(n4704) );
  OR4_X1 U35670 ( .A1(n2321), .A2(IR_REG_30__SCAN_IN), .A3(n2760), .A4(U3149), 
        .ZN(n2761) );
  OAI21_X1 U35680 ( .B1(STATE_REG_SCAN_IN), .B2(n4704), .A(n2761), .ZN(U3321)
         );
  INV_X1 U35690 ( .A(DATAI_30_), .ZN(n4568) );
  NAND2_X1 U35700 ( .A1(n2325), .A2(STATE_REG_SCAN_IN), .ZN(n2762) );
  OAI21_X1 U35710 ( .B1(STATE_REG_SCAN_IN), .B2(n4568), .A(n2762), .ZN(U3322)
         );
  INV_X1 U35720 ( .A(DATAI_28_), .ZN(n4717) );
  NAND2_X1 U35730 ( .A1(n2883), .A2(STATE_REG_SCAN_IN), .ZN(n2763) );
  OAI21_X1 U35740 ( .B1(STATE_REG_SCAN_IN), .B2(n4717), .A(n2763), .ZN(U3324)
         );
  NAND2_X1 U35750 ( .A1(n3885), .A2(DATAO_REG_30__SCAN_IN), .ZN(n2764) );
  OAI21_X1 U35760 ( .B1(n3885), .B2(n3756), .A(n2764), .ZN(U3580) );
  INV_X1 U35770 ( .A(n2928), .ZN(n2765) );
  INV_X1 U35780 ( .A(D_REG_1__SCAN_IN), .ZN(n2768) );
  INV_X1 U35790 ( .A(n2820), .ZN(n2767) );
  AOI22_X1 U35800 ( .A1(n4514), .A2(n2768), .B1(n2767), .B2(n4515), .ZN(U3459)
         );
  INV_X1 U35810 ( .A(D_REG_0__SCAN_IN), .ZN(n2772) );
  AND2_X1 U3582 ( .A1(n4515), .A2(n2769), .ZN(n2771) );
  AOI22_X1 U3583 ( .A1(n4514), .A2(n2772), .B1(n2771), .B2(n2770), .ZN(U3458)
         );
  OR2_X1 U3584 ( .A1(n2773), .A2(U3149), .ZN(n3881) );
  NAND2_X1 U3585 ( .A1(n2928), .A2(n3881), .ZN(n2782) );
  AOI21_X1 U3586 ( .B1(n2774), .B2(n2773), .A(n3742), .ZN(n2781) );
  INV_X1 U3587 ( .A(n2781), .ZN(n2775) );
  NOR2_X1 U3588 ( .A1(n4486), .A2(U4043), .ZN(U3148) );
  XNOR2_X1 U3589 ( .A(n4388), .B(n4557), .ZN(n3915) );
  AND2_X1 U3590 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3914)
         );
  NAND2_X1 U3591 ( .A1(n3915), .A2(n3914), .ZN(n3913) );
  NAND2_X1 U3592 ( .A1(n4388), .A2(REG1_REG_1__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U3593 ( .A1(n3913), .A2(n2776), .ZN(n2892) );
  INV_X1 U3594 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3016) );
  XNOR2_X1 U3595 ( .A(n4387), .B(n3016), .ZN(n2893) );
  NAND2_X1 U3596 ( .A1(n2892), .A2(n2893), .ZN(n2891) );
  NAND2_X1 U3597 ( .A1(n4387), .A2(REG1_REG_2__SCAN_IN), .ZN(n2777) );
  XNOR2_X1 U3598 ( .A(n2778), .B(n2787), .ZN(n3922) );
  NAND2_X1 U3599 ( .A1(n3922), .A2(REG1_REG_3__SCAN_IN), .ZN(n3921) );
  NAND2_X1 U3600 ( .A1(n2778), .A2(n4386), .ZN(n2779) );
  INV_X1 U3601 ( .A(n4385), .ZN(n2920) );
  XNOR2_X1 U3602 ( .A(n2780), .B(n2920), .ZN(n2916) );
  XOR2_X1 U3603 ( .A(REG1_REG_5__SCAN_IN), .B(n2796), .Z(n2783) );
  INV_X1 U3604 ( .A(n4488), .ZN(n2800) );
  AOI211_X1 U3605 ( .C1(n2784), .C2(n2783), .A(n2799), .B(n2800), .ZN(n2795)
         );
  AND2_X1 U3606 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2786)
         );
  NAND2_X1 U3607 ( .A1(n3912), .A2(n2786), .ZN(n3911) );
  NAND2_X1 U3608 ( .A1(n4388), .A2(REG2_REG_1__SCAN_IN), .ZN(n2896) );
  MUX2_X1 U3609 ( .A(n2362), .B(REG2_REG_2__SCAN_IN), .S(n4387), .Z(n2895) );
  AOI21_X1 U3610 ( .B1(n3911), .B2(n2896), .A(n2895), .ZN(n2894) );
  AOI21_X1 U3611 ( .B1(n4387), .B2(REG2_REG_2__SCAN_IN), .A(n2894), .ZN(n2788)
         );
  XNOR2_X1 U3612 ( .A(n2788), .B(n2787), .ZN(n3923) );
  MUX2_X1 U3613 ( .A(REG2_REG_5__SCAN_IN), .B(n2395), .S(n2796), .Z(n2790) );
  NOR2_X1 U3614 ( .A1(n2886), .A2(n3902), .ZN(n3876) );
  AOI211_X1 U3615 ( .C1(n2791), .C2(n2790), .A(n2797), .B(n4482), .ZN(n2794)
         );
  NAND2_X1 U3616 ( .A1(n3906), .A2(n2886), .ZN(n4493) );
  NOR2_X1 U3617 ( .A1(STATE_REG_SCAN_IN), .A2(n2089), .ZN(n3134) );
  AOI21_X1 U3618 ( .B1(n4486), .B2(ADDR_REG_5__SCAN_IN), .A(n3134), .ZN(n2792)
         );
  OAI21_X1 U3619 ( .B1(n4493), .B2(n2796), .A(n2792), .ZN(n2793) );
  OR3_X1 U3620 ( .A1(n2795), .A2(n2794), .A3(n2793), .ZN(U3245) );
  INV_X1 U3621 ( .A(n2796), .ZN(n4384) );
  XNOR2_X1 U3622 ( .A(n2813), .B(REG2_REG_6__SCAN_IN), .ZN(n2805) );
  INV_X1 U3623 ( .A(n4493), .ZN(n3920) );
  NAND2_X1 U3624 ( .A1(n4486), .A2(ADDR_REG_6__SCAN_IN), .ZN(n2798) );
  NAND2_X1 U3625 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U3626 ( .A1(n2798), .A2(n3150), .ZN(n2803) );
  INV_X1 U3627 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3094) );
  AOI211_X1 U3628 ( .C1(n2801), .C2(n3094), .A(n2800), .B(n2807), .ZN(n2802)
         );
  AOI211_X1 U3629 ( .C1(n3920), .C2(n4383), .A(n2803), .B(n2802), .ZN(n2804)
         );
  OAI21_X1 U3630 ( .B1(n2805), .B2(n4482), .A(n2804), .ZN(U3246) );
  INV_X1 U3631 ( .A(n2806), .ZN(n2808) );
  INV_X1 U3632 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4562) );
  MUX2_X1 U3633 ( .A(REG1_REG_7__SCAN_IN), .B(n4562), .S(n4382), .Z(n2809) );
  XNOR2_X1 U3634 ( .A(n2905), .B(n2809), .ZN(n2818) );
  INV_X1 U3635 ( .A(n4382), .ZN(n2903) );
  AND2_X1 U3636 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3172) );
  AOI21_X1 U3637 ( .B1(n4486), .B2(ADDR_REG_7__SCAN_IN), .A(n3172), .ZN(n2810)
         );
  OAI21_X1 U3638 ( .B1(n4493), .B2(n2903), .A(n2810), .ZN(n2817) );
  INV_X1 U3639 ( .A(n2811), .ZN(n2812) );
  AOI22_X1 U3640 ( .A1(n2813), .A2(REG2_REG_6__SCAN_IN), .B1(n4383), .B2(n2812), .ZN(n2815) );
  MUX2_X1 U3641 ( .A(n2421), .B(REG2_REG_7__SCAN_IN), .S(n4382), .Z(n2814) );
  NOR2_X1 U3642 ( .A1(n2815), .A2(n2814), .ZN(n2907) );
  AOI211_X1 U3643 ( .C1(n2815), .C2(n2814), .A(n4482), .B(n2907), .ZN(n2816)
         );
  AOI211_X1 U3644 ( .C1(n4488), .C2(n2818), .A(n2817), .B(n2816), .ZN(n2819)
         );
  INV_X1 U3645 ( .A(n2819), .ZN(U3247) );
  NAND3_X1 U3646 ( .A1(n2931), .A2(n2822), .A3(n2929), .ZN(n2851) );
  INV_X1 U3647 ( .A(n2856), .ZN(n2824) );
  NAND2_X1 U3648 ( .A1(n4515), .A2(n2824), .ZN(n2825) );
  NOR2_X1 U3649 ( .A1(n2049), .A2(n2825), .ZN(n3877) );
  NAND2_X1 U3650 ( .A1(n2851), .A2(n3877), .ZN(n2954) );
  INV_X1 U3651 ( .A(n2954), .ZN(n2832) );
  OR2_X1 U3652 ( .A1(n2827), .A2(n2826), .ZN(n2829) );
  NAND2_X1 U3653 ( .A1(n2829), .A2(n2828), .ZN(n2844) );
  NAND2_X1 U3654 ( .A1(n2844), .A2(n4168), .ZN(n2830) );
  NAND2_X1 U3655 ( .A1(n2851), .A2(n2830), .ZN(n2831) );
  NAND2_X1 U3656 ( .A1(n2831), .A2(n2926), .ZN(n2953) );
  NOR3_X1 U3657 ( .A1(n2832), .A2(n2953), .A3(n2928), .ZN(n2878) );
  OR2_X1 U3658 ( .A1(n2928), .A2(n4168), .ZN(n2833) );
  OR2_X1 U3659 ( .A1(n2851), .A2(n2833), .ZN(n2835) );
  AND2_X2 U3660 ( .A1(n2835), .A2(n4494), .ZN(n3675) );
  INV_X1 U3661 ( .A(n3675), .ZN(n3590) );
  INV_X1 U3662 ( .A(n2836), .ZN(n2952) );
  NAND2_X1 U3663 ( .A1(n2952), .A2(REG1_REG_0__SCAN_IN), .ZN(n2837) );
  NAND2_X1 U3664 ( .A1(n3901), .A2(n3542), .ZN(n2838) );
  NAND2_X1 U3665 ( .A1(n2839), .A2(n2838), .ZN(n2843) );
  NAND2_X1 U3666 ( .A1(n3023), .A2(n3901), .ZN(n2841) );
  AOI22_X1 U3667 ( .A1(n3542), .A2(n3071), .B1(n2952), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2840) );
  NAND2_X1 U3668 ( .A1(n2841), .A2(n2840), .ZN(n2842) );
  OAI21_X1 U3669 ( .B1(n2843), .B2(n2842), .A(n2861), .ZN(n2884) );
  OR2_X1 U3670 ( .A1(n2928), .A2(n2844), .ZN(n2845) );
  NAND2_X1 U3671 ( .A1(n3877), .A2(n2886), .ZN(n2846) );
  OAI22_X1 U3672 ( .A1(n2884), .A2(n3716), .B1(n3700), .B2(n2854), .ZN(n2847)
         );
  AOI21_X1 U3673 ( .B1(n3071), .B2(n3590), .A(n2847), .ZN(n2848) );
  OAI21_X1 U3674 ( .B1(n2878), .B2(n2849), .A(n2848), .ZN(U3229) );
  NAND2_X1 U3675 ( .A1(n3877), .A2(n2883), .ZN(n2850) );
  OAI22_X1 U3676 ( .A1(n2852), .A2(n3699), .B1(n3700), .B2(n2867), .ZN(n2853)
         );
  AOI21_X1 U3677 ( .B1(n3070), .B2(n3590), .A(n2853), .ZN(n2866) );
  NOR2_X1 U3678 ( .A1(n3499), .A2(n3078), .ZN(n2858) );
  XNOR2_X1 U3679 ( .A(n2870), .B(n2871), .ZN(n2863) );
  INV_X1 U3680 ( .A(n2860), .ZN(n2862) );
  OAI21_X1 U3681 ( .B1(n2862), .B2(n2050), .A(n2861), .ZN(n2864) );
  NAND2_X1 U3682 ( .A1(n2863), .A2(n2864), .ZN(n2874) );
  OAI211_X1 U3683 ( .C1(n2863), .C2(n2864), .A(n2874), .B(n3685), .ZN(n2865)
         );
  OAI211_X1 U3684 ( .C1(n2878), .C2(n3075), .A(n2866), .B(n2865), .ZN(U3219)
         );
  AOI21_X1 U3685 ( .B1(n2876), .B2(n2875), .A(n2944), .ZN(n2882) );
  OAI22_X1 U3686 ( .A1(n3036), .A2(n3700), .B1(n3699), .B2(n2854), .ZN(n2880)
         );
  NOR2_X1 U3687 ( .A1(n2878), .A2(n2877), .ZN(n2879) );
  AOI211_X1 U3688 ( .C1(n3013), .C2(n3590), .A(n2880), .B(n2879), .ZN(n2881)
         );
  OAI21_X1 U3689 ( .B1(n2882), .B2(n3716), .A(n2881), .ZN(U3234) );
  OAI21_X1 U3690 ( .B1(REG2_REG_0__SCAN_IN), .B2(n3902), .A(n2883), .ZN(n3904)
         );
  NAND2_X1 U3691 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3910) );
  NOR2_X1 U3692 ( .A1(n2884), .A2(n2887), .ZN(n2885) );
  AOI211_X1 U3693 ( .C1(n2887), .C2(n3910), .A(n2886), .B(n2885), .ZN(n2888)
         );
  INV_X1 U3694 ( .A(n4387), .ZN(n2890) );
  AOI22_X1 U3695 ( .A1(n4486), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2889) );
  OAI21_X1 U3696 ( .B1(n4493), .B2(n2890), .A(n2889), .ZN(n2902) );
  OAI211_X1 U3697 ( .C1(n2893), .C2(n2892), .A(n4488), .B(n2891), .ZN(n2900)
         );
  INV_X1 U3698 ( .A(n2894), .ZN(n2898) );
  NAND3_X1 U3699 ( .A1(n3911), .A2(n2896), .A3(n2895), .ZN(n2897) );
  NAND3_X1 U3700 ( .A1(n4435), .A2(n2898), .A3(n2897), .ZN(n2899) );
  NAND2_X1 U3701 ( .A1(n2900), .A2(n2899), .ZN(n2901) );
  OR3_X1 U3702 ( .A1(n2921), .A2(n2902), .A3(n2901), .ZN(U3242) );
  NOR2_X1 U3703 ( .A1(n4382), .A2(REG1_REG_7__SCAN_IN), .ZN(n2904) );
  XOR2_X1 U3704 ( .A(REG1_REG_8__SCAN_IN), .B(n3954), .Z(n2906) );
  NAND2_X1 U3705 ( .A1(n2906), .A2(n4488), .ZN(n2912) );
  XNOR2_X1 U3706 ( .A(REG2_REG_8__SCAN_IN), .B(n3932), .ZN(n2908) );
  NAND2_X1 U3707 ( .A1(n4435), .A2(n2908), .ZN(n2909) );
  NAND2_X1 U3708 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3214) );
  NAND2_X1 U3709 ( .A1(n2909), .A2(n3214), .ZN(n2910) );
  AOI21_X1 U3710 ( .B1(n4486), .B2(ADDR_REG_8__SCAN_IN), .A(n2910), .ZN(n2911)
         );
  OAI211_X1 U3711 ( .C1(n4493), .C2(n3952), .A(n2912), .B(n2911), .ZN(U3248)
         );
  XOR2_X1 U3712 ( .A(REG2_REG_4__SCAN_IN), .B(n2913), .Z(n2923) );
  INV_X1 U3713 ( .A(n2914), .ZN(n2915) );
  OAI211_X1 U3714 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2916), .A(n4488), .B(n2915), 
        .ZN(n2919) );
  NAND2_X1 U3715 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3037) );
  INV_X1 U3716 ( .A(n3037), .ZN(n2917) );
  AOI21_X1 U3717 ( .B1(n4486), .B2(ADDR_REG_4__SCAN_IN), .A(n2917), .ZN(n2918)
         );
  OAI211_X1 U3718 ( .C1(n4493), .C2(n2920), .A(n2919), .B(n2918), .ZN(n2922)
         );
  AOI211_X1 U3719 ( .C1(n4435), .C2(n2923), .A(n2922), .B(n2921), .ZN(n2924)
         );
  INV_X1 U3720 ( .A(n2924), .ZN(U3244) );
  NAND2_X1 U3721 ( .A1(n3901), .A2(n2925), .ZN(n3809) );
  AND2_X1 U3722 ( .A1(n3807), .A2(n3809), .ZN(n4529) );
  INV_X1 U3723 ( .A(n2926), .ZN(n2927) );
  NOR2_X1 U3724 ( .A1(n2928), .A2(n2927), .ZN(n2930) );
  NAND4_X1 U3725 ( .A1(n2932), .A2(n2931), .A3(n2930), .A4(n2929), .ZN(n2933)
         );
  NAND2_X1 U3726 ( .A1(n2934), .A2(n4380), .ZN(n2990) );
  INV_X1 U3727 ( .A(n2990), .ZN(n2935) );
  NAND2_X1 U3728 ( .A1(n4200), .A2(n2935), .ZN(n4156) );
  NAND2_X1 U3729 ( .A1(n3071), .A2(n2936), .ZN(n4527) );
  AOI21_X1 U3730 ( .B1(n4172), .B2(n4147), .A(n4529), .ZN(n2937) );
  AOI21_X1 U3731 ( .B1(n4319), .B2(n3900), .A(n2937), .ZN(n4528) );
  OAI21_X1 U3732 ( .B1(n2938), .B2(n4527), .A(n4528), .ZN(n2939) );
  INV_X1 U3733 ( .A(n4494), .ZN(n4504) );
  AOI22_X1 U3734 ( .A1(n2939), .A2(n4200), .B1(REG3_REG_0__SCAN_IN), .B2(n4504), .ZN(n2941) );
  INV_X1 U3735 ( .A(n4200), .ZN(n4227) );
  NAND2_X1 U3736 ( .A1(n4227), .A2(REG2_REG_0__SCAN_IN), .ZN(n2940) );
  OAI211_X1 U3737 ( .C1(n4529), .C2(n4156), .A(n2941), .B(n2940), .ZN(U3290)
         );
  INV_X1 U3738 ( .A(n2942), .ZN(n2946) );
  INV_X1 U3739 ( .A(n2943), .ZN(n2945) );
  NAND2_X1 U3740 ( .A1(n3898), .A2(n2047), .ZN(n2949) );
  NAND2_X1 U3741 ( .A1(n2045), .A2(n2963), .ZN(n2948) );
  NAND2_X1 U3742 ( .A1(n2949), .A2(n2948), .ZN(n2950) );
  XNOR2_X1 U3743 ( .A(n2950), .B(n2050), .ZN(n3029) );
  OAI22_X1 U3744 ( .A1(n3036), .A2(n2048), .B1(n3554), .B2(n2968), .ZN(n3028)
         );
  XNOR2_X1 U3745 ( .A(n3029), .B(n3028), .ZN(n3031) );
  XOR2_X1 U3746 ( .A(n3032), .B(n3031), .Z(n2960) );
  OAI22_X1 U3747 ( .A1(n2867), .A2(n3699), .B1(n3700), .B2(n2982), .ZN(n2958)
         );
  OAI21_X1 U3748 ( .B1(n2953), .B2(n2952), .A(STATE_REG_SCAN_IN), .ZN(n2956)
         );
  AND2_X1 U3749 ( .A1(n2954), .A2(n3881), .ZN(n2955) );
  MUX2_X1 U3750 ( .A(n3713), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2957) );
  AOI211_X1 U3751 ( .C1(n2963), .C2(n3590), .A(n2958), .B(n2957), .ZN(n2959)
         );
  OAI21_X1 U3752 ( .B1(n2960), .B2(n3716), .A(n2959), .ZN(U3215) );
  XNOR2_X1 U3753 ( .A(n2961), .B(n3770), .ZN(n3060) );
  XNOR2_X1 U3754 ( .A(n2962), .B(n3770), .ZN(n2967) );
  AOI22_X1 U3755 ( .A1(n3899), .A2(n4278), .B1(n4318), .B2(n2963), .ZN(n2964)
         );
  OAI21_X1 U3756 ( .B1(n2982), .B2(n4282), .A(n2964), .ZN(n2966) );
  NOR2_X1 U3757 ( .A1(n3060), .A2(n4147), .ZN(n2965) );
  AOI211_X1 U3758 ( .C1(n2967), .C2(n4206), .A(n2966), .B(n2965), .ZN(n3067)
         );
  OAI21_X1 U3759 ( .B1(n3060), .B2(n4532), .A(n3067), .ZN(n2975) );
  OR2_X1 U3760 ( .A1(n3012), .A2(n2968), .ZN(n2969) );
  NAND2_X1 U3761 ( .A1(n3052), .A2(n2969), .ZN(n3063) );
  INV_X1 U3762 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2970) );
  OAI22_X1 U3763 ( .A1(n4328), .A2(n3063), .B1(n4564), .B2(n2970), .ZN(n2971)
         );
  AOI21_X1 U3764 ( .B1(n2975), .B2(n4564), .A(n2971), .ZN(n2972) );
  INV_X1 U3765 ( .A(n2972), .ZN(U3521) );
  INV_X1 U3766 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2973) );
  OAI22_X1 U3767 ( .A1(n4378), .A2(n3063), .B1(n4554), .B2(n2973), .ZN(n2974)
         );
  AOI21_X1 U3768 ( .B1(n2975), .B2(n4554), .A(n2974), .ZN(n2976) );
  INV_X1 U3769 ( .A(n2976), .ZN(U3473) );
  INV_X1 U3770 ( .A(n2977), .ZN(n3820) );
  NAND2_X1 U3771 ( .A1(n3820), .A2(n3825), .ZN(n3789) );
  XOR2_X1 U3772 ( .A(n2978), .B(n3789), .Z(n3108) );
  XNOR2_X1 U3773 ( .A(n2979), .B(n3789), .ZN(n2980) );
  NAND2_X1 U3774 ( .A1(n2980), .A2(n4206), .ZN(n3105) );
  AOI22_X1 U3775 ( .A1(n3895), .A2(n4319), .B1(n4318), .B2(n2984), .ZN(n2981)
         );
  OAI211_X1 U3776 ( .C1(n2982), .C2(n4323), .A(n3105), .B(n2981), .ZN(n2983)
         );
  AOI21_X1 U3777 ( .B1(n3108), .B2(n4546), .A(n2983), .ZN(n2988) );
  AND2_X1 U3778 ( .A1(n3053), .A2(n2984), .ZN(n2985) );
  NOR2_X1 U3779 ( .A1(n2993), .A2(n2985), .ZN(n3099) );
  AOI22_X1 U3780 ( .A1(n2740), .A2(n3099), .B1(REG1_REG_5__SCAN_IN), .B2(n4561), .ZN(n2986) );
  OAI21_X1 U3781 ( .B1(n2988), .B2(n4561), .A(n2986), .ZN(U3523) );
  AOI22_X1 U3782 ( .A1(n2726), .A2(n3099), .B1(REG0_REG_5__SCAN_IN), .B2(n4552), .ZN(n2987) );
  OAI21_X1 U3783 ( .B1(n2988), .B2(n4552), .A(n2987), .ZN(U3477) );
  AND2_X1 U3784 ( .A1(n3827), .A2(n3823), .ZN(n3784) );
  XOR2_X1 U3785 ( .A(n2989), .B(n3784), .Z(n3090) );
  NAND2_X1 U3786 ( .A1(n4147), .A2(n2990), .ZN(n2991) );
  NAND2_X1 U3787 ( .A1(n4200), .A2(n2991), .ZN(n4203) );
  XNOR2_X1 U3788 ( .A(n2992), .B(n3784), .ZN(n3088) );
  NAND2_X1 U3789 ( .A1(n4200), .A2(n4206), .ZN(n3388) );
  INV_X1 U3790 ( .A(n3388), .ZN(n3001) );
  NAND2_X1 U3791 ( .A1(n4200), .A2(n3981), .ZN(n4196) );
  INV_X1 U3792 ( .A(n4537), .ZN(n3114) );
  OR2_X1 U3793 ( .A1(n2993), .A2(n3149), .ZN(n2994) );
  NAND2_X1 U3794 ( .A1(n3116), .A2(n2994), .ZN(n3095) );
  AND2_X1 U3795 ( .A1(n4200), .A2(n4278), .ZN(n4027) );
  OAI22_X1 U3796 ( .A1(n4200), .A2(n2995), .B1(n3155), .B2(n4494), .ZN(n2996)
         );
  AOI21_X1 U3797 ( .B1(n4027), .B2(n3896), .A(n2996), .ZN(n2999) );
  NAND2_X1 U3798 ( .A1(n4200), .A2(n4319), .ZN(n4220) );
  NAND2_X1 U3799 ( .A1(n4200), .A2(n4318), .ZN(n4219) );
  OAI22_X1 U3800 ( .A1(n3215), .A2(n4220), .B1(n4219), .B2(n3149), .ZN(n2997)
         );
  INV_X1 U3801 ( .A(n2997), .ZN(n2998) );
  OAI211_X1 U3802 ( .C1(n4179), .C2(n3095), .A(n2999), .B(n2998), .ZN(n3000)
         );
  AOI21_X1 U3803 ( .B1(n3088), .B2(n3001), .A(n3000), .ZN(n3002) );
  OAI21_X1 U3804 ( .B1(n3090), .B2(n4203), .A(n3002), .ZN(U3284) );
  INV_X1 U3805 ( .A(n3003), .ZN(n3004) );
  AOI21_X1 U3806 ( .B1(n2224), .B2(n3005), .A(n3004), .ZN(n4505) );
  OAI21_X1 U3807 ( .B1(n2224), .B2(n3007), .A(n3006), .ZN(n3011) );
  AOI22_X1 U3808 ( .A1(n3900), .A2(n4278), .B1(n3013), .B2(n4318), .ZN(n3008)
         );
  OAI21_X1 U3809 ( .B1(n3036), .B2(n4282), .A(n3008), .ZN(n3010) );
  NOR2_X1 U3810 ( .A1(n4505), .A2(n4147), .ZN(n3009) );
  AOI211_X1 U3811 ( .C1(n4206), .C2(n3011), .A(n3010), .B(n3009), .ZN(n4513)
         );
  OAI21_X1 U3812 ( .B1(n4505), .B2(n4532), .A(n4513), .ZN(n3021) );
  INV_X1 U3813 ( .A(n3012), .ZN(n3015) );
  NAND2_X1 U3814 ( .A1(n3068), .A2(n3013), .ZN(n3014) );
  NAND2_X1 U3815 ( .A1(n3015), .A2(n3014), .ZN(n4506) );
  OAI22_X1 U3816 ( .A1(n4328), .A2(n4506), .B1(n4564), .B2(n3016), .ZN(n3017)
         );
  AOI21_X1 U3817 ( .B1(n3021), .B2(n4564), .A(n3017), .ZN(n3018) );
  INV_X1 U3818 ( .A(n3018), .ZN(U3520) );
  INV_X1 U3819 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3019) );
  OAI22_X1 U3820 ( .A1(n4378), .A2(n4506), .B1(n4554), .B2(n3019), .ZN(n3020)
         );
  AOI21_X1 U3821 ( .B1(n3021), .B2(n4554), .A(n3020), .ZN(n3022) );
  INV_X1 U3822 ( .A(n3022), .ZN(U3471) );
  NOR2_X1 U3823 ( .A1(n3554), .A2(n3054), .ZN(n3024) );
  AOI21_X1 U3824 ( .B1(n3547), .B2(n3897), .A(n3024), .ZN(n3124) );
  NAND2_X1 U3825 ( .A1(n3897), .A2(n2047), .ZN(n3026) );
  NAND2_X1 U3826 ( .A1(n2045), .A2(n3046), .ZN(n3025) );
  NAND2_X1 U3827 ( .A1(n3026), .A2(n3025), .ZN(n3027) );
  XNOR2_X1 U3828 ( .A(n3027), .B(n2050), .ZN(n3126) );
  XOR2_X1 U3829 ( .A(n3124), .B(n3126), .Z(n3034) );
  OR2_X1 U3830 ( .A1(n3029), .A2(n3028), .ZN(n3030) );
  AOI211_X1 U3831 ( .C1(n3034), .C2(n3033), .A(n3716), .B(n3127), .ZN(n3035)
         );
  INV_X1 U3832 ( .A(n3035), .ZN(n3041) );
  OAI22_X1 U3833 ( .A1(n3675), .A2(n3054), .B1(n3036), .B2(n3699), .ZN(n3039)
         );
  OAI21_X1 U3834 ( .B1(n3700), .B2(n3148), .A(n3037), .ZN(n3038) );
  NOR2_X1 U3835 ( .A1(n3039), .A2(n3038), .ZN(n3040) );
  OAI211_X1 U3836 ( .C1(n3692), .C2(n3056), .A(n3041), .B(n3040), .ZN(U3227)
         );
  NAND2_X1 U3837 ( .A1(n3043), .A2(n3772), .ZN(n3044) );
  NAND2_X1 U3838 ( .A1(n3042), .A2(n3044), .ZN(n4539) );
  XNOR2_X1 U3839 ( .A(n3772), .B(n3045), .ZN(n3050) );
  AOI22_X1 U3840 ( .A1(n3898), .A2(n4278), .B1(n3046), .B2(n4318), .ZN(n3048)
         );
  NAND2_X1 U3841 ( .A1(n3896), .A2(n4319), .ZN(n3047) );
  OAI211_X1 U3842 ( .C1(n4539), .C2(n4147), .A(n3048), .B(n3047), .ZN(n3049)
         );
  AOI21_X1 U3843 ( .B1(n3050), .B2(n4206), .A(n3049), .ZN(n3051) );
  INV_X1 U3844 ( .A(n3051), .ZN(n4541) );
  INV_X1 U3845 ( .A(n3052), .ZN(n3055) );
  OAI211_X1 U3846 ( .C1(n3055), .C2(n3054), .A(n4537), .B(n3053), .ZN(n4540)
         );
  OAI22_X1 U3847 ( .A1(n4540), .A2(n4380), .B1(n4494), .B2(n3056), .ZN(n3057)
         );
  OAI21_X1 U3848 ( .B1(n4541), .B2(n3057), .A(n4200), .ZN(n3059) );
  NAND2_X1 U3849 ( .A1(n4227), .A2(REG2_REG_4__SCAN_IN), .ZN(n3058) );
  OAI211_X1 U3850 ( .C1(n4539), .C2(n4156), .A(n3059), .B(n3058), .ZN(U3286)
         );
  INV_X1 U3851 ( .A(n3060), .ZN(n3065) );
  INV_X1 U3852 ( .A(n4156), .ZN(n4509) );
  INV_X1 U3853 ( .A(n4200), .ZN(n4215) );
  AOI22_X1 U3854 ( .A1(n4215), .A2(REG2_REG_3__SCAN_IN), .B1(n4504), .B2(n3061), .ZN(n3062) );
  OAI21_X1 U3855 ( .B1(n4179), .B2(n3063), .A(n3062), .ZN(n3064) );
  AOI21_X1 U3856 ( .B1(n3065), .B2(n4509), .A(n3064), .ZN(n3066) );
  OAI21_X1 U3857 ( .B1(n3067), .B2(n4227), .A(n3066), .ZN(U3287) );
  INV_X1 U3858 ( .A(n3068), .ZN(n3069) );
  AOI21_X1 U3859 ( .B1(n3071), .B2(n3070), .A(n3069), .ZN(n4536) );
  OR2_X1 U3860 ( .A1(n3768), .A2(n3072), .ZN(n3073) );
  NAND2_X1 U3861 ( .A1(n3074), .A2(n3073), .ZN(n4533) );
  OAI22_X1 U3862 ( .A1(n4156), .A2(n4533), .B1(n3075), .B2(n4494), .ZN(n3084)
         );
  NAND2_X1 U3863 ( .A1(n3901), .A2(n4278), .ZN(n3077) );
  NAND2_X1 U3864 ( .A1(n3899), .A2(n4319), .ZN(n3076) );
  OAI211_X1 U3865 ( .C1(n4168), .C2(n3078), .A(n3077), .B(n3076), .ZN(n3079)
         );
  INV_X1 U3866 ( .A(n3079), .ZN(n3082) );
  XNOR2_X1 U3867 ( .A(n3768), .B(n3807), .ZN(n3080) );
  NAND2_X1 U3868 ( .A1(n3080), .A2(n4206), .ZN(n3081) );
  OAI211_X1 U3869 ( .C1(n4533), .C2(n4147), .A(n3082), .B(n3081), .ZN(n4534)
         );
  MUX2_X1 U3870 ( .A(n4534), .B(REG2_REG_1__SCAN_IN), .S(n4227), .Z(n3083) );
  AOI211_X1 U3871 ( .C1(n4508), .C2(n4536), .A(n3084), .B(n3083), .ZN(n3085)
         );
  INV_X1 U3872 ( .A(n3085), .ZN(U3289) );
  INV_X1 U3873 ( .A(n4546), .ZN(n4315) );
  AOI22_X1 U3874 ( .A1(n3894), .A2(n4319), .B1(n3145), .B2(n4318), .ZN(n3086)
         );
  OAI21_X1 U3875 ( .B1(n3148), .B2(n4323), .A(n3086), .ZN(n3087) );
  AOI21_X1 U3876 ( .B1(n3088), .B2(n4206), .A(n3087), .ZN(n3089) );
  OAI21_X1 U3877 ( .B1(n3090), .B2(n4315), .A(n3089), .ZN(n3097) );
  INV_X1 U3878 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3091) );
  OAI22_X1 U3879 ( .A1(n4378), .A2(n3095), .B1(n4554), .B2(n3091), .ZN(n3092)
         );
  AOI21_X1 U3880 ( .B1(n3097), .B2(n4554), .A(n3092), .ZN(n3093) );
  INV_X1 U3881 ( .A(n3093), .ZN(U3479) );
  OAI22_X1 U3882 ( .A1(n4328), .A2(n3095), .B1(n4564), .B2(n3094), .ZN(n3096)
         );
  AOI21_X1 U3883 ( .B1(n3097), .B2(n4564), .A(n3096), .ZN(n3098) );
  INV_X1 U3884 ( .A(n3098), .ZN(U3524) );
  INV_X1 U3885 ( .A(n3099), .ZN(n3104) );
  OAI22_X1 U3886 ( .A1(n4200), .A2(n2395), .B1(n3137), .B2(n4494), .ZN(n3100)
         );
  AOI21_X1 U3887 ( .B1(n4027), .B2(n3897), .A(n3100), .ZN(n3103) );
  OAI22_X1 U3888 ( .A1(n3143), .A2(n4220), .B1(n4219), .B2(n3132), .ZN(n3101)
         );
  INV_X1 U3889 ( .A(n3101), .ZN(n3102) );
  OAI211_X1 U3890 ( .C1(n4179), .C2(n3104), .A(n3103), .B(n3102), .ZN(n3107)
         );
  NOR2_X1 U3891 ( .A1(n3105), .A2(n4215), .ZN(n3106) );
  AOI211_X1 U3892 ( .C1(n3108), .C2(n4210), .A(n3107), .B(n3106), .ZN(n3109)
         );
  INV_X1 U3893 ( .A(n3109), .ZN(U3285) );
  XNOR2_X1 U3894 ( .A(n3110), .B(n3773), .ZN(n3113) );
  AOI22_X1 U3895 ( .A1(n3893), .A2(n4319), .B1(n4318), .B2(n3115), .ZN(n3111)
         );
  OAI21_X1 U3896 ( .B1(n3143), .B2(n4323), .A(n3111), .ZN(n3112) );
  AOI21_X1 U3897 ( .B1(n3113), .B2(n4206), .A(n3112), .ZN(n4551) );
  AOI21_X1 U3898 ( .B1(n3116), .B2(n3115), .A(n3114), .ZN(n3117) );
  NAND2_X1 U3899 ( .A1(n3117), .A2(n3227), .ZN(n4550) );
  INV_X1 U3900 ( .A(n4550), .ZN(n3120) );
  INV_X1 U3901 ( .A(n4196), .ZN(n3119) );
  OAI22_X1 U3902 ( .A1(n4200), .A2(n2421), .B1(n3171), .B2(n4494), .ZN(n3118)
         );
  AOI21_X1 U3903 ( .B1(n3120), .B2(n3119), .A(n3118), .ZN(n3123) );
  NAND2_X1 U3904 ( .A1(n3121), .A2(n3773), .ZN(n4547) );
  NAND3_X1 U3905 ( .A1(n4548), .A2(n4547), .A3(n4210), .ZN(n3122) );
  OAI211_X1 U3906 ( .C1(n4551), .C2(n4215), .A(n3123), .B(n3122), .ZN(U3283)
         );
  INV_X1 U3907 ( .A(n3124), .ZN(n3125) );
  INV_X2 U3908 ( .A(n2047), .ZN(n3554) );
  NOR2_X1 U3909 ( .A1(n3554), .A2(n3132), .ZN(n3128) );
  AOI21_X1 U3910 ( .B1(n3547), .B2(n3896), .A(n3128), .ZN(n3138) );
  OAI22_X1 U3911 ( .A1(n3148), .A2(n3554), .B1(n3553), .B2(n3132), .ZN(n3129)
         );
  XNOR2_X1 U3912 ( .A(n3129), .B(n2050), .ZN(n3140) );
  XOR2_X1 U3913 ( .A(n3138), .B(n3140), .Z(n3130) );
  AOI211_X1 U3914 ( .C1(n2086), .C2(n3130), .A(n3716), .B(n3142), .ZN(n3131)
         );
  INV_X1 U3915 ( .A(n3131), .ZN(n3136) );
  OAI22_X1 U3916 ( .A1(n3675), .A2(n3132), .B1(n3143), .B2(n3700), .ZN(n3133)
         );
  AOI211_X1 U3917 ( .C1(n3708), .C2(n3897), .A(n3134), .B(n3133), .ZN(n3135)
         );
  OAI211_X1 U3918 ( .C1(n3692), .C2(n3137), .A(n3136), .B(n3135), .ZN(U3224)
         );
  INV_X1 U3919 ( .A(n3138), .ZN(n3139) );
  AND2_X1 U3920 ( .A1(n3140), .A2(n3139), .ZN(n3141) );
  OAI22_X1 U3921 ( .A1(n3143), .A2(n3554), .B1(n3553), .B2(n3149), .ZN(n3144)
         );
  XNOR2_X1 U3922 ( .A(n3144), .B(n2050), .ZN(n3168) );
  AOI22_X1 U3923 ( .A1(n3547), .A2(n3895), .B1(n2047), .B2(n3145), .ZN(n3167)
         );
  XNOR2_X1 U3924 ( .A(n3168), .B(n3167), .ZN(n3146) );
  XNOR2_X1 U3925 ( .A(n3166), .B(n3146), .ZN(n3147) );
  NAND2_X1 U3926 ( .A1(n3147), .A2(n3685), .ZN(n3154) );
  OAI22_X1 U3927 ( .A1(n3675), .A2(n3149), .B1(n3148), .B2(n3699), .ZN(n3152)
         );
  OAI21_X1 U3928 ( .B1(n3700), .B2(n3215), .A(n3150), .ZN(n3151) );
  NOR2_X1 U3929 ( .A1(n3152), .A2(n3151), .ZN(n3153) );
  OAI211_X1 U3930 ( .C1(n3692), .C2(n3155), .A(n3154), .B(n3153), .ZN(U3236)
         );
  INV_X1 U3931 ( .A(n3156), .ZN(n3836) );
  AND2_X1 U3932 ( .A1(n3836), .A2(n3834), .ZN(n3787) );
  XOR2_X1 U3933 ( .A(n3787), .B(n3157), .Z(n3158) );
  NAND2_X1 U3934 ( .A1(n3158), .A2(n4206), .ZN(n3181) );
  INV_X1 U3935 ( .A(n3226), .ZN(n3159) );
  AOI21_X1 U3936 ( .B1(n3248), .B2(n3159), .A(n3191), .ZN(n3186) );
  OAI22_X1 U3937 ( .A1(n3252), .A2(n4494), .B1(n2449), .B2(n4200), .ZN(n3162)
         );
  INV_X1 U3938 ( .A(n4220), .ZN(n4034) );
  AOI22_X1 U3939 ( .A1(n4034), .A2(n3891), .B1(n4027), .B2(n3893), .ZN(n3160)
         );
  OAI21_X1 U3940 ( .B1(n3255), .B2(n4219), .A(n3160), .ZN(n3161) );
  AOI211_X1 U3941 ( .C1(n3186), .C2(n4508), .A(n3162), .B(n3161), .ZN(n3165)
         );
  XNOR2_X1 U3942 ( .A(n3163), .B(n3787), .ZN(n3184) );
  NAND2_X1 U3943 ( .A1(n3184), .A2(n4210), .ZN(n3164) );
  OAI211_X1 U3944 ( .C1(n3181), .C2(n4215), .A(n3165), .B(n3164), .ZN(U3281)
         );
  NOR2_X1 U3945 ( .A1(n3554), .A2(n3175), .ZN(n3169) );
  AOI21_X1 U3946 ( .B1(n3547), .B2(n3894), .A(n3169), .ZN(n3201) );
  OAI22_X1 U3947 ( .A1(n3215), .A2(n3554), .B1(n3553), .B2(n3175), .ZN(n3170)
         );
  XNOR2_X1 U3948 ( .A(n3170), .B(n2050), .ZN(n3199) );
  XOR2_X1 U3949 ( .A(n3201), .B(n3199), .Z(n3202) );
  XNOR2_X1 U3950 ( .A(n3203), .B(n3202), .ZN(n3179) );
  INV_X1 U3951 ( .A(n3171), .ZN(n3177) );
  AOI21_X1 U3952 ( .B1(n3708), .B2(n3895), .A(n3172), .ZN(n3174) );
  NAND2_X1 U3953 ( .A1(n3707), .A2(n3893), .ZN(n3173) );
  OAI211_X1 U3954 ( .C1(n3675), .C2(n3175), .A(n3174), .B(n3173), .ZN(n3176)
         );
  AOI21_X1 U3955 ( .B1(n3177), .B2(n3713), .A(n3176), .ZN(n3178) );
  OAI21_X1 U3956 ( .B1(n3179), .B2(n3716), .A(n3178), .ZN(U3210) );
  AOI22_X1 U3957 ( .A1(n3891), .A2(n4319), .B1(n4318), .B2(n3248), .ZN(n3180)
         );
  OAI211_X1 U3958 ( .C1(n3182), .C2(n4323), .A(n3181), .B(n3180), .ZN(n3183)
         );
  AOI21_X1 U3959 ( .B1(n3184), .B2(n4546), .A(n3183), .ZN(n3188) );
  AOI22_X1 U3960 ( .A1(n3186), .A2(n2740), .B1(REG1_REG_9__SCAN_IN), .B2(n4561), .ZN(n3185) );
  OAI21_X1 U3961 ( .B1(n3188), .B2(n4561), .A(n3185), .ZN(U3527) );
  AOI22_X1 U3962 ( .A1(n3186), .A2(n2726), .B1(REG0_REG_9__SCAN_IN), .B2(n4552), .ZN(n3187) );
  OAI21_X1 U3963 ( .B1(n3188), .B2(n4552), .A(n3187), .ZN(U3485) );
  AND2_X1 U3964 ( .A1(n3842), .A2(n3838), .ZN(n3785) );
  XOR2_X1 U3965 ( .A(n3785), .B(n3189), .Z(n3238) );
  XOR2_X1 U3966 ( .A(n3785), .B(n3190), .Z(n3240) );
  NAND2_X1 U3967 ( .A1(n3240), .A2(n4210), .ZN(n3198) );
  INV_X1 U3968 ( .A(n3191), .ZN(n3192) );
  AOI21_X1 U3969 ( .B1(n3284), .B2(n3192), .A(n2085), .ZN(n3242) );
  INV_X1 U3970 ( .A(n4027), .ZN(n4217) );
  INV_X1 U3971 ( .A(n4219), .ZN(n3439) );
  AOI22_X1 U3972 ( .A1(n3439), .A2(n3284), .B1(n4034), .B2(n3890), .ZN(n3195)
         );
  INV_X1 U3973 ( .A(n3298), .ZN(n3193) );
  AOI22_X1 U3974 ( .A1(n4215), .A2(REG2_REG_10__SCAN_IN), .B1(n3193), .B2(
        n4504), .ZN(n3194) );
  OAI211_X1 U3975 ( .C1(n3293), .C2(n4217), .A(n3195), .B(n3194), .ZN(n3196)
         );
  AOI21_X1 U3976 ( .B1(n3242), .B2(n4508), .A(n3196), .ZN(n3197) );
  OAI211_X1 U3977 ( .C1(n3238), .C2(n3388), .A(n3198), .B(n3197), .ZN(U3280)
         );
  INV_X1 U3978 ( .A(n3199), .ZN(n3200) );
  NAND2_X1 U3979 ( .A1(n3893), .A2(n2047), .ZN(n3205) );
  NAND2_X1 U3980 ( .A1(n2045), .A2(n3228), .ZN(n3204) );
  NAND2_X1 U3981 ( .A1(n3205), .A2(n3204), .ZN(n3206) );
  XNOR2_X1 U3982 ( .A(n3206), .B(n2074), .ZN(n3209) );
  NOR2_X1 U3983 ( .A1(n2049), .A2(n3213), .ZN(n3207) );
  AOI21_X1 U3984 ( .B1(n3547), .B2(n3893), .A(n3207), .ZN(n3208) );
  NOR2_X1 U3985 ( .A1(n3209), .A2(n3208), .ZN(n3246) );
  INV_X1 U3986 ( .A(n3246), .ZN(n3210) );
  NAND2_X1 U3987 ( .A1(n3209), .A2(n3208), .ZN(n3247) );
  NAND2_X1 U3988 ( .A1(n3210), .A2(n3247), .ZN(n3211) );
  XNOR2_X1 U3989 ( .A(n3245), .B(n3211), .ZN(n3212) );
  NAND2_X1 U3990 ( .A1(n3212), .A2(n3685), .ZN(n3219) );
  OAI22_X1 U3991 ( .A1(n3675), .A2(n3213), .B1(n3293), .B2(n3700), .ZN(n3217)
         );
  OAI21_X1 U3992 ( .B1(n3699), .B2(n3215), .A(n3214), .ZN(n3216) );
  NOR2_X1 U3993 ( .A1(n3217), .A2(n3216), .ZN(n3218) );
  OAI211_X1 U3994 ( .C1(n3692), .C2(n4495), .A(n3219), .B(n3218), .ZN(U3218)
         );
  INV_X1 U3995 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U3996 ( .A1(n3833), .A2(n3829), .ZN(n3788) );
  XNOR2_X1 U3997 ( .A(n3220), .B(n3788), .ZN(n4498) );
  XNOR2_X1 U3998 ( .A(n3221), .B(n3788), .ZN(n3225) );
  AOI22_X1 U3999 ( .A1(n3894), .A2(n4278), .B1(n3228), .B2(n4318), .ZN(n3222)
         );
  OAI21_X1 U4000 ( .B1(n3293), .B2(n4282), .A(n3222), .ZN(n3224) );
  NOR2_X1 U4001 ( .A1(n4498), .A2(n4147), .ZN(n3223) );
  AOI211_X1 U4002 ( .C1(n4206), .C2(n3225), .A(n3224), .B(n3223), .ZN(n4503)
         );
  OAI21_X1 U4003 ( .B1(n4532), .B2(n4498), .A(n4503), .ZN(n3232) );
  NAND2_X1 U4004 ( .A1(n3232), .A2(n4564), .ZN(n3230) );
  AOI21_X1 U4005 ( .B1(n3228), .B2(n3227), .A(n3226), .ZN(n4499) );
  NAND2_X1 U4006 ( .A1(n4499), .A2(n2740), .ZN(n3229) );
  OAI211_X1 U4007 ( .C1(n4564), .C2(n3231), .A(n3230), .B(n3229), .ZN(U3526)
         );
  INV_X1 U4008 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4009 ( .A1(n3232), .A2(n4554), .ZN(n3234) );
  NAND2_X1 U4010 ( .A1(n4499), .A2(n2726), .ZN(n3233) );
  OAI211_X1 U4011 ( .C1(n4554), .C2(n3235), .A(n3234), .B(n3233), .ZN(U3483)
         );
  OAI22_X1 U4012 ( .A1(n3405), .A2(n4282), .B1(n4168), .B2(n3292), .ZN(n3236)
         );
  AOI21_X1 U4013 ( .B1(n4278), .B2(n3892), .A(n3236), .ZN(n3237) );
  OAI21_X1 U4014 ( .B1(n3238), .B2(n4172), .A(n3237), .ZN(n3239) );
  AOI21_X1 U4015 ( .B1(n4546), .B2(n3240), .A(n3239), .ZN(n3244) );
  AOI22_X1 U4016 ( .A1(n3242), .A2(n2740), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4561), .ZN(n3241) );
  OAI21_X1 U4017 ( .B1(n3244), .B2(n4561), .A(n3241), .ZN(U3528) );
  AOI22_X1 U4018 ( .A1(n3242), .A2(n2726), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4552), .ZN(n3243) );
  OAI21_X1 U4019 ( .B1(n3244), .B2(n4552), .A(n3243), .ZN(U3487) );
  OAI22_X1 U4020 ( .A1(n3293), .A2(n2048), .B1(n2049), .B2(n3255), .ZN(n3279)
         );
  NAND2_X1 U4021 ( .A1(n3892), .A2(n2047), .ZN(n3250) );
  NAND2_X1 U4022 ( .A1(n2045), .A2(n3248), .ZN(n3249) );
  NAND2_X1 U4023 ( .A1(n3250), .A2(n3249), .ZN(n3251) );
  XNOR2_X1 U4024 ( .A(n3251), .B(n2050), .ZN(n3278) );
  XOR2_X1 U4025 ( .A(n3279), .B(n3278), .Z(n3276) );
  XOR2_X1 U4026 ( .A(n3277), .B(n3276), .Z(n3259) );
  INV_X1 U4027 ( .A(n3252), .ZN(n3257) );
  NOR2_X1 U4028 ( .A1(STATE_REG_SCAN_IN), .A2(n2446), .ZN(n4401) );
  AOI21_X1 U4029 ( .B1(n3707), .B2(n3891), .A(n4401), .ZN(n3254) );
  NAND2_X1 U4030 ( .A1(n3708), .A2(n3893), .ZN(n3253) );
  OAI211_X1 U4031 ( .C1(n3675), .C2(n3255), .A(n3254), .B(n3253), .ZN(n3256)
         );
  AOI21_X1 U4032 ( .B1(n3257), .B2(n3713), .A(n3256), .ZN(n3258) );
  OAI21_X1 U4033 ( .B1(n3259), .B2(n3716), .A(n3258), .ZN(U3228) );
  AND2_X1 U4034 ( .A1(n3305), .A2(n3303), .ZN(n3786) );
  INV_X1 U4035 ( .A(n3786), .ZN(n3271) );
  XNOR2_X1 U4036 ( .A(n3260), .B(n3271), .ZN(n3368) );
  AND2_X1 U4037 ( .A1(n3341), .A2(n3395), .ZN(n3261) );
  NOR2_X1 U4038 ( .A1(n3311), .A2(n3261), .ZN(n3375) );
  NAND2_X1 U4039 ( .A1(n3375), .A2(n4508), .ZN(n3267) );
  OAI22_X1 U4040 ( .A1(n4200), .A2(n3262), .B1(n3410), .B2(n4494), .ZN(n3263)
         );
  AOI21_X1 U4041 ( .B1(n4027), .B2(n3890), .A(n3263), .ZN(n3266) );
  INV_X1 U4042 ( .A(n3888), .ZN(n3579) );
  OAI22_X1 U40430 ( .A1(n3579), .A2(n4220), .B1(n4219), .B2(n3404), .ZN(n3264)
         );
  INV_X1 U4044 ( .A(n3264), .ZN(n3265) );
  NAND3_X1 U4045 ( .A1(n3267), .A2(n3266), .A3(n3265), .ZN(n3274) );
  INV_X1 U4046 ( .A(n3268), .ZN(n3269) );
  AOI21_X1 U4047 ( .B1(n3335), .B2(n3270), .A(n3269), .ZN(n3306) );
  XNOR2_X1 U4048 ( .A(n3306), .B(n3271), .ZN(n3272) );
  NAND2_X1 U4049 ( .A1(n3272), .A2(n4206), .ZN(n3366) );
  NOR2_X1 U4050 ( .A1(n3366), .A2(n4227), .ZN(n3273) );
  AOI211_X1 U4051 ( .C1(n4210), .C2(n3368), .A(n3274), .B(n3273), .ZN(n3275)
         );
  INV_X1 U4052 ( .A(n3275), .ZN(U3278) );
  INV_X1 U4053 ( .A(n3278), .ZN(n3281) );
  INV_X1 U4054 ( .A(n3279), .ZN(n3280) );
  NAND2_X1 U4055 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  NOR2_X1 U4056 ( .A1(n3554), .A2(n3292), .ZN(n3283) );
  AOI21_X1 U4057 ( .B1(n3547), .B2(n3891), .A(n3283), .ZN(n3318) );
  NAND2_X1 U4058 ( .A1(n3891), .A2(n2047), .ZN(n3286) );
  NAND2_X1 U4059 ( .A1(n2045), .A2(n3284), .ZN(n3285) );
  NAND2_X1 U4060 ( .A1(n3286), .A2(n3285), .ZN(n3287) );
  XNOR2_X1 U4061 ( .A(n3287), .B(n2050), .ZN(n3320) );
  XOR2_X1 U4062 ( .A(n3318), .B(n3320), .Z(n3289) );
  AOI21_X1 U4063 ( .B1(n3288), .B2(n3289), .A(n3716), .ZN(n3291) );
  NAND2_X1 U4064 ( .A1(n3291), .A2(n3322), .ZN(n3297) );
  OAI22_X1 U4065 ( .A1(n3675), .A2(n3292), .B1(n3405), .B2(n3700), .ZN(n3295)
         );
  NAND2_X1 U4066 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4405) );
  OAI21_X1 U4067 ( .B1(n3699), .B2(n3293), .A(n4405), .ZN(n3294) );
  NOR2_X1 U4068 ( .A1(n3295), .A2(n3294), .ZN(n3296) );
  OAI211_X1 U4069 ( .C1(n3692), .C2(n3298), .A(n3297), .B(n3296), .ZN(U3214)
         );
  INV_X1 U4070 ( .A(n3300), .ZN(n3302) );
  OR2_X1 U4071 ( .A1(n3302), .A2(n3301), .ZN(n3794) );
  XNOR2_X1 U4072 ( .A(n3299), .B(n3794), .ZN(n3348) );
  INV_X1 U4073 ( .A(n3348), .ZN(n3317) );
  INV_X1 U4074 ( .A(n3303), .ZN(n3304) );
  AOI21_X1 U4075 ( .B1(n3306), .B2(n3305), .A(n3304), .ZN(n3307) );
  XNOR2_X1 U4076 ( .A(n3307), .B(n3794), .ZN(n3310) );
  OAI22_X1 U4077 ( .A1(n4324), .A2(n4282), .B1(n4168), .B2(n3456), .ZN(n3308)
         );
  AOI21_X1 U4078 ( .B1(n4278), .B2(n3889), .A(n3308), .ZN(n3309) );
  OAI21_X1 U4079 ( .B1(n3310), .B2(n4172), .A(n3309), .ZN(n3347) );
  NOR2_X1 U4080 ( .A1(n3311), .A2(n3456), .ZN(n3312) );
  OR2_X1 U4081 ( .A1(n3380), .A2(n3312), .ZN(n3354) );
  INV_X1 U4082 ( .A(n3313), .ZN(n3458) );
  AOI22_X1 U4083 ( .A1(n4215), .A2(REG2_REG_13__SCAN_IN), .B1(n3458), .B2(
        n4504), .ZN(n3314) );
  OAI21_X1 U4084 ( .B1(n3354), .B2(n4179), .A(n3314), .ZN(n3315) );
  AOI21_X1 U4085 ( .B1(n3347), .B2(n4200), .A(n3315), .ZN(n3316) );
  OAI21_X1 U4086 ( .B1(n3317), .B2(n4203), .A(n3316), .ZN(U3277) );
  INV_X1 U4087 ( .A(n3318), .ZN(n3319) );
  NAND2_X1 U4088 ( .A1(n3320), .A2(n3319), .ZN(n3321) );
  OAI22_X1 U4089 ( .A1(n3405), .A2(n2049), .B1(n3553), .B2(n3342), .ZN(n3323)
         );
  XNOR2_X1 U4090 ( .A(n3323), .B(n2050), .ZN(n3389) );
  OAI22_X1 U4091 ( .A1(n3405), .A2(n2048), .B1(n2049), .B2(n3342), .ZN(n3390)
         );
  INV_X1 U4092 ( .A(n3390), .ZN(n3393) );
  XNOR2_X1 U4093 ( .A(n3389), .B(n3393), .ZN(n3324) );
  XNOR2_X1 U4094 ( .A(n3391), .B(n3324), .ZN(n3330) );
  INV_X1 U4095 ( .A(n3339), .ZN(n3328) );
  AND2_X1 U4096 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4422) );
  AOI21_X1 U4097 ( .B1(n3707), .B2(n3889), .A(n4422), .ZN(n3326) );
  NAND2_X1 U4098 ( .A1(n3708), .A2(n3891), .ZN(n3325) );
  OAI211_X1 U4099 ( .C1(n3675), .C2(n3342), .A(n3326), .B(n3325), .ZN(n3327)
         );
  AOI21_X1 U4100 ( .B1(n3328), .B2(n3713), .A(n3327), .ZN(n3329) );
  OAI21_X1 U4101 ( .B1(n3330), .B2(n3716), .A(n3329), .ZN(U3233) );
  INV_X1 U4102 ( .A(n3331), .ZN(n3332) );
  AOI21_X1 U4103 ( .B1(n3774), .B2(n3333), .A(n3332), .ZN(n3356) );
  AOI22_X1 U4104 ( .A1(n3889), .A2(n4319), .B1(n4318), .B2(n3334), .ZN(n3338)
         );
  XNOR2_X1 U4105 ( .A(n3335), .B(n3774), .ZN(n3336) );
  NAND2_X1 U4106 ( .A1(n3336), .A2(n4206), .ZN(n3337) );
  OAI211_X1 U4107 ( .C1(n3356), .C2(n4147), .A(n3338), .B(n3337), .ZN(n3358)
         );
  NAND2_X1 U4108 ( .A1(n3358), .A2(n4200), .ZN(n3346) );
  OAI22_X1 U4109 ( .A1(n4200), .A2(n3340), .B1(n3339), .B2(n4494), .ZN(n3344)
         );
  OAI21_X1 U4110 ( .B1(n2085), .B2(n3342), .A(n3341), .ZN(n3364) );
  NOR2_X1 U4111 ( .A1(n3364), .A2(n4179), .ZN(n3343) );
  AOI211_X1 U4112 ( .C1(n4027), .C2(n3891), .A(n3344), .B(n3343), .ZN(n3345)
         );
  OAI211_X1 U4113 ( .C1(n3356), .C2(n4156), .A(n3346), .B(n3345), .ZN(U3279)
         );
  INV_X1 U4114 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3349) );
  AOI21_X1 U4115 ( .B1(n4546), .B2(n3348), .A(n3347), .ZN(n3351) );
  MUX2_X1 U4116 ( .A(n3349), .B(n3351), .S(n4564), .Z(n3350) );
  OAI21_X1 U4117 ( .B1(n4328), .B2(n3354), .A(n3350), .ZN(U3531) );
  INV_X1 U4118 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3352) );
  MUX2_X1 U4119 ( .A(n3352), .B(n3351), .S(n4554), .Z(n3353) );
  OAI21_X1 U4120 ( .B1(n3354), .B2(n4378), .A(n3353), .ZN(U3493) );
  INV_X1 U4121 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3359) );
  OAI22_X1 U4122 ( .A1(n3356), .A2(n4532), .B1(n3355), .B2(n4323), .ZN(n3357)
         );
  NOR2_X1 U4123 ( .A1(n3358), .A2(n3357), .ZN(n3361) );
  MUX2_X1 U4124 ( .A(n3359), .B(n3361), .S(n4564), .Z(n3360) );
  OAI21_X1 U4125 ( .B1(n4328), .B2(n3364), .A(n3360), .ZN(U3529) );
  INV_X1 U4126 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3362) );
  MUX2_X1 U4127 ( .A(n3362), .B(n3361), .S(n4554), .Z(n3363) );
  OAI21_X1 U4128 ( .B1(n3364), .B2(n4378), .A(n3363), .ZN(U3489) );
  AOI22_X1 U4129 ( .A1(n3888), .A2(n4319), .B1(n4318), .B2(n3395), .ZN(n3365)
         );
  OAI211_X1 U4130 ( .C1(n3405), .C2(n4323), .A(n3366), .B(n3365), .ZN(n3367)
         );
  INV_X1 U4131 ( .A(n3367), .ZN(n3370) );
  NAND2_X1 U4132 ( .A1(n3368), .A2(n4546), .ZN(n3369) );
  NAND2_X1 U4133 ( .A1(n3370), .A2(n3369), .ZN(n3373) );
  MUX2_X1 U4134 ( .A(REG1_REG_12__SCAN_IN), .B(n3373), .S(n4564), .Z(n3371) );
  AOI21_X1 U4135 ( .B1(n2740), .B2(n3375), .A(n3371), .ZN(n3372) );
  INV_X1 U4136 ( .A(n3372), .ZN(U3530) );
  MUX2_X1 U4137 ( .A(REG0_REG_12__SCAN_IN), .B(n3373), .S(n4554), .Z(n3374) );
  AOI21_X1 U4138 ( .B1(n3375), .B2(n2726), .A(n3374), .ZN(n3376) );
  INV_X1 U4139 ( .A(n3376), .ZN(U3491) );
  XNOR2_X1 U4140 ( .A(n3719), .B(n3378), .ZN(n3426) );
  OAI21_X1 U4141 ( .B1(n3379), .B2(n3378), .A(n3377), .ZN(n3428) );
  NAND2_X1 U4142 ( .A1(n3428), .A2(n4210), .ZN(n3387) );
  OAI21_X1 U4143 ( .B1(n3380), .B2(n3577), .A(n3415), .ZN(n3434) );
  INV_X1 U4144 ( .A(n3434), .ZN(n3385) );
  AOI22_X1 U4145 ( .A1(n3439), .A2(n3464), .B1(n4034), .B2(n3886), .ZN(n3383)
         );
  INV_X1 U4146 ( .A(n3584), .ZN(n3381) );
  AOI22_X1 U4147 ( .A1(n4215), .A2(REG2_REG_14__SCAN_IN), .B1(n3381), .B2(
        n4504), .ZN(n3382) );
  OAI211_X1 U4148 ( .C1(n3579), .C2(n4217), .A(n3383), .B(n3382), .ZN(n3384)
         );
  AOI21_X1 U4149 ( .B1(n3385), .B2(n4508), .A(n3384), .ZN(n3386) );
  OAI211_X1 U4150 ( .C1(n3426), .C2(n3388), .A(n3387), .B(n3386), .ZN(U3276)
         );
  INV_X1 U4151 ( .A(n3391), .ZN(n3394) );
  OAI21_X1 U4152 ( .B1(n3394), .B2(n3393), .A(n3392), .ZN(n3450) );
  NAND2_X1 U4153 ( .A1(n3889), .A2(n2047), .ZN(n3397) );
  NAND2_X1 U4154 ( .A1(n2045), .A2(n3395), .ZN(n3396) );
  NAND2_X1 U4155 ( .A1(n3397), .A2(n3396), .ZN(n3398) );
  XNOR2_X1 U4156 ( .A(n3398), .B(n2074), .ZN(n3401) );
  NOR2_X1 U4157 ( .A1(n2049), .A2(n3404), .ZN(n3399) );
  AOI21_X1 U4158 ( .B1(n3547), .B2(n3889), .A(n3399), .ZN(n3400) );
  NOR2_X1 U4159 ( .A1(n3401), .A2(n3400), .ZN(n3449) );
  NAND2_X1 U4160 ( .A1(n3401), .A2(n3400), .ZN(n3448) );
  NAND2_X1 U4161 ( .A1(n2184), .A2(n3448), .ZN(n3402) );
  XNOR2_X1 U4162 ( .A(n3450), .B(n3402), .ZN(n3403) );
  NAND2_X1 U4163 ( .A1(n3403), .A2(n3685), .ZN(n3409) );
  OAI22_X1 U4164 ( .A1(n3675), .A2(n3404), .B1(n3579), .B2(n3700), .ZN(n3407)
         );
  NAND2_X1 U4165 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4426) );
  OAI21_X1 U4166 ( .B1(n3699), .B2(n3405), .A(n4426), .ZN(n3406) );
  NOR2_X1 U4167 ( .A1(n3407), .A2(n3406), .ZN(n3408) );
  OAI211_X1 U4168 ( .C1(n3692), .C2(n3410), .A(n3409), .B(n3408), .ZN(U3221)
         );
  AOI21_X1 U4169 ( .B1(n3411), .B2(n3769), .A(n4172), .ZN(n3413) );
  NAND2_X1 U4170 ( .A1(n3413), .A2(n3412), .ZN(n4322) );
  XNOR2_X1 U4171 ( .A(n3414), .B(n3769), .ZN(n4326) );
  NAND2_X1 U4172 ( .A1(n4326), .A2(n4210), .ZN(n3423) );
  INV_X1 U4173 ( .A(n3415), .ZN(n3416) );
  OAI21_X1 U4174 ( .B1(n3416), .B2(n3711), .A(n3438), .ZN(n4379) );
  INV_X1 U4175 ( .A(n4379), .ZN(n3421) );
  AOI22_X1 U4176 ( .A1(n3439), .A2(n4317), .B1(n4034), .B2(n4320), .ZN(n3419)
         );
  INV_X1 U4177 ( .A(n3417), .ZN(n3714) );
  AOI22_X1 U4178 ( .A1(n4215), .A2(REG2_REG_15__SCAN_IN), .B1(n3714), .B2(
        n4504), .ZN(n3418) );
  OAI211_X1 U4179 ( .C1(n4324), .C2(n4217), .A(n3419), .B(n3418), .ZN(n3420)
         );
  AOI21_X1 U4180 ( .B1(n3421), .B2(n4508), .A(n3420), .ZN(n3422) );
  OAI211_X1 U4181 ( .C1(n4227), .C2(n4322), .A(n3423), .B(n3422), .ZN(U3275)
         );
  OAI22_X1 U4182 ( .A1(n4310), .A2(n4282), .B1(n4168), .B2(n3577), .ZN(n3424)
         );
  AOI21_X1 U4183 ( .B1(n4278), .B2(n3888), .A(n3424), .ZN(n3425) );
  OAI21_X1 U4184 ( .B1(n3426), .B2(n4172), .A(n3425), .ZN(n3427) );
  AOI21_X1 U4185 ( .B1(n3428), .B2(n4546), .A(n3427), .ZN(n3432) );
  INV_X1 U4186 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3429) );
  MUX2_X1 U4187 ( .A(n3432), .B(n3429), .S(n4561), .Z(n3430) );
  OAI21_X1 U4188 ( .B1(n4328), .B2(n3434), .A(n3430), .ZN(U3532) );
  INV_X1 U4189 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3431) );
  MUX2_X1 U4190 ( .A(n3432), .B(n3431), .S(n4552), .Z(n3433) );
  OAI21_X1 U4191 ( .B1(n3434), .B2(n4378), .A(n3433), .ZN(U3495) );
  OAI21_X1 U4192 ( .B1(n3435), .B2(n2534), .A(n3436), .ZN(n4316) );
  INV_X1 U4193 ( .A(n3437), .ZN(n4213) );
  AOI21_X1 U4194 ( .B1(n4307), .B2(n3438), .A(n4213), .ZN(n4312) );
  AOI22_X1 U4195 ( .A1(n3439), .A2(n4307), .B1(n4034), .B2(n4308), .ZN(n3442)
         );
  INV_X1 U4196 ( .A(n3440), .ZN(n3636) );
  AOI22_X1 U4197 ( .A1(n4215), .A2(REG2_REG_16__SCAN_IN), .B1(n3636), .B2(
        n4504), .ZN(n3441) );
  OAI211_X1 U4198 ( .C1(n4310), .C2(n4217), .A(n3442), .B(n3441), .ZN(n3446)
         );
  OAI211_X1 U4199 ( .C1(n3444), .C2(n3793), .A(n3443), .B(n4206), .ZN(n4313)
         );
  NOR2_X1 U4200 ( .A1(n4313), .A2(n4227), .ZN(n3445) );
  AOI211_X1 U4201 ( .C1(n4312), .C2(n4508), .A(n3446), .B(n3445), .ZN(n3447)
         );
  OAI21_X1 U4202 ( .B1(n4316), .B2(n4203), .A(n3447), .ZN(U3274) );
  AOI22_X1 U4203 ( .A1(n3888), .A2(n2047), .B1(n2045), .B2(n3451), .ZN(n3452)
         );
  XNOR2_X1 U4204 ( .A(n2183), .B(n3461), .ZN(n3453) );
  XNOR2_X1 U4205 ( .A(n3463), .B(n3453), .ZN(n3460) );
  NOR2_X1 U4206 ( .A1(STATE_REG_SCAN_IN), .A2(n2488), .ZN(n4439) );
  AOI21_X1 U4207 ( .B1(n3707), .B2(n3887), .A(n4439), .ZN(n3455) );
  NAND2_X1 U4208 ( .A1(n3708), .A2(n3889), .ZN(n3454) );
  OAI211_X1 U4209 ( .C1(n3675), .C2(n3456), .A(n3455), .B(n3454), .ZN(n3457)
         );
  AOI21_X1 U4210 ( .B1(n3458), .B2(n3713), .A(n3457), .ZN(n3459) );
  OAI21_X1 U4211 ( .B1(n3460), .B2(n3716), .A(n3459), .ZN(U3231) );
  NAND2_X1 U4212 ( .A1(n3887), .A2(n2047), .ZN(n3466) );
  NAND2_X1 U4213 ( .A1(n2045), .A2(n3464), .ZN(n3465) );
  NAND2_X1 U4214 ( .A1(n3466), .A2(n3465), .ZN(n3467) );
  XNOR2_X1 U4215 ( .A(n3467), .B(n2074), .ZN(n3470) );
  NOR2_X1 U4216 ( .A1(n2049), .A2(n3577), .ZN(n3468) );
  AOI21_X1 U4217 ( .B1(n3547), .B2(n3887), .A(n3468), .ZN(n3469) );
  NOR2_X1 U4218 ( .A1(n3470), .A2(n3469), .ZN(n3572) );
  NAND2_X1 U4219 ( .A1(n3470), .A2(n3469), .ZN(n3573) );
  OAI21_X2 U4220 ( .B1(n3571), .B2(n3572), .A(n3573), .ZN(n3475) );
  OAI22_X1 U4221 ( .A1(n4310), .A2(n2049), .B1(n3553), .B2(n3711), .ZN(n3471)
         );
  XOR2_X1 U4222 ( .A(n2050), .B(n3471), .Z(n3474) );
  INV_X1 U4223 ( .A(n3473), .ZN(n3628) );
  NAND2_X1 U4224 ( .A1(n3475), .A2(n3474), .ZN(n3629) );
  NAND2_X1 U4225 ( .A1(n3547), .A2(n3886), .ZN(n3477) );
  NAND2_X1 U4226 ( .A1(n2047), .A2(n4317), .ZN(n3476) );
  NAND2_X1 U4227 ( .A1(n3477), .A2(n3476), .ZN(n3706) );
  NAND2_X1 U4228 ( .A1(n3629), .A2(n3706), .ZN(n3481) );
  OAI22_X1 U4229 ( .A1(n4303), .A2(n2049), .B1(n3553), .B2(n3634), .ZN(n3478)
         );
  XNOR2_X1 U4230 ( .A(n3478), .B(n2050), .ZN(n3480) );
  OAI22_X1 U4231 ( .A1(n4303), .A2(n2048), .B1(n2049), .B2(n3634), .ZN(n3479)
         );
  NOR2_X1 U4232 ( .A1(n3480), .A2(n3479), .ZN(n3482) );
  AOI21_X1 U4233 ( .B1(n3480), .B2(n3479), .A(n3482), .ZN(n3631) );
  INV_X1 U4234 ( .A(n3482), .ZN(n3483) );
  NAND2_X1 U4235 ( .A1(n4308), .A2(n2047), .ZN(n3485) );
  NAND2_X1 U4236 ( .A1(n2045), .A2(n4299), .ZN(n3484) );
  NAND2_X1 U4237 ( .A1(n3485), .A2(n3484), .ZN(n3486) );
  XNOR2_X1 U4238 ( .A(n3486), .B(n2050), .ZN(n3489) );
  NAND2_X1 U4239 ( .A1(n3547), .A2(n4308), .ZN(n3488) );
  NAND2_X1 U4240 ( .A1(n2047), .A2(n4299), .ZN(n3487) );
  NAND2_X1 U4241 ( .A1(n3488), .A2(n3487), .ZN(n3490) );
  NAND2_X1 U4242 ( .A1(n3489), .A2(n3490), .ZN(n3641) );
  INV_X1 U4243 ( .A(n3489), .ZN(n3492) );
  INV_X1 U4244 ( .A(n3490), .ZN(n3491) );
  NAND2_X1 U4245 ( .A1(n3492), .A2(n3491), .ZN(n3640) );
  AOI22_X1 U4246 ( .A1(n4300), .A2(n3547), .B1(n2047), .B2(n4189), .ZN(n3683)
         );
  AOI22_X1 U4247 ( .A1(n4300), .A2(n2047), .B1(n2045), .B2(n4189), .ZN(n3493)
         );
  XNOR2_X1 U4248 ( .A(n3493), .B(n2050), .ZN(n3682) );
  NOR2_X1 U4249 ( .A1(n3681), .A2(n3683), .ZN(n3494) );
  NOR2_X1 U4250 ( .A1(n3495), .A2(n3494), .ZN(n3596) );
  NAND2_X1 U4251 ( .A1(n4142), .A2(n2047), .ZN(n3497) );
  NAND2_X1 U4252 ( .A1(n2045), .A2(n4174), .ZN(n3496) );
  NAND2_X1 U4253 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  XNOR2_X1 U4254 ( .A(n3498), .B(n2074), .ZN(n3502) );
  NOR2_X1 U4255 ( .A1(n2049), .A2(n4169), .ZN(n3500) );
  AOI21_X1 U4256 ( .B1(n4142), .B2(n3547), .A(n3500), .ZN(n3501) );
  NAND2_X1 U4257 ( .A1(n3502), .A2(n3501), .ZN(n3504) );
  OAI21_X1 U4258 ( .B1(n3502), .B2(n3501), .A(n3504), .ZN(n3600) );
  NAND2_X1 U4259 ( .A1(n3596), .A2(n3503), .ZN(n3597) );
  OAI22_X1 U4260 ( .A1(n4132), .A2(n2049), .B1(n3553), .B2(n3665), .ZN(n3505)
         );
  XNOR2_X1 U4261 ( .A(n3505), .B(n2050), .ZN(n3506) );
  OAI22_X1 U4262 ( .A1(n4132), .A2(n2048), .B1(n2049), .B2(n3665), .ZN(n3507)
         );
  NAND2_X1 U4263 ( .A1(n3506), .A2(n3507), .ZN(n3662) );
  INV_X1 U4264 ( .A(n3506), .ZN(n3509) );
  INV_X1 U4265 ( .A(n3507), .ZN(n3508) );
  NAND2_X1 U4266 ( .A1(n3509), .A2(n3508), .ZN(n3661) );
  NAND2_X1 U4267 ( .A1(n4109), .A2(n2047), .ZN(n3511) );
  NAND2_X1 U4268 ( .A1(n2045), .A2(n4277), .ZN(n3510) );
  NAND2_X1 U4269 ( .A1(n3511), .A2(n3510), .ZN(n3512) );
  XNOR2_X1 U4270 ( .A(n3512), .B(n2050), .ZN(n3516) );
  NAND2_X1 U4271 ( .A1(n4109), .A2(n3547), .ZN(n3514) );
  NAND2_X1 U4272 ( .A1(n2047), .A2(n4277), .ZN(n3513) );
  NAND2_X1 U4273 ( .A1(n3514), .A2(n3513), .ZN(n3515) );
  NOR2_X1 U4274 ( .A1(n3516), .A2(n3515), .ZN(n3607) );
  NAND2_X1 U4275 ( .A1(n3516), .A2(n3515), .ZN(n3608) );
  OAI22_X1 U4276 ( .A1(n4283), .A2(n2049), .B1(n3553), .B2(n4112), .ZN(n3517)
         );
  XNOR2_X1 U4277 ( .A(n3517), .B(n2050), .ZN(n3522) );
  OAI22_X1 U4278 ( .A1(n4283), .A2(n2048), .B1(n2049), .B2(n4112), .ZN(n3523)
         );
  XNOR2_X1 U4279 ( .A(n3522), .B(n3523), .ZN(n3673) );
  NAND2_X1 U4280 ( .A1(n4259), .A2(n2047), .ZN(n3519) );
  NAND2_X1 U4281 ( .A1(n2045), .A2(n4098), .ZN(n3518) );
  NAND2_X1 U4282 ( .A1(n3519), .A2(n3518), .ZN(n3520) );
  XNOR2_X1 U4283 ( .A(n3520), .B(n2050), .ZN(n3528) );
  NOR2_X1 U4284 ( .A1(n2049), .A2(n4093), .ZN(n3521) );
  AOI21_X1 U4285 ( .B1(n4259), .B2(n3547), .A(n3521), .ZN(n3526) );
  XNOR2_X1 U4286 ( .A(n3528), .B(n3526), .ZN(n3588) );
  INV_X1 U4287 ( .A(n3522), .ZN(n3525) );
  INV_X1 U4288 ( .A(n3523), .ZN(n3524) );
  NAND2_X1 U4289 ( .A1(n3525), .A2(n3524), .ZN(n3586) );
  NAND2_X1 U4290 ( .A1(n3585), .A2(n3534), .ZN(n3532) );
  INV_X1 U4291 ( .A(n3526), .ZN(n3527) );
  NOR2_X1 U4292 ( .A1(n2049), .A2(n4079), .ZN(n3529) );
  AOI21_X1 U4293 ( .B1(n4095), .B2(n3547), .A(n3529), .ZN(n3535) );
  NAND2_X1 U4294 ( .A1(n3532), .A2(n3531), .ZN(n3650) );
  OAI22_X1 U4295 ( .A1(n4058), .A2(n2049), .B1(n3553), .B2(n4079), .ZN(n3533)
         );
  XNOR2_X1 U4296 ( .A(n3533), .B(n2050), .ZN(n3652) );
  NAND2_X1 U4297 ( .A1(n3650), .A2(n3652), .ZN(n3537) );
  OAI22_X1 U4298 ( .A1(n4262), .A2(n2049), .B1(n3553), .B2(n4062), .ZN(n3538)
         );
  XNOR2_X1 U4299 ( .A(n3538), .B(n2050), .ZN(n3540) );
  OAI22_X1 U4300 ( .A1(n4262), .A2(n2048), .B1(n2049), .B2(n4062), .ZN(n3539)
         );
  OR2_X1 U4301 ( .A1(n3540), .A2(n3539), .ZN(n3619) );
  NAND2_X1 U4302 ( .A1(n3540), .A2(n3539), .ZN(n3618) );
  NAND2_X1 U4303 ( .A1(n4237), .A2(n2047), .ZN(n3544) );
  NAND2_X1 U4304 ( .A1(n2045), .A2(n4245), .ZN(n3543) );
  NAND2_X1 U4305 ( .A1(n3544), .A2(n3543), .ZN(n3545) );
  XNOR2_X1 U4306 ( .A(n3545), .B(n2074), .ZN(n3549) );
  NOR2_X1 U4307 ( .A1(n2049), .A2(n4048), .ZN(n3546) );
  AOI21_X1 U4308 ( .B1(n4237), .B2(n3547), .A(n3546), .ZN(n3548) );
  NOR2_X1 U4309 ( .A1(n3549), .A2(n3548), .ZN(n3696) );
  NAND2_X1 U4310 ( .A1(n3549), .A2(n3548), .ZN(n3694) );
  OAI22_X1 U4311 ( .A1(n4249), .A2(n2049), .B1(n4029), .B2(n3553), .ZN(n3550)
         );
  XNOR2_X1 U4312 ( .A(n3550), .B(n2050), .ZN(n3552) );
  OAI22_X1 U4313 ( .A1(n4249), .A2(n2048), .B1(n4029), .B2(n2049), .ZN(n3551)
         );
  XNOR2_X1 U4314 ( .A(n3552), .B(n3551), .ZN(n3564) );
  OAI22_X1 U4315 ( .A1(n4240), .A2(n2048), .B1(n2049), .B2(n4008), .ZN(n3557)
         );
  OAI22_X1 U4316 ( .A1(n4240), .A2(n2049), .B1(n3553), .B2(n4008), .ZN(n3555)
         );
  XNOR2_X1 U4317 ( .A(n3555), .B(n2050), .ZN(n3556) );
  XOR2_X1 U4318 ( .A(n3557), .B(n3556), .Z(n3558) );
  INV_X1 U4319 ( .A(n3883), .ZN(n4009) );
  INV_X1 U4320 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3559) );
  OAI22_X1 U4321 ( .A1(n4009), .A2(n3700), .B1(STATE_REG_SCAN_IN), .B2(n3559), 
        .ZN(n3561) );
  OAI22_X1 U4322 ( .A1(n4249), .A2(n3699), .B1(n3675), .B2(n4008), .ZN(n3560)
         );
  AOI211_X1 U4323 ( .C1(n4005), .C2(n3713), .A(n3561), .B(n3560), .ZN(n3562)
         );
  OAI21_X1 U4324 ( .B1(n3563), .B2(n3716), .A(n3562), .ZN(U3217) );
  XNOR2_X1 U4325 ( .A(n3565), .B(n3564), .ZN(n3570) );
  NOR2_X1 U4326 ( .A1(n4025), .A2(n3692), .ZN(n3568) );
  AOI22_X1 U4327 ( .A1(n4237), .A2(n3708), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3566) );
  OAI21_X1 U4328 ( .B1(n3675), .B2(n4029), .A(n3566), .ZN(n3567) );
  AOI211_X1 U4329 ( .C1(n4033), .C2(n3707), .A(n3568), .B(n3567), .ZN(n3569)
         );
  OAI21_X1 U4330 ( .B1(n3570), .B2(n3716), .A(n3569), .ZN(U3211) );
  INV_X1 U4331 ( .A(n3572), .ZN(n3574) );
  NAND2_X1 U4332 ( .A1(n3574), .A2(n3573), .ZN(n3575) );
  XNOR2_X1 U4333 ( .A(n3571), .B(n3575), .ZN(n3576) );
  NAND2_X1 U4334 ( .A1(n3576), .A2(n3685), .ZN(n3583) );
  OAI22_X1 U4335 ( .A1(n3675), .A2(n3577), .B1(n4310), .B2(n3700), .ZN(n3581)
         );
  NOR2_X1 U4336 ( .A1(n4693), .A2(STATE_REG_SCAN_IN), .ZN(n4449) );
  INV_X1 U4337 ( .A(n4449), .ZN(n3578) );
  OAI21_X1 U4338 ( .B1(n3699), .B2(n3579), .A(n3578), .ZN(n3580) );
  NOR2_X1 U4339 ( .A1(n3581), .A2(n3580), .ZN(n3582) );
  OAI211_X1 U4340 ( .C1(n3692), .C2(n3584), .A(n3583), .B(n3582), .ZN(U3212)
         );
  INV_X1 U4341 ( .A(n3585), .ZN(n3671) );
  OAI211_X1 U4342 ( .C1(n3589), .C2(n3588), .A(n3685), .B(n3587), .ZN(n3595)
         );
  AOI22_X1 U4343 ( .A1(n4095), .A2(n3707), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3594) );
  AOI22_X1 U4344 ( .A1(n3590), .A2(n4098), .B1(n3708), .B2(n3884), .ZN(n3593)
         );
  INV_X1 U4345 ( .A(n3591), .ZN(n4101) );
  NAND2_X1 U4346 ( .A1(n3713), .A2(n4101), .ZN(n3592) );
  NAND4_X1 U4347 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(U3213)
         );
  INV_X1 U4348 ( .A(n3596), .ZN(n3599) );
  INV_X1 U4349 ( .A(n3597), .ZN(n3598) );
  AOI21_X1 U4350 ( .B1(n3600), .B2(n3599), .A(n3598), .ZN(n3606) );
  INV_X1 U4351 ( .A(n4300), .ZN(n4221) );
  OAI22_X1 U4352 ( .A1(n3675), .A2(n4169), .B1(n4221), .B2(n3699), .ZN(n3602)
         );
  NAND2_X1 U4353 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3980) );
  OAI21_X1 U4354 ( .B1(n3700), .B2(n4132), .A(n3980), .ZN(n3601) );
  NOR2_X1 U4355 ( .A1(n3602), .A2(n3601), .ZN(n3605) );
  INV_X1 U4356 ( .A(n3603), .ZN(n4177) );
  NAND2_X1 U4357 ( .A1(n3713), .A2(n4177), .ZN(n3604) );
  OAI211_X1 U4358 ( .C1(n3606), .C2(n3716), .A(n3605), .B(n3604), .ZN(U3216)
         );
  INV_X1 U4359 ( .A(n3607), .ZN(n3609) );
  NAND2_X1 U4360 ( .A1(n3609), .A2(n3608), .ZN(n3611) );
  OAI211_X1 U4361 ( .C1(n3660), .C2(n2295), .A(n3662), .B(n3611), .ZN(n3610)
         );
  OAI211_X1 U4362 ( .C1(n3612), .C2(n3611), .A(n3685), .B(n3610), .ZN(n3617)
         );
  AOI22_X1 U4363 ( .A1(n3707), .A2(n3884), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3616) );
  OAI22_X1 U4364 ( .A1(n3675), .A2(n4133), .B1(n4132), .B2(n3699), .ZN(n3613)
         );
  INV_X1 U4365 ( .A(n3613), .ZN(n3615) );
  NAND2_X1 U4366 ( .A1(n3713), .A2(n4130), .ZN(n3614) );
  NAND4_X1 U4367 ( .A1(n3617), .A2(n3616), .A3(n3615), .A4(n3614), .ZN(U3220)
         );
  NAND2_X1 U4368 ( .A1(n3619), .A2(n3618), .ZN(n3621) );
  XOR2_X1 U4369 ( .A(n3621), .B(n3620), .Z(n3627) );
  INV_X1 U4370 ( .A(n3622), .ZN(n4065) );
  OAI22_X1 U4371 ( .A1(n4058), .A2(n3699), .B1(n3675), .B2(n4062), .ZN(n3625)
         );
  INV_X1 U4372 ( .A(n4237), .ZN(n3623) );
  OAI22_X1 U4373 ( .A1(n3623), .A2(n3700), .B1(STATE_REG_SCAN_IN), .B2(n4690), 
        .ZN(n3624) );
  AOI211_X1 U4374 ( .C1(n4065), .C2(n3713), .A(n3625), .B(n3624), .ZN(n3626)
         );
  OAI21_X1 U4375 ( .B1(n3627), .B2(n3716), .A(n3626), .ZN(U3222) );
  OAI21_X1 U4376 ( .B1(n3473), .B2(n3706), .A(n3629), .ZN(n3630) );
  XOR2_X1 U4377 ( .A(n3631), .B(n3630), .Z(n3638) );
  AND2_X1 U4378 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4466) );
  AOI21_X1 U4379 ( .B1(n3707), .B2(n4308), .A(n4466), .ZN(n3633) );
  NAND2_X1 U4380 ( .A1(n3708), .A2(n3886), .ZN(n3632) );
  OAI211_X1 U4381 ( .C1(n3675), .C2(n3634), .A(n3633), .B(n3632), .ZN(n3635)
         );
  AOI21_X1 U4382 ( .B1(n3636), .B2(n3713), .A(n3635), .ZN(n3637) );
  OAI21_X1 U4383 ( .B1(n3638), .B2(n3716), .A(n3637), .ZN(U3223) );
  NAND2_X1 U4384 ( .A1(n3641), .A2(n3640), .ZN(n3642) );
  XNOR2_X1 U4385 ( .A(n3639), .B(n3642), .ZN(n3648) );
  INV_X1 U4386 ( .A(n3643), .ZN(n4214) );
  NOR2_X1 U4387 ( .A1(STATE_REG_SCAN_IN), .A2(n2536), .ZN(n4475) );
  AOI21_X1 U4388 ( .B1(n3707), .B2(n4300), .A(n4475), .ZN(n3645) );
  NAND2_X1 U4389 ( .A1(n3708), .A2(n4320), .ZN(n3644) );
  OAI211_X1 U4390 ( .C1(n3675), .C2(n4218), .A(n3645), .B(n3644), .ZN(n3646)
         );
  AOI21_X1 U4391 ( .B1(n4214), .B2(n3713), .A(n3646), .ZN(n3647) );
  OAI21_X1 U4392 ( .B1(n3648), .B2(n3716), .A(n3647), .ZN(U3225) );
  NAND2_X1 U4393 ( .A1(n3649), .A2(n3650), .ZN(n3651) );
  XOR2_X1 U4394 ( .A(n3652), .B(n3651), .Z(n3658) );
  INV_X1 U4395 ( .A(n3653), .ZN(n4077) );
  OAI22_X1 U4396 ( .A1(n4107), .A2(n3699), .B1(n3675), .B2(n4079), .ZN(n3656)
         );
  INV_X1 U4397 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3654) );
  OAI22_X1 U4398 ( .A1(n4262), .A2(n3700), .B1(STATE_REG_SCAN_IN), .B2(n3654), 
        .ZN(n3655) );
  AOI211_X1 U4399 ( .C1(n4077), .C2(n3713), .A(n3656), .B(n3655), .ZN(n3657)
         );
  OAI21_X1 U4400 ( .B1(n3658), .B2(n3716), .A(n3657), .ZN(U3226) );
  NOR2_X1 U4401 ( .A1(n3659), .A2(n2295), .ZN(n3664) );
  AOI21_X1 U4402 ( .B1(n3662), .B2(n3661), .A(n3660), .ZN(n3663) );
  OAI21_X1 U4403 ( .B1(n3664), .B2(n3663), .A(n3685), .ZN(n3670) );
  AOI22_X1 U4404 ( .A1(n3707), .A2(n4109), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3669) );
  INV_X1 U4405 ( .A(n4142), .ZN(n4191) );
  OAI22_X1 U4406 ( .A1(n3675), .A2(n3665), .B1(n4191), .B2(n3699), .ZN(n3666)
         );
  INV_X1 U4407 ( .A(n3666), .ZN(n3668) );
  NAND2_X1 U4408 ( .A1(n3713), .A2(n4151), .ZN(n3667) );
  NAND4_X1 U4409 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), .ZN(U3230)
         );
  AOI21_X1 U4410 ( .B1(n3673), .B2(n3672), .A(n3671), .ZN(n3680) );
  INV_X1 U4411 ( .A(n3674), .ZN(n4115) );
  OAI22_X1 U4412 ( .A1(n3675), .A2(n4112), .B1(n4144), .B2(n3699), .ZN(n3678)
         );
  OAI22_X1 U4413 ( .A1(n4107), .A2(n3700), .B1(STATE_REG_SCAN_IN), .B2(n3676), 
        .ZN(n3677) );
  AOI211_X1 U4414 ( .C1(n4115), .C2(n3713), .A(n3678), .B(n3677), .ZN(n3679)
         );
  OAI21_X1 U4415 ( .B1(n3680), .B2(n3716), .A(n3679), .ZN(U3232) );
  XOR2_X1 U4416 ( .A(n3683), .B(n3682), .Z(n3684) );
  XNOR2_X1 U4417 ( .A(n3681), .B(n3684), .ZN(n3686) );
  NAND2_X1 U4418 ( .A1(n3686), .A2(n3685), .ZN(n3691) );
  OAI22_X1 U4419 ( .A1(n3675), .A2(n4195), .B1(n3687), .B2(n3699), .ZN(n3689)
         );
  NAND2_X1 U4420 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4481) );
  OAI21_X1 U4421 ( .B1(n3700), .B2(n4191), .A(n4481), .ZN(n3688) );
  NOR2_X1 U4422 ( .A1(n3689), .A2(n3688), .ZN(n3690) );
  OAI211_X1 U4423 ( .C1(n3692), .C2(n4197), .A(n3691), .B(n3690), .ZN(U3235)
         );
  INV_X1 U4424 ( .A(n3694), .ZN(n3695) );
  NOR2_X1 U4425 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  XNOR2_X1 U4426 ( .A(n3693), .B(n3697), .ZN(n3704) );
  OAI22_X1 U4427 ( .A1(n4262), .A2(n3699), .B1(STATE_REG_SCAN_IN), .B2(n3698), 
        .ZN(n3702) );
  OAI22_X1 U4428 ( .A1(n4249), .A2(n3700), .B1(n3675), .B2(n4048), .ZN(n3701)
         );
  AOI211_X1 U4429 ( .C1(n4046), .C2(n3713), .A(n3702), .B(n3701), .ZN(n3703)
         );
  OAI21_X1 U4430 ( .B1(n3704), .B2(n3716), .A(n3703), .ZN(U3237) );
  NAND2_X1 U4431 ( .A1(n3628), .A2(n3629), .ZN(n3705) );
  XOR2_X1 U4432 ( .A(n3706), .B(n3705), .Z(n3717) );
  AND2_X1 U4433 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4457) );
  AOI21_X1 U4434 ( .B1(n3707), .B2(n4320), .A(n4457), .ZN(n3710) );
  NAND2_X1 U4435 ( .A1(n3708), .A2(n3887), .ZN(n3709) );
  OAI211_X1 U4436 ( .C1(n3675), .C2(n3711), .A(n3710), .B(n3709), .ZN(n3712)
         );
  AOI21_X1 U4437 ( .B1(n3714), .B2(n3713), .A(n3712), .ZN(n3715) );
  OAI21_X1 U4438 ( .B1(n3717), .B2(n3716), .A(n3715), .ZN(U3238) );
  INV_X1 U4439 ( .A(n3848), .ZN(n3723) );
  NAND2_X1 U4440 ( .A1(n3722), .A2(n3718), .ZN(n3846) );
  NOR3_X1 U4441 ( .A1(n3719), .A2(n3723), .A3(n3846), .ZN(n3721) );
  INV_X1 U4442 ( .A(n3720), .ZN(n3850) );
  OAI21_X1 U4443 ( .B1(n3721), .B2(n3850), .A(n3849), .ZN(n3731) );
  INV_X1 U4444 ( .A(n3722), .ZN(n3724) );
  AOI211_X1 U4445 ( .C1(n3726), .C2(n3725), .A(n3724), .B(n3723), .ZN(n3728)
         );
  OAI21_X1 U4446 ( .B1(n3728), .B2(n3727), .A(n3849), .ZN(n3730) );
  AND2_X1 U4447 ( .A1(n3730), .A2(n3729), .ZN(n3853) );
  NAND2_X1 U4448 ( .A1(n3731), .A2(n3853), .ZN(n3733) );
  INV_X1 U4449 ( .A(n3766), .ZN(n3732) );
  NOR2_X1 U4450 ( .A1(n3780), .A2(n3732), .ZN(n3857) );
  OAI221_X1 U4451 ( .B1(n3734), .B2(n3856), .C1(n3734), .C2(n3733), .A(n3857), 
        .ZN(n3745) );
  OR2_X1 U4452 ( .A1(n3736), .A2(n3735), .ZN(n3750) );
  NAND2_X1 U4453 ( .A1(n3737), .A2(REG1_REG_31__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U4454 ( .A1(n2558), .A2(REG0_REG_31__SCAN_IN), .ZN(n3740) );
  INV_X1 U4455 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3990) );
  OR2_X1 U4456 ( .A1(n3738), .A2(n3990), .ZN(n3739) );
  AND3_X1 U4457 ( .A1(n3741), .A2(n3740), .A3(n3739), .ZN(n3988) );
  INV_X1 U4458 ( .A(n3988), .ZN(n3882) );
  NOR2_X1 U4459 ( .A1(n2487), .A2(n4704), .ZN(n3989) );
  INV_X1 U4460 ( .A(n3989), .ZN(n3986) );
  AND2_X1 U4461 ( .A1(n3882), .A2(n3986), .ZN(n3868) );
  INV_X1 U4462 ( .A(n3868), .ZN(n3744) );
  NOR2_X1 U4463 ( .A1(n3742), .A2(n4568), .ZN(n4233) );
  NAND2_X1 U4464 ( .A1(n3756), .A2(n4233), .ZN(n3743) );
  AND2_X1 U4465 ( .A1(n3744), .A2(n3743), .ZN(n3797) );
  OAI21_X1 U4466 ( .B1(n3883), .B2(n3995), .A(n3797), .ZN(n3749) );
  AOI211_X1 U4467 ( .C1(n4037), .C2(n3745), .A(n3750), .B(n3749), .ZN(n3753)
         );
  NAND2_X1 U4468 ( .A1(n3883), .A2(n3995), .ZN(n3746) );
  AND2_X1 U4469 ( .A1(n3747), .A2(n3746), .ZN(n3862) );
  NAND3_X1 U4470 ( .A1(n4022), .A2(n3862), .A3(n3748), .ZN(n3751) );
  AOI21_X1 U4471 ( .B1(n3862), .B2(n3750), .A(n3749), .ZN(n3867) );
  AOI22_X1 U4472 ( .A1(n3753), .A2(n3752), .B1(n3751), .B2(n3867), .ZN(n3760)
         );
  INV_X1 U4473 ( .A(n4233), .ZN(n3754) );
  NOR2_X1 U4474 ( .A1(n3882), .A2(n3754), .ZN(n3759) );
  INV_X1 U4475 ( .A(n3755), .ZN(n3758) );
  NOR2_X1 U4476 ( .A1(n3756), .A2(n4233), .ZN(n3796) );
  OAI21_X1 U4477 ( .B1(n3796), .B2(n3988), .A(n3989), .ZN(n3757) );
  OAI211_X1 U4478 ( .C1(n3760), .C2(n3759), .A(n3758), .B(n3757), .ZN(n3875)
         );
  INV_X1 U4479 ( .A(n3761), .ZN(n3763) );
  OR2_X1 U4480 ( .A1(n3763), .A2(n3762), .ZN(n4043) );
  INV_X1 U4481 ( .A(n4043), .ZN(n3805) );
  NAND2_X1 U4482 ( .A1(n3764), .A2(n4038), .ZN(n4056) );
  NAND2_X1 U4483 ( .A1(n3766), .A2(n3765), .ZN(n4092) );
  INV_X1 U4484 ( .A(n4092), .ZN(n3778) );
  INV_X1 U4485 ( .A(n4087), .ZN(n3852) );
  AND2_X1 U4486 ( .A1(n3852), .A2(n4086), .ZN(n4127) );
  INV_X1 U4487 ( .A(n4162), .ZN(n3767) );
  AND2_X1 U4488 ( .A1(n3767), .A2(n4161), .ZN(n4208) );
  INV_X1 U4489 ( .A(n3768), .ZN(n3771) );
  NAND4_X1 U4490 ( .A1(n4208), .A2(n3771), .A3(n3770), .A4(n2133), .ZN(n3776)
         );
  NAND4_X1 U4491 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n2224), .ZN(n3775)
         );
  NOR2_X1 U4492 ( .A1(n3776), .A2(n3775), .ZN(n3777) );
  NAND3_X1 U4493 ( .A1(n3778), .A2(n4127), .A3(n3777), .ZN(n3803) );
  INV_X1 U4494 ( .A(n3779), .ZN(n4055) );
  NOR2_X1 U4495 ( .A1(n3780), .A2(n4055), .ZN(n4073) );
  INV_X1 U4496 ( .A(n4117), .ZN(n4090) );
  XNOR2_X1 U4497 ( .A(n4142), .B(n4169), .ZN(n4159) );
  INV_X1 U4498 ( .A(n4159), .ZN(n4166) );
  INV_X1 U4499 ( .A(n3781), .ZN(n3783) );
  AND2_X1 U4500 ( .A1(n3783), .A2(n3782), .ZN(n4146) );
  INV_X1 U4501 ( .A(n4184), .ZN(n4187) );
  AND4_X1 U4502 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3792)
         );
  NOR2_X1 U4503 ( .A1(n3789), .A2(n3788), .ZN(n3790) );
  NAND4_X1 U4504 ( .A1(n4187), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3801)
         );
  NAND2_X1 U4505 ( .A1(n3793), .A2(n4529), .ZN(n3800) );
  INV_X1 U4506 ( .A(n3794), .ZN(n3799) );
  NOR2_X1 U4507 ( .A1(n3882), .A2(n3986), .ZN(n3795) );
  NOR2_X1 U4508 ( .A1(n3796), .A2(n3795), .ZN(n3869) );
  OR3_X1 U4509 ( .A1(n4056), .A2(n3803), .A3(n3802), .ZN(n3804) );
  OR3_X1 U4510 ( .A1(n3806), .A2(n3805), .A3(n3804), .ZN(n3874) );
  NOR2_X1 U4511 ( .A1(n4249), .A2(n4236), .ZN(n3866) );
  INV_X1 U4512 ( .A(n3807), .ZN(n3810) );
  OAI211_X1 U4513 ( .C1(n3810), .C2(n2667), .A(n3809), .B(n3808), .ZN(n3813)
         );
  NAND3_X1 U4514 ( .A1(n3813), .A2(n3812), .A3(n3811), .ZN(n3816) );
  NAND3_X1 U4515 ( .A1(n3816), .A2(n3815), .A3(n3814), .ZN(n3819) );
  NAND3_X1 U4516 ( .A1(n3819), .A2(n3818), .A3(n3817), .ZN(n3822) );
  NAND3_X1 U4517 ( .A1(n3822), .A2(n3821), .A3(n3820), .ZN(n3826) );
  INV_X1 U4518 ( .A(n3823), .ZN(n3824) );
  AOI21_X1 U4519 ( .B1(n3826), .B2(n3825), .A(n3824), .ZN(n3832) );
  NAND2_X1 U4520 ( .A1(n3828), .A2(n3827), .ZN(n3831) );
  OAI211_X1 U4521 ( .C1(n3832), .C2(n3831), .A(n3830), .B(n3829), .ZN(n3835)
         );
  NAND3_X1 U4522 ( .A1(n3835), .A2(n3834), .A3(n3833), .ZN(n3837) );
  NAND2_X1 U4523 ( .A1(n3837), .A2(n3836), .ZN(n3843) );
  INV_X1 U4524 ( .A(n3838), .ZN(n3841) );
  INV_X1 U4525 ( .A(n3839), .ZN(n3840) );
  AOI211_X1 U4526 ( .C1(n3843), .C2(n3842), .A(n3841), .B(n3840), .ZN(n3847)
         );
  INV_X1 U4527 ( .A(n3844), .ZN(n3845) );
  NOR3_X1 U4528 ( .A1(n3847), .A2(n3846), .A3(n3845), .ZN(n3851) );
  OAI211_X1 U4529 ( .C1(n3851), .C2(n3850), .A(n3849), .B(n3848), .ZN(n3854)
         );
  NAND3_X1 U4530 ( .A1(n3854), .A2(n3853), .A3(n3852), .ZN(n3855) );
  NAND2_X1 U4531 ( .A1(n3856), .A2(n3855), .ZN(n3860) );
  INV_X1 U4532 ( .A(n3857), .ZN(n3858) );
  AOI211_X1 U4533 ( .C1(n3861), .C2(n3860), .A(n3859), .B(n3858), .ZN(n3865)
         );
  INV_X1 U4534 ( .A(n3862), .ZN(n3863) );
  NOR4_X1 U4535 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3871)
         );
  INV_X1 U4536 ( .A(n3867), .ZN(n3870) );
  OAI22_X1 U4537 ( .A1(n3871), .A2(n3870), .B1(n3869), .B2(n3868), .ZN(n3873)
         );
  NAND2_X1 U4538 ( .A1(n3877), .A2(n3876), .ZN(n3878) );
  OAI211_X1 U4539 ( .C1(n3879), .C2(n3881), .A(n3878), .B(B_REG_SCAN_IN), .ZN(
        n3880) );
  MUX2_X1 U4540 ( .A(DATAO_REG_31__SCAN_IN), .B(n3882), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4541 ( .A(DATAO_REG_29__SCAN_IN), .B(n3883), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4542 ( .A(DATAO_REG_28__SCAN_IN), .B(n4033), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4543 ( .A(DATAO_REG_27__SCAN_IN), .B(n4012), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4544 ( .A(DATAO_REG_26__SCAN_IN), .B(n4237), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4545 ( .A(DATAO_REG_25__SCAN_IN), .B(n4246), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4546 ( .A(DATAO_REG_24__SCAN_IN), .B(n4095), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4547 ( .A(DATAO_REG_23__SCAN_IN), .B(n4259), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4548 ( .A(n3884), .B(DATAO_REG_22__SCAN_IN), .S(n3885), .Z(U3572)
         );
  MUX2_X1 U4549 ( .A(DATAO_REG_21__SCAN_IN), .B(n4109), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4550 ( .A(DATAO_REG_20__SCAN_IN), .B(n4279), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4551 ( .A(n4142), .B(DATAO_REG_19__SCAN_IN), .S(n3885), .Z(U3569)
         );
  MUX2_X1 U4552 ( .A(n4300), .B(DATAO_REG_18__SCAN_IN), .S(n3885), .Z(U3568)
         );
  MUX2_X1 U4553 ( .A(DATAO_REG_17__SCAN_IN), .B(n4308), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4554 ( .A(n4320), .B(DATAO_REG_16__SCAN_IN), .S(n3885), .Z(U3566)
         );
  MUX2_X1 U4555 ( .A(DATAO_REG_15__SCAN_IN), .B(n3886), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4556 ( .A(DATAO_REG_14__SCAN_IN), .B(n3887), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4557 ( .A(DATAO_REG_13__SCAN_IN), .B(n3888), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4558 ( .A(DATAO_REG_12__SCAN_IN), .B(n3889), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4559 ( .A(DATAO_REG_11__SCAN_IN), .B(n3890), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4560 ( .A(DATAO_REG_10__SCAN_IN), .B(n3891), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4561 ( .A(DATAO_REG_9__SCAN_IN), .B(n3892), .S(U4043), .Z(U3559) );
  MUX2_X1 U4562 ( .A(DATAO_REG_8__SCAN_IN), .B(n3893), .S(U4043), .Z(U3558) );
  MUX2_X1 U4563 ( .A(DATAO_REG_7__SCAN_IN), .B(n3894), .S(U4043), .Z(U3557) );
  MUX2_X1 U4564 ( .A(DATAO_REG_6__SCAN_IN), .B(n3895), .S(U4043), .Z(U3556) );
  MUX2_X1 U4565 ( .A(DATAO_REG_5__SCAN_IN), .B(n3896), .S(U4043), .Z(U3555) );
  MUX2_X1 U4566 ( .A(DATAO_REG_4__SCAN_IN), .B(n3897), .S(U4043), .Z(U3554) );
  MUX2_X1 U4567 ( .A(DATAO_REG_3__SCAN_IN), .B(n3898), .S(U4043), .Z(U3553) );
  MUX2_X1 U4568 ( .A(DATAO_REG_2__SCAN_IN), .B(n3899), .S(U4043), .Z(U3552) );
  MUX2_X1 U4569 ( .A(DATAO_REG_1__SCAN_IN), .B(n3900), .S(U4043), .Z(U3551) );
  MUX2_X1 U4570 ( .A(DATAO_REG_0__SCAN_IN), .B(n3901), .S(U4043), .Z(U3550) );
  INV_X1 U4571 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4555) );
  NAND3_X1 U4572 ( .A1(n4488), .A2(IR_REG_0__SCAN_IN), .A3(n4555), .ZN(n3909)
         );
  AOI21_X1 U4573 ( .B1(n4555), .B2(n3902), .A(n3904), .ZN(n3903) );
  MUX2_X1 U4574 ( .A(n3904), .B(n3903), .S(n2273), .Z(n3905) );
  AOI22_X1 U4575 ( .A1(n3906), .A2(n3905), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3908) );
  NAND2_X1 U4576 ( .A1(n4486), .A2(ADDR_REG_0__SCAN_IN), .ZN(n3907) );
  NAND3_X1 U4577 ( .A1(n3909), .A2(n3908), .A3(n3907), .ZN(U3240) );
  NAND2_X1 U4578 ( .A1(n3920), .A2(n4388), .ZN(n3919) );
  OAI211_X1 U4579 ( .C1(n2786), .C2(n3912), .A(n4435), .B(n3911), .ZN(n3918)
         );
  OAI211_X1 U4580 ( .C1(n3915), .C2(n3914), .A(n4488), .B(n3913), .ZN(n3917)
         );
  AOI22_X1 U4581 ( .A1(n4486), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3916) );
  NAND4_X1 U4582 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(U3241)
         );
  NAND2_X1 U4583 ( .A1(n3920), .A2(n4386), .ZN(n3928) );
  OAI211_X1 U4584 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3922), .A(n4488), .B(n3921), 
        .ZN(n3927) );
  AOI22_X1 U4585 ( .A1(n4486), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3926) );
  XNOR2_X1 U4586 ( .A(n3923), .B(REG2_REG_3__SCAN_IN), .ZN(n3924) );
  NAND2_X1 U4587 ( .A1(n4435), .A2(n3924), .ZN(n3925) );
  NAND4_X1 U4588 ( .A1(n3928), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(U3243)
         );
  INV_X1 U4589 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3929) );
  MUX2_X1 U4590 ( .A(REG2_REG_19__SCAN_IN), .B(n3929), .S(n4380), .Z(n3945) );
  INV_X1 U4591 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4592 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4516), .B1(n3946), .B2(
        n3930), .ZN(n4484) );
  NOR2_X1 U4593 ( .A1(n3973), .A2(REG2_REG_17__SCAN_IN), .ZN(n3931) );
  AOI21_X1 U4594 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3973), .A(n3931), .ZN(n4473) );
  INV_X1 U4595 ( .A(n3965), .ZN(n4520) );
  INV_X1 U4596 ( .A(n3949), .ZN(n4521) );
  NOR2_X1 U4597 ( .A1(n4434), .A2(n4521), .ZN(n4433) );
  NAND2_X1 U4598 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4523), .ZN(n3936) );
  INV_X1 U4599 ( .A(n4523), .ZN(n4420) );
  AOI22_X1 U4600 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4523), .B1(n4420), .B2(
        n3340), .ZN(n4417) );
  NAND2_X1 U4601 ( .A1(n3951), .A2(REG2_REG_9__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4602 ( .A1(n3951), .A2(REG2_REG_9__SCAN_IN), .B1(n2449), .B2(n4526), .ZN(n4397) );
  NAND2_X1 U4603 ( .A1(n3933), .A2(n4395), .ZN(n3934) );
  NAND2_X1 U4604 ( .A1(n3957), .A2(n3934), .ZN(n3935) );
  INV_X1 U4605 ( .A(n3957), .ZN(n4525) );
  XNOR2_X1 U4606 ( .A(n3934), .B(n4525), .ZN(n4404) );
  NAND2_X1 U4607 ( .A1(n3961), .A2(n3937), .ZN(n3938) );
  INV_X1 U4608 ( .A(n3961), .ZN(n4522) );
  XNOR2_X1 U4609 ( .A(n3937), .B(n4522), .ZN(n4425) );
  NOR2_X1 U4610 ( .A1(n4520), .A2(n3939), .ZN(n3940) );
  NOR2_X1 U4611 ( .A1(n2500), .A2(n4447), .ZN(n4446) );
  NAND2_X1 U4612 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3948), .ZN(n3941) );
  OAI21_X1 U4613 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3948), .A(n3941), .ZN(n4454) );
  INV_X1 U4614 ( .A(n3969), .ZN(n4518) );
  NAND2_X1 U4615 ( .A1(n3942), .A2(n4518), .ZN(n3943) );
  XOR2_X1 U4616 ( .A(n3945), .B(n3944), .Z(n3985) );
  INV_X1 U4617 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4618 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3946), .B1(n4516), .B2(
        n3975), .ZN(n4490) );
  NOR2_X1 U4619 ( .A1(n3973), .A2(REG1_REG_17__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U4620 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3948), .ZN(n3968) );
  INV_X1 U4621 ( .A(n3948), .ZN(n4519) );
  INV_X1 U4622 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4623 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3948), .B1(n4519), .B2(
        n3947), .ZN(n4460) );
  NAND2_X1 U4624 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3949), .ZN(n3964) );
  AOI22_X1 U4625 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3949), .B1(n4521), .B2(
        n3349), .ZN(n4443) );
  NAND2_X1 U4626 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4523), .ZN(n3960) );
  AOI22_X1 U4627 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4523), .B1(n4420), .B2(
        n3359), .ZN(n4414) );
  NAND2_X1 U4628 ( .A1(n3951), .A2(REG1_REG_9__SCAN_IN), .ZN(n3956) );
  INV_X1 U4629 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4630 ( .A1(n3951), .A2(REG1_REG_9__SCAN_IN), .B1(n3950), .B2(n4526), .ZN(n4394) );
  INV_X1 U4631 ( .A(n3952), .ZN(n4381) );
  AOI22_X1 U4632 ( .A1(n3954), .A2(REG1_REG_8__SCAN_IN), .B1(n4381), .B2(n3953), .ZN(n3955) );
  INV_X1 U4633 ( .A(n3955), .ZN(n4393) );
  NAND2_X1 U4634 ( .A1(n4394), .A2(n4393), .ZN(n4392) );
  NAND2_X1 U4635 ( .A1(n3956), .A2(n4392), .ZN(n3958) );
  NAND2_X1 U4636 ( .A1(n3957), .A2(n3958), .ZN(n3959) );
  NAND2_X1 U4637 ( .A1(n3961), .A2(n3962), .ZN(n3963) );
  XNOR2_X1 U4638 ( .A(n3962), .B(n4522), .ZN(n4430) );
  NAND2_X1 U4639 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4430), .ZN(n4429) );
  NAND2_X1 U4640 ( .A1(n3963), .A2(n4429), .ZN(n4442) );
  NAND2_X1 U4641 ( .A1(n4443), .A2(n4442), .ZN(n4441) );
  NAND2_X1 U4642 ( .A1(n3964), .A2(n4441), .ZN(n3966) );
  NAND2_X1 U4643 ( .A1(n3965), .A2(n3966), .ZN(n3967) );
  XNOR2_X1 U4644 ( .A(n3966), .B(n4520), .ZN(n4451) );
  NAND2_X1 U4645 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4451), .ZN(n4450) );
  NAND2_X1 U4646 ( .A1(n3967), .A2(n4450), .ZN(n4459) );
  NAND2_X1 U4647 ( .A1(n4460), .A2(n4459), .ZN(n4458) );
  NOR2_X1 U4648 ( .A1(n3969), .A2(n3970), .ZN(n3971) );
  INV_X1 U4649 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4650 ( .A1(n3973), .A2(n3972), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4517), .ZN(n4476) );
  NAND2_X1 U4651 ( .A1(n4490), .A2(n4489), .ZN(n4487) );
  OAI21_X1 U4652 ( .B1(n3975), .B2(n4516), .A(n4487), .ZN(n3978) );
  INV_X1 U4653 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3976) );
  MUX2_X1 U4654 ( .A(n3976), .B(REG1_REG_19__SCAN_IN), .S(n4380), .Z(n3977) );
  XNOR2_X1 U4655 ( .A(n3978), .B(n3977), .ZN(n3983) );
  NAND2_X1 U4656 ( .A1(n4486), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3979) );
  OAI211_X1 U4657 ( .C1(n4493), .C2(n3981), .A(n3980), .B(n3979), .ZN(n3982)
         );
  OAI21_X1 U4658 ( .B1(n3985), .B2(n4482), .A(n3984), .ZN(U3259) );
  NOR2_X2 U4659 ( .A1(n4231), .A2(n4233), .ZN(n4230) );
  XNOR2_X1 U4660 ( .A(n4230), .B(n3986), .ZN(n4332) );
  NOR2_X1 U4661 ( .A1(n3988), .A2(n3987), .ZN(n4232) );
  AOI21_X1 U4662 ( .B1(n3989), .B2(n4318), .A(n4232), .ZN(n4329) );
  MUX2_X1 U4663 ( .A(n3990), .B(n4329), .S(n4200), .Z(n3991) );
  OAI21_X1 U4664 ( .B1(n4332), .B2(n4179), .A(n3991), .ZN(U3260) );
  XNOR2_X1 U4665 ( .A(n3993), .B(n3992), .ZN(n4003) );
  OAI22_X1 U4666 ( .A1(n4219), .A2(n3995), .B1(n3994), .B2(n4200), .ZN(n3996)
         );
  AOI21_X1 U4667 ( .B1(n4033), .B2(n4027), .A(n3996), .ZN(n4002) );
  OAI22_X1 U4668 ( .A1(n3998), .A2(n4179), .B1(n3997), .B2(n4494), .ZN(n3999)
         );
  OAI21_X1 U4669 ( .B1(n4000), .B2(n3999), .A(n4200), .ZN(n4001) );
  OAI211_X1 U4670 ( .C1(n4003), .C2(n4203), .A(n4002), .B(n4001), .ZN(U3354)
         );
  INV_X1 U4671 ( .A(n4004), .ZN(n4018) );
  NAND2_X1 U4672 ( .A1(n4005), .A2(n4504), .ZN(n4006) );
  OAI21_X1 U4673 ( .B1(n4200), .B2(n4007), .A(n4006), .ZN(n4011) );
  OAI22_X1 U4674 ( .A1(n4009), .A2(n4220), .B1(n4008), .B2(n4219), .ZN(n4010)
         );
  AOI211_X1 U4675 ( .C1(n4027), .C2(n4012), .A(n4011), .B(n4010), .ZN(n4013)
         );
  OAI21_X1 U4676 ( .B1(n4014), .B2(n4179), .A(n4013), .ZN(n4015) );
  AOI21_X1 U4677 ( .B1(n4016), .B2(n4200), .A(n4015), .ZN(n4017) );
  OAI21_X1 U4678 ( .B1(n4018), .B2(n4203), .A(n4017), .ZN(U3262) );
  OAI21_X1 U4679 ( .B1(n4022), .B2(n4020), .A(n4019), .ZN(n4021) );
  NAND2_X1 U4680 ( .A1(n4021), .A2(n4206), .ZN(n4239) );
  XNOR2_X1 U4681 ( .A(n4023), .B(n4022), .ZN(n4242) );
  NAND2_X1 U4682 ( .A1(n4242), .A2(n4210), .ZN(n4036) );
  OAI22_X1 U4683 ( .A1(n4025), .A2(n4494), .B1(n4024), .B2(n4200), .ZN(n4026)
         );
  AOI21_X1 U4684 ( .B1(n4027), .B2(n4237), .A(n4026), .ZN(n4028) );
  OAI21_X1 U4685 ( .B1(n4029), .B2(n4219), .A(n4028), .ZN(n4032) );
  NAND2_X1 U4686 ( .A1(n4045), .A2(n4236), .ZN(n4030) );
  NAND2_X1 U4687 ( .A1(n2059), .A2(n4030), .ZN(n4339) );
  NOR2_X1 U4688 ( .A1(n4339), .A2(n4179), .ZN(n4031) );
  AOI211_X1 U4689 ( .C1(n4034), .C2(n4033), .A(n4032), .B(n4031), .ZN(n4035)
         );
  OAI211_X1 U4690 ( .C1(n4227), .C2(n4239), .A(n4036), .B(n4035), .ZN(U3263)
         );
  INV_X1 U4691 ( .A(n4037), .ZN(n4039) );
  OAI21_X1 U4692 ( .B1(n2062), .B2(n4039), .A(n4038), .ZN(n4040) );
  XNOR2_X1 U4693 ( .A(n4040), .B(n4043), .ZN(n4041) );
  NAND2_X1 U4694 ( .A1(n4041), .A2(n4206), .ZN(n4248) );
  XOR2_X1 U4695 ( .A(n4043), .B(n4042), .Z(n4251) );
  NAND2_X1 U4696 ( .A1(n4251), .A2(n4210), .ZN(n4053) );
  OR2_X1 U4697 ( .A1(n4064), .A2(n4048), .ZN(n4044) );
  NAND2_X1 U4698 ( .A1(n4045), .A2(n4044), .ZN(n4343) );
  INV_X1 U4699 ( .A(n4343), .ZN(n4051) );
  AOI22_X1 U4700 ( .A1(n4046), .A2(n4504), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4227), .ZN(n4047) );
  OAI21_X1 U4701 ( .B1(n4262), .B2(n4217), .A(n4047), .ZN(n4050) );
  OAI22_X1 U4702 ( .A1(n4249), .A2(n4220), .B1(n4219), .B2(n4048), .ZN(n4049)
         );
  AOI211_X1 U4703 ( .C1(n4051), .C2(n4508), .A(n4050), .B(n4049), .ZN(n4052)
         );
  OAI211_X1 U4704 ( .C1(n4227), .C2(n4248), .A(n4053), .B(n4052), .ZN(U3264)
         );
  XNOR2_X1 U4705 ( .A(n4054), .B(n4056), .ZN(n4255) );
  INV_X1 U4706 ( .A(n4255), .ZN(n4069) );
  NOR2_X1 U4707 ( .A1(n2062), .A2(n4055), .ZN(n4057) );
  XNOR2_X1 U4708 ( .A(n4057), .B(n4056), .ZN(n4061) );
  OAI22_X1 U4709 ( .A1(n4058), .A2(n4323), .B1(n4062), .B2(n4168), .ZN(n4059)
         );
  AOI21_X1 U4710 ( .B1(n4319), .B2(n4237), .A(n4059), .ZN(n4060) );
  OAI21_X1 U4711 ( .B1(n4061), .B2(n4172), .A(n4060), .ZN(n4254) );
  NOR2_X1 U4712 ( .A1(n4074), .A2(n4062), .ZN(n4063) );
  OR2_X1 U4713 ( .A1(n4064), .A2(n4063), .ZN(n4347) );
  AOI22_X1 U4714 ( .A1(n4065), .A2(n4504), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4227), .ZN(n4066) );
  OAI21_X1 U4715 ( .B1(n4347), .B2(n4179), .A(n4066), .ZN(n4067) );
  AOI21_X1 U4716 ( .B1(n4254), .B2(n4200), .A(n4067), .ZN(n4068) );
  OAI21_X1 U4717 ( .B1(n4069), .B2(n4203), .A(n4068), .ZN(U3265) );
  XNOR2_X1 U4718 ( .A(n4070), .B(n4073), .ZN(n4071) );
  NAND2_X1 U4719 ( .A1(n4071), .A2(n4206), .ZN(n4261) );
  XOR2_X1 U4720 ( .A(n4073), .B(n4072), .Z(n4264) );
  NAND2_X1 U4721 ( .A1(n4264), .A2(n4210), .ZN(n4084) );
  INV_X1 U4722 ( .A(n4100), .ZN(n4076) );
  INV_X1 U4723 ( .A(n4074), .ZN(n4075) );
  OAI21_X1 U4724 ( .B1(n4076), .B2(n4079), .A(n4075), .ZN(n4351) );
  INV_X1 U4725 ( .A(n4351), .ZN(n4082) );
  AOI22_X1 U4726 ( .A1(n4077), .A2(n4504), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4227), .ZN(n4078) );
  OAI21_X1 U4727 ( .B1(n4107), .B2(n4217), .A(n4078), .ZN(n4081) );
  OAI22_X1 U4728 ( .A1(n4262), .A2(n4220), .B1(n4219), .B2(n4079), .ZN(n4080)
         );
  AOI211_X1 U4729 ( .C1(n4082), .C2(n4508), .A(n4081), .B(n4080), .ZN(n4083)
         );
  OAI211_X1 U4730 ( .C1(n4227), .C2(n4261), .A(n4084), .B(n4083), .ZN(U3266)
         );
  XOR2_X1 U4731 ( .A(n4092), .B(n4085), .Z(n4268) );
  INV_X1 U4732 ( .A(n4268), .ZN(n4105) );
  OAI21_X1 U4733 ( .B1(n4124), .B2(n4087), .A(n4086), .ZN(n4106) );
  INV_X1 U4734 ( .A(n4088), .ZN(n4089) );
  AOI21_X1 U4735 ( .B1(n4106), .B2(n4090), .A(n4089), .ZN(n4091) );
  XOR2_X1 U4736 ( .A(n4092), .B(n4091), .Z(n4097) );
  OAI22_X1 U4737 ( .A1(n4283), .A2(n4323), .B1(n4168), .B2(n4093), .ZN(n4094)
         );
  AOI21_X1 U4738 ( .B1(n4319), .B2(n4095), .A(n4094), .ZN(n4096) );
  OAI21_X1 U4739 ( .B1(n4097), .B2(n4172), .A(n4096), .ZN(n4267) );
  NAND2_X1 U4740 ( .A1(n4114), .A2(n4098), .ZN(n4099) );
  NAND2_X1 U4741 ( .A1(n4100), .A2(n4099), .ZN(n4355) );
  AOI22_X1 U4742 ( .A1(n4101), .A2(n4504), .B1(n4227), .B2(
        REG2_REG_23__SCAN_IN), .ZN(n4102) );
  OAI21_X1 U4743 ( .B1(n4355), .B2(n4179), .A(n4102), .ZN(n4103) );
  AOI21_X1 U4744 ( .B1(n4267), .B2(n4200), .A(n4103), .ZN(n4104) );
  OAI21_X1 U4745 ( .B1(n4105), .B2(n4203), .A(n4104), .ZN(U3267) );
  XNOR2_X1 U4746 ( .A(n4106), .B(n4117), .ZN(n4111) );
  OAI22_X1 U4747 ( .A1(n4107), .A2(n4282), .B1(n4112), .B2(n4168), .ZN(n4108)
         );
  AOI21_X1 U4748 ( .B1(n4278), .B2(n4109), .A(n4108), .ZN(n4110) );
  OAI21_X1 U4749 ( .B1(n4111), .B2(n4172), .A(n4110), .ZN(n4272) );
  OR2_X1 U4750 ( .A1(n4128), .A2(n4112), .ZN(n4113) );
  NAND2_X1 U4751 ( .A1(n4114), .A2(n4113), .ZN(n4359) );
  AOI22_X1 U4752 ( .A1(n4227), .A2(REG2_REG_22__SCAN_IN), .B1(n4115), .B2(
        n4504), .ZN(n4116) );
  OAI21_X1 U4753 ( .B1(n4359), .B2(n4179), .A(n4116), .ZN(n4121) );
  NOR2_X1 U4754 ( .A1(n4118), .A2(n4117), .ZN(n4271) );
  INV_X1 U4755 ( .A(n4273), .ZN(n4119) );
  NOR3_X1 U4756 ( .A1(n4271), .A2(n4119), .A3(n4203), .ZN(n4120) );
  AOI211_X1 U4757 ( .C1(n4200), .C2(n4272), .A(n4121), .B(n4120), .ZN(n4122)
         );
  INV_X1 U4758 ( .A(n4122), .ZN(U3268) );
  INV_X1 U4759 ( .A(n4127), .ZN(n4123) );
  XNOR2_X1 U4760 ( .A(n4124), .B(n4123), .ZN(n4125) );
  NAND2_X1 U4761 ( .A1(n4125), .A2(n4206), .ZN(n4281) );
  XOR2_X1 U4762 ( .A(n4127), .B(n4126), .Z(n4285) );
  NAND2_X1 U4763 ( .A1(n4285), .A2(n4210), .ZN(n4138) );
  INV_X1 U4764 ( .A(n4128), .ZN(n4129) );
  OAI21_X1 U4765 ( .B1(n4152), .B2(n4133), .A(n4129), .ZN(n4363) );
  INV_X1 U4766 ( .A(n4363), .ZN(n4136) );
  AOI22_X1 U4767 ( .A1(n4227), .A2(REG2_REG_21__SCAN_IN), .B1(n4130), .B2(
        n4504), .ZN(n4131) );
  OAI21_X1 U4768 ( .B1(n4217), .B2(n4132), .A(n4131), .ZN(n4135) );
  OAI22_X1 U4769 ( .A1(n4283), .A2(n4220), .B1(n4219), .B2(n4133), .ZN(n4134)
         );
  AOI211_X1 U4770 ( .C1(n4136), .C2(n4508), .A(n4135), .B(n4134), .ZN(n4137)
         );
  OAI211_X1 U4771 ( .C1(n4227), .C2(n4281), .A(n4138), .B(n4137), .ZN(U3269)
         );
  NAND2_X1 U4772 ( .A1(n4140), .A2(n4139), .ZN(n4141) );
  XNOR2_X1 U4773 ( .A(n4141), .B(n2094), .ZN(n4150) );
  AOI22_X1 U4774 ( .A1(n4142), .A2(n4278), .B1(n4153), .B2(n4318), .ZN(n4143)
         );
  OAI21_X1 U4775 ( .B1(n4144), .B2(n4282), .A(n4143), .ZN(n4149) );
  XNOR2_X1 U4776 ( .A(n4145), .B(n4146), .ZN(n4292) );
  NOR2_X1 U4777 ( .A1(n4292), .A2(n4147), .ZN(n4148) );
  AOI211_X1 U4778 ( .C1(n4206), .C2(n4150), .A(n4149), .B(n4148), .ZN(n4291)
         );
  AOI22_X1 U4779 ( .A1(n4227), .A2(REG2_REG_20__SCAN_IN), .B1(n4151), .B2(
        n4504), .ZN(n4155) );
  INV_X1 U4780 ( .A(n4152), .ZN(n4289) );
  NAND2_X1 U4781 ( .A1(n4176), .A2(n4153), .ZN(n4288) );
  NAND3_X1 U4782 ( .A1(n4289), .A2(n4508), .A3(n4288), .ZN(n4154) );
  OAI211_X1 U4783 ( .C1(n4292), .C2(n4156), .A(n4155), .B(n4154), .ZN(n4157)
         );
  INV_X1 U4784 ( .A(n4157), .ZN(n4158) );
  OAI21_X1 U4785 ( .B1(n4291), .B2(n4215), .A(n4158), .ZN(U3270) );
  XNOR2_X1 U4786 ( .A(n4160), .B(n4159), .ZN(n4294) );
  INV_X1 U4787 ( .A(n4294), .ZN(n4182) );
  OAI21_X1 U4788 ( .B1(n4205), .B2(n4162), .A(n4161), .ZN(n4188) );
  INV_X1 U4789 ( .A(n4163), .ZN(n4165) );
  OAI21_X1 U4790 ( .B1(n4188), .B2(n4165), .A(n4164), .ZN(n4167) );
  XNOR2_X1 U4791 ( .A(n4167), .B(n4166), .ZN(n4173) );
  OAI22_X1 U4792 ( .A1(n4221), .A2(n4323), .B1(n4169), .B2(n4168), .ZN(n4170)
         );
  AOI21_X1 U4793 ( .B1(n4279), .B2(n4319), .A(n4170), .ZN(n4171) );
  OAI21_X1 U4794 ( .B1(n4173), .B2(n4172), .A(n4171), .ZN(n4293) );
  NAND2_X1 U4795 ( .A1(n4194), .A2(n4174), .ZN(n4175) );
  NAND2_X1 U4796 ( .A1(n4176), .A2(n4175), .ZN(n4368) );
  AOI22_X1 U4797 ( .A1(n4215), .A2(REG2_REG_19__SCAN_IN), .B1(n4177), .B2(
        n4504), .ZN(n4178) );
  OAI21_X1 U4798 ( .B1(n4368), .B2(n4179), .A(n4178), .ZN(n4180) );
  AOI21_X1 U4799 ( .B1(n4293), .B2(n4200), .A(n4180), .ZN(n4181) );
  OAI21_X1 U4800 ( .B1(n4182), .B2(n4203), .A(n4181), .ZN(U3271) );
  OAI21_X1 U4801 ( .B1(n4185), .B2(n4184), .A(n4183), .ZN(n4186) );
  INV_X1 U4802 ( .A(n4186), .ZN(n4298) );
  XNOR2_X1 U4803 ( .A(n4188), .B(n4187), .ZN(n4193) );
  AOI22_X1 U4804 ( .A1(n4308), .A2(n4278), .B1(n4318), .B2(n4189), .ZN(n4190)
         );
  OAI21_X1 U4805 ( .B1(n4191), .B2(n4282), .A(n4190), .ZN(n4192) );
  AOI21_X1 U4806 ( .B1(n4193), .B2(n4206), .A(n4192), .ZN(n4297) );
  INV_X1 U4807 ( .A(n4297), .ZN(n4201) );
  OAI211_X1 U4808 ( .C1(n4211), .C2(n4195), .A(n4194), .B(n4537), .ZN(n4296)
         );
  NOR2_X1 U4809 ( .A1(n4296), .A2(n4196), .ZN(n4199) );
  OAI22_X1 U4810 ( .A1(n4200), .A2(n3930), .B1(n4197), .B2(n4494), .ZN(n4198)
         );
  AOI211_X1 U4811 ( .C1(n4201), .C2(n4200), .A(n4199), .B(n4198), .ZN(n4202)
         );
  OAI21_X1 U4812 ( .B1(n4298), .B2(n4203), .A(n4202), .ZN(U3272) );
  INV_X1 U4813 ( .A(n4208), .ZN(n4204) );
  XNOR2_X1 U4814 ( .A(n4205), .B(n4204), .ZN(n4207) );
  NAND2_X1 U4815 ( .A1(n4207), .A2(n4206), .ZN(n4302) );
  XNOR2_X1 U4816 ( .A(n4209), .B(n4208), .ZN(n4305) );
  NAND2_X1 U4817 ( .A1(n4305), .A2(n4210), .ZN(n4226) );
  INV_X1 U4818 ( .A(n4211), .ZN(n4212) );
  OAI21_X1 U4819 ( .B1(n4213), .B2(n4218), .A(n4212), .ZN(n4373) );
  INV_X1 U4820 ( .A(n4373), .ZN(n4224) );
  AOI22_X1 U4821 ( .A1(n4215), .A2(REG2_REG_17__SCAN_IN), .B1(n4214), .B2(
        n4504), .ZN(n4216) );
  OAI21_X1 U4822 ( .B1(n4217), .B2(n4303), .A(n4216), .ZN(n4223) );
  OAI22_X1 U4823 ( .A1(n4221), .A2(n4220), .B1(n4219), .B2(n4218), .ZN(n4222)
         );
  AOI211_X1 U4824 ( .C1(n4224), .C2(n4508), .A(n4223), .B(n4222), .ZN(n4225)
         );
  OAI211_X1 U4825 ( .C1(n4227), .C2(n4302), .A(n4226), .B(n4225), .ZN(U3273)
         );
  NOR2_X1 U4826 ( .A1(n4561), .A2(n4329), .ZN(n4228) );
  AOI21_X1 U4827 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4561), .A(n4228), .ZN(n4229) );
  OAI21_X1 U4828 ( .B1(n4332), .B2(n4328), .A(n4229), .ZN(U3549) );
  AOI21_X1 U4829 ( .B1(n4233), .B2(n4231), .A(n4230), .ZN(n4389) );
  INV_X1 U4830 ( .A(n4389), .ZN(n4335) );
  INV_X1 U4831 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4234) );
  AOI21_X1 U4832 ( .B1(n4233), .B2(n4318), .A(n4232), .ZN(n4391) );
  MUX2_X1 U4833 ( .A(n4234), .B(n4391), .S(n4564), .Z(n4235) );
  OAI21_X1 U4834 ( .B1(n4335), .B2(n4328), .A(n4235), .ZN(U3548) );
  INV_X1 U4835 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U4836 ( .A1(n4237), .A2(n4278), .B1(n4236), .B2(n4318), .ZN(n4238)
         );
  OAI211_X1 U4837 ( .C1(n4240), .C2(n4282), .A(n4239), .B(n4238), .ZN(n4241)
         );
  AOI21_X1 U4838 ( .B1(n4242), .B2(n4546), .A(n4241), .ZN(n4336) );
  MUX2_X1 U4839 ( .A(n4243), .B(n4336), .S(n4564), .Z(n4244) );
  OAI21_X1 U4840 ( .B1(n4328), .B2(n4339), .A(n4244), .ZN(U3545) );
  INV_X1 U4841 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U4842 ( .A1(n4246), .A2(n4278), .B1(n4245), .B2(n4318), .ZN(n4247)
         );
  OAI211_X1 U4843 ( .C1(n4249), .C2(n4282), .A(n4248), .B(n4247), .ZN(n4250)
         );
  AOI21_X1 U4844 ( .B1(n4251), .B2(n4546), .A(n4250), .ZN(n4340) );
  MUX2_X1 U4845 ( .A(n4252), .B(n4340), .S(n4564), .Z(n4253) );
  OAI21_X1 U4846 ( .B1(n4328), .B2(n4343), .A(n4253), .ZN(U3544) );
  INV_X1 U4847 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4256) );
  AOI21_X1 U4848 ( .B1(n4255), .B2(n4546), .A(n4254), .ZN(n4344) );
  MUX2_X1 U4849 ( .A(n4256), .B(n4344), .S(n4564), .Z(n4257) );
  OAI21_X1 U4850 ( .B1(n4328), .B2(n4347), .A(n4257), .ZN(U3543) );
  INV_X1 U4851 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4265) );
  AOI22_X1 U4852 ( .A1(n4259), .A2(n4278), .B1(n4318), .B2(n4258), .ZN(n4260)
         );
  OAI211_X1 U4853 ( .C1(n4262), .C2(n4282), .A(n4261), .B(n4260), .ZN(n4263)
         );
  AOI21_X1 U4854 ( .B1(n4264), .B2(n4546), .A(n4263), .ZN(n4348) );
  MUX2_X1 U4855 ( .A(n4265), .B(n4348), .S(n4564), .Z(n4266) );
  OAI21_X1 U4856 ( .B1(n4328), .B2(n4351), .A(n4266), .ZN(U3542) );
  INV_X1 U4857 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4269) );
  AOI21_X1 U4858 ( .B1(n4268), .B2(n4546), .A(n4267), .ZN(n4352) );
  MUX2_X1 U4859 ( .A(n4269), .B(n4352), .S(n4564), .Z(n4270) );
  OAI21_X1 U4860 ( .B1(n4328), .B2(n4355), .A(n4270), .ZN(U3541) );
  INV_X1 U4861 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4275) );
  NOR2_X1 U4862 ( .A1(n4271), .A2(n4315), .ZN(n4274) );
  AOI21_X1 U4863 ( .B1(n4274), .B2(n4273), .A(n4272), .ZN(n4356) );
  MUX2_X1 U4864 ( .A(n4275), .B(n4356), .S(n4564), .Z(n4276) );
  OAI21_X1 U4865 ( .B1(n4328), .B2(n4359), .A(n4276), .ZN(U3540) );
  INV_X1 U4866 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4286) );
  AOI22_X1 U4867 ( .A1(n4279), .A2(n4278), .B1(n4277), .B2(n4318), .ZN(n4280)
         );
  OAI211_X1 U4868 ( .C1(n4283), .C2(n4282), .A(n4281), .B(n4280), .ZN(n4284)
         );
  AOI21_X1 U4869 ( .B1(n4285), .B2(n4546), .A(n4284), .ZN(n4360) );
  MUX2_X1 U4870 ( .A(n4286), .B(n4360), .S(n4564), .Z(n4287) );
  OAI21_X1 U4871 ( .B1(n4328), .B2(n4363), .A(n4287), .ZN(U3539) );
  NAND3_X1 U4872 ( .A1(n4289), .A2(n4288), .A3(n4537), .ZN(n4290) );
  OAI211_X1 U4873 ( .C1(n4292), .C2(n4532), .A(n4291), .B(n4290), .ZN(n4364)
         );
  MUX2_X1 U4874 ( .A(REG1_REG_20__SCAN_IN), .B(n4364), .S(n4564), .Z(U3538) );
  AOI21_X1 U4875 ( .B1(n4294), .B2(n4546), .A(n4293), .ZN(n4365) );
  MUX2_X1 U4876 ( .A(n3976), .B(n4365), .S(n4564), .Z(n4295) );
  OAI21_X1 U4877 ( .B1(n4328), .B2(n4368), .A(n4295), .ZN(U3537) );
  OAI211_X1 U4878 ( .C1(n4298), .C2(n4315), .A(n4297), .B(n4296), .ZN(n4369)
         );
  MUX2_X1 U4879 ( .A(REG1_REG_18__SCAN_IN), .B(n4369), .S(n4564), .Z(U3536) );
  AOI22_X1 U4880 ( .A1(n4300), .A2(n4319), .B1(n4299), .B2(n4318), .ZN(n4301)
         );
  OAI211_X1 U4881 ( .C1(n4303), .C2(n4323), .A(n4302), .B(n4301), .ZN(n4304)
         );
  AOI21_X1 U4882 ( .B1(n4305), .B2(n4546), .A(n4304), .ZN(n4371) );
  MUX2_X1 U4883 ( .A(n4371), .B(n3972), .S(n4561), .Z(n4306) );
  OAI21_X1 U4884 ( .B1(n4328), .B2(n4373), .A(n4306), .ZN(U3535) );
  AOI22_X1 U4885 ( .A1(n4308), .A2(n4319), .B1(n4318), .B2(n4307), .ZN(n4309)
         );
  OAI21_X1 U4886 ( .B1(n4310), .B2(n4323), .A(n4309), .ZN(n4311) );
  AOI21_X1 U4887 ( .B1(n4312), .B2(n4537), .A(n4311), .ZN(n4314) );
  OAI211_X1 U4888 ( .C1(n4316), .C2(n4315), .A(n4314), .B(n4313), .ZN(n4374)
         );
  MUX2_X1 U4889 ( .A(REG1_REG_16__SCAN_IN), .B(n4374), .S(n4564), .Z(U3534) );
  AOI22_X1 U4890 ( .A1(n4320), .A2(n4319), .B1(n4318), .B2(n4317), .ZN(n4321)
         );
  OAI211_X1 U4891 ( .C1(n4324), .C2(n4323), .A(n4322), .B(n4321), .ZN(n4325)
         );
  AOI21_X1 U4892 ( .B1(n4326), .B2(n4546), .A(n4325), .ZN(n4376) );
  MUX2_X1 U4893 ( .A(n4376), .B(n3947), .S(n4561), .Z(n4327) );
  OAI21_X1 U4894 ( .B1(n4328), .B2(n4379), .A(n4327), .ZN(U3533) );
  NOR2_X1 U4895 ( .A1(n4552), .A2(n4329), .ZN(n4330) );
  AOI21_X1 U4896 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4552), .A(n4330), .ZN(n4331) );
  OAI21_X1 U4897 ( .B1(n4332), .B2(n4378), .A(n4331), .ZN(U3517) );
  INV_X1 U4898 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4333) );
  MUX2_X1 U4899 ( .A(n4333), .B(n4391), .S(n4554), .Z(n4334) );
  OAI21_X1 U4900 ( .B1(n4335), .B2(n4378), .A(n4334), .ZN(U3516) );
  INV_X1 U4901 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4337) );
  MUX2_X1 U4902 ( .A(n4337), .B(n4336), .S(n4554), .Z(n4338) );
  OAI21_X1 U4903 ( .B1(n4339), .B2(n4378), .A(n4338), .ZN(U3513) );
  INV_X1 U4904 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4341) );
  MUX2_X1 U4905 ( .A(n4341), .B(n4340), .S(n4554), .Z(n4342) );
  OAI21_X1 U4906 ( .B1(n4343), .B2(n4378), .A(n4342), .ZN(U3512) );
  INV_X1 U4907 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4345) );
  MUX2_X1 U4908 ( .A(n4345), .B(n4344), .S(n4554), .Z(n4346) );
  OAI21_X1 U4909 ( .B1(n4347), .B2(n4378), .A(n4346), .ZN(U3511) );
  INV_X1 U4910 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4349) );
  MUX2_X1 U4911 ( .A(n4349), .B(n4348), .S(n4554), .Z(n4350) );
  OAI21_X1 U4912 ( .B1(n4351), .B2(n4378), .A(n4350), .ZN(U3510) );
  INV_X1 U4913 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4353) );
  MUX2_X1 U4914 ( .A(n4353), .B(n4352), .S(n4554), .Z(n4354) );
  OAI21_X1 U4915 ( .B1(n4355), .B2(n4378), .A(n4354), .ZN(U3509) );
  INV_X1 U4916 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4357) );
  MUX2_X1 U4917 ( .A(n4357), .B(n4356), .S(n4554), .Z(n4358) );
  OAI21_X1 U4918 ( .B1(n4359), .B2(n4378), .A(n4358), .ZN(U3508) );
  INV_X1 U4919 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4361) );
  MUX2_X1 U4920 ( .A(n4361), .B(n4360), .S(n4554), .Z(n4362) );
  OAI21_X1 U4921 ( .B1(n4363), .B2(n4378), .A(n4362), .ZN(U3507) );
  MUX2_X1 U4922 ( .A(REG0_REG_20__SCAN_IN), .B(n4364), .S(n4554), .Z(U3506) );
  INV_X1 U4923 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4366) );
  MUX2_X1 U4924 ( .A(n4366), .B(n4365), .S(n4554), .Z(n4367) );
  OAI21_X1 U4925 ( .B1(n4368), .B2(n4378), .A(n4367), .ZN(U3505) );
  MUX2_X1 U4926 ( .A(REG0_REG_18__SCAN_IN), .B(n4369), .S(n4554), .Z(U3503) );
  INV_X1 U4927 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4370) );
  MUX2_X1 U4928 ( .A(n4371), .B(n4370), .S(n4552), .Z(n4372) );
  OAI21_X1 U4929 ( .B1(n4373), .B2(n4378), .A(n4372), .ZN(U3501) );
  MUX2_X1 U4930 ( .A(REG0_REG_16__SCAN_IN), .B(n4374), .S(n4554), .Z(U3499) );
  INV_X1 U4931 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4375) );
  MUX2_X1 U4932 ( .A(n4376), .B(n4375), .S(n4552), .Z(n4377) );
  OAI21_X1 U4933 ( .B1(n4379), .B2(n4378), .A(n4377), .ZN(U3497) );
  MUX2_X1 U4934 ( .A(DATAI_21_), .B(n2667), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U4935 ( .A(n4380), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4936 ( .A(DATAI_8_), .B(n4381), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4937 ( .A(n4382), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4938 ( .A(n4383), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4939 ( .A(n4384), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4940 ( .A(DATAI_4_), .B(n4385), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4941 ( .A(n4386), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4942 ( .A(n4387), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4943 ( .A(n4388), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4944 ( .A1(n4389), .A2(n4508), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4215), .ZN(n4390) );
  OAI21_X1 U4945 ( .B1(n4227), .B2(n4391), .A(n4390), .ZN(U3261) );
  OAI211_X1 U4946 ( .C1(n4394), .C2(n4393), .A(n4488), .B(n4392), .ZN(n4399)
         );
  OAI211_X1 U4947 ( .C1(n4397), .C2(n4396), .A(n4435), .B(n4395), .ZN(n4398)
         );
  OAI211_X1 U4948 ( .C1(n4493), .C2(n4526), .A(n4399), .B(n4398), .ZN(n4400)
         );
  AOI211_X1 U4949 ( .C1(n4486), .C2(ADDR_REG_9__SCAN_IN), .A(n4401), .B(n4400), 
        .ZN(n4402) );
  INV_X1 U4950 ( .A(n4402), .ZN(U3249) );
  OAI211_X1 U4951 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4404), .A(n4435), .B(n4403), .ZN(n4406) );
  NAND2_X1 U4952 ( .A1(n4406), .A2(n4405), .ZN(n4407) );
  AOI21_X1 U4953 ( .B1(n4486), .B2(ADDR_REG_10__SCAN_IN), .A(n4407), .ZN(n4411) );
  OAI211_X1 U4954 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4409), .A(n4488), .B(n4408), .ZN(n4410) );
  OAI211_X1 U4955 ( .C1(n4493), .C2(n4525), .A(n4411), .B(n4410), .ZN(U3250)
         );
  OAI211_X1 U4956 ( .C1(n4414), .C2(n4413), .A(n4488), .B(n4412), .ZN(n4419)
         );
  OAI211_X1 U4957 ( .C1(n4417), .C2(n4416), .A(n4435), .B(n4415), .ZN(n4418)
         );
  OAI211_X1 U4958 ( .C1(n4493), .C2(n4420), .A(n4419), .B(n4418), .ZN(n4421)
         );
  AOI211_X1 U4959 ( .C1(n4486), .C2(ADDR_REG_11__SCAN_IN), .A(n4422), .B(n4421), .ZN(n4423) );
  INV_X1 U4960 ( .A(n4423), .ZN(U3251) );
  OAI211_X1 U4961 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4425), .A(n4435), .B(n4424), .ZN(n4427) );
  NAND2_X1 U4962 ( .A1(n4427), .A2(n4426), .ZN(n4428) );
  AOI21_X1 U4963 ( .B1(n4486), .B2(ADDR_REG_12__SCAN_IN), .A(n4428), .ZN(n4432) );
  OAI211_X1 U4964 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4430), .A(n4488), .B(n4429), .ZN(n4431) );
  OAI211_X1 U4965 ( .C1(n4493), .C2(n4522), .A(n4432), .B(n4431), .ZN(U3252)
         );
  AOI21_X1 U4966 ( .B1(n4434), .B2(n4521), .A(n4433), .ZN(n4438) );
  OAI21_X1 U4967 ( .B1(n4438), .B2(n4437), .A(n4435), .ZN(n4436) );
  AOI21_X1 U4968 ( .B1(n4438), .B2(n4437), .A(n4436), .ZN(n4440) );
  AOI211_X1 U4969 ( .C1(n4486), .C2(ADDR_REG_13__SCAN_IN), .A(n4440), .B(n4439), .ZN(n4445) );
  OAI211_X1 U4970 ( .C1(n4443), .C2(n4442), .A(n4488), .B(n4441), .ZN(n4444)
         );
  OAI211_X1 U4971 ( .C1(n4493), .C2(n4521), .A(n4445), .B(n4444), .ZN(U3253)
         );
  AOI211_X1 U4972 ( .C1(n2500), .C2(n4447), .A(n4446), .B(n4482), .ZN(n4448)
         );
  AOI211_X1 U4973 ( .C1(n4486), .C2(ADDR_REG_14__SCAN_IN), .A(n4449), .B(n4448), .ZN(n4453) );
  OAI211_X1 U4974 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4451), .A(n4488), .B(n4450), .ZN(n4452) );
  OAI211_X1 U4975 ( .C1(n4493), .C2(n4520), .A(n4453), .B(n4452), .ZN(U3254)
         );
  AOI211_X1 U4976 ( .C1(n4455), .C2(n4454), .A(n2068), .B(n4482), .ZN(n4456)
         );
  AOI211_X1 U4977 ( .C1(n4486), .C2(ADDR_REG_15__SCAN_IN), .A(n4457), .B(n4456), .ZN(n4462) );
  OAI211_X1 U4978 ( .C1(n4460), .C2(n4459), .A(n4488), .B(n4458), .ZN(n4461)
         );
  OAI211_X1 U4979 ( .C1(n4493), .C2(n4519), .A(n4462), .B(n4461), .ZN(U3255)
         );
  AOI221_X1 U4980 ( .B1(n4464), .B2(n4463), .C1(n2525), .C2(n4463), .A(n4482), 
        .ZN(n4465) );
  AOI211_X1 U4981 ( .C1(n4486), .C2(ADDR_REG_16__SCAN_IN), .A(n4466), .B(n4465), .ZN(n4470) );
  OAI221_X1 U4982 ( .B1(n4468), .B2(REG1_REG_16__SCAN_IN), .C1(n4468), .C2(
        n4467), .A(n4488), .ZN(n4469) );
  OAI211_X1 U4983 ( .C1(n4493), .C2(n4518), .A(n4470), .B(n4469), .ZN(U3256)
         );
  AOI221_X1 U4984 ( .B1(n4473), .B2(n4472), .C1(n4471), .C2(n4472), .A(n4482), 
        .ZN(n4474) );
  AOI211_X1 U4985 ( .C1(n4486), .C2(ADDR_REG_17__SCAN_IN), .A(n4475), .B(n4474), .ZN(n4480) );
  OAI221_X1 U4986 ( .B1(n4478), .B2(n4477), .C1(n4478), .C2(n4476), .A(n4488), 
        .ZN(n4479) );
  OAI211_X1 U4987 ( .C1(n4493), .C2(n4517), .A(n4480), .B(n4479), .ZN(U3257)
         );
  INV_X1 U4988 ( .A(n4481), .ZN(n4485) );
  OAI211_X1 U4989 ( .C1(n4490), .C2(n4489), .A(n4488), .B(n4487), .ZN(n4491)
         );
  OAI211_X1 U4990 ( .C1(n4493), .C2(n4516), .A(n4492), .B(n4491), .ZN(U3258)
         );
  OAI22_X1 U4991 ( .A1(n4200), .A2(n4496), .B1(n4495), .B2(n4494), .ZN(n4497)
         );
  INV_X1 U4992 ( .A(n4497), .ZN(n4502) );
  INV_X1 U4993 ( .A(n4498), .ZN(n4500) );
  AOI22_X1 U4994 ( .A1(n4500), .A2(n4509), .B1(n4508), .B2(n4499), .ZN(n4501)
         );
  OAI211_X1 U4995 ( .C1(n4215), .C2(n4503), .A(n4502), .B(n4501), .ZN(U3282)
         );
  AOI22_X1 U4996 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4227), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4504), .ZN(n4512) );
  INV_X1 U4997 ( .A(n4505), .ZN(n4510) );
  INV_X1 U4998 ( .A(n4506), .ZN(n4507) );
  AOI22_X1 U4999 ( .A1(n4510), .A2(n4509), .B1(n4508), .B2(n4507), .ZN(n4511)
         );
  OAI211_X1 U5000 ( .C1(n4227), .C2(n4513), .A(n4512), .B(n4511), .ZN(U3288)
         );
  AND2_X1 U5001 ( .A1(D_REG_31__SCAN_IN), .A2(n4514), .ZN(U3291) );
  AND2_X1 U5002 ( .A1(D_REG_30__SCAN_IN), .A2(n4514), .ZN(U3292) );
  AND2_X1 U5003 ( .A1(D_REG_29__SCAN_IN), .A2(n4514), .ZN(U3293) );
  AND2_X1 U5004 ( .A1(D_REG_28__SCAN_IN), .A2(n4514), .ZN(U3294) );
  AND2_X1 U5005 ( .A1(D_REG_27__SCAN_IN), .A2(n4514), .ZN(U3295) );
  AND2_X1 U5006 ( .A1(D_REG_26__SCAN_IN), .A2(n4514), .ZN(U3296) );
  AND2_X1 U5007 ( .A1(D_REG_25__SCAN_IN), .A2(n4514), .ZN(U3297) );
  AND2_X1 U5008 ( .A1(D_REG_24__SCAN_IN), .A2(n4514), .ZN(U3298) );
  AND2_X1 U5009 ( .A1(D_REG_23__SCAN_IN), .A2(n4514), .ZN(U3299) );
  AND2_X1 U5010 ( .A1(D_REG_22__SCAN_IN), .A2(n4514), .ZN(U3300) );
  AND2_X1 U5011 ( .A1(D_REG_21__SCAN_IN), .A2(n4514), .ZN(U3301) );
  AND2_X1 U5012 ( .A1(D_REG_20__SCAN_IN), .A2(n4514), .ZN(U3302) );
  AND2_X1 U5013 ( .A1(D_REG_19__SCAN_IN), .A2(n4514), .ZN(U3303) );
  AND2_X1 U5014 ( .A1(D_REG_18__SCAN_IN), .A2(n4514), .ZN(U3304) );
  AND2_X1 U5015 ( .A1(D_REG_17__SCAN_IN), .A2(n4514), .ZN(U3305) );
  AND2_X1 U5016 ( .A1(D_REG_16__SCAN_IN), .A2(n4514), .ZN(U3306) );
  AND2_X1 U5017 ( .A1(D_REG_15__SCAN_IN), .A2(n4514), .ZN(U3307) );
  AND2_X1 U5018 ( .A1(D_REG_14__SCAN_IN), .A2(n4514), .ZN(U3308) );
  AND2_X1 U5019 ( .A1(D_REG_13__SCAN_IN), .A2(n4514), .ZN(U3309) );
  AND2_X1 U5020 ( .A1(D_REG_12__SCAN_IN), .A2(n4514), .ZN(U3310) );
  AND2_X1 U5021 ( .A1(D_REG_11__SCAN_IN), .A2(n4514), .ZN(U3311) );
  AND2_X1 U5022 ( .A1(D_REG_10__SCAN_IN), .A2(n4514), .ZN(U3312) );
  AND2_X1 U5023 ( .A1(D_REG_9__SCAN_IN), .A2(n4514), .ZN(U3313) );
  AND2_X1 U5024 ( .A1(D_REG_8__SCAN_IN), .A2(n4514), .ZN(U3314) );
  AND2_X1 U5025 ( .A1(D_REG_7__SCAN_IN), .A2(n4514), .ZN(U3315) );
  AND2_X1 U5026 ( .A1(D_REG_6__SCAN_IN), .A2(n4514), .ZN(U3316) );
  AND2_X1 U5027 ( .A1(D_REG_5__SCAN_IN), .A2(n4514), .ZN(U3317) );
  AND2_X1 U5028 ( .A1(D_REG_4__SCAN_IN), .A2(n4514), .ZN(U3318) );
  AND2_X1 U5029 ( .A1(D_REG_3__SCAN_IN), .A2(n4514), .ZN(U3319) );
  AND2_X1 U5030 ( .A1(D_REG_2__SCAN_IN), .A2(n4514), .ZN(U3320) );
  INV_X1 U5031 ( .A(DATAI_23_), .ZN(n4707) );
  AOI21_X1 U5032 ( .B1(U3149), .B2(n4707), .A(n4515), .ZN(U3329) );
  AOI22_X1 U5033 ( .A1(STATE_REG_SCAN_IN), .A2(n4516), .B1(n2554), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5034 ( .A1(STATE_REG_SCAN_IN), .A2(n4517), .B1(n4734), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5035 ( .A(DATAI_16_), .ZN(n4592) );
  AOI22_X1 U5036 ( .A1(STATE_REG_SCAN_IN), .A2(n4518), .B1(n4592), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5037 ( .A(DATAI_15_), .ZN(n4566) );
  AOI22_X1 U5038 ( .A1(STATE_REG_SCAN_IN), .A2(n4519), .B1(n4566), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5039 ( .A(DATAI_14_), .ZN(n4731) );
  AOI22_X1 U5040 ( .A1(STATE_REG_SCAN_IN), .A2(n4520), .B1(n4731), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5041 ( .A(DATAI_13_), .ZN(n4729) );
  AOI22_X1 U5042 ( .A1(STATE_REG_SCAN_IN), .A2(n4521), .B1(n4729), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5043 ( .A(DATAI_12_), .ZN(n4709) );
  AOI22_X1 U5044 ( .A1(STATE_REG_SCAN_IN), .A2(n4522), .B1(n4709), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5045 ( .A1(U3149), .A2(n4523), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4524) );
  INV_X1 U5046 ( .A(n4524), .ZN(U3341) );
  INV_X1 U5047 ( .A(DATAI_10_), .ZN(n4695) );
  AOI22_X1 U5048 ( .A1(STATE_REG_SCAN_IN), .A2(n4525), .B1(n4695), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5049 ( .A(DATAI_9_), .ZN(n4694) );
  AOI22_X1 U5050 ( .A1(STATE_REG_SCAN_IN), .A2(n4526), .B1(n4694), .B2(U3149), 
        .ZN(U3343) );
  OAI211_X1 U5051 ( .C1(n4529), .C2(n4532), .A(n4528), .B(n4527), .ZN(n4530)
         );
  INV_X1 U5052 ( .A(n4530), .ZN(n4556) );
  INV_X1 U5053 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4531) );
  AOI22_X1 U5054 ( .A1(n4554), .A2(n4556), .B1(n4531), .B2(n4552), .ZN(U3467)
         );
  NOR2_X1 U5055 ( .A1(n4533), .A2(n4532), .ZN(n4535) );
  AOI211_X1 U5056 ( .C1(n4537), .C2(n4536), .A(n4535), .B(n4534), .ZN(n4558)
         );
  INV_X1 U5057 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5058 ( .A1(n4554), .A2(n4558), .B1(n4538), .B2(n4552), .ZN(U3469)
         );
  INV_X1 U5059 ( .A(n4539), .ZN(n4544) );
  INV_X1 U5060 ( .A(n4540), .ZN(n4542) );
  AOI211_X1 U5061 ( .C1(n4544), .C2(n4543), .A(n4542), .B(n4541), .ZN(n4560)
         );
  INV_X1 U5062 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5063 ( .A1(n4554), .A2(n4560), .B1(n4545), .B2(n4552), .ZN(U3475)
         );
  NAND3_X1 U5064 ( .A1(n4548), .A2(n4547), .A3(n4546), .ZN(n4549) );
  AND3_X1 U5065 ( .A1(n4551), .A2(n4550), .A3(n4549), .ZN(n4563) );
  INV_X1 U5066 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4553) );
  AOI22_X1 U5067 ( .A1(n4554), .A2(n4563), .B1(n4553), .B2(n4552), .ZN(U3481)
         );
  AOI22_X1 U5068 ( .A1(n4564), .A2(n4556), .B1(n4555), .B2(n4561), .ZN(U3518)
         );
  INV_X1 U5069 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4557) );
  AOI22_X1 U5070 ( .A1(n4564), .A2(n4558), .B1(n4557), .B2(n4561), .ZN(U3519)
         );
  INV_X1 U5071 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4559) );
  AOI22_X1 U5072 ( .A1(n4564), .A2(n4560), .B1(n4559), .B2(n4561), .ZN(U3522)
         );
  AOI22_X1 U5073 ( .A1(n4564), .A2(n4563), .B1(n4562), .B2(n4561), .ZN(U3525)
         );
  AOI22_X1 U5074 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4755) );
  AOI22_X1 U5075 ( .A1(n4566), .A2(keyinput_g16), .B1(keyinput_g17), .B2(n4731), .ZN(n4565) );
  OAI221_X1 U5076 ( .B1(n4566), .B2(keyinput_g16), .C1(n4731), .C2(
        keyinput_g17), .A(n4565), .ZN(n4576) );
  AOI22_X1 U5077 ( .A1(n4695), .A2(keyinput_g21), .B1(keyinput_g1), .B2(n4568), 
        .ZN(n4567) );
  OAI221_X1 U5078 ( .B1(n4695), .B2(keyinput_g21), .C1(n4568), .C2(keyinput_g1), .A(n4567), .ZN(n4575) );
  INV_X1 U5079 ( .A(DATAI_6_), .ZN(n4570) );
  AOI22_X1 U5080 ( .A1(n4728), .A2(keyinput_g7), .B1(n4570), .B2(keyinput_g25), 
        .ZN(n4569) );
  OAI221_X1 U5081 ( .B1(n4728), .B2(keyinput_g7), .C1(n4570), .C2(keyinput_g25), .A(n4569), .ZN(n4574) );
  XOR2_X1 U5082 ( .A(n2317), .B(keyinput_g4), .Z(n4572) );
  XNOR2_X1 U5083 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_g42), .ZN(n4571) );
  NAND2_X1 U5084 ( .A1(n4572), .A2(n4571), .ZN(n4573) );
  NOR4_X1 U5085 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(n4614)
         );
  AOI22_X1 U5086 ( .A1(n4578), .A2(keyinput_g5), .B1(keyinput_g13), .B2(n2554), 
        .ZN(n4577) );
  OAI221_X1 U5087 ( .B1(n4578), .B2(keyinput_g5), .C1(n2554), .C2(keyinput_g13), .A(n4577), .ZN(n4587) );
  AOI22_X1 U5088 ( .A1(n4690), .A2(keyinput_g45), .B1(n4580), .B2(keyinput_g34), .ZN(n4579) );
  OAI221_X1 U5089 ( .B1(n4690), .B2(keyinput_g45), .C1(n4580), .C2(
        keyinput_g34), .A(n4579), .ZN(n4586) );
  XNOR2_X1 U5090 ( .A(DATAI_1_), .B(keyinput_g30), .ZN(n4584) );
  XNOR2_X1 U5091 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_g50), .ZN(n4583) );
  XNOR2_X1 U5092 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_g59), .ZN(n4582) );
  XNOR2_X1 U5093 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_g44), .ZN(n4581) );
  NAND4_X1 U5094 ( .A1(n4584), .A2(n4583), .A3(n4582), .A4(n4581), .ZN(n4585)
         );
  NOR3_X1 U5095 ( .A1(n4587), .A2(n4586), .A3(n4585), .ZN(n4613) );
  AOI22_X1 U5096 ( .A1(n4590), .A2(keyinput_g6), .B1(keyinput_g9), .B2(n4589), 
        .ZN(n4588) );
  OAI221_X1 U5097 ( .B1(n4590), .B2(keyinput_g6), .C1(n4589), .C2(keyinput_g9), 
        .A(n4588), .ZN(n4599) );
  INV_X1 U5098 ( .A(DATAI_21_), .ZN(n4719) );
  AOI22_X1 U5099 ( .A1(n4592), .A2(keyinput_g15), .B1(n4719), .B2(keyinput_g10), .ZN(n4591) );
  OAI221_X1 U5100 ( .B1(n4592), .B2(keyinput_g15), .C1(n4719), .C2(
        keyinput_g10), .A(n4591), .ZN(n4598) );
  XOR2_X1 U5101 ( .A(n2536), .B(keyinput_g48), .Z(n4596) );
  XNOR2_X1 U5102 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_g60), .ZN(n4595) );
  XNOR2_X1 U5103 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_g35), .ZN(n4594) );
  XNOR2_X1 U5104 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_g55), .ZN(n4593) );
  NAND4_X1 U5105 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(n4593), .ZN(n4597)
         );
  NOR3_X1 U5106 ( .A1(n4599), .A2(n4598), .A3(n4597), .ZN(n4612) );
  AOI22_X1 U5107 ( .A1(n2488), .A2(keyinput_g54), .B1(keyinput_g2), .B2(n4601), 
        .ZN(n4600) );
  OAI221_X1 U5108 ( .B1(n2488), .B2(keyinput_g54), .C1(n4601), .C2(keyinput_g2), .A(n4600), .ZN(n4610) );
  AOI22_X1 U5109 ( .A1(U3149), .A2(keyinput_g32), .B1(keyinput_g36), .B2(n4603), .ZN(n4602) );
  OAI221_X1 U5110 ( .B1(U3149), .B2(keyinput_g32), .C1(n4603), .C2(
        keyinput_g36), .A(n4602), .ZN(n4609) );
  XNOR2_X1 U5111 ( .A(DATAI_0_), .B(keyinput_g31), .ZN(n4607) );
  XNOR2_X1 U5112 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .ZN(n4606) );
  XNOR2_X1 U5113 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n4605) );
  XNOR2_X1 U5114 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_g57), .ZN(n4604) );
  NAND4_X1 U5115 ( .A1(n4607), .A2(n4606), .A3(n4605), .A4(n4604), .ZN(n4608)
         );
  NOR3_X1 U5116 ( .A1(n4610), .A2(n4609), .A3(n4608), .ZN(n4611) );
  NAND4_X1 U5117 ( .A1(n4614), .A2(n4613), .A3(n4612), .A4(n4611), .ZN(n4753)
         );
  AOI22_X1 U5118 ( .A1(DATAI_17_), .A2(keyinput_g14), .B1(DATAI_19_), .B2(
        keyinput_g12), .ZN(n4615) );
  OAI221_X1 U5119 ( .B1(DATAI_17_), .B2(keyinput_g14), .C1(DATAI_19_), .C2(
        keyinput_g12), .A(n4615), .ZN(n4622) );
  AOI22_X1 U5120 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(DATAI_28_), .B2(
        keyinput_g3), .ZN(n4616) );
  OAI221_X1 U5121 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(DATAI_28_), .C2(
        keyinput_g3), .A(n4616), .ZN(n4621) );
  AOI22_X1 U5122 ( .A1(DATAI_11_), .A2(keyinput_g20), .B1(DATAI_12_), .B2(
        keyinput_g19), .ZN(n4617) );
  OAI221_X1 U5123 ( .B1(DATAI_11_), .B2(keyinput_g20), .C1(DATAI_12_), .C2(
        keyinput_g19), .A(n4617), .ZN(n4620) );
  AOI22_X1 U5124 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput_g38), .B1(
        REG3_REG_7__SCAN_IN), .B2(keyinput_g33), .ZN(n4618) );
  OAI221_X1 U5125 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_g38), .C1(
        REG3_REG_7__SCAN_IN), .C2(keyinput_g33), .A(n4618), .ZN(n4619) );
  NOR4_X1 U5126 ( .A1(n4622), .A2(n4621), .A3(n4620), .A4(n4619), .ZN(n4652)
         );
  INV_X1 U5127 ( .A(DATAI_4_), .ZN(n4623) );
  XOR2_X1 U5128 ( .A(n4623), .B(keyinput_g27), .Z(n4630) );
  AOI22_X1 U5129 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput_g40), .B1(n2443), 
        .B2(keyinput_g23), .ZN(n4624) );
  OAI221_X1 U5130 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_g40), .C1(n2443), 
        .C2(keyinput_g23), .A(n4624), .ZN(n4629) );
  AOI22_X1 U5131 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_g53), .B1(
        REG3_REG_24__SCAN_IN), .B2(keyinput_g49), .ZN(n4625) );
  OAI221_X1 U5132 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_g53), .C1(
        REG3_REG_24__SCAN_IN), .C2(keyinput_g49), .A(n4625), .ZN(n4628) );
  AOI22_X1 U5133 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_g39), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput_g43), .ZN(n4626) );
  OAI221_X1 U5134 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_g39), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput_g43), .A(n4626), .ZN(n4627) );
  NOR4_X1 U5135 ( .A1(n4630), .A2(n4629), .A3(n4628), .A4(n4627), .ZN(n4651)
         );
  INV_X1 U5136 ( .A(DATAI_2_), .ZN(n4705) );
  AOI22_X1 U5137 ( .A1(n4707), .A2(keyinput_g8), .B1(keyinput_g29), .B2(n4705), 
        .ZN(n4631) );
  OAI221_X1 U5138 ( .B1(n4707), .B2(keyinput_g8), .C1(n4705), .C2(keyinput_g29), .A(n4631), .ZN(n4640) );
  AOI22_X1 U5139 ( .A1(n4704), .A2(keyinput_g0), .B1(n4633), .B2(keyinput_g26), 
        .ZN(n4632) );
  OAI221_X1 U5140 ( .B1(n4704), .B2(keyinput_g0), .C1(n4633), .C2(keyinput_g26), .A(n4632), .ZN(n4639) );
  AOI22_X1 U5141 ( .A1(DATAI_13_), .A2(keyinput_g18), .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .ZN(n4634) );
  OAI221_X1 U5142 ( .B1(DATAI_13_), .B2(keyinput_g18), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput_g46), .A(n4634), .ZN(n4638) );
  XNOR2_X1 U5143 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_g62), .ZN(n4636) );
  XNOR2_X1 U5144 ( .A(DATAI_3_), .B(keyinput_g28), .ZN(n4635) );
  NAND2_X1 U5145 ( .A1(n4636), .A2(n4635), .ZN(n4637) );
  NOR4_X1 U5146 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4650)
         );
  AOI22_X1 U5147 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_g47), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput_g58), .ZN(n4641) );
  OAI221_X1 U5148 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_g47), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput_g58), .A(n4641), .ZN(n4648) );
  AOI22_X1 U5149 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(IR_REG_1__SCAN_IN), 
        .B2(keyinput_g56), .ZN(n4642) );
  OAI221_X1 U5150 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(IR_REG_1__SCAN_IN), 
        .C2(keyinput_g56), .A(n4642), .ZN(n4647) );
  AOI22_X1 U5151 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(REG3_REG_8__SCAN_IN), 
        .B2(keyinput_g41), .ZN(n4643) );
  OAI221_X1 U5152 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(REG3_REG_8__SCAN_IN), 
        .C2(keyinput_g41), .A(n4643), .ZN(n4646) );
  AOI22_X1 U5153 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_g51), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .ZN(n4644) );
  OAI221_X1 U5154 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_g51), .C1(
        REG3_REG_10__SCAN_IN), .C2(keyinput_g37), .A(n4644), .ZN(n4645) );
  NOR4_X1 U5155 ( .A1(n4648), .A2(n4647), .A3(n4646), .A4(n4645), .ZN(n4649)
         );
  NAND4_X1 U5156 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4752)
         );
  AOI22_X1 U5157 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f38), .ZN(n4653) );
  OAI221_X1 U5158 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(REG3_REG_3__SCAN_IN), .C2(keyinput_f38), .A(n4653), .ZN(n4660) );
  AOI22_X1 U5159 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(DATAI_25_), .B2(
        keyinput_f6), .ZN(n4654) );
  OAI221_X1 U5160 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(DATAI_25_), .C2(
        keyinput_f6), .A(n4654), .ZN(n4659) );
  AOI22_X1 U5161 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_f33), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_f55), .ZN(n4655) );
  OAI221_X1 U5162 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_f33), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_f55), .A(n4655), .ZN(n4658) );
  AOI22_X1 U5163 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_f42), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .ZN(n4656) );
  OAI221_X1 U5164 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_f42), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_f44), .A(n4656), .ZN(n4657) );
  NOR4_X1 U5165 ( .A1(n4660), .A2(n4659), .A3(n4658), .A4(n4657), .ZN(n4688)
         );
  XOR2_X1 U5166 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_f53), .Z(n4667) );
  AOI22_X1 U5167 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(REG3_REG_19__SCAN_IN), 
        .B2(keyinput_f39), .ZN(n4661) );
  OAI221_X1 U5168 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(REG3_REG_19__SCAN_IN), .C2(keyinput_f39), .A(n4661), .ZN(n4666) );
  AOI22_X1 U5169 ( .A1(DATAI_26_), .A2(keyinput_f5), .B1(DATAI_27_), .B2(
        keyinput_f4), .ZN(n4662) );
  OAI221_X1 U5170 ( .B1(DATAI_26_), .B2(keyinput_f5), .C1(DATAI_27_), .C2(
        keyinput_f4), .A(n4662), .ZN(n4665) );
  AOI22_X1 U5171 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_f43), .B1(
        REG3_REG_24__SCAN_IN), .B2(keyinput_f49), .ZN(n4663) );
  OAI221_X1 U5172 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_f43), .C1(
        REG3_REG_24__SCAN_IN), .C2(keyinput_f49), .A(n4663), .ZN(n4664) );
  NOR4_X1 U5173 ( .A1(n4667), .A2(n4666), .A3(n4665), .A4(n4664), .ZN(n4687)
         );
  AOI22_X1 U5174 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(REG3_REG_27__SCAN_IN), 
        .B2(keyinput_f34), .ZN(n4668) );
  OAI221_X1 U5175 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(REG3_REG_27__SCAN_IN), .C2(keyinput_f34), .A(n4668), .ZN(n4676) );
  AOI22_X1 U5176 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_f37), .ZN(n4669) );
  OAI221_X1 U5177 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(
        REG3_REG_10__SCAN_IN), .C2(keyinput_f37), .A(n4669), .ZN(n4675) );
  AOI22_X1 U5178 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(REG3_REG_23__SCAN_IN), 
        .B2(keyinput_f36), .ZN(n4670) );
  OAI221_X1 U5179 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(REG3_REG_23__SCAN_IN), .C2(keyinput_f36), .A(n4670), .ZN(n4674) );
  XNOR2_X1 U5180 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_f60), .ZN(n4672) );
  XNOR2_X1 U5181 ( .A(DATAI_15_), .B(keyinput_f16), .ZN(n4671) );
  NAND2_X1 U5182 ( .A1(n4672), .A2(n4671), .ZN(n4673) );
  NOR4_X1 U5183 ( .A1(n4676), .A2(n4675), .A3(n4674), .A4(n4673), .ZN(n4686)
         );
  AOI22_X1 U5184 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(IR_REG_1__SCAN_IN), 
        .B2(keyinput_f56), .ZN(n4677) );
  OAI221_X1 U5185 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(IR_REG_1__SCAN_IN), 
        .C2(keyinput_f56), .A(n4677), .ZN(n4684) );
  AOI22_X1 U5186 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(IR_REG_7__SCAN_IN), 
        .B2(keyinput_f62), .ZN(n4678) );
  OAI221_X1 U5187 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(IR_REG_7__SCAN_IN), 
        .C2(keyinput_f62), .A(n4678), .ZN(n4683) );
  AOI22_X1 U5188 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(DATAI_8_), .B2(
        keyinput_f23), .ZN(n4679) );
  OAI221_X1 U5189 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(DATAI_8_), .C2(
        keyinput_f23), .A(n4679), .ZN(n4682) );
  AOI22_X1 U5190 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_f57), .B1(
        IR_REG_4__SCAN_IN), .B2(keyinput_f59), .ZN(n4680) );
  OAI221_X1 U5191 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_f57), .C1(
        IR_REG_4__SCAN_IN), .C2(keyinput_f59), .A(n4680), .ZN(n4681) );
  NOR4_X1 U5192 ( .A1(n4684), .A2(n4683), .A3(n4682), .A4(n4681), .ZN(n4685)
         );
  NAND4_X1 U5193 ( .A1(n4688), .A2(n4687), .A3(n4686), .A4(n4685), .ZN(n4746)
         );
  INV_X1 U5194 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4691) );
  AOI22_X1 U5195 ( .A1(n4691), .A2(keyinput_f46), .B1(n4690), .B2(keyinput_f45), .ZN(n4689) );
  OAI221_X1 U5196 ( .B1(n4691), .B2(keyinput_f46), .C1(n4690), .C2(
        keyinput_f45), .A(n4689), .ZN(n4702) );
  AOI22_X1 U5197 ( .A1(n4694), .A2(keyinput_f22), .B1(n4693), .B2(keyinput_f35), .ZN(n4692) );
  OAI221_X1 U5198 ( .B1(n4694), .B2(keyinput_f22), .C1(n4693), .C2(
        keyinput_f35), .A(n4692), .ZN(n4701) );
  XOR2_X1 U5199 ( .A(n4695), .B(keyinput_f21), .Z(n4699) );
  XNOR2_X1 U5200 ( .A(DATAI_3_), .B(keyinput_f28), .ZN(n4698) );
  XNOR2_X1 U5201 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_f41), .ZN(n4697) );
  XNOR2_X1 U5202 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n4696) );
  NAND4_X1 U5203 ( .A1(n4699), .A2(n4698), .A3(n4697), .A4(n4696), .ZN(n4700)
         );
  NOR3_X1 U5204 ( .A1(n4702), .A2(n4701), .A3(n4700), .ZN(n4744) );
  AOI22_X1 U5205 ( .A1(n4705), .A2(keyinput_f29), .B1(keyinput_f0), .B2(n4704), 
        .ZN(n4703) );
  OAI221_X1 U5206 ( .B1(n4705), .B2(keyinput_f29), .C1(n4704), .C2(keyinput_f0), .A(n4703), .ZN(n4714) );
  AOI22_X1 U5207 ( .A1(n2536), .A2(keyinput_f48), .B1(keyinput_f8), .B2(n4707), 
        .ZN(n4706) );
  OAI221_X1 U5208 ( .B1(n2536), .B2(keyinput_f48), .C1(n4707), .C2(keyinput_f8), .A(n4706), .ZN(n4713) );
  AOI22_X1 U5209 ( .A1(n2488), .A2(keyinput_f54), .B1(keyinput_f19), .B2(n4709), .ZN(n4708) );
  OAI221_X1 U5210 ( .B1(n2488), .B2(keyinput_f54), .C1(n4709), .C2(
        keyinput_f19), .A(n4708), .ZN(n4712) );
  AOI22_X1 U5211 ( .A1(n2446), .A2(keyinput_f51), .B1(n3559), .B2(keyinput_f40), .ZN(n4710) );
  OAI221_X1 U5212 ( .B1(n2446), .B2(keyinput_f51), .C1(n3559), .C2(
        keyinput_f40), .A(n4710), .ZN(n4711) );
  NOR4_X1 U5213 ( .A1(n4714), .A2(n4713), .A3(n4712), .A4(n4711), .ZN(n4743)
         );
  AOI22_X1 U5214 ( .A1(n4717), .A2(keyinput_f3), .B1(keyinput_f11), .B2(n4716), 
        .ZN(n4715) );
  OAI221_X1 U5215 ( .B1(n4717), .B2(keyinput_f3), .C1(n4716), .C2(keyinput_f11), .A(n4715), .ZN(n4726) );
  AOI22_X1 U5216 ( .A1(n2089), .A2(keyinput_f47), .B1(keyinput_f10), .B2(n4719), .ZN(n4718) );
  OAI221_X1 U5217 ( .B1(n2089), .B2(keyinput_f47), .C1(n4719), .C2(
        keyinput_f10), .A(n4718), .ZN(n4725) );
  XNOR2_X1 U5218 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_f52), .ZN(n4723) );
  XNOR2_X1 U5219 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n4722) );
  XNOR2_X1 U5220 ( .A(DATAI_0_), .B(keyinput_f31), .ZN(n4721) );
  XNOR2_X1 U5221 ( .A(DATAI_7_), .B(keyinput_f24), .ZN(n4720) );
  NAND4_X1 U5222 ( .A1(n4723), .A2(n4722), .A3(n4721), .A4(n4720), .ZN(n4724)
         );
  NOR3_X1 U5223 ( .A1(n4726), .A2(n4725), .A3(n4724), .ZN(n4742) );
  AOI22_X1 U5224 ( .A1(n4729), .A2(keyinput_f18), .B1(keyinput_f7), .B2(n4728), 
        .ZN(n4727) );
  OAI221_X1 U5225 ( .B1(n4729), .B2(keyinput_f18), .C1(n4728), .C2(keyinput_f7), .A(n4727), .ZN(n4740) );
  INV_X1 U5226 ( .A(DATAI_19_), .ZN(n4732) );
  AOI22_X1 U5227 ( .A1(n4732), .A2(keyinput_f12), .B1(keyinput_f17), .B2(n4731), .ZN(n4730) );
  OAI221_X1 U5228 ( .B1(n4732), .B2(keyinput_f12), .C1(n4731), .C2(
        keyinput_f17), .A(n4730), .ZN(n4739) );
  AOI22_X1 U5229 ( .A1(n4734), .A2(keyinput_f14), .B1(U3149), .B2(keyinput_f32), .ZN(n4733) );
  OAI221_X1 U5230 ( .B1(n4734), .B2(keyinput_f14), .C1(U3149), .C2(
        keyinput_f32), .A(n4733), .ZN(n4738) );
  XNOR2_X1 U5231 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_f58), .ZN(n4736) );
  XNOR2_X1 U5232 ( .A(keyinput_f25), .B(DATAI_6_), .ZN(n4735) );
  NAND2_X1 U5233 ( .A1(n4736), .A2(n4735), .ZN(n4737) );
  NOR4_X1 U5234 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n4741)
         );
  NAND4_X1 U5235 ( .A1(n4744), .A2(n4743), .A3(n4742), .A4(n4741), .ZN(n4745)
         );
  OAI22_X1 U5236 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput_f63), .B1(n4746), .B2(
        n4745), .ZN(n4748) );
  INV_X1 U5237 ( .A(keyinput_g63), .ZN(n4747) );
  NAND2_X1 U5238 ( .A1(n4748), .A2(n4747), .ZN(n4750) );
  OAI211_X1 U5239 ( .C1(n4748), .C2(keyinput_f63), .A(IR_REG_8__SCAN_IN), .B(
        keyinput_g63), .ZN(n4749) );
  OAI21_X1 U5240 ( .B1(IR_REG_8__SCAN_IN), .B2(n4750), .A(n4749), .ZN(n4751)
         );
  OAI21_X1 U5241 ( .B1(n4753), .B2(n4752), .A(n4751), .ZN(n4754) );
  XOR2_X1 U5242 ( .A(n4755), .B(n4754), .Z(U3352) );
  BUF_X2 U2310 ( .A(n3542), .Z(n2047) );
  BUF_X1 U2318 ( .A(n3023), .Z(n3547) );
  OR2_X1 U2865 ( .A1(n2944), .A2(n2072), .ZN(n2172) );
  CLKBUF_X1 U2297 ( .A(n2951), .Z(n2048) );
  AOI21_X1 U2313 ( .B1(n4383), .B2(n2808), .A(n2807), .ZN(n2905) );
endmodule

