

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2957, n2958, n2959, n2960, n2961, n2963, n2964, n2969, n2970, n2971,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782;

  AOI21_X1 U3405 ( .B1(n5697), .B2(n5516), .A(n5505), .ZN(n5741) );
  INV_X1 U3406 ( .A(n6254), .ZN(n6266) );
  INV_X1 U3407 ( .A(n5655), .ZN(n2989) );
  INV_X2 U3408 ( .A(n5655), .ZN(n5674) );
  NAND2_X2 U3410 ( .A1(n4560), .A2(n4546), .ZN(n6277) );
  XNOR2_X1 U3411 ( .A(n4008), .B(n4630), .ZN(n4461) );
  NAND2_X2 U3412 ( .A1(n4685), .A2(n4537), .ZN(n4005) );
  CLKBUF_X3 U3413 ( .A(n4164), .Z(n2959) );
  NAND2_X1 U3414 ( .A1(n3397), .A2(n3396), .ZN(n4726) );
  CLKBUF_X2 U3415 ( .A(n3470), .Z(n2971) );
  CLKBUF_X2 U3416 ( .A(n3400), .Z(n2979) );
  CLKBUF_X2 U3417 ( .A(n3373), .Z(n2984) );
  INV_X2 U3418 ( .A(n3810), .ZN(n2961) );
  CLKBUF_X2 U3419 ( .A(n3372), .Z(n2973) );
  BUF_X1 U3420 ( .A(n3402), .Z(n2969) );
  AND2_X2 U3421 ( .A1(n2981), .A2(n4707), .ZN(n2983) );
  AND2_X2 U3422 ( .A1(n3227), .A2(n4711), .ZN(n3416) );
  AND2_X2 U3423 ( .A1(n4436), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3225)
         );
  INV_X1 U3425 ( .A(n3374), .ZN(n3848) );
  AND2_X1 U3426 ( .A1(n4003), .A2(n4021), .ZN(n3158) );
  NAND2_X1 U3427 ( .A1(n4164), .A2(n4002), .ZN(n4021) );
  AND2_X1 U3429 ( .A1(n5322), .A2(n5308), .ZN(n5442) );
  NOR2_X1 U3430 ( .A1(n3160), .A2(n5104), .ZN(n3159) );
  XNOR2_X1 U3431 ( .A(n4726), .B(n4727), .ZN(n4653) );
  NAND2_X1 U3432 ( .A1(n5371), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4343) );
  INV_X1 U3433 ( .A(n3340), .ZN(n3345) );
  NAND2_X1 U3434 ( .A1(n5598), .A2(n4323), .ZN(n3197) );
  NAND2_X1 U3435 ( .A1(n4624), .A2(n3159), .ZN(n5107) );
  INV_X1 U3436 ( .A(n6155), .ZN(n6174) );
  AND2_X2 U3437 ( .A1(n3219), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5147)
         );
  INV_X1 U3438 ( .A(n6152), .ZN(n6095) );
  INV_X1 U3439 ( .A(n3003), .ZN(n4164) );
  OAI21_X2 U3443 ( .B1(n4195), .B2(n5181), .A(n4192), .ZN(n4163) );
  NAND3_X2 U3444 ( .A1(n3992), .A2(n3370), .A3(n3369), .ZN(n3387) );
  AND2_X2 U34460 ( .A1(n3227), .A2(n4711), .ZN(n2957) );
  NAND2_X2 U34470 ( .A1(n3272), .A2(n3271), .ZN(n3359) );
  AND2_X2 U34480 ( .A1(n3367), .A2(n3366), .ZN(n3370) );
  INV_X1 U3449 ( .A(n2976), .ZN(n2958) );
  AOI21_X2 U34510 ( .B1(n3074), .B2(n5680), .A(n3026), .ZN(n3073) );
  XNOR2_X2 U34520 ( .A(n4308), .B(n4307), .ZN(n5680) );
  AOI21_X2 U34530 ( .B1(n4739), .B2(n3177), .A(n3020), .ZN(n3176) );
  BUF_X4 U3454 ( .A(n4164), .Z(n2960) );
  INV_X1 U34560 ( .A(n3810), .ZN(n3049) );
  NOR2_X2 U3457 ( .A1(n6098), .A2(n4172), .ZN(n6093) );
  AND2_X1 U34590 ( .A1(n2980), .A2(n4707), .ZN(n2964) );
  AND2_X1 U34610 ( .A1(n2980), .A2(n4707), .ZN(n3402) );
  OR2_X1 U34620 ( .A1(n5598), .A2(n3151), .ZN(n3147) );
  CLKBUF_X1 U34630 ( .A(n5237), .Z(n5238) );
  NOR2_X1 U34640 ( .A1(n5747), .A2(n3103), .ZN(n5727) );
  OR2_X1 U34650 ( .A1(n5787), .A2(n5708), .ZN(n5763) );
  AND2_X1 U3466 ( .A1(n4281), .A2(n4280), .ZN(n4302) );
  OAI21_X1 U3467 ( .B1(n4239), .B2(n3675), .A(n3508), .ZN(n4621) );
  AND2_X1 U34680 ( .A1(n4246), .A2(n4247), .ZN(n5920) );
  INV_X1 U34690 ( .A(n4246), .ZN(n3132) );
  NAND2_X1 U34700 ( .A1(n3141), .A2(n3079), .ZN(n4246) );
  OR2_X1 U34710 ( .A1(n3141), .A2(n3079), .ZN(n4247) );
  OR2_X1 U34720 ( .A1(n4476), .A2(n4477), .ZN(n4478) );
  AND2_X1 U34730 ( .A1(n3187), .A2(n3186), .ZN(n3388) );
  CLKBUF_X1 U34740 ( .A(n4138), .Z(n4419) );
  CLKBUF_X2 U3475 ( .A(n3339), .Z(n4223) );
  INV_X1 U3476 ( .A(n3981), .ZN(n4001) );
  NAND2_X1 U3477 ( .A1(n3330), .A2(n4250), .ZN(n3358) );
  NAND2_X1 U3478 ( .A1(n4250), .A2(n3332), .ZN(n3981) );
  AND4_X1 U3480 ( .A1(n3290), .A2(n3289), .A3(n3288), .A4(n3287), .ZN(n3297)
         );
  AND4_X1 U3481 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3260)
         );
  CLKBUF_X2 U3482 ( .A(n3298), .Z(n4119) );
  CLKBUF_X2 U3483 ( .A(n3465), .Z(n3489) );
  BUF_X1 U3484 ( .A(n3509), .Z(n2977) );
  CLKBUF_X2 U3485 ( .A(n3421), .Z(n4120) );
  CLKBUF_X2 U3486 ( .A(n3313), .Z(n3537) );
  AND2_X1 U3487 ( .A1(n3936), .A2(n3935), .ZN(n5506) );
  OR2_X1 U3488 ( .A1(n5532), .A2(n5523), .ZN(n5515) );
  OAI21_X1 U3489 ( .B1(n5197), .B2(n5198), .A(n3933), .ZN(n5521) );
  OAI21_X1 U3490 ( .B1(n4112), .B2(n5179), .A(n5178), .ZN(n5499) );
  XNOR2_X1 U3491 ( .A(n4137), .B(n4136), .ZN(n4232) );
  OR2_X1 U3492 ( .A1(n5624), .A2(n5620), .ZN(n5610) );
  AND2_X1 U3493 ( .A1(n5197), .A2(n3042), .ZN(n4137) );
  NOR2_X2 U3494 ( .A1(n5237), .A2(n3044), .ZN(n5197) );
  OR2_X1 U3495 ( .A1(n3155), .A2(n3008), .ZN(n3153) );
  OAI21_X1 U3496 ( .B1(n5597), .B2(n3157), .A(n5544), .ZN(n3156) );
  AOI21_X1 U3497 ( .B1(n3185), .B2(n4318), .A(n3023), .ZN(n3184) );
  AND2_X1 U3498 ( .A1(n2993), .A2(n3012), .ZN(n2994) );
  NAND2_X1 U3499 ( .A1(n4292), .A2(n4291), .ZN(n5131) );
  OR2_X1 U3500 ( .A1(n3216), .A2(n3029), .ZN(n3185) );
  AND2_X1 U3501 ( .A1(n4208), .A2(n4179), .ZN(n5186) );
  NOR2_X1 U3502 ( .A1(n5224), .A2(n4184), .ZN(n5208) );
  OR2_X1 U3503 ( .A1(n4309), .A2(n6297), .ZN(n5663) );
  OR2_X1 U3504 ( .A1(n4295), .A2(n4294), .ZN(n4298) );
  NAND2_X2 U3505 ( .A1(n4302), .A2(n4304), .ZN(n4309) );
  NOR3_X1 U3506 ( .A1(n6084), .A2(n5572), .A3(n3056), .ZN(n5255) );
  OR2_X1 U3507 ( .A1(n5287), .A2(n4175), .ZN(n5254) );
  NAND2_X1 U3508 ( .A1(n5293), .A2(n4183), .ZN(n6084) );
  XNOR2_X1 U3509 ( .A(n4281), .B(n3566), .ZN(n4293) );
  NOR2_X1 U3510 ( .A1(n5307), .A2(n5306), .ZN(n5293) );
  NOR2_X2 U3511 ( .A1(n5355), .A2(n5354), .ZN(n5339) );
  OR2_X2 U3512 ( .A1(n3062), .A2(n3061), .ZN(n5355) );
  NAND2_X1 U3513 ( .A1(n3091), .A2(n5905), .ZN(n5913) );
  NAND2_X1 U3514 ( .A1(n6277), .A2(n4572), .ZN(n3091) );
  NOR2_X1 U3516 ( .A1(n4697), .A2(n4679), .ZN(n6498) );
  NOR2_X1 U3517 ( .A1(n4697), .A2(n4672), .ZN(n6530) );
  NOR2_X1 U3518 ( .A1(n4697), .A2(n3343), .ZN(n6516) );
  NOR2_X1 U3519 ( .A1(n4697), .A2(n4691), .ZN(n6492) );
  NOR2_X1 U3520 ( .A1(n4697), .A2(n3362), .ZN(n6522) );
  NOR2_X1 U3521 ( .A1(n4697), .A2(n4554), .ZN(n6510) );
  INV_X1 U3522 ( .A(n4343), .ZN(n4332) );
  INV_X2 U3523 ( .A(n6193), .ZN(n2970) );
  NAND2_X1 U3524 ( .A1(n4553), .A2(n4552), .ZN(n4586) );
  NAND2_X1 U3525 ( .A1(n4542), .A2(n4541), .ZN(n4560) );
  OR2_X1 U3526 ( .A1(n4566), .A2(n4540), .ZN(n4541) );
  OR2_X1 U3527 ( .A1(n4662), .A2(n4294), .ZN(n4257) );
  AOI21_X1 U3528 ( .B1(n3007), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3395), 
        .ZN(n3398) );
  NOR2_X1 U3529 ( .A1(n4014), .A2(n3162), .ZN(n3161) );
  OAI21_X1 U3530 ( .B1(n3954), .B2(n3099), .A(n2998), .ZN(n3100) );
  NAND2_X1 U3531 ( .A1(n3323), .A2(n4406), .ZN(n3357) );
  MUX2_X1 U3532 ( .A(n4085), .B(n4005), .S(EBX_REG_1__SCAN_IN), .Z(n4004) );
  AND2_X1 U3533 ( .A1(n3335), .A2(n3354), .ZN(n3188) );
  NAND2_X1 U3534 ( .A1(n4005), .A2(n3981), .ZN(n4629) );
  AND2_X1 U3535 ( .A1(n4261), .A2(n3343), .ZN(n3344) );
  OR2_X1 U3536 ( .A1(n3339), .A2(n2974), .ZN(n4440) );
  NOR2_X1 U3537 ( .A1(n3328), .A2(n4544), .ZN(n3986) );
  CLKBUF_X1 U3538 ( .A(n3330), .Z(n3987) );
  NAND2_X1 U3539 ( .A1(n4554), .A2(n3324), .ZN(n3339) );
  BUF_X2 U3540 ( .A(n3325), .Z(n4691) );
  INV_X1 U3541 ( .A(n3361), .ZN(n3347) );
  CLKBUF_X2 U3542 ( .A(n3360), .Z(n4544) );
  NAND3_X1 U3543 ( .A1(n3297), .A2(n3296), .A3(n3295), .ZN(n3340) );
  NAND2_X2 U3544 ( .A1(n3260), .A2(n3218), .ZN(n3360) );
  AND4_X1 U3545 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3250)
         );
  AND4_X1 U3546 ( .A1(n3231), .A2(n3230), .A3(n3229), .A4(n3228), .ZN(n3232)
         );
  AND4_X1 U3547 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3271)
         );
  AND4_X1 U3548 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(n3233)
         );
  CLKBUF_X1 U3549 ( .A(n3291), .Z(n4121) );
  AND4_X1 U3550 ( .A1(n3311), .A2(n3310), .A3(n3309), .A4(n3308), .ZN(n3320)
         );
  AND4_X1 U3551 ( .A1(n3234), .A2(n3240), .A3(n3237), .A4(n3235), .ZN(n3140)
         );
  AND4_X1 U3552 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3218)
         );
  AND4_X1 U3553 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n3321)
         );
  AND3_X1 U3554 ( .A1(n3294), .A2(n3293), .A3(n3292), .ZN(n3295) );
  AND4_X1 U3555 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3251)
         );
  AND4_X1 U3556 ( .A1(n3266), .A2(n3265), .A3(n3264), .A4(n3263), .ZN(n3272)
         );
  AND4_X1 U3557 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3319)
         );
  AND4_X1 U3558 ( .A1(n3302), .A2(n3301), .A3(n3300), .A4(n3299), .ZN(n3322)
         );
  AND4_X1 U3559 ( .A1(n3236), .A2(n3241), .A3(n3239), .A4(n3238), .ZN(n3139)
         );
  AND2_X2 U3560 ( .A1(n3220), .A2(n4415), .ZN(n3407) );
  INV_X2 U3561 ( .A(n6021), .ZN(n4375) );
  AND2_X2 U3563 ( .A1(n4707), .A2(n4415), .ZN(n3314) );
  AND2_X2 U3565 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4415) );
  AND2_X2 U3566 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4707) );
  NOR2_X2 U3567 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4706) );
  NOR2_X4 U3568 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4723) );
  BUF_X2 U3569 ( .A(n4723), .Z(n2980) );
  AND2_X1 U3570 ( .A1(n4785), .A2(n3500), .ZN(n3131) );
  NAND2_X1 U3571 ( .A1(n3132), .A2(n4785), .ZN(n3502) );
  INV_X2 U3572 ( .A(n3360), .ZN(n4554) );
  NAND2_X1 U3573 ( .A1(n3433), .A2(n6566), .ZN(n3431) );
  INV_X1 U3574 ( .A(n3387), .ZN(n3386) );
  AND2_X1 U3576 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4711) );
  AND4_X2 U3577 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3325)
         );
  NAND2_X1 U3578 ( .A1(n4250), .A2(n3332), .ZN(n2974) );
  NAND2_X1 U3579 ( .A1(n4250), .A2(n3332), .ZN(n2975) );
  AND2_X2 U3580 ( .A1(n5147), .A2(n3220), .ZN(n2976) );
  AND2_X2 U3581 ( .A1(n4586), .A2(n4267), .ZN(n4570) );
  BUF_X8 U3582 ( .A(n3509), .Z(n2978) );
  AND2_X2 U3583 ( .A1(n3226), .A2(n4707), .ZN(n3509) );
  AND2_X2 U3584 ( .A1(n3226), .A2(n4706), .ZN(n3400) );
  AND2_X2 U3585 ( .A1(n2980), .A2(n4706), .ZN(n3373) );
  INV_X4 U3586 ( .A(n3325), .ZN(n3332) );
  NOR2_X2 U3587 ( .A1(n3286), .A2(n3285), .ZN(n3342) );
  XNOR2_X2 U3588 ( .A(n5911), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4553)
         );
  AND2_X1 U3589 ( .A1(n2980), .A2(n4707), .ZN(n2982) );
  NAND2_X4 U3590 ( .A1(n3251), .A2(n3250), .ZN(n3324) );
  INV_X1 U3591 ( .A(n5655), .ZN(n2988) );
  AND2_X2 U3592 ( .A1(n3225), .A2(n4415), .ZN(n3421) );
  NOR2_X1 U3593 ( .A1(n3170), .A2(n5421), .ZN(n3169) );
  INV_X1 U3594 ( .A(n3217), .ZN(n3170) );
  INV_X1 U3595 ( .A(n3501), .ZN(n3500) );
  OR2_X1 U3596 ( .A1(n3385), .A2(n3384), .ZN(n4259) );
  OR2_X1 U3597 ( .A1(n3413), .A2(n3412), .ZN(n4233) );
  OAI21_X1 U3598 ( .B1(n3347), .B2(n3360), .A(n3359), .ZN(n3273) );
  AND2_X2 U3599 ( .A1(n5147), .A2(n4707), .ZN(n3465) );
  NOR2_X1 U3600 ( .A1(n3203), .A2(n3034), .ZN(n3202) );
  INV_X1 U3601 ( .A(n5245), .ZN(n3203) );
  NAND2_X1 U3602 ( .A1(n3130), .A2(n3128), .ZN(n3127) );
  INV_X1 U3603 ( .A(n5738), .ZN(n3128) );
  INV_X1 U3604 ( .A(n5543), .ZN(n3157) );
  NAND2_X1 U3605 ( .A1(n3150), .A2(n5580), .ZN(n3149) );
  INV_X1 U3606 ( .A(n3153), .ZN(n3150) );
  AND3_X1 U3607 ( .A1(n3343), .A2(n4679), .A3(n4685), .ZN(n4438) );
  NAND2_X1 U3608 ( .A1(n5142), .A2(n3345), .ZN(n4217) );
  INV_X1 U3609 ( .A(n3346), .ZN(n4406) );
  INV_X1 U3610 ( .A(n5371), .ZN(n6135) );
  NAND2_X1 U3611 ( .A1(n3050), .A2(n3021), .ZN(n4528) );
  NAND2_X1 U3612 ( .A1(n3051), .A2(n3017), .ZN(n3050) );
  OR2_X2 U3613 ( .A1(n4528), .A2(n6573), .ZN(n4566) );
  INV_X1 U3614 ( .A(n4326), .ZN(n3196) );
  AND2_X1 U3615 ( .A1(n5707), .A2(n5708), .ZN(n3104) );
  AND2_X1 U3616 ( .A1(n3168), .A2(n3167), .ZN(n3166) );
  INV_X1 U3617 ( .A(n5270), .ZN(n3167) );
  INV_X1 U3618 ( .A(n5347), .ZN(n4041) );
  NAND2_X1 U3619 ( .A1(n5915), .A2(n4662), .ZN(n5967) );
  AND2_X1 U3620 ( .A1(n4230), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4205) );
  AOI21_X1 U3621 ( .B1(n4223), .B2(n3945), .A(n3345), .ZN(n3938) );
  OAI21_X1 U3622 ( .B1(n3361), .B2(n3324), .A(n3359), .ZN(n3328) );
  INV_X1 U3623 ( .A(n3349), .ZN(n3124) );
  NAND2_X1 U3624 ( .A1(n3100), .A2(n2990), .ZN(n3054) );
  NAND2_X1 U3625 ( .A1(n3963), .A2(n3102), .ZN(n3101) );
  NAND2_X1 U3626 ( .A1(n3970), .A2(n4280), .ZN(n3976) );
  OR2_X1 U3627 ( .A1(n3499), .A2(n3498), .ZN(n4236) );
  NAND2_X1 U3628 ( .A1(n3345), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3441) );
  OAI21_X1 U3629 ( .B1(n3433), .B2(n3066), .A(n6566), .ZN(n3065) );
  INV_X1 U3630 ( .A(n3447), .ZN(n3068) );
  OR2_X1 U3631 ( .A1(n3476), .A2(n3475), .ZN(n4241) );
  NAND2_X1 U3632 ( .A1(n3361), .A2(n3324), .ZN(n3330) );
  AOI22_X1 U3633 ( .A1(n3470), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U3634 ( .A1(n3372), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3049), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3231) );
  MUX2_X1 U3635 ( .A(n3994), .B(n4225), .S(n6309), .Z(n3354) );
  NOR2_X1 U3636 ( .A1(n4443), .A2(n3993), .ZN(n4547) );
  NAND2_X2 U3637 ( .A1(n3441), .A2(n3055), .ZN(n3979) );
  NAND2_X1 U3638 ( .A1(n3502), .A2(n3501), .ZN(n3144) );
  NAND2_X1 U3639 ( .A1(n3724), .A2(n3045), .ZN(n3762) );
  NOR2_X1 U3640 ( .A1(n3207), .A2(n3082), .ZN(n3081) );
  INV_X1 U3641 ( .A(n5427), .ZN(n3082) );
  NOR2_X1 U3642 ( .A1(n3725), .A2(n5625), .ZN(n3107) );
  INV_X1 U3643 ( .A(n4132), .ZN(n4106) );
  NOR2_X1 U3644 ( .A1(n5142), .A2(n6566), .ZN(n4132) );
  NOR2_X1 U3645 ( .A1(n5291), .A2(n5439), .ZN(n3208) );
  NAND2_X1 U3646 ( .A1(n3086), .A2(n5332), .ZN(n3085) );
  INV_X1 U3647 ( .A(n3087), .ZN(n3086) );
  NAND2_X1 U3648 ( .A1(n5121), .A2(n3200), .ZN(n3199) );
  INV_X1 U3649 ( .A(n5123), .ZN(n3200) );
  OR2_X1 U3650 ( .A1(n5164), .A2(n5978), .ZN(n3032) );
  NOR2_X2 U3651 ( .A1(n3996), .A2(n5978), .ZN(n3685) );
  AND2_X1 U3652 ( .A1(n3195), .A2(n4321), .ZN(n3075) );
  INV_X1 U3653 ( .A(n4323), .ZN(n3194) );
  AND2_X1 U3654 ( .A1(n2994), .A2(n3146), .ZN(n4315) );
  INV_X1 U3655 ( .A(n4627), .ZN(n3162) );
  NAND2_X1 U3656 ( .A1(n3182), .A2(n4252), .ZN(n4268) );
  NAND2_X1 U3657 ( .A1(n5920), .A2(n4280), .ZN(n3182) );
  NOR2_X1 U3658 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n4916), .ZN(n5972)
         );
  AOI21_X1 U3659 ( .B1(n3298), .B2(INSTQUEUE_REG_1__4__SCAN_IN), .A(n3019), 
        .ZN(n3253) );
  INV_X1 U3660 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4916) );
  INV_X1 U3661 ( .A(n6394), .ZN(n4869) );
  OAI21_X1 U3662 ( .B1(n6615), .B2(n4651), .A(n6567), .ZN(n4656) );
  CLKBUF_X1 U3663 ( .A(n3480), .Z(n3481) );
  NAND2_X1 U3664 ( .A1(n5978), .A2(n6059), .ZN(n3819) );
  INV_X1 U3665 ( .A(n4213), .ZN(n4543) );
  NAND2_X1 U3666 ( .A1(n4332), .A2(n4169), .ZN(n6159) );
  NAND2_X1 U3667 ( .A1(n3389), .A2(n3391), .ZN(n3440) );
  OR2_X2 U3668 ( .A1(n3063), .A2(n2997), .ZN(n5371) );
  INV_X1 U3669 ( .A(n3706), .ZN(n4135) );
  OR2_X1 U3670 ( .A1(n3843), .A2(n5246), .ZN(n3878) );
  NAND2_X1 U3671 ( .A1(n3794), .A2(n3105), .ZN(n3798) );
  INV_X1 U3672 ( .A(n3762), .ZN(n3794) );
  AND2_X1 U3673 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n3705), .ZN(n3724)
         );
  INV_X1 U3674 ( .A(n3704), .ZN(n3705) );
  NOR2_X1 U3675 ( .A1(n3604), .A2(n3111), .ZN(n3110) );
  AND2_X1 U3676 ( .A1(n3588), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3603)
         );
  NOR2_X1 U3677 ( .A1(n3567), .A2(n6263), .ZN(n3588) );
  NOR2_X1 U3678 ( .A1(n3522), .A2(n6272), .ZN(n3544) );
  NAND2_X1 U3679 ( .A1(n3544), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3567)
         );
  NAND2_X1 U3680 ( .A1(n4478), .A2(n3439), .ZN(n4335) );
  NAND2_X1 U3681 ( .A1(n4477), .A2(n3438), .ZN(n3439) );
  NOR2_X1 U3682 ( .A1(n3127), .A2(n3048), .ZN(n3126) );
  NOR2_X1 U3683 ( .A1(n3174), .A2(n3172), .ZN(n3171) );
  OR2_X1 U3684 ( .A1(n4161), .A2(n3173), .ZN(n3172) );
  INV_X1 U3685 ( .A(n5213), .ZN(n3173) );
  INV_X1 U3686 ( .A(n3127), .ZN(n3125) );
  NAND2_X1 U3687 ( .A1(n3197), .A2(n3195), .ZN(n5532) );
  OR2_X1 U3688 ( .A1(n3008), .A2(n3157), .ZN(n3154) );
  INV_X1 U3689 ( .A(n3156), .ZN(n3155) );
  NAND2_X1 U3690 ( .A1(n2995), .A2(n5362), .ZN(n3163) );
  NAND2_X1 U3691 ( .A1(n5609), .A2(n6297), .ZN(n3138) );
  NAND2_X1 U3692 ( .A1(n5609), .A2(n6307), .ZN(n4310) );
  INV_X1 U3693 ( .A(n4301), .ZN(n3074) );
  NAND2_X1 U3694 ( .A1(n3072), .A2(n5680), .ZN(n3071) );
  INV_X1 U3695 ( .A(n3142), .ZN(n3072) );
  INV_X1 U3696 ( .A(n3091), .ZN(n5870) );
  OR2_X1 U3697 ( .A1(n4845), .A2(n6059), .ZN(n5043) );
  AND2_X1 U3698 ( .A1(n4419), .A2(n3332), .ZN(n5144) );
  INV_X1 U3699 ( .A(n4866), .ZN(n4914) );
  OAI21_X1 U3700 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6588), .A(n4869), 
        .ZN(n4840) );
  AND2_X1 U3701 ( .A1(n4994), .A2(n4959), .ZN(n4964) );
  INV_X1 U3702 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6059) );
  INV_X1 U3703 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5241) );
  INV_X1 U3704 ( .A(n3114), .ZN(n3113) );
  AOI21_X1 U3705 ( .B1(n5254), .B2(REIP_REG_24__SCAN_IN), .A(n3115), .ZN(n3114) );
  OAI21_X1 U3706 ( .B1(n5769), .B2(n6172), .A(n3116), .ZN(n3115) );
  OAI21_X1 U3707 ( .B1(n6186), .B2(n5274), .A(n3120), .ZN(n3119) );
  AND2_X1 U3708 ( .A1(n5371), .A2(n3121), .ZN(n3118) );
  INV_X1 U3709 ( .A(n5581), .ZN(n3121) );
  AND2_X1 U3710 ( .A1(n5371), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6142) );
  AND2_X1 U3711 ( .A1(n4167), .A2(n4165), .ZN(n6161) );
  INV_X1 U3712 ( .A(n6161), .ZN(n6172) );
  NAND2_X1 U3713 ( .A1(n4205), .A2(n5371), .ZN(n6155) );
  INV_X1 U3714 ( .A(n6182), .ZN(n5405) );
  OR2_X1 U3715 ( .A1(n5734), .A2(n5428), .ZN(n4089) );
  NAND2_X1 U3716 ( .A1(n4054), .A2(n3168), .ZN(n5271) );
  OR2_X1 U3717 ( .A1(n4566), .A2(n4444), .ZN(n4218) );
  INV_X1 U3718 ( .A(n5491), .ZN(n5486) );
  INV_X1 U3719 ( .A(n6233), .ZN(n6212) );
  XNOR2_X1 U3720 ( .A(n4152), .B(n4151), .ZN(n4230) );
  NAND2_X1 U3721 ( .A1(n4150), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4152)
         );
  INV_X1 U3722 ( .A(n4149), .ZN(n4150) );
  NAND2_X1 U3723 ( .A1(n3933), .A2(n3934), .ZN(n3935) );
  NAND2_X1 U3724 ( .A1(n5772), .A2(n3014), .ZN(n5747) );
  NOR2_X2 U3725 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6419) );
  INV_X1 U3726 ( .A(n6419), .ZN(n6476) );
  INV_X1 U3727 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U3728 ( .A1(n3979), .A2(n3332), .ZN(n3944) );
  NAND2_X1 U3729 ( .A1(n3098), .A2(n4140), .ZN(n3097) );
  NAND2_X1 U3730 ( .A1(n3976), .A2(n3016), .ZN(n3095) );
  NAND2_X1 U3731 ( .A1(n3944), .A2(n3324), .ZN(n3947) );
  XNOR2_X1 U3732 ( .A(n3481), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3965)
         );
  NAND2_X1 U3733 ( .A1(n3961), .A2(n3960), .ZN(n3967) );
  AND2_X1 U3734 ( .A1(n6309), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3941)
         );
  XNOR2_X1 U3735 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3942) );
  NAND2_X1 U3736 ( .A1(n3225), .A2(n5147), .ZN(n3810) );
  NAND2_X1 U3737 ( .A1(n3152), .A2(n5580), .ZN(n3151) );
  INV_X1 U3738 ( .A(n3154), .ZN(n3152) );
  AND2_X1 U3739 ( .A1(n4318), .A2(n4319), .ZN(n3136) );
  AND2_X1 U3740 ( .A1(n3345), .A2(n4250), .ZN(n4253) );
  NAND2_X1 U3741 ( .A1(n3421), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3310)
         );
  AOI22_X1 U3742 ( .A1(n3372), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U3743 ( .A1(n2977), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3248) );
  OR2_X1 U3744 ( .A1(n3351), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3352)
         );
  INV_X1 U3745 ( .A(n3351), .ZN(n3077) );
  NAND2_X1 U3746 ( .A1(n3189), .A2(n3039), .ZN(n3078) );
  NAND2_X1 U3747 ( .A1(n3975), .A2(n3974), .ZN(n4143) );
  OR2_X1 U3748 ( .A1(n3973), .A2(n3972), .ZN(n3975) );
  AND2_X1 U3749 ( .A1(n6662), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3972)
         );
  NAND2_X1 U3750 ( .A1(n3052), .A2(n3977), .ZN(n3051) );
  INV_X1 U3751 ( .A(n3934), .ZN(n3212) );
  NOR2_X1 U3752 ( .A1(n5211), .A2(n3089), .ZN(n3088) );
  INV_X1 U3753 ( .A(n5223), .ZN(n3089) );
  INV_X1 U3754 ( .A(n5259), .ZN(n3204) );
  NOR2_X1 U3755 ( .A1(n5274), .A2(n3106), .ZN(n3105) );
  AND2_X1 U3756 ( .A1(n5269), .A2(n3206), .ZN(n3205) );
  INV_X1 U3757 ( .A(n5280), .ZN(n3206) );
  NAND2_X1 U3758 ( .A1(n5430), .A2(n3208), .ZN(n3207) );
  OR2_X1 U3759 ( .A1(n3198), .A2(n5343), .ZN(n3087) );
  OR2_X1 U3760 ( .A1(n3199), .A2(n5359), .ZN(n3198) );
  XNOR2_X1 U3761 ( .A(n3530), .B(n3531), .ZN(n4273) );
  OR2_X1 U3762 ( .A1(n5199), .A2(n4086), .ZN(n3174) );
  INV_X1 U3763 ( .A(n5126), .ZN(n3165) );
  NAND2_X1 U3764 ( .A1(n3143), .A2(n4238), .ZN(n4272) );
  AND2_X2 U3765 ( .A1(n4679), .A2(n4250), .ZN(n4261) );
  OAI21_X1 U3766 ( .B1(n3963), .B2(n4806), .A(n3025), .ZN(n3444) );
  NAND2_X1 U3767 ( .A1(n3191), .A2(n3414), .ZN(n3141) );
  AOI22_X1 U3768 ( .A1(n3979), .A2(n4233), .B1(INSTQUEUE_REG_0__2__SCAN_IN), 
        .B2(n3970), .ZN(n3414) );
  NAND2_X1 U3769 ( .A1(n3069), .A2(n3067), .ZN(n3079) );
  NAND2_X1 U3770 ( .A1(n4341), .A2(n3064), .ZN(n3069) );
  NAND2_X1 U3771 ( .A1(n3070), .A2(n3068), .ZN(n3067) );
  AND2_X1 U3772 ( .A1(n5041), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4751) );
  AND2_X2 U3773 ( .A1(n3233), .A2(n3232), .ZN(n3361) );
  AOI22_X1 U3774 ( .A1(n3465), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3230) );
  AND2_X1 U3775 ( .A1(n3460), .A2(n5039), .ZN(n6388) );
  AND2_X1 U3776 ( .A1(n3394), .A2(n6423), .ZN(n4791) );
  NAND2_X1 U3777 ( .A1(n3478), .A2(n3477), .ZN(n4785) );
  INV_X1 U3778 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6547) );
  AND2_X1 U3779 ( .A1(n4419), .A2(n4146), .ZN(n4404) );
  NAND2_X1 U3780 ( .A1(n4213), .A2(n4537), .ZN(n4408) );
  NAND2_X1 U3781 ( .A1(n3058), .A2(n3057), .ZN(n3056) );
  INV_X1 U3782 ( .A(n6025), .ZN(n3058) );
  NOR2_X1 U3783 ( .A1(n3059), .A2(n5588), .ZN(n3057) );
  NAND2_X1 U3784 ( .A1(n4332), .A2(n3038), .ZN(n3062) );
  INV_X1 U3785 ( .A(n4182), .ZN(n3060) );
  OAI21_X1 U3786 ( .B1(n3368), .B2(n4685), .A(n3332), .ZN(n3369) );
  AND3_X1 U3787 ( .A1(n3365), .A2(n3364), .A3(n4712), .ZN(n3366) );
  NAND2_X1 U3788 ( .A1(n3354), .A2(n3040), .ZN(n3186) );
  AND2_X1 U3789 ( .A1(n3169), .A2(n4064), .ZN(n3168) );
  NAND2_X1 U3790 ( .A1(n3530), .A2(n3144), .ZN(n4239) );
  NOR2_X1 U3791 ( .A1(n3213), .A2(n3211), .ZN(n3210) );
  INV_X1 U3792 ( .A(n5179), .ZN(n3213) );
  INV_X1 U3793 ( .A(n4191), .ZN(n3209) );
  OR2_X1 U3794 ( .A1(n4109), .A2(n5180), .ZN(n4149) );
  NAND2_X1 U3795 ( .A1(n3879), .A2(n2991), .ZN(n3931) );
  NOR2_X1 U3796 ( .A1(n3878), .A2(n5241), .ZN(n3879) );
  NAND2_X1 U3797 ( .A1(n3879), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3914)
         );
  NAND2_X1 U3798 ( .A1(n3724), .A2(n3000), .ZN(n3745) );
  AOI21_X1 U3799 ( .B1(n3744), .B2(n3743), .A(n3742), .ZN(n5427) );
  AND2_X1 U3800 ( .A1(n3709), .A2(n3708), .ZN(n5291) );
  NAND2_X1 U3801 ( .A1(n3688), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3704)
         );
  NOR2_X1 U3802 ( .A1(n3672), .A2(n5325), .ZN(n3688) );
  CLKBUF_X1 U3803 ( .A(n5303), .Z(n5304) );
  NAND2_X1 U3804 ( .A1(n3603), .A2(n3109), .ZN(n3672) );
  AND2_X1 U3805 ( .A1(n3001), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3109)
         );
  NAND2_X1 U3806 ( .A1(n3084), .A2(n5317), .ZN(n3083) );
  INV_X1 U3807 ( .A(n3085), .ZN(n3084) );
  AND3_X1 U3808 ( .A1(n3587), .A2(n3586), .A3(n3585), .ZN(n5123) );
  CLKBUF_X1 U3809 ( .A(n4903), .Z(n4904) );
  AOI21_X1 U3810 ( .B1(n4282), .B2(n3685), .A(n3547), .ZN(n4832) );
  NAND2_X1 U3811 ( .A1(n3503), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3522)
         );
  NOR2_X1 U3812 ( .A1(n3483), .A2(n3482), .ZN(n3503) );
  INV_X1 U3813 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3482) );
  AOI21_X1 U3814 ( .B1(n6590), .B2(n3685), .A(n3488), .ZN(n4622) );
  NAND2_X1 U3815 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3483) );
  AND2_X1 U3816 ( .A1(n3456), .A2(n3455), .ZN(n4492) );
  AOI21_X1 U3817 ( .B1(n3195), .B2(n3194), .A(n3018), .ZN(n3193) );
  NOR2_X1 U3818 ( .A1(n5578), .A2(n5569), .ZN(n5563) );
  AND2_X1 U3819 ( .A1(n4051), .A2(n4050), .ZN(n5432) );
  NAND2_X1 U3820 ( .A1(n3137), .A2(n3184), .ZN(n5558) );
  OR2_X1 U3821 ( .A1(n4315), .A2(n3185), .ZN(n3183) );
  AND2_X1 U3822 ( .A1(n4037), .A2(n4036), .ZN(n5348) );
  NAND2_X1 U3823 ( .A1(n5346), .A2(n5348), .ZN(n5347) );
  NAND2_X1 U3824 ( .A1(n3145), .A2(n2993), .ZN(n5652) );
  NAND2_X1 U3825 ( .A1(n6049), .A2(n6566), .ZN(n4225) );
  NAND2_X1 U3826 ( .A1(n3165), .A2(n4030), .ZN(n6106) );
  AND2_X1 U3827 ( .A1(n4027), .A2(n4026), .ZN(n4907) );
  INV_X1 U3828 ( .A(n3161), .ZN(n3160) );
  NAND2_X1 U3829 ( .A1(n4624), .A2(n3161), .ZN(n5105) );
  INV_X1 U3830 ( .A(n6277), .ZN(n5114) );
  INV_X1 U3831 ( .A(n4268), .ZN(n3181) );
  OR2_X1 U3832 ( .A1(n3427), .A2(n3426), .ZN(n4260) );
  OR2_X1 U3833 ( .A1(n3987), .A2(n3701), .ZN(n5142) );
  AND2_X1 U3834 ( .A1(n4433), .A2(n4432), .ZN(n6540) );
  CLKBUF_X3 U3835 ( .A(n3340), .Z(n4537) );
  NAND2_X1 U3836 ( .A1(n4652), .A2(n4656), .ZN(n4697) );
  INV_X1 U3837 ( .A(n4840), .ZN(n6426) );
  INV_X1 U3838 ( .A(n4528), .ZN(n4431) );
  AND2_X1 U3839 ( .A1(n5170), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3994) );
  INV_X1 U3840 ( .A(n4734), .ZN(n4651) );
  INV_X1 U3841 ( .A(n6573), .ZN(n6559) );
  NAND2_X1 U3842 ( .A1(n5173), .A2(n5171), .ZN(n6609) );
  NOR2_X1 U3843 ( .A1(n6135), .A2(n6057), .ZN(n6167) );
  CLKBUF_X1 U3844 ( .A(n3433), .Z(n6421) );
  XNOR2_X1 U3845 ( .A(n4163), .B(n4162), .ZN(n5687) );
  AND2_X1 U3846 ( .A1(n4054), .A2(n3169), .ZN(n5281) );
  INV_X1 U3847 ( .A(n5506), .ZN(n5461) );
  NOR2_X1 U3848 ( .A1(n6779), .A2(n4482), .ZN(n6197) );
  INV_X2 U3849 ( .A(n6197), .ZN(n6776) );
  OR2_X1 U3850 ( .A1(n6779), .A2(n4483), .ZN(n5491) );
  OR2_X1 U3851 ( .A1(n4566), .A2(n4565), .ZN(n6233) );
  OR2_X1 U3853 ( .A1(n4566), .A2(n4417), .ZN(n4497) );
  NOR2_X1 U3854 ( .A1(n5173), .A2(n3332), .ZN(n6241) );
  NAND2_X1 U3855 ( .A1(n3794), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3795)
         );
  NAND2_X1 U3856 ( .A1(n3724), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3726)
         );
  NAND2_X1 U3857 ( .A1(n3603), .A2(n3110), .ZN(n3634) );
  NAND2_X1 U3858 ( .A1(n3603), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3619)
         );
  INV_X1 U3859 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6272) );
  OR2_X1 U3860 ( .A1(n4566), .A2(n6552), .ZN(n6256) );
  NAND2_X1 U3861 ( .A1(n6271), .A2(n4484), .ZN(n6254) );
  XNOR2_X1 U3862 ( .A(n4328), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5686)
         );
  AND2_X1 U3863 ( .A1(n3197), .A2(n3028), .ZN(n3129) );
  AOI21_X1 U3864 ( .B1(n2992), .B2(n5726), .A(n5155), .ZN(n5156) );
  AND2_X1 U3865 ( .A1(n6286), .A2(n5737), .ZN(n3103) );
  NAND2_X1 U3866 ( .A1(n3197), .A2(n4326), .ZN(n5534) );
  NAND2_X1 U3867 ( .A1(n5800), .A2(n3013), .ZN(n5784) );
  NAND2_X1 U3868 ( .A1(n3148), .A2(n3153), .ZN(n5579) );
  OR2_X1 U3869 ( .A1(n5598), .A2(n3154), .ZN(n3148) );
  NAND2_X1 U3870 ( .A1(n5826), .A2(n5543), .ZN(n5587) );
  NAND2_X1 U3871 ( .A1(n5598), .A2(n5597), .ZN(n5826) );
  INV_X1 U3872 ( .A(n5872), .ZN(n6039) );
  NAND2_X1 U3873 ( .A1(n3145), .A2(n4310), .ZN(n5667) );
  INV_X1 U3874 ( .A(n3138), .ZN(n5664) );
  NAND2_X1 U3875 ( .A1(n3071), .A2(n3073), .ZN(n5676) );
  NAND2_X1 U3876 ( .A1(n3142), .A2(n4301), .ZN(n5681) );
  AND2_X1 U3877 ( .A1(n4560), .A2(n4545), .ZN(n6300) );
  INV_X1 U3878 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6309) );
  INV_X1 U3879 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6662) );
  OAI21_X1 U3880 ( .B1(n4733), .B2(n6586), .A(n6394), .ZN(n6599) );
  INV_X1 U3881 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5153) );
  INV_X1 U3882 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5170) );
  INV_X1 U3883 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6053) );
  NOR2_X1 U3884 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6049) );
  NAND2_X1 U3885 ( .A1(n4914), .A2(n4757), .ZN(n4824) );
  OAI21_X1 U3886 ( .B1(n4872), .B2(n4871), .A(n5977), .ZN(n4896) );
  INV_X1 U3887 ( .A(n5057), .ZN(n5081) );
  INV_X1 U3888 ( .A(n6418), .ZN(n6391) );
  NOR2_X2 U3889 ( .A1(n6428), .A2(n4920), .ZN(n6414) );
  INV_X1 U3890 ( .A(n6536), .ZN(n6477) );
  INV_X1 U3891 ( .A(n5006), .ZN(n6475) );
  NOR2_X1 U3892 ( .A1(n6713), .A2(n6394), .ZN(n6474) );
  NOR2_X1 U3893 ( .A1(n4692), .A2(n6394), .ZN(n6491) );
  NOR2_X1 U3894 ( .A1(n4680), .A2(n6394), .ZN(n6497) );
  NOR2_X1 U3895 ( .A1(n4667), .A2(n6394), .ZN(n6509) );
  NOR2_X1 U3896 ( .A1(n6675), .A2(n6394), .ZN(n6515) );
  NOR2_X1 U3897 ( .A1(n4837), .A2(n6394), .ZN(n6521) );
  OAI21_X1 U3898 ( .B1(n4843), .B2(n4842), .A(n4841), .ZN(n4862) );
  AND2_X1 U3899 ( .A1(n4846), .A2(n4662), .ZN(n6531) );
  OAI211_X1 U3900 ( .C1(n4963), .C2(n6588), .A(n4962), .B(n4961), .ZN(n4987)
         );
  INV_X1 U3901 ( .A(n6491), .ZN(n6363) );
  INV_X1 U3902 ( .A(n6497), .ZN(n6366) );
  INV_X1 U3903 ( .A(n6503), .ZN(n6369) );
  INV_X1 U3904 ( .A(n6509), .ZN(n6372) );
  INV_X1 U3905 ( .A(n6521), .ZN(n6378) );
  NAND2_X1 U3906 ( .A1(n4994), .A2(n6429), .ZN(n5032) );
  INV_X1 U3907 ( .A(n4964), .ZN(n5033) );
  INV_X1 U3908 ( .A(n6528), .ZN(n6384) );
  NAND2_X1 U3909 ( .A1(n4431), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U3910 ( .A1(n3994), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6573) );
  INV_X1 U3911 ( .A(n6568), .ZN(n6615) );
  INV_X1 U3912 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6588) );
  AND2_X1 U3913 ( .A1(n6014), .A2(STATE_REG_1__SCAN_IN), .ZN(n6021) );
  OAI211_X1 U3914 ( .C1(n5471), .C2(n6095), .A(n3117), .B(n3024), .ZN(U2803)
         );
  INV_X1 U3915 ( .A(n5242), .ZN(n3117) );
  AOI21_X1 U3916 ( .B1(n4205), .B2(n3118), .A(n3119), .ZN(n5275) );
  OR4_X1 U3917 ( .A1(n4346), .A2(n4345), .A3(n4344), .A4(n5391), .ZN(U2826) );
  NAND2_X1 U3918 ( .A1(n4091), .A2(n4090), .ZN(U2831) );
  AND2_X1 U3919 ( .A1(n4089), .A2(n4088), .ZN(n4090) );
  NAND2_X1 U3920 ( .A1(n5506), .A2(n6193), .ZN(n4091) );
  AND2_X2 U3921 ( .A1(n5147), .A2(n4706), .ZN(n3298) );
  NAND2_X1 U3922 ( .A1(n3201), .A2(n3205), .ZN(n5258) );
  OR2_X1 U3923 ( .A1(n3976), .A2(n4141), .ZN(n2990) );
  INV_X1 U3924 ( .A(n5303), .ZN(n3080) );
  INV_X1 U3925 ( .A(n2973), .ZN(n3808) );
  AND3_X1 U3926 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .A3(PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n2991) );
  AND2_X2 U3927 ( .A1(n3197), .A2(n3015), .ZN(n2992) );
  NOR2_X1 U3928 ( .A1(n5237), .A2(n3041), .ZN(n4112) );
  OR2_X1 U3929 ( .A1(n4544), .A2(n6566), .ZN(n3055) );
  AND2_X2 U3930 ( .A1(n4537), .A2(n3332), .ZN(n3003) );
  NAND2_X1 U3931 ( .A1(n5222), .A2(n5223), .ZN(n5210) );
  OR2_X1 U3932 ( .A1(n4903), .A2(n3199), .ZN(n5120) );
  OR2_X1 U3933 ( .A1(n4903), .A2(n3085), .ZN(n5315) );
  NOR2_X1 U3934 ( .A1(n5303), .A2(n3207), .ZN(n5426) );
  AND2_X1 U3935 ( .A1(n3138), .A2(n4310), .ZN(n2993) );
  NAND2_X1 U3936 ( .A1(n3190), .A2(n3192), .ZN(n4437) );
  NOR2_X1 U3937 ( .A1(n3164), .A2(n6107), .ZN(n2995) );
  OR3_X1 U3938 ( .A1(n3973), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6662), 
        .ZN(n4144) );
  INV_X1 U3939 ( .A(n4144), .ZN(n3102) );
  OR3_X1 U3940 ( .A1(n5187), .A2(REIP_REG_30__SCAN_IN), .A3(n5493), .ZN(n2996)
         );
  NAND2_X1 U3941 ( .A1(n5171), .A2(n3037), .ZN(n2997) );
  NOR2_X1 U3942 ( .A1(n5279), .A2(n3034), .ZN(n5244) );
  NAND2_X1 U3943 ( .A1(n3963), .A2(n3962), .ZN(n2998) );
  AND2_X1 U3944 ( .A1(n3949), .A2(n3948), .ZN(n2999) );
  NOR2_X1 U3945 ( .A1(n4566), .A2(n4408), .ZN(n3063) );
  AND2_X1 U3946 ( .A1(n3107), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3000)
         );
  AND2_X1 U3947 ( .A1(n3110), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3001)
         );
  AND2_X1 U3948 ( .A1(n3081), .A2(n3761), .ZN(n3002) );
  NAND2_X2 U3949 ( .A1(n3431), .A2(n3430), .ZN(n4662) );
  NAND2_X1 U3951 ( .A1(n5442), .A2(n5441), .ZN(n5297) );
  INV_X1 U3952 ( .A(n3314), .ZN(n3374) );
  NAND2_X1 U3953 ( .A1(n3183), .A2(n4318), .ZN(n5602) );
  NOR2_X1 U3954 ( .A1(n5279), .A2(n5280), .ZN(n5268) );
  NAND2_X1 U3955 ( .A1(n3080), .A2(n3081), .ZN(n5413) );
  NOR2_X1 U3956 ( .A1(n4315), .A2(n3216), .ZN(n3004) );
  OR2_X1 U3957 ( .A1(n2989), .A2(n6307), .ZN(n3005) );
  NOR2_X1 U3958 ( .A1(n4903), .A2(n3083), .ZN(n5302) );
  OR2_X1 U3959 ( .A1(n4903), .A2(n3198), .ZN(n5342) );
  AND2_X1 U3960 ( .A1(n3080), .A2(n3208), .ZN(n3006) );
  NAND2_X1 U3961 ( .A1(n3080), .A2(n3692), .ZN(n5290) );
  AND2_X2 U3962 ( .A1(n4706), .A2(n4415), .ZN(n3313) );
  AND2_X1 U3963 ( .A1(n3189), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3007) );
  AND2_X1 U3964 ( .A1(n3986), .A2(n3344), .ZN(n4213) );
  NAND2_X1 U3965 ( .A1(n4054), .A2(n3217), .ZN(n5416) );
  NOR2_X1 U3966 ( .A1(n5674), .A2(n6736), .ZN(n3008) );
  NOR2_X1 U3967 ( .A1(n4903), .A2(n5123), .ZN(n3009) );
  OR2_X1 U3968 ( .A1(n3330), .A2(n3360), .ZN(n3010) );
  AND2_X1 U3969 ( .A1(n3073), .A2(n3005), .ZN(n3011) );
  NOR2_X1 U3970 ( .A1(n5535), .A2(n3196), .ZN(n3195) );
  INV_X2 U3971 ( .A(n3379), .ZN(n3291) );
  AND2_X1 U3972 ( .A1(n5887), .A2(n5653), .ZN(n3012) );
  OR2_X1 U3973 ( .A1(n5820), .A2(n5790), .ZN(n3013) );
  OR2_X1 U3974 ( .A1(n5820), .A2(n5753), .ZN(n3014) );
  AND2_X1 U3975 ( .A1(n3125), .A2(n3195), .ZN(n3015) );
  INV_X1 U3976 ( .A(n3175), .ZN(n5201) );
  NOR2_X1 U3977 ( .A1(n5215), .A2(n5199), .ZN(n3175) );
  AND2_X1 U3978 ( .A1(n3324), .A2(n3096), .ZN(n3016) );
  OR2_X1 U3979 ( .A1(n3976), .A2(n4143), .ZN(n3017) );
  AND2_X1 U3980 ( .A1(n5674), .A2(n5764), .ZN(n3018) );
  AND3_X1 U3981 ( .A1(n3225), .A2(n5147), .A3(INSTQUEUE_REG_9__4__SCAN_IN), 
        .ZN(n3019) );
  AND2_X1 U3982 ( .A1(n4272), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3020)
         );
  NAND2_X1 U3983 ( .A1(n3979), .A2(n3978), .ZN(n3021) );
  NOR2_X1 U3984 ( .A1(n4903), .A2(n3087), .ZN(n3022) );
  NOR2_X1 U3985 ( .A1(n5609), .A2(n5864), .ZN(n3023) );
  NOR2_X1 U3986 ( .A1(n5243), .A2(n3113), .ZN(n3024) );
  AND2_X1 U3987 ( .A1(n3443), .A2(n3055), .ZN(n3025) );
  NAND2_X1 U3988 ( .A1(n3080), .A2(n3002), .ZN(n5279) );
  AND2_X1 U3989 ( .A1(n4308), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3026)
         );
  AND2_X1 U3990 ( .A1(n3329), .A2(n3010), .ZN(n3980) );
  AND3_X1 U3991 ( .A1(n4537), .A2(n4544), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3970) );
  INV_X1 U3992 ( .A(n3970), .ZN(n3963) );
  NOR2_X1 U3993 ( .A1(n6084), .A2(n6025), .ZN(n3027) );
  AND2_X1 U3994 ( .A1(n3195), .A2(n3126), .ZN(n3028) );
  NOR2_X1 U3995 ( .A1(n2988), .A2(n4316), .ZN(n3029) );
  INV_X1 U3996 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6566) );
  OR2_X1 U3997 ( .A1(n6084), .A2(n3056), .ZN(n3030) );
  INV_X1 U3998 ( .A(n3964), .ZN(n3099) );
  INV_X1 U3999 ( .A(n5523), .ZN(n3130) );
  OR2_X1 U4000 ( .A1(n2989), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5523)
         );
  NOR2_X2 U4001 ( .A1(n6779), .A2(n4536), .ZN(n3031) );
  AND2_X1 U4002 ( .A1(n3724), .A2(n3107), .ZN(n3033) );
  NAND2_X1 U4003 ( .A1(n3204), .A2(n3205), .ZN(n3034) );
  NOR2_X1 U4004 ( .A1(n5126), .A2(n3163), .ZN(n5346) );
  INV_X1 U4005 ( .A(n3090), .ZN(n6201) );
  NOR2_X1 U4006 ( .A1(n6233), .A2(n3345), .ZN(n3090) );
  AND2_X1 U4007 ( .A1(n3603), .A2(n3001), .ZN(n3035) );
  AND2_X1 U4008 ( .A1(n5371), .A2(n4153), .ZN(n6152) );
  AND2_X1 U4009 ( .A1(n4624), .A2(n4623), .ZN(n3036) );
  NOR2_X1 U4010 ( .A1(n6564), .A2(n4148), .ZN(n3037) );
  INV_X1 U4011 ( .A(n3063), .ZN(n5173) );
  AND2_X1 U4012 ( .A1(n4169), .A2(n3060), .ZN(n3038) );
  OR2_X1 U4013 ( .A1(n3563), .A2(n3562), .ZN(n4304) );
  AND2_X1 U4014 ( .A1(STATE2_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3039) );
  NAND2_X1 U4015 ( .A1(STATE2_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3040) );
  INV_X1 U4016 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U4017 ( .A1(n3212), .A2(n5198), .ZN(n3211) );
  INV_X1 U4018 ( .A(n5414), .ZN(n3761) );
  OR2_X1 U4019 ( .A1(n3211), .A2(n3044), .ZN(n3041) );
  NAND2_X1 U4020 ( .A1(n3415), .A2(n3706), .ZN(n4490) );
  AND2_X1 U4021 ( .A1(n3210), .A2(n3209), .ZN(n3042) );
  AND2_X1 U4022 ( .A1(n3332), .A2(n3324), .ZN(n4280) );
  AND2_X1 U4023 ( .A1(n3165), .A2(n2995), .ZN(n3043) );
  NAND2_X1 U4024 ( .A1(n3088), .A2(n3863), .ZN(n3044) );
  INV_X1 U4025 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5978) );
  INV_X1 U4026 ( .A(n6258), .ZN(n6265) );
  INV_X1 U4027 ( .A(n4030), .ZN(n3164) );
  INV_X1 U4028 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6678) );
  AND2_X1 U4029 ( .A1(n3000), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3045)
         );
  AND2_X1 U4030 ( .A1(n3105), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3046)
         );
  AND2_X1 U4031 ( .A1(n2991), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3047)
         );
  INV_X1 U4032 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4457) );
  INV_X1 U4033 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3112) );
  INV_X1 U4034 ( .A(REIP_REG_21__SCAN_IN), .ZN(n3059) );
  INV_X1 U4035 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4436) );
  INV_X1 U4036 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3106) );
  INV_X1 U4037 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3180) );
  INV_X1 U4038 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3111) );
  OR2_X1 U4039 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3048) );
  NAND2_X1 U4040 ( .A1(n6143), .A2(EBX_REG_21__SCAN_IN), .ZN(n3120) );
  NAND2_X1 U4041 ( .A1(n6143), .A2(EBX_REG_24__SCAN_IN), .ZN(n3116) );
  NAND2_X1 U4042 ( .A1(n3553), .A2(n3552), .ZN(n4281) );
  INV_X2 U4043 ( .A(n4309), .ZN(n5655) );
  AND2_X1 U4044 ( .A1(n3342), .A2(n3341), .ZN(n4138) );
  NAND2_X1 U4045 ( .A1(n3353), .A2(n3352), .ZN(n3389) );
  NAND2_X1 U4046 ( .A1(n3134), .A2(n4319), .ZN(n3133) );
  INV_X1 U4047 ( .A(n3184), .ZN(n3134) );
  INV_X1 U4048 ( .A(n3350), .ZN(n3353) );
  AND2_X2 U4049 ( .A1(n3135), .A2(n3133), .ZN(n4322) );
  NAND2_X2 U4050 ( .A1(n4322), .A2(n4321), .ZN(n5598) );
  AOI22_X1 U4051 ( .A1(n3421), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3049), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4052 ( .A1(n3312), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3049), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4053 ( .A1(n3470), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3049), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4054 ( .A1(n3372), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3049), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4055 ( .A1(n3372), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3049), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3290) );
  NAND3_X1 U4056 ( .A1(n3054), .A2(n3101), .A3(n3053), .ZN(n3052) );
  NAND3_X1 U4057 ( .A1(n2999), .A2(n2990), .A3(n3964), .ZN(n3053) );
  INV_X1 U4058 ( .A(n3055), .ZN(n3066) );
  NAND2_X1 U4059 ( .A1(n3055), .A2(n4537), .ZN(n3428) );
  NOR2_X1 U4060 ( .A1(n3997), .A2(n3055), .ZN(n3998) );
  NAND2_X1 U4061 ( .A1(n3431), .A2(n3055), .ZN(n3070) );
  INV_X1 U4062 ( .A(n3062), .ZN(n5364) );
  NAND2_X1 U4063 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n3061) );
  INV_X1 U4064 ( .A(n3065), .ZN(n3064) );
  NAND2_X2 U4066 ( .A1(n3071), .A2(n3011), .ZN(n3146) );
  NAND3_X1 U4067 ( .A1(n3530), .A2(n4280), .A3(n3144), .ZN(n3143) );
  NAND2_X1 U4068 ( .A1(n4322), .A2(n3075), .ZN(n3076) );
  AND2_X2 U4070 ( .A1(n3076), .A2(n3193), .ZN(n5525) );
  NAND3_X1 U4071 ( .A1(n3078), .A2(n3350), .A3(n3077), .ZN(n3391) );
  NAND3_X1 U4072 ( .A1(n4247), .A2(n3685), .A3(n4246), .ZN(n3415) );
  NOR2_X1 U4073 ( .A1(n5237), .A2(n5239), .ZN(n5222) );
  NAND3_X1 U4074 ( .A1(n3225), .A2(n5147), .A3(INSTQUEUE_REG_9__1__SCAN_IN), 
        .ZN(n3317) );
  NAND2_X1 U4075 ( .A1(n5913), .A2(n5906), .ZN(n5133) );
  OAI211_X1 U4076 ( .C1(n3095), .C2(n3094), .A(n3097), .B(n3092), .ZN(n3949)
         );
  NAND2_X1 U4077 ( .A1(n3093), .A2(n3976), .ZN(n3092) );
  NAND3_X1 U4078 ( .A1(n3946), .A2(n3945), .A3(n3979), .ZN(n3093) );
  INV_X1 U4079 ( .A(n3944), .ZN(n3094) );
  INV_X1 U4080 ( .A(n4140), .ZN(n3096) );
  INV_X1 U4081 ( .A(n3946), .ZN(n3098) );
  NOR2_X2 U4082 ( .A1(n5784), .A2(n3104), .ZN(n5772) );
  NAND2_X1 U4083 ( .A1(n3794), .A2(n3046), .ZN(n3843) );
  INV_X1 U4084 ( .A(n3798), .ZN(n3842) );
  INV_X1 U4085 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U4086 ( .A1(n3879), .A2(n3047), .ZN(n4109) );
  INV_X1 U4087 ( .A(n4109), .ZN(n4108) );
  NAND2_X1 U4088 ( .A1(n3122), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3350) );
  NAND3_X1 U4089 ( .A1(n6048), .A2(n3123), .A3(n4555), .ZN(n3122) );
  NAND2_X2 U4090 ( .A1(n4138), .A2(n4691), .ZN(n6048) );
  NAND3_X1 U4091 ( .A1(n4213), .A2(n4537), .A3(n3124), .ZN(n3123) );
  NAND2_X1 U4092 ( .A1(n3348), .A2(n4438), .ZN(n4555) );
  AOI21_X1 U4093 ( .B1(n5155), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n3129), 
        .ZN(n4328) );
  NAND3_X1 U4095 ( .A1(n2994), .A2(n3146), .A3(n3136), .ZN(n3135) );
  NAND3_X1 U4096 ( .A1(n2994), .A2(n3146), .A3(n4318), .ZN(n3137) );
  NAND2_X2 U4097 ( .A1(n3140), .A2(n3139), .ZN(n4529) );
  NAND2_X1 U4098 ( .A1(n5131), .A2(n5130), .ZN(n3142) );
  XNOR2_X2 U4099 ( .A(n4272), .B(n4240), .ZN(n4739) );
  CLKBUF_X1 U4100 ( .A(n3146), .Z(n3145) );
  NAND2_X1 U4101 ( .A1(n3147), .A2(n3149), .ZN(n5546) );
  NAND2_X1 U4102 ( .A1(n4004), .A2(n3158), .ZN(n4008) );
  NAND2_X2 U4103 ( .A1(n4054), .A2(n3166), .ZN(n5273) );
  NAND2_X1 U4104 ( .A1(n5228), .A2(n3171), .ZN(n4197) );
  NAND2_X1 U4105 ( .A1(n5228), .A2(n5213), .ZN(n5215) );
  NOR2_X2 U4106 ( .A1(n5215), .A2(n3174), .ZN(n5183) );
  NAND2_X1 U4107 ( .A1(n3179), .A2(n4271), .ZN(n4738) );
  OAI21_X2 U4108 ( .B1(n3179), .B2(n3178), .A(n3176), .ZN(n5102) );
  INV_X1 U4109 ( .A(n4271), .ZN(n3177) );
  INV_X1 U4110 ( .A(n4739), .ZN(n3178) );
  NAND2_X1 U4111 ( .A1(n4634), .A2(n4633), .ZN(n3179) );
  NAND2_X1 U4112 ( .A1(n3181), .A2(n3180), .ZN(n4569) );
  NAND4_X1 U4113 ( .A1(n3367), .A2(n3357), .A3(n3336), .A4(n3335), .ZN(n3189)
         );
  NAND4_X1 U4114 ( .A1(n3188), .A2(n3336), .A3(n3367), .A4(n3357), .ZN(n3187)
         );
  CLKBUF_X1 U4115 ( .A(n4726), .Z(n3190) );
  NAND3_X1 U4116 ( .A1(n4726), .A2(n3192), .A3(n6566), .ZN(n3191) );
  NAND2_X1 U4117 ( .A1(n3399), .A2(n3398), .ZN(n3192) );
  AND2_X2 U4118 ( .A1(n3502), .A2(n3479), .ZN(n6590) );
  INV_X1 U4119 ( .A(n5279), .ZN(n3201) );
  NAND2_X1 U4120 ( .A1(n3201), .A2(n3202), .ZN(n5237) );
  NAND2_X1 U4121 ( .A1(n5197), .A2(n3210), .ZN(n5178) );
  NAND2_X1 U4122 ( .A1(n5197), .A2(n5198), .ZN(n3933) );
  INV_X1 U4123 ( .A(n4112), .ZN(n3936) );
  XNOR2_X2 U4124 ( .A(n5565), .B(n5564), .ZN(n5780) );
  OR2_X2 U4125 ( .A1(n5563), .A2(n5562), .ZN(n5565) );
  AOI22_X1 U4126 ( .A1(n3312), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4127 ( .A1(n3312), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3223) );
  INV_X1 U4128 ( .A(n3334), .ZN(n3335) );
  AND2_X2 U4129 ( .A1(n3480), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3220)
         );
  AOI22_X1 U4130 ( .A1(n3400), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4131 ( .A1(n3303), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3224) );
  INV_X1 U4132 ( .A(n4440), .ZN(n3326) );
  NAND2_X1 U4133 ( .A1(n6590), .A2(n5044), .ZN(n6428) );
  NAND2_X1 U4134 ( .A1(n6590), .A2(n4280), .ZN(n4245) );
  NAND2_X1 U4135 ( .A1(n5920), .A2(n4912), .ZN(n6352) );
  AND2_X1 U4136 ( .A1(n5920), .A2(n4785), .ZN(n4994) );
  OR2_X1 U4137 ( .A1(n6590), .A2(n5920), .ZN(n4866) );
  INV_X1 U4138 ( .A(n5920), .ZN(n5044) );
  NAND2_X1 U4139 ( .A1(n4653), .A2(n6566), .ZN(n3478) );
  CLKBUF_X1 U4140 ( .A(n4653), .Z(n4654) );
  NAND2_X1 U4141 ( .A1(n5686), .A2(n4329), .ZN(n4330) );
  INV_X1 U4142 ( .A(n5169), .ZN(n5157) );
  INV_X2 U4143 ( .A(n5452), .ZN(n6195) );
  AND2_X1 U4144 ( .A1(n4000), .A2(n3999), .ZN(n5452) );
  AND2_X1 U4145 ( .A1(n5489), .A2(n4672), .ZN(n3214) );
  AND2_X1 U4146 ( .A1(n5706), .A2(n6286), .ZN(n3215) );
  INV_X1 U4147 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3725) );
  INV_X1 U4148 ( .A(n5428), .ZN(n6192) );
  NAND2_X1 U4149 ( .A1(n6195), .A2(n4672), .ZN(n5428) );
  NAND2_X1 U4150 ( .A1(n5663), .A2(n4314), .ZN(n3216) );
  NOR2_X1 U4151 ( .A1(n5432), .A2(n5431), .ZN(n3217) );
  INV_X1 U4152 ( .A(n3819), .ZN(n3859) );
  NAND2_X1 U4153 ( .A1(n3980), .A2(n3331), .ZN(n3368) );
  INV_X1 U4154 ( .A(n4261), .ZN(n3982) );
  INV_X1 U4155 ( .A(n3537), .ZN(n3593) );
  OR2_X1 U4156 ( .A1(n3519), .A2(n3518), .ZN(n4283) );
  OR2_X1 U4157 ( .A1(n3893), .A2(n3892), .ZN(n3900) );
  INV_X1 U4158 ( .A(n4832), .ZN(n3548) );
  INV_X1 U4159 ( .A(n4648), .ZN(n3528) );
  INV_X1 U4160 ( .A(n3398), .ZN(n3396) );
  OR2_X1 U4161 ( .A1(n3875), .A2(n3874), .ZN(n3894) );
  INV_X1 U4162 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5274) );
  INV_X1 U4163 ( .A(n5439), .ZN(n3692) );
  OR2_X1 U4164 ( .A1(n3543), .A2(n3542), .ZN(n4286) );
  INV_X1 U4165 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U4166 ( .A1(n4041), .A2(n4040), .ZN(n5321) );
  AND2_X1 U4167 ( .A1(n3388), .A2(n3387), .ZN(n3371) );
  AND2_X1 U4168 ( .A1(n4047), .A2(n4046), .ZN(n5441) );
  OR2_X1 U4169 ( .A1(n2989), .A2(n4320), .ZN(n4321) );
  NAND2_X1 U4170 ( .A1(n3464), .A2(n3463), .ZN(n4727) );
  INV_X1 U4171 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5246) );
  INV_X1 U4172 ( .A(n3863), .ZN(n5239) );
  INV_X1 U4173 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5594) );
  AND3_X1 U4174 ( .A1(n3691), .A2(n3690), .A3(n3689), .ZN(n5439) );
  AND3_X1 U4175 ( .A1(n3980), .A2(n4261), .A3(n4217), .ZN(n4421) );
  INV_X1 U4176 ( .A(n5522), .ZN(n4327) );
  OR2_X1 U4177 ( .A1(n5674), .A2(n4325), .ZN(n4326) );
  INV_X1 U4178 ( .A(n6300), .ZN(n6288) );
  INV_X1 U4179 ( .A(n4867), .ZN(n4898) );
  NAND2_X1 U4180 ( .A1(n4914), .A2(n6429), .ZN(n5080) );
  OR2_X1 U4181 ( .A1(n6352), .A2(n5929), .ZN(n5961) );
  INV_X1 U4182 ( .A(n6462), .ZN(n6009) );
  INV_X1 U4183 ( .A(n4654), .ZN(n6592) );
  NAND2_X1 U4184 ( .A1(n4994), .A2(n5041), .ZN(n4845) );
  NAND2_X1 U4185 ( .A1(n4404), .A2(n6559), .ZN(n5171) );
  NAND2_X1 U4186 ( .A1(n5452), .A2(EBX_REG_28__SCAN_IN), .ZN(n4088) );
  AND2_X1 U4187 ( .A1(n6195), .A2(n5164), .ZN(n6193) );
  NOR2_X2 U4188 ( .A1(n6779), .A2(n5165), .ZN(n6774) );
  AND3_X2 U4189 ( .A1(n4497), .A2(n4219), .A3(n4218), .ZN(n6779) );
  INV_X1 U4190 ( .A(n6214), .ZN(n6229) );
  OR2_X1 U4191 ( .A1(n4557), .A2(READY_N), .ZN(n4417) );
  OAI21_X1 U4192 ( .B1(n4464), .B2(n6611), .A(n3063), .ZN(n4495) );
  INV_X1 U4193 ( .A(n4497), .ZN(n6243) );
  INV_X1 U4194 ( .A(n4499), .ZN(n6242) );
  INV_X1 U4195 ( .A(n6271), .ZN(n6246) );
  AND2_X1 U4196 ( .A1(n4560), .A2(n5144), .ZN(n5872) );
  INV_X1 U4197 ( .A(n5903), .ZN(n6304) );
  NAND2_X1 U4198 ( .A1(n6566), .A2(n4656), .ZN(n6394) );
  AOI21_X1 U4199 ( .B1(n4914), .B2(n4751), .A(n6476), .ZN(n4790) );
  NOR2_X1 U4200 ( .A1(n4866), .A2(n5967), .ZN(n5057) );
  OAI211_X1 U4201 ( .C1(n5055), .C2(n5054), .A(n6426), .B(n5053), .ZN(n5079)
         );
  INV_X1 U4202 ( .A(n5961), .ZN(n6341) );
  OAI21_X1 U4203 ( .B1(n6389), .B2(n5978), .A(n4869), .ZN(n5933) );
  NOR2_X2 U4204 ( .A1(n6352), .A2(n5967), .ZN(n6380) );
  OR2_X1 U4205 ( .A1(n4662), .A2(n5041), .ZN(n6351) );
  NOR2_X2 U4206 ( .A1(n6428), .A2(n5929), .ZN(n6007) );
  AND2_X1 U4207 ( .A1(n5970), .A2(n4654), .ZN(n6422) );
  NOR2_X1 U4208 ( .A1(n6428), .A2(n5967), .ZN(n6462) );
  INV_X1 U4209 ( .A(n6351), .ZN(n6429) );
  NOR2_X1 U4210 ( .A1(n4686), .A2(n6394), .ZN(n6503) );
  NOR2_X1 U4211 ( .A1(n5040), .A2(n6394), .ZN(n6528) );
  NOR2_X2 U4212 ( .A1(n4845), .A2(n4662), .ZN(n4990) );
  AND2_X1 U4213 ( .A1(n6566), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4222) );
  INV_X1 U4214 ( .A(n4387), .ZN(n4398) );
  NOR2_X1 U4215 ( .A1(n4188), .A2(n4187), .ZN(n4189) );
  INV_X1 U4216 ( .A(n6143), .ZN(n6179) );
  INV_X1 U4217 ( .A(n6142), .ZN(n6186) );
  INV_X1 U4218 ( .A(n6779), .ZN(n5489) );
  INV_X1 U4219 ( .A(n4495), .ZN(n4499) );
  INV_X2 U4220 ( .A(n6241), .ZN(n4526) );
  OR2_X1 U4221 ( .A1(n5302), .A2(n5318), .ZN(n5651) );
  INV_X1 U4222 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U4223 ( .A1(n6256), .A2(n4226), .ZN(n6271) );
  INV_X1 U4224 ( .A(n5686), .ZN(n5715) );
  OR2_X1 U4225 ( .A1(n5807), .A2(n5695), .ZN(n5787) );
  NAND2_X1 U4226 ( .A1(n4560), .A2(n4559), .ZN(n5903) );
  AOI21_X1 U4227 ( .B1(n4790), .B2(n4789), .A(n4788), .ZN(n4830) );
  AOI22_X1 U4228 ( .A1(n5051), .A2(n5054), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5050), .ZN(n5086) );
  NOR2_X1 U4229 ( .A1(n4919), .A2(n4918), .ZN(n4957) );
  AOI22_X1 U4230 ( .A1(n6313), .A2(n6314), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6317), .ZN(n6337) );
  OR2_X1 U4231 ( .A1(n6352), .A2(n6351), .ZN(n6418) );
  INV_X1 U4232 ( .A(n6474), .ZN(n6360) );
  INV_X1 U4233 ( .A(n6515), .ZN(n6375) );
  AOI21_X1 U4234 ( .B1(n6476), .B2(n6432), .A(n6427), .ZN(n6458) );
  NAND2_X1 U4235 ( .A1(n6430), .A2(n6429), .ZN(n6536) );
  INV_X1 U4236 ( .A(n6492), .ZN(n5010) );
  INV_X1 U4237 ( .A(n6530), .ZN(n5018) );
  NAND2_X1 U4238 ( .A1(n4375), .A2(n4402), .ZN(n6582) );
  INV_X1 U4239 ( .A(n4385), .ZN(n4400) );
  OAI211_X1 U4240 ( .C1(n5169), .C2(n6095), .A(n2996), .B(n4212), .ZN(U2797)
         );
  INV_X1 U4241 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3219) );
  INV_X1 U4242 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3480) );
  AND2_X4 U4243 ( .A1(n2981), .A2(n3220), .ZN(n3312) );
  AOI22_X1 U4244 ( .A1(n3421), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3222) );
  AND2_X2 U4245 ( .A1(n4457), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3226)
         );
  AOI22_X1 U4246 ( .A1(n2977), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3229) );
  NOR2_X2 U4247 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4248 ( .A1(n3400), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4249 ( .A1(n3465), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4250 ( .A1(n3400), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4251 ( .A1(n3470), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n2982), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4252 ( .A1(n3303), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4253 ( .A1(n2978), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4254 ( .A1(n3421), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4255 ( .A1(n3312), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3238) );
  INV_X2 U4256 ( .A(n4529), .ZN(n4679) );
  AOI22_X1 U4257 ( .A1(n2963), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4258 ( .A1(n3407), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4259 ( .A1(n3421), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4260 ( .A1(n3373), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3246) );
  NAND3_X1 U4261 ( .A1(n3347), .A2(n4679), .A3(n3324), .ZN(n3262) );
  AOI22_X1 U4262 ( .A1(n3372), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4263 ( .A1(n3303), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4264 ( .A1(n3400), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4265 ( .A1(n3407), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4266 ( .A1(n2977), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4267 ( .A1(n3373), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3257) );
  NAND2_X1 U4268 ( .A1(n3339), .A2(n4529), .ZN(n3261) );
  NAND2_X1 U4269 ( .A1(n3262), .A2(n3261), .ZN(n3286) );
  AOI22_X1 U4270 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n3372), .B1(n3298), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4271 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n3465), .B1(n3373), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4272 ( .A1(n2983), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4273 ( .A1(n3400), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4274 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n3303), .B1(n3312), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4275 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n3407), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4276 ( .A1(n2978), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3267) );
  INV_X1 U4277 ( .A(n3273), .ZN(n3284) );
  AOI22_X1 U4278 ( .A1(n2978), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4279 ( .A1(n3400), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4280 ( .A1(n3407), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3274) );
  NAND4_X1 U4281 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3283)
         );
  AOI22_X1 U4282 ( .A1(n3298), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4283 ( .A1(n3465), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4284 ( .A1(n3372), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4285 ( .A1(n3303), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3278) );
  NAND4_X1 U4286 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3282)
         );
  OR2_X2 U4287 ( .A1(n3283), .A2(n3282), .ZN(n4250) );
  NAND2_X1 U4288 ( .A1(n3284), .A2(n3358), .ZN(n3285) );
  INV_X1 U4289 ( .A(n3342), .ZN(n3323) );
  AOI22_X1 U4290 ( .A1(n3465), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4291 ( .A1(n2977), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4292 ( .A1(n3400), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3287) );
  INV_X1 U4293 ( .A(n3312), .ZN(n3379) );
  AOI22_X1 U4294 ( .A1(n3291), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4295 ( .A1(n3303), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4296 ( .A1(n3470), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4297 ( .A1(n3421), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3292) );
  NAND2_X1 U4298 ( .A1(n3400), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3302) );
  NAND2_X1 U4299 ( .A1(n3465), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3301)
         );
  NAND2_X1 U4300 ( .A1(n3298), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3300) );
  NAND2_X1 U4301 ( .A1(n3407), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U4302 ( .A1(n2977), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3307)
         );
  NAND2_X1 U4303 ( .A1(n3303), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4304 ( .A1(n3470), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4305 ( .A1(n2983), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3304)
         );
  NAND2_X1 U4306 ( .A1(n3372), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3311)
         );
  NAND2_X1 U4307 ( .A1(n3373), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3309) );
  NAND2_X1 U4308 ( .A1(n3416), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4309 ( .A1(n3312), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U4310 ( .A1(n3313), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4311 ( .A1(n3314), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3315)
         );
  NAND2_X2 U4312 ( .A1(n3345), .A2(n4691), .ZN(n3346) );
  INV_X1 U4313 ( .A(n3986), .ZN(n3327) );
  AND2_X2 U4314 ( .A1(n3325), .A2(n3340), .ZN(n4464) );
  AOI21_X2 U4315 ( .B1(n3327), .B2(n4464), .A(n3326), .ZN(n3367) );
  INV_X1 U4316 ( .A(n3328), .ZN(n3329) );
  NAND2_X1 U4317 ( .A1(n3987), .A2(n4544), .ZN(n3331) );
  INV_X1 U4318 ( .A(n3368), .ZN(n3336) );
  NAND2_X1 U4319 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n4380) );
  OAI21_X1 U4320 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n4380), .ZN(n4166) );
  INV_X1 U4321 ( .A(n4166), .ZN(n3333) );
  NOR2_X1 U4322 ( .A1(n3332), .A2(n3333), .ZN(n3349) );
  NAND2_X1 U4323 ( .A1(n3345), .A2(n3332), .ZN(n4342) );
  OAI211_X1 U4324 ( .C1(n3349), .C2(n3324), .A(n4261), .B(n4342), .ZN(n3334)
         );
  INV_X1 U4325 ( .A(n4225), .ZN(n3462) );
  XNOR2_X1 U4326 ( .A(n6309), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6389)
         );
  NAND2_X1 U4327 ( .A1(n3462), .A2(n6389), .ZN(n3338) );
  INV_X1 U4328 ( .A(n3994), .ZN(n3461) );
  NAND2_X1 U4329 ( .A1(n3461), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U4330 ( .A1(n3338), .A2(n3337), .ZN(n3351) );
  NOR2_X1 U4331 ( .A1(n4223), .A2(n4537), .ZN(n3341) );
  INV_X1 U4332 ( .A(n3324), .ZN(n3343) );
  NAND2_X1 U4333 ( .A1(n5164), .A2(n3996), .ZN(n4536) );
  NOR2_X1 U4334 ( .A1(n3346), .A2(n4536), .ZN(n3348) );
  INV_X2 U4335 ( .A(n4250), .ZN(n4685) );
  INV_X1 U4336 ( .A(n4342), .ZN(n3355) );
  NAND2_X1 U4337 ( .A1(n3355), .A2(n4223), .ZN(n3356) );
  AND2_X2 U4338 ( .A1(n3357), .A2(n3356), .ZN(n3992) );
  NAND2_X1 U4339 ( .A1(n3358), .A2(n4464), .ZN(n3365) );
  NAND2_X1 U4340 ( .A1(n6049), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6574) );
  AOI21_X1 U4341 ( .B1(n4537), .B2(n4529), .A(n6574), .ZN(n3364) );
  NAND2_X1 U4342 ( .A1(n3360), .A2(n3359), .ZN(n3701) );
  INV_X1 U4343 ( .A(n3701), .ZN(n3363) );
  BUF_X1 U4344 ( .A(n3361), .Z(n3362) );
  NAND4_X1 U4345 ( .A1(n3363), .A2(n3362), .A3(n4679), .A4(n4685), .ZN(n4712)
         );
  AOI22_X1 U4346 ( .A1(n2961), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4347 ( .A1(n2973), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3377) );
  INV_X1 U4348 ( .A(n2984), .ZN(n3401) );
  AOI22_X1 U4349 ( .A1(n2978), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4350 ( .A1(n2976), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3375) );
  NAND4_X1 U4351 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3385)
         );
  INV_X1 U4352 ( .A(n2979), .ZN(n3772) );
  AOI22_X1 U4353 ( .A1(n3400), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3421), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4354 ( .A1(n4092), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4355 ( .A1(n3291), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4356 ( .A1(n3298), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3380) );
  NAND4_X1 U4357 ( .A1(n3383), .A2(n3382), .A3(n3381), .A4(n3380), .ZN(n3384)
         );
  NAND2_X1 U4358 ( .A1(n3066), .A2(n4259), .ZN(n3447) );
  XNOR2_X2 U4359 ( .A(n3388), .B(n3386), .ZN(n3433) );
  NAND2_X1 U4360 ( .A1(n3388), .A2(n3387), .ZN(n3390) );
  NAND2_X1 U4361 ( .A1(n3390), .A2(n3389), .ZN(n3392) );
  NAND2_X1 U4362 ( .A1(n3392), .A2(n3391), .ZN(n3399) );
  INV_X1 U4363 ( .A(n3399), .ZN(n3397) );
  NAND2_X1 U4364 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4365 ( .A1(n3393), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4366 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5972), .ZN(n6423) );
  OAI22_X1 U4367 ( .A1(n4225), .A2(n4791), .B1(n3994), .B2(n6547), .ZN(n3395)
         );
  AOI22_X1 U4368 ( .A1(n2973), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4369 ( .A1(n2979), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4370 ( .A1(n2984), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4371 ( .A1(n3291), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3403) );
  NAND4_X1 U4372 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3413)
         );
  AOI22_X1 U4373 ( .A1(n2961), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4374 ( .A1(n3489), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4375 ( .A1(n2978), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4377 ( .A1(n4092), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3408) );
  NAND4_X1 U4378 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(n3412)
         );
  NAND2_X1 U4379 ( .A1(n5978), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3706) );
  INV_X1 U4380 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4810) );
  AOI22_X1 U4381 ( .A1(n2973), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4382 ( .A1(n3489), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4383 ( .A1(n2978), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3373), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4384 ( .A1(n3400), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3417) );
  NAND4_X1 U4385 ( .A1(n3420), .A2(n3419), .A3(n3418), .A4(n3417), .ZN(n3427)
         );
  AOI22_X1 U4386 ( .A1(n2971), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4387 ( .A1(n3421), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4388 ( .A1(n2976), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2982), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4389 ( .A1(n3291), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3422) );
  NAND4_X1 U4390 ( .A1(n3425), .A2(n3424), .A3(n3423), .A4(n3422), .ZN(n3426)
         );
  NAND2_X1 U4391 ( .A1(n3428), .A2(n4260), .ZN(n3429) );
  OAI211_X1 U4392 ( .C1(n4810), .C2(n3963), .A(n3429), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3430) );
  NAND2_X1 U4393 ( .A1(n4662), .A2(n3362), .ZN(n3432) );
  NAND2_X1 U4394 ( .A1(n3432), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4476) );
  INV_X1 U4395 ( .A(n4536), .ZN(n3434) );
  NAND2_X1 U4396 ( .A1(n3434), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3506) );
  INV_X2 U4397 ( .A(n3032), .ZN(n3721) );
  NAND2_X1 U4398 ( .A1(n3721), .A2(EAX_REG_0__SCAN_IN), .ZN(n3436) );
  NAND2_X1 U4399 ( .A1(n5978), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3435)
         );
  OAI211_X1 U4400 ( .C1(n3506), .C2(n4457), .A(n3436), .B(n3435), .ZN(n3437)
         );
  AOI21_X1 U4401 ( .B1(n3433), .B2(n3685), .A(n3437), .ZN(n4477) );
  INV_X1 U4402 ( .A(n3819), .ZN(n3438) );
  NAND2_X1 U4403 ( .A1(n3440), .A2(n6566), .ZN(n3446) );
  INV_X1 U4404 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4806) );
  INV_X1 U4405 ( .A(n3441), .ZN(n3442) );
  NAND2_X1 U4406 ( .A1(n3442), .A2(n4259), .ZN(n3443) );
  INV_X1 U4407 ( .A(n3444), .ZN(n3445) );
  NAND2_X1 U4408 ( .A1(n3446), .A2(n3445), .ZN(n3448) );
  INV_X1 U4410 ( .A(n3685), .ZN(n3675) );
  OR2_X1 U4411 ( .A1(n5041), .A2(n3675), .ZN(n3450) );
  AOI22_X1 U4412 ( .A1(n3721), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5978), .ZN(n3449) );
  OAI211_X1 U4413 ( .C1(n3506), .C2(n5153), .A(n3450), .B(n3449), .ZN(n4336)
         );
  AND2_X2 U4414 ( .A1(n4335), .A2(n4336), .ZN(n4334) );
  NAND2_X1 U4415 ( .A1(n4490), .A2(n4334), .ZN(n3457) );
  INV_X1 U4416 ( .A(n3506), .ZN(n3451) );
  NAND2_X1 U4417 ( .A1(n3451), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3456) );
  INV_X1 U4418 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3453) );
  OAI21_X1 U4419 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3483), .ZN(n5384) );
  NAND2_X1 U4420 ( .A1(n3859), .A2(n5384), .ZN(n3452) );
  OAI21_X1 U4421 ( .B1(n3706), .B2(n3453), .A(n3452), .ZN(n3454) );
  AOI21_X1 U4422 ( .B1(n3721), .B2(EAX_REG_2__SCAN_IN), .A(n3454), .ZN(n3455)
         );
  NAND2_X1 U4423 ( .A1(n3457), .A2(n4492), .ZN(n3459) );
  OR2_X1 U4424 ( .A1(n4490), .A2(n4334), .ZN(n3458) );
  NAND2_X1 U4425 ( .A1(n3459), .A2(n3458), .ZN(n4489) );
  NAND2_X1 U4426 ( .A1(n3007), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3464) );
  NOR3_X1 U4427 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6547), .A3(n4916), 
        .ZN(n6353) );
  NAND2_X1 U4428 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6353), .ZN(n6350) );
  NAND2_X1 U4429 ( .A1(n6598), .A2(n6350), .ZN(n3460) );
  NAND3_X1 U4430 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4958) );
  INV_X1 U4431 ( .A(n4958), .ZN(n5001) );
  NAND2_X1 U4432 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5001), .ZN(n5039) );
  AOI22_X1 U4433 ( .A1(n3462), .A2(n6388), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3461), .ZN(n3463) );
  INV_X1 U4434 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6624) );
  AOI22_X1 U4435 ( .A1(n2973), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4436 ( .A1(n3489), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4437 ( .A1(n2978), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4438 ( .A1(n2979), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4439 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3476)
         );
  AOI22_X1 U4440 ( .A1(n2971), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4441 ( .A1(n4120), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4442 ( .A1(n2976), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4443 ( .A1(n3291), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3471) );
  NAND4_X1 U4444 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3475)
         );
  AOI22_X1 U4445 ( .A1(n3979), .A2(n4241), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3970), .ZN(n3477) );
  AND2_X1 U4446 ( .A1(n3478), .A2(n3477), .ZN(n4912) );
  NAND2_X1 U4447 ( .A1(n4912), .A2(n4246), .ZN(n3479) );
  INV_X1 U4448 ( .A(n3483), .ZN(n3485) );
  INV_X1 U4449 ( .A(n3503), .ZN(n3484) );
  OAI21_X1 U4450 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3485), .A(n3484), 
        .ZN(n5374) );
  AOI22_X1 U4451 ( .A1(n3859), .A2(n5374), .B1(n4135), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3487) );
  NAND2_X1 U4452 ( .A1(n3721), .A2(EAX_REG_3__SCAN_IN), .ZN(n3486) );
  OAI211_X1 U4453 ( .C1(n3506), .C2(n3481), .A(n3487), .B(n3486), .ZN(n3488)
         );
  NOR2_X2 U4454 ( .A1(n4489), .A2(n4622), .ZN(n4619) );
  AOI22_X1 U4455 ( .A1(n2973), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4456 ( .A1(n3489), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4457 ( .A1(n2978), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4458 ( .A1(n2979), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3490) );
  NAND4_X1 U4459 ( .A1(n3493), .A2(n3492), .A3(n3491), .A4(n3490), .ZN(n3499)
         );
  AOI22_X1 U4460 ( .A1(n2971), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U4461 ( .A1(n4120), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4462 ( .A1(n2976), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4463 ( .A1(n3291), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3494) );
  NAND4_X1 U4464 ( .A1(n3497), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n3498)
         );
  AOI22_X1 U4465 ( .A1(n3979), .A2(n4236), .B1(INSTQUEUE_REG_0__4__SCAN_IN), 
        .B2(n3970), .ZN(n3501) );
  OAI21_X1 U4466 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3503), .A(n3522), 
        .ZN(n6173) );
  OAI21_X1 U4467 ( .B1(n6059), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5978), 
        .ZN(n3505) );
  NAND2_X1 U4468 ( .A1(n3721), .A2(EAX_REG_4__SCAN_IN), .ZN(n3504) );
  OAI211_X1 U4469 ( .C1(n3506), .C2(n6053), .A(n3505), .B(n3504), .ZN(n3507)
         );
  OAI21_X1 U4470 ( .B1(n3819), .B2(n6173), .A(n3507), .ZN(n3508) );
  NAND2_X1 U4471 ( .A1(n4619), .A2(n4621), .ZN(n4620) );
  INV_X1 U4472 ( .A(n4620), .ZN(n3529) );
  AOI22_X1 U4473 ( .A1(n2973), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4474 ( .A1(n3489), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4475 ( .A1(n2978), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3511) );
  INV_X1 U4476 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6672) );
  AOI22_X1 U4477 ( .A1(n2979), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3510) );
  NAND4_X1 U4478 ( .A1(n3513), .A2(n3512), .A3(n3511), .A4(n3510), .ZN(n3519)
         );
  AOI22_X1 U4479 ( .A1(n2971), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4480 ( .A1(n4120), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4481 ( .A1(n2976), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n2982), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4482 ( .A1(n3291), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3514) );
  NAND4_X1 U4483 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3518)
         );
  NAND2_X1 U4484 ( .A1(n3979), .A2(n4283), .ZN(n3521) );
  NAND2_X1 U4485 ( .A1(n3970), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4486 ( .A1(n3521), .A2(n3520), .ZN(n3531) );
  INV_X1 U4487 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3526) );
  INV_X1 U4488 ( .A(n3522), .ZN(n3524) );
  INV_X1 U4489 ( .A(n3544), .ZN(n3523) );
  OAI21_X1 U4490 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3524), .A(n3523), 
        .ZN(n6162) );
  AOI22_X1 U4491 ( .A1(n3438), .A2(n6162), .B1(n4135), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3525) );
  OAI21_X1 U4492 ( .B1(n3032), .B2(n3526), .A(n3525), .ZN(n3527) );
  AOI21_X1 U4493 ( .B1(n4273), .B2(n3685), .A(n3527), .ZN(n4648) );
  NAND2_X1 U4494 ( .A1(n3529), .A2(n3528), .ZN(n4647) );
  INV_X1 U4495 ( .A(n4647), .ZN(n3549) );
  INV_X1 U4496 ( .A(n3530), .ZN(n3532) );
  NAND2_X1 U4497 ( .A1(n3532), .A2(n3531), .ZN(n3550) );
  AOI22_X1 U4498 ( .A1(n2973), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4499 ( .A1(n2978), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4500 ( .A1(n2961), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4501 ( .A1(n2971), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3533) );
  NAND4_X1 U4502 ( .A1(n3536), .A2(n3535), .A3(n3534), .A4(n3533), .ZN(n3543)
         );
  AOI22_X1 U4503 ( .A1(n2979), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4504 ( .A1(n2976), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4505 ( .A1(n4121), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4506 ( .A1(n4119), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3538) );
  NAND4_X1 U4507 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3542)
         );
  AOI22_X1 U4508 ( .A1(n3979), .A2(n4286), .B1(n3970), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U4509 ( .A1(n3550), .A2(n3551), .ZN(n4282) );
  OAI21_X1 U4510 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n3544), .A(n3567), 
        .ZN(n6156) );
  INV_X1 U4511 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3545) );
  INV_X1 U4512 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6659) );
  OAI22_X1 U4513 ( .A1(n3032), .A2(n3545), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6659), .ZN(n3546) );
  MUX2_X1 U4514 ( .A(n6156), .B(n3546), .S(n3819), .Z(n3547) );
  NAND2_X1 U4515 ( .A1(n3549), .A2(n3548), .ZN(n4831) );
  INV_X1 U4516 ( .A(n4831), .ZN(n3574) );
  INV_X1 U4517 ( .A(n3550), .ZN(n3553) );
  INV_X1 U4518 ( .A(n3551), .ZN(n3552) );
  AOI22_X1 U4519 ( .A1(n2978), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4520 ( .A1(n4120), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4521 ( .A1(n2973), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4522 ( .A1(n2984), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3554) );
  NAND4_X1 U4523 ( .A1(n3557), .A2(n3556), .A3(n3555), .A4(n3554), .ZN(n3563)
         );
  AOI22_X1 U4524 ( .A1(n3489), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4525 ( .A1(n2979), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4526 ( .A1(n2976), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4527 ( .A1(n2971), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4528 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3562)
         );
  NAND2_X1 U4529 ( .A1(n3979), .A2(n4304), .ZN(n3565) );
  NAND2_X1 U4530 ( .A1(n3970), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3564) );
  NAND2_X1 U4531 ( .A1(n3565), .A2(n3564), .ZN(n3566) );
  INV_X1 U4532 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3571) );
  INV_X1 U4533 ( .A(n3567), .ZN(n3569) );
  INV_X1 U4534 ( .A(n3588), .ZN(n3568) );
  OAI21_X1 U4535 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3569), .A(n3568), 
        .ZN(n6255) );
  AOI22_X1 U4536 ( .A1(n3438), .A2(n6255), .B1(n4135), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3570) );
  OAI21_X1 U4537 ( .B1(n3032), .B2(n3571), .A(n3570), .ZN(n3572) );
  AOI21_X1 U4538 ( .B1(n4293), .B2(n3685), .A(n3572), .ZN(n4905) );
  INV_X1 U4539 ( .A(n4905), .ZN(n3573) );
  NAND2_X1 U4540 ( .A1(n3574), .A2(n3573), .ZN(n4903) );
  AOI22_X1 U4541 ( .A1(n2973), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4542 ( .A1(n4121), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4543 ( .A1(n4120), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4544 ( .A1(n2979), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3575) );
  NAND4_X1 U4545 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(n3584)
         );
  AOI22_X1 U4546 ( .A1(n2961), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4547 ( .A1(n2978), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4548 ( .A1(n2976), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n2982), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4549 ( .A1(n2971), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4550 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3583)
         );
  OAI21_X1 U4551 ( .B1(n3584), .B2(n3583), .A(n3685), .ZN(n3587) );
  NAND2_X1 U4552 ( .A1(n3721), .A2(EAX_REG_8__SCAN_IN), .ZN(n3586) );
  XNOR2_X1 U4553 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3588), .ZN(n6121) );
  AOI22_X1 U4554 ( .A1(n3859), .A2(n6121), .B1(n4135), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3585) );
  XOR2_X1 U4555 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3603), .Z(n6112) );
  AOI22_X1 U4556 ( .A1(n2973), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4557 ( .A1(n2978), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4558 ( .A1(n2971), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4559 ( .A1(n2976), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3589) );
  NAND4_X1 U4560 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3599)
         );
  AOI22_X1 U4561 ( .A1(n3489), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4562 ( .A1(n2961), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4563 ( .A1(n2979), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4564 ( .A1(n2984), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3594) );
  NAND4_X1 U4565 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .ZN(n3598)
         );
  OR2_X1 U4566 ( .A1(n3599), .A2(n3598), .ZN(n3600) );
  AOI22_X1 U4567 ( .A1(n3685), .A2(n3600), .B1(n4135), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3602) );
  NAND2_X1 U4568 ( .A1(n3721), .A2(EAX_REG_9__SCAN_IN), .ZN(n3601) );
  OAI211_X1 U4569 ( .C1(n6112), .C2(n3819), .A(n3602), .B(n3601), .ZN(n5121)
         );
  INV_X1 U4570 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3604) );
  XNOR2_X1 U4571 ( .A(n3619), .B(n3604), .ZN(n5669) );
  AOI22_X1 U4572 ( .A1(n2973), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4573 ( .A1(n4119), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4574 ( .A1(n2961), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4575 ( .A1(n2976), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3605) );
  NAND4_X1 U4576 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(n3614)
         );
  AOI22_X1 U4577 ( .A1(n2978), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4578 ( .A1(n2971), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4579 ( .A1(n4120), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4580 ( .A1(n3291), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3609) );
  NAND4_X1 U4581 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3613)
         );
  OAI21_X1 U4582 ( .B1(n3614), .B2(n3613), .A(n3685), .ZN(n3617) );
  NAND2_X1 U4583 ( .A1(n3721), .A2(EAX_REG_10__SCAN_IN), .ZN(n3616) );
  NAND2_X1 U4584 ( .A1(n4135), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3615)
         );
  NAND3_X1 U4585 ( .A1(n3617), .A2(n3616), .A3(n3615), .ZN(n3618) );
  AOI21_X1 U4586 ( .B1(n5669), .B2(n3859), .A(n3618), .ZN(n5359) );
  XNOR2_X1 U4587 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3634), .ZN(n6249)
         );
  INV_X1 U4588 ( .A(n6249), .ZN(n5345) );
  AOI22_X1 U4589 ( .A1(n2978), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4590 ( .A1(n2973), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4591 ( .A1(n4120), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4592 ( .A1(n2979), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3620) );
  NAND4_X1 U4593 ( .A1(n3623), .A2(n3622), .A3(n3621), .A4(n3620), .ZN(n3629)
         );
  AOI22_X1 U4594 ( .A1(n4119), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4595 ( .A1(n2961), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4596 ( .A1(n2983), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4597 ( .A1(n2971), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3624) );
  NAND4_X1 U4598 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n3628)
         );
  OAI21_X1 U4599 ( .B1(n3629), .B2(n3628), .A(n3685), .ZN(n3632) );
  NAND2_X1 U4600 ( .A1(n3721), .A2(EAX_REG_11__SCAN_IN), .ZN(n3631) );
  NAND2_X1 U4601 ( .A1(n4135), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3630)
         );
  NAND3_X1 U4602 ( .A1(n3632), .A2(n3631), .A3(n3630), .ZN(n3633) );
  AOI21_X1 U4603 ( .B1(n5345), .B2(n3438), .A(n3633), .ZN(n5343) );
  XNOR2_X1 U4604 ( .A(n3035), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5658)
         );
  AOI21_X1 U4605 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3112), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3636) );
  AND2_X1 U4606 ( .A1(n3721), .A2(EAX_REG_12__SCAN_IN), .ZN(n3635) );
  OAI22_X1 U4607 ( .A1(n5658), .A2(n3819), .B1(n3636), .B2(n3635), .ZN(n3648)
         );
  AOI22_X1 U4608 ( .A1(n2973), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4609 ( .A1(n2961), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4610 ( .A1(n2976), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4611 ( .A1(n4121), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3637) );
  NAND4_X1 U4612 ( .A1(n3640), .A2(n3639), .A3(n3638), .A4(n3637), .ZN(n3646)
         );
  AOI22_X1 U4613 ( .A1(n3489), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4614 ( .A1(n2971), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4615 ( .A1(n2978), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4616 ( .A1(n4120), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3641) );
  NAND4_X1 U4617 ( .A1(n3644), .A2(n3643), .A3(n3642), .A4(n3641), .ZN(n3645)
         );
  OAI21_X1 U4618 ( .B1(n3646), .B2(n3645), .A(n3685), .ZN(n3647) );
  NAND2_X1 U4619 ( .A1(n3648), .A2(n3647), .ZN(n5332) );
  XNOR2_X1 U4620 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3672), .ZN(n5648)
         );
  AOI22_X1 U4621 ( .A1(n2973), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4622 ( .A1(n2971), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4623 ( .A1(n2978), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4624 ( .A1(n4119), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3649) );
  NAND4_X1 U4625 ( .A1(n3652), .A2(n3651), .A3(n3650), .A4(n3649), .ZN(n3658)
         );
  AOI22_X1 U4626 ( .A1(n2979), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4627 ( .A1(n4120), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4628 ( .A1(n2976), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4629 ( .A1(n4092), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3653) );
  NAND4_X1 U4630 ( .A1(n3656), .A2(n3655), .A3(n3654), .A4(n3653), .ZN(n3657)
         );
  OR2_X1 U4631 ( .A1(n3658), .A2(n3657), .ZN(n3659) );
  AOI22_X1 U4632 ( .A1(n3685), .A2(n3659), .B1(n4135), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U4633 ( .A1(n3721), .A2(EAX_REG_13__SCAN_IN), .ZN(n3660) );
  OAI211_X1 U4634 ( .C1(n5648), .C2(n3819), .A(n3661), .B(n3660), .ZN(n5317)
         );
  AOI22_X1 U4635 ( .A1(n3489), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4636 ( .A1(n2978), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4637 ( .A1(n2976), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4638 ( .A1(n2971), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4639 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3671)
         );
  AOI22_X1 U4640 ( .A1(n2973), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4641 ( .A1(n2984), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4642 ( .A1(n3312), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n2982), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4643 ( .A1(n2961), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4644 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3670)
         );
  NOR2_X1 U4645 ( .A1(n3671), .A2(n3670), .ZN(n3676) );
  XNOR2_X1 U4646 ( .A(n3688), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5639)
         );
  NAND2_X1 U4647 ( .A1(n5639), .A2(n3859), .ZN(n3674) );
  AOI22_X1 U4648 ( .A1(n3721), .A2(EAX_REG_14__SCAN_IN), .B1(n4135), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3673) );
  OAI211_X1 U4649 ( .C1(n3676), .C2(n3675), .A(n3674), .B(n3673), .ZN(n5305)
         );
  NAND2_X1 U4650 ( .A1(n5302), .A2(n5305), .ZN(n5303) );
  AOI22_X1 U4651 ( .A1(n2978), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4652 ( .A1(n2961), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4653 ( .A1(n2984), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4654 ( .A1(n3407), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3677) );
  NAND4_X1 U4655 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(n3687)
         );
  AOI22_X1 U4656 ( .A1(n2973), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4657 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4120), .B1(n4119), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4658 ( .A1(n2979), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4659 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n2976), .B1(n2982), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3681) );
  NAND4_X1 U4660 ( .A1(n3684), .A2(n3683), .A3(n3682), .A4(n3681), .ZN(n3686)
         );
  OAI21_X1 U4661 ( .B1(n3687), .B2(n3686), .A(n3685), .ZN(n3691) );
  NAND2_X1 U4662 ( .A1(n3721), .A2(EAX_REG_15__SCAN_IN), .ZN(n3690) );
  XNOR2_X1 U4663 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3704), .ZN(n5633)
         );
  INV_X1 U4664 ( .A(n5633), .ZN(n6094) );
  AOI22_X1 U4665 ( .A1(n4135), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n3859), 
        .B2(n6094), .ZN(n3689) );
  AOI22_X1 U4666 ( .A1(n2978), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4667 ( .A1(n4119), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4668 ( .A1(n3407), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4669 ( .A1(n4121), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3693) );
  NAND4_X1 U4670 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3703)
         );
  AOI22_X1 U4671 ( .A1(n2961), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4672 ( .A1(n2976), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4673 ( .A1(n2973), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4674 ( .A1(n4120), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3697) );
  NAND4_X1 U4675 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3702)
         );
  OAI21_X1 U4676 ( .B1(n3703), .B2(n3702), .A(n4132), .ZN(n3709) );
  INV_X1 U4677 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5625) );
  XNOR2_X1 U4678 ( .A(n3724), .B(n5625), .ZN(n5629) );
  OAI22_X1 U4679 ( .A1(n5629), .A2(n3819), .B1(n3706), .B2(n5625), .ZN(n3707)
         );
  AOI21_X1 U4680 ( .B1(n3721), .B2(EAX_REG_16__SCAN_IN), .A(n3707), .ZN(n3708)
         );
  AOI22_X1 U4681 ( .A1(n2973), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4682 ( .A1(n2961), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4683 ( .A1(n2979), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4684 ( .A1(n2978), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3710) );
  NAND4_X1 U4685 ( .A1(n3713), .A2(n3712), .A3(n3711), .A4(n3710), .ZN(n3719)
         );
  AOI22_X1 U4686 ( .A1(n2976), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4687 ( .A1(n2971), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4688 ( .A1(n4120), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4689 ( .A1(n3407), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3714) );
  NAND4_X1 U4690 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3718)
         );
  NOR2_X1 U4691 ( .A1(n3719), .A2(n3718), .ZN(n3723) );
  NOR2_X1 U4692 ( .A1(n3725), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3720) );
  AOI21_X1 U4693 ( .B1(n3721), .B2(EAX_REG_17__SCAN_IN), .A(n3720), .ZN(n3722)
         );
  OAI21_X1 U4694 ( .B1(n4106), .B2(n3723), .A(n3722), .ZN(n3728) );
  AND2_X1 U4695 ( .A1(n3726), .A2(n3725), .ZN(n3727) );
  OR2_X1 U4696 ( .A1(n3727), .A2(n3033), .ZN(n6086) );
  MUX2_X1 U4697 ( .A(n3728), .B(n6086), .S(n3859), .Z(n5430) );
  NAND2_X1 U4698 ( .A1(n4106), .A2(n3819), .ZN(n3763) );
  AOI22_X1 U4699 ( .A1(n2979), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4700 ( .A1(n2978), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4701 ( .A1(n2984), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3732) );
  AOI21_X1 U4702 ( .B1(n2957), .B2(INSTQUEUE_REG_9__2__SCAN_IN), .A(n3859), 
        .ZN(n3730) );
  NAND2_X1 U4703 ( .A1(n2963), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3729)
         );
  AND2_X1 U4704 ( .A1(n3730), .A2(n3729), .ZN(n3731) );
  NAND4_X1 U4705 ( .A1(n3734), .A2(n3733), .A3(n3732), .A4(n3731), .ZN(n3740)
         );
  AOI22_X1 U4706 ( .A1(n2961), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4707 ( .A1(n2973), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4708 ( .A1(n2971), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4709 ( .A1(n4121), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3735) );
  NAND4_X1 U4710 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(n3739)
         );
  OR2_X1 U4711 ( .A1(n3740), .A2(n3739), .ZN(n3741) );
  NAND2_X1 U4712 ( .A1(n3763), .A2(n3741), .ZN(n3744) );
  AOI22_X1 U4713 ( .A1(n3721), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5978), .ZN(n3743) );
  XNOR2_X1 U4714 ( .A(n3033), .B(n3108), .ZN(n6075) );
  AND2_X1 U4715 ( .A1(n6075), .A2(n3438), .ZN(n3742) );
  NAND2_X1 U4716 ( .A1(n3745), .A2(n5594), .ZN(n3746) );
  NAND2_X1 U4717 ( .A1(n3762), .A2(n3746), .ZN(n6022) );
  INV_X1 U4718 ( .A(n6022), .ZN(n5596) );
  AOI22_X1 U4719 ( .A1(n3489), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4720 ( .A1(n2976), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4721 ( .A1(n2979), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4722 ( .A1(n2961), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3747) );
  NAND4_X1 U4723 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3756)
         );
  AOI22_X1 U4724 ( .A1(n2978), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4725 ( .A1(n2973), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4726 ( .A1(n4092), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2982), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4727 ( .A1(n4121), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3751) );
  NAND4_X1 U4728 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(n3755)
         );
  OR2_X1 U4729 ( .A1(n3756), .A2(n3755), .ZN(n3759) );
  INV_X1 U4730 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3757) );
  OAI22_X1 U4731 ( .A1(n3032), .A2(n3757), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5594), .ZN(n3758) );
  AOI21_X1 U4732 ( .B1(n4132), .B2(n3759), .A(n3758), .ZN(n3760) );
  MUX2_X1 U4733 ( .A(n5596), .B(n3760), .S(n3819), .Z(n5414) );
  XNOR2_X1 U4734 ( .A(n3794), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5590)
         );
  INV_X1 U4735 ( .A(n3763), .ZN(n3817) );
  AOI22_X1 U4736 ( .A1(n2961), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4737 ( .A1(n2976), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4738 ( .A1(n4119), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4739 ( .A1(n3312), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4740 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3778)
         );
  INV_X1 U4741 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4742 ( .A1(n2978), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3769) );
  AOI21_X1 U4743 ( .B1(n3416), .B2(INSTQUEUE_REG_9__4__SCAN_IN), .A(n3859), 
        .ZN(n3768) );
  OAI211_X1 U4744 ( .C1(n3374), .C2(n3770), .A(n3769), .B(n3768), .ZN(n3777)
         );
  INV_X1 U4745 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3773) );
  INV_X1 U4746 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3771) );
  OAI22_X1 U4747 ( .A1(n3808), .A2(n3773), .B1(n3772), .B2(n3771), .ZN(n3776)
         );
  INV_X1 U4748 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3774) );
  INV_X1 U4749 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5952) );
  OAI22_X1 U4750 ( .A1(n3401), .A2(n3774), .B1(n3593), .B2(n5952), .ZN(n3775)
         );
  NOR4_X1 U4751 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3780)
         );
  AOI22_X1 U4752 ( .A1(n3721), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5978), .ZN(n3779) );
  OAI21_X1 U4753 ( .B1(n3817), .B2(n3780), .A(n3779), .ZN(n3781) );
  OAI21_X1 U4754 ( .B1(n3819), .B2(n5590), .A(n3781), .ZN(n5280) );
  AOI22_X1 U4755 ( .A1(n2978), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4756 ( .A1(n2979), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4757 ( .A1(n2961), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4758 ( .A1(n2971), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3782) );
  NAND4_X1 U4759 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3791)
         );
  AOI22_X1 U4760 ( .A1(n2973), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4761 ( .A1(n4119), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4762 ( .A1(n2984), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4763 ( .A1(n4121), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4764 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3790)
         );
  OAI21_X1 U4765 ( .B1(n3791), .B2(n3790), .A(n4132), .ZN(n3793) );
  AOI22_X1 U4766 ( .A1(n3721), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5978), .ZN(n3792) );
  NAND2_X1 U4767 ( .A1(n3793), .A2(n3792), .ZN(n3797) );
  NAND2_X1 U4768 ( .A1(n3795), .A2(n5274), .ZN(n3796) );
  NAND2_X1 U4769 ( .A1(n3798), .A2(n3796), .ZN(n5581) );
  MUX2_X1 U4770 ( .A(n3797), .B(n5581), .S(n3859), .Z(n5269) );
  XNOR2_X1 U4771 ( .A(n3842), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5574)
         );
  AOI22_X1 U4772 ( .A1(n2979), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4773 ( .A1(n4119), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4774 ( .A1(n4120), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4775 ( .A1(n2978), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3799) );
  NAND4_X1 U4776 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n3814)
         );
  INV_X1 U4777 ( .A(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4778 ( .A1(n4092), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3804) );
  AOI21_X1 U4779 ( .B1(n2957), .B2(INSTQUEUE_REG_9__6__SCAN_IN), .A(n3859), 
        .ZN(n3803) );
  OAI211_X1 U4780 ( .C1(n3379), .C2(n3805), .A(n3804), .B(n3803), .ZN(n3813)
         );
  INV_X1 U4781 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3807) );
  INV_X1 U4782 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3806) );
  OAI22_X1 U4783 ( .A1(n3808), .A2(n3807), .B1(n2958), .B2(n3806), .ZN(n3812)
         );
  INV_X1 U4784 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3809) );
  INV_X1 U4785 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5960) );
  OAI22_X1 U4786 ( .A1(n3810), .A2(n3809), .B1(n3593), .B2(n5960), .ZN(n3811)
         );
  NOR4_X1 U4787 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3816)
         );
  AOI22_X1 U4788 ( .A1(n3721), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5978), .ZN(n3815) );
  OAI21_X1 U4789 ( .B1(n3817), .B2(n3816), .A(n3815), .ZN(n3818) );
  OAI21_X1 U4790 ( .B1(n3819), .B2(n5574), .A(n3818), .ZN(n5259) );
  AOI22_X1 U4791 ( .A1(n2978), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4792 ( .A1(n2971), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4793 ( .A1(n4120), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4794 ( .A1(n2973), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4795 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4796 ( .A1(n2979), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4797 ( .A1(n4119), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4798 ( .A1(n2976), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4799 ( .A1(n3291), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4800 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  NOR2_X1 U4801 ( .A1(n3829), .A2(n3828), .ZN(n3846) );
  AOI22_X1 U4802 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n2979), .B1(n2961), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4803 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n2978), .B1(n2984), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4804 ( .A1(n4120), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4805 ( .A1(n4121), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4806 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3839)
         );
  AOI22_X1 U4807 ( .A1(n2973), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4808 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n2971), .B1(n4092), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4809 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n2976), .B1(n3537), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4810 ( .A1(n4119), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4811 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3838)
         );
  NOR2_X1 U4812 ( .A1(n3839), .A2(n3838), .ZN(n3847) );
  XNOR2_X1 U4813 ( .A(n3846), .B(n3847), .ZN(n3841) );
  AOI22_X1 U4814 ( .A1(n3721), .A2(EAX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5978), .ZN(n3840) );
  OAI21_X1 U4815 ( .B1(n4106), .B2(n3841), .A(n3840), .ZN(n3845) );
  INV_X1 U4816 ( .A(n3843), .ZN(n3844) );
  OAI21_X1 U4817 ( .B1(n3844), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n3878), 
        .ZN(n5555) );
  MUX2_X1 U4818 ( .A(n3845), .B(n5555), .S(n3438), .Z(n5245) );
  OR2_X1 U4819 ( .A1(n3847), .A2(n3846), .ZN(n3875) );
  INV_X1 U4820 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U4821 ( .A1(n2961), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4822 ( .A1(n3312), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4823 ( .A1(n2971), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4824 ( .A1(n3489), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4825 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3858)
         );
  AOI22_X1 U4826 ( .A1(n2979), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4827 ( .A1(n2973), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4828 ( .A1(n2978), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4829 ( .A1(n2976), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4830 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3857)
         );
  NOR2_X1 U4831 ( .A1(n3858), .A2(n3857), .ZN(n3874) );
  XNOR2_X1 U4832 ( .A(n3875), .B(n3874), .ZN(n3862) );
  AOI22_X1 U4833 ( .A1(n3721), .A2(EAX_REG_24__SCAN_IN), .B1(n4135), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3861) );
  XNOR2_X1 U4834 ( .A(n3878), .B(n5241), .ZN(n5550) );
  NAND2_X1 U4835 ( .A1(n5550), .A2(n3859), .ZN(n3860) );
  OAI211_X1 U4836 ( .C1(n3862), .C2(n4106), .A(n3861), .B(n3860), .ZN(n3863)
         );
  AOI22_X1 U4837 ( .A1(n2973), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4838 ( .A1(n3489), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4839 ( .A1(n2978), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4840 ( .A1(n2979), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3864) );
  NAND4_X1 U4841 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(n3873)
         );
  AOI22_X1 U4842 ( .A1(n2971), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4843 ( .A1(n4120), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4844 ( .A1(n2976), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n2982), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4845 ( .A1(n4121), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3868) );
  NAND4_X1 U4846 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3872)
         );
  NOR2_X1 U4847 ( .A1(n3873), .A2(n3872), .ZN(n3895) );
  XNOR2_X1 U4848 ( .A(n3895), .B(n3894), .ZN(n3877) );
  AOI22_X1 U4849 ( .A1(n3721), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5978), .ZN(n3876) );
  OAI21_X1 U4850 ( .B1(n3877), .B2(n4106), .A(n3876), .ZN(n3883) );
  INV_X1 U4851 ( .A(n3879), .ZN(n3881) );
  INV_X1 U4852 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3880) );
  NAND2_X1 U4853 ( .A1(n3881), .A2(n3880), .ZN(n3882) );
  NAND2_X1 U4854 ( .A1(n3914), .A2(n3882), .ZN(n5539) );
  MUX2_X1 U4855 ( .A(n3883), .B(n5539), .S(n3859), .Z(n5223) );
  AOI22_X1 U4856 ( .A1(n2971), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4857 ( .A1(n4120), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4858 ( .A1(n2976), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4859 ( .A1(n3312), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3884) );
  NAND4_X1 U4860 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3893)
         );
  AOI22_X1 U4861 ( .A1(n2973), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4862 ( .A1(n3489), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4863 ( .A1(n2978), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4864 ( .A1(n2979), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3888) );
  NAND4_X1 U4865 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3892)
         );
  NOR2_X1 U4866 ( .A1(n3895), .A2(n3894), .ZN(n3901) );
  XOR2_X1 U4867 ( .A(n3900), .B(n3901), .Z(n3898) );
  INV_X1 U4868 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3896) );
  INV_X1 U4869 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5528) );
  OAI22_X1 U4870 ( .A1(n3032), .A2(n3896), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5528), .ZN(n3897) );
  AOI21_X1 U4871 ( .B1(n3898), .B2(n4132), .A(n3897), .ZN(n3899) );
  XNOR2_X1 U4872 ( .A(n3914), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5526)
         );
  MUX2_X1 U4873 ( .A(n3899), .B(n5526), .S(n3859), .Z(n5211) );
  NAND2_X1 U4874 ( .A1(n3901), .A2(n3900), .ZN(n3927) );
  AOI22_X1 U4875 ( .A1(n2973), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4876 ( .A1(n3489), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4877 ( .A1(n2971), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4878 ( .A1(n2979), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4879 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3911)
         );
  AOI22_X1 U4880 ( .A1(n2978), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4881 ( .A1(n2976), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4882 ( .A1(n4120), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4883 ( .A1(n3312), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4884 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3910)
         );
  NOR2_X1 U4885 ( .A1(n3911), .A2(n3910), .ZN(n3928) );
  XNOR2_X1 U4886 ( .A(n3927), .B(n3928), .ZN(n3913) );
  AOI22_X1 U4887 ( .A1(n3721), .A2(EAX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5978), .ZN(n3912) );
  OAI21_X1 U4888 ( .B1(n3913), .B2(n4106), .A(n3912), .ZN(n3916) );
  NOR2_X1 U4889 ( .A1(n3914), .A2(n5528), .ZN(n3915) );
  INV_X1 U4890 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5203) );
  OAI21_X1 U4891 ( .B1(n3915), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n3931), 
        .ZN(n5513) );
  MUX2_X1 U4892 ( .A(n3916), .B(n5513), .S(n3438), .Z(n5198) );
  AOI22_X1 U4893 ( .A1(n2973), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4894 ( .A1(n3489), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4895 ( .A1(n2978), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4896 ( .A1(n2979), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4897 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3926)
         );
  AOI22_X1 U4898 ( .A1(n2971), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4899 ( .A1(n3421), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4900 ( .A1(n2976), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4901 ( .A1(n4121), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3921) );
  NAND4_X1 U4902 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3925)
         );
  OR2_X1 U4903 ( .A1(n3926), .A2(n3925), .ZN(n4103) );
  NOR2_X1 U4904 ( .A1(n3928), .A2(n3927), .ZN(n4104) );
  XOR2_X1 U4905 ( .A(n4103), .B(n4104), .Z(n3930) );
  INV_X1 U4906 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4496) );
  OAI22_X1 U4907 ( .A1(n3032), .A2(n4496), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6678), .ZN(n3929) );
  AOI21_X1 U4908 ( .B1(n3930), .B2(n4132), .A(n3929), .ZN(n3932) );
  AOI21_X1 U4909 ( .B1(n6678), .B2(n3931), .A(n4108), .ZN(n5509) );
  MUX2_X1 U4910 ( .A(n3932), .B(n5509), .S(n3859), .Z(n3934) );
  XNOR2_X1 U4911 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3945) );
  NAND2_X1 U4912 ( .A1(n4691), .A2(n3324), .ZN(n3937) );
  NAND2_X1 U4913 ( .A1(n3346), .A2(n3937), .ZN(n3956) );
  OR2_X1 U4914 ( .A1(n3938), .A2(n3956), .ZN(n3946) );
  INV_X1 U4915 ( .A(n3941), .ZN(n3940) );
  INV_X1 U4916 ( .A(n3942), .ZN(n3939) );
  NAND2_X1 U4917 ( .A1(n3940), .A2(n3939), .ZN(n3943) );
  NAND2_X1 U4918 ( .A1(n3942), .A2(n3941), .ZN(n3951) );
  AND2_X1 U4919 ( .A1(n3943), .A2(n3951), .ZN(n4140) );
  NAND3_X1 U4920 ( .A1(n3947), .A2(STATE2_REG_0__SCAN_IN), .A3(n4140), .ZN(
        n3948) );
  NAND2_X1 U4921 ( .A1(n4916), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3950) );
  NAND2_X1 U4922 ( .A1(n3951), .A2(n3950), .ZN(n3959) );
  XNOR2_X1 U4923 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3958) );
  INV_X1 U4924 ( .A(n3958), .ZN(n3952) );
  XNOR2_X1 U4925 ( .A(n3959), .B(n3952), .ZN(n4139) );
  NAND2_X1 U4926 ( .A1(n3979), .A2(n4139), .ZN(n3955) );
  INV_X1 U4927 ( .A(n3956), .ZN(n3953) );
  OAI211_X1 U4928 ( .C1(n4139), .C2(n3963), .A(n3955), .B(n3953), .ZN(n3954)
         );
  INV_X1 U4929 ( .A(n3955), .ZN(n3957) );
  NAND2_X1 U4930 ( .A1(n3957), .A2(n3956), .ZN(n3964) );
  NAND2_X1 U4931 ( .A1(n3959), .A2(n3958), .ZN(n3961) );
  NAND2_X1 U4932 ( .A1(n6547), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3960) );
  XNOR2_X1 U4933 ( .A(n3967), .B(n3965), .ZN(n4141) );
  INV_X1 U4934 ( .A(n4141), .ZN(n3962) );
  INV_X1 U4935 ( .A(n3965), .ZN(n3966) );
  NAND2_X1 U4936 ( .A1(n3967), .A2(n3966), .ZN(n3969) );
  NAND2_X1 U4937 ( .A1(n6598), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3968) );
  NAND2_X1 U4938 ( .A1(n3969), .A2(n3968), .ZN(n3973) );
  INV_X1 U4939 ( .A(n3976), .ZN(n3971) );
  AOI22_X1 U4940 ( .A1(n3971), .A2(n3102), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6566), .ZN(n3977) );
  NAND2_X1 U4941 ( .A1(n6053), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3974) );
  INV_X1 U4942 ( .A(n4143), .ZN(n3978) );
  NOR2_X1 U4943 ( .A1(n4342), .A2(n4529), .ZN(n4425) );
  OAI21_X1 U4944 ( .B1(n4425), .B2(n4629), .A(n3982), .ZN(n3984) );
  OAI21_X1 U4945 ( .B1(n4536), .B2(n4537), .A(n4529), .ZN(n3983) );
  OAI211_X1 U4946 ( .C1(n3980), .C2(n2975), .A(n3984), .B(n3983), .ZN(n3990)
         );
  NAND2_X1 U4947 ( .A1(n3987), .A2(n4537), .ZN(n3985) );
  OR2_X1 U4948 ( .A1(n3986), .A2(n3985), .ZN(n3989) );
  INV_X1 U4949 ( .A(n3987), .ZN(n4481) );
  NAND2_X1 U4950 ( .A1(n4481), .A2(n4464), .ZN(n3988) );
  NAND2_X1 U4951 ( .A1(n3989), .A2(n3988), .ZN(n4420) );
  NOR2_X1 U4952 ( .A1(n3990), .A2(n4420), .ZN(n3991) );
  NAND2_X1 U4953 ( .A1(n3992), .A2(n3991), .ZN(n4443) );
  OAI21_X1 U4954 ( .B1(n4440), .B2(n4537), .A(n4712), .ZN(n3993) );
  NOR2_X1 U4955 ( .A1(n5142), .A2(n4691), .ZN(n4527) );
  NAND2_X1 U4956 ( .A1(n4547), .A2(n4527), .ZN(n4445) );
  NOR2_X1 U4957 ( .A1(n4445), .A2(n6573), .ZN(n3995) );
  NAND2_X1 U4958 ( .A1(n4528), .A2(n3995), .ZN(n4000) );
  NAND2_X1 U4959 ( .A1(n3996), .A2(n5170), .ZN(n3997) );
  NAND3_X1 U4960 ( .A1(n4438), .A2(n3721), .A3(n3998), .ZN(n4215) );
  OR2_X1 U4961 ( .A1(n4215), .A2(n2959), .ZN(n3999) );
  NAND2_X2 U4962 ( .A1(n3003), .A2(n4001), .ZN(n4085) );
  INV_X1 U4963 ( .A(n4005), .ZN(n4002) );
  NAND2_X1 U4964 ( .A1(n2960), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4003)
         );
  NAND2_X1 U4965 ( .A1(n4005), .A2(EBX_REG_0__SCAN_IN), .ZN(n4007) );
  INV_X1 U4966 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U4967 ( .A1(n2975), .A2(n4632), .ZN(n4006) );
  NAND2_X1 U4968 ( .A1(n4007), .A2(n4006), .ZN(n4630) );
  NAND2_X1 U4969 ( .A1(n4461), .A2(n3003), .ZN(n4009) );
  AND2_X2 U4970 ( .A1(n4009), .A2(n4008), .ZN(n4577) );
  MUX2_X1 U4971 ( .A(n4085), .B(n4005), .S(EBX_REG_2__SCAN_IN), .Z(n4012) );
  NAND2_X1 U4972 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n2960), .ZN(n4010)
         );
  AND2_X1 U4973 ( .A1(n4021), .A2(n4010), .ZN(n4011) );
  NAND2_X1 U4974 ( .A1(n4012), .A2(n4011), .ZN(n4576) );
  AND2_X2 U4975 ( .A1(n4577), .A2(n4576), .ZN(n4624) );
  OR2_X2 U4976 ( .A1(n2959), .A2(n4001), .ZN(n4081) );
  MUX2_X1 U4977 ( .A(n4081), .B(n3981), .S(EBX_REG_3__SCAN_IN), .Z(n4013) );
  OAI21_X1 U4978 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4629), .A(n4013), 
        .ZN(n4014) );
  INV_X1 U4979 ( .A(n4014), .ZN(n4623) );
  MUX2_X1 U4980 ( .A(n4085), .B(n4005), .S(EBX_REG_4__SCAN_IN), .Z(n4017) );
  NAND2_X1 U4981 ( .A1(n2959), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4015)
         );
  AND2_X1 U4982 ( .A1(n4021), .A2(n4015), .ZN(n4016) );
  NAND2_X1 U4983 ( .A1(n4017), .A2(n4016), .ZN(n4627) );
  NAND2_X1 U4984 ( .A1(n2975), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4018)
         );
  OAI211_X1 U4985 ( .C1(n2959), .C2(EBX_REG_5__SCAN_IN), .A(n4005), .B(n4018), 
        .ZN(n4019) );
  OAI21_X1 U4986 ( .B1(n4081), .B2(EBX_REG_5__SCAN_IN), .A(n4019), .ZN(n5104)
         );
  MUX2_X1 U4987 ( .A(n4085), .B(n4005), .S(EBX_REG_6__SCAN_IN), .Z(n4023) );
  NAND2_X1 U4988 ( .A1(n2960), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4020)
         );
  AND2_X1 U4989 ( .A1(n4021), .A2(n4020), .ZN(n4022) );
  NAND2_X1 U4990 ( .A1(n4023), .A2(n4022), .ZN(n4834) );
  INV_X1 U4991 ( .A(n4834), .ZN(n4024) );
  NOR2_X2 U4992 ( .A1(n5107), .A2(n4024), .ZN(n4908) );
  INV_X1 U4993 ( .A(n4081), .ZN(n4159) );
  INV_X1 U4994 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U4995 ( .A1(n4159), .A2(n6129), .ZN(n4027) );
  NAND2_X1 U4996 ( .A1(n2975), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4025)
         );
  OAI211_X1 U4997 ( .C1(n2960), .C2(EBX_REG_7__SCAN_IN), .A(n4005), .B(n4025), 
        .ZN(n4026) );
  NAND2_X1 U4998 ( .A1(n4908), .A2(n4907), .ZN(n5126) );
  INV_X1 U4999 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4307) );
  NAND2_X1 U5000 ( .A1(n4005), .A2(n4307), .ZN(n4028) );
  OAI211_X1 U5001 ( .C1(n2959), .C2(EBX_REG_8__SCAN_IN), .A(n2975), .B(n4028), 
        .ZN(n4029) );
  OAI21_X1 U5002 ( .B1(n4085), .B2(EBX_REG_8__SCAN_IN), .A(n4029), .ZN(n4030)
         );
  NAND2_X1 U5003 ( .A1(n2975), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4031)
         );
  OAI211_X1 U5004 ( .C1(n2960), .C2(EBX_REG_9__SCAN_IN), .A(n4005), .B(n4031), 
        .ZN(n4032) );
  OAI21_X1 U5005 ( .B1(n4081), .B2(EBX_REG_9__SCAN_IN), .A(n4032), .ZN(n6107)
         );
  INV_X1 U5006 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U5007 ( .A1(n4005), .A2(n6297), .ZN(n4033) );
  OAI211_X1 U5008 ( .C1(n2960), .C2(EBX_REG_10__SCAN_IN), .A(n2975), .B(n4033), 
        .ZN(n4034) );
  OAI21_X1 U5009 ( .B1(n4085), .B2(EBX_REG_10__SCAN_IN), .A(n4034), .ZN(n5362)
         );
  INV_X1 U5010 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U5011 ( .A1(n4159), .A2(n6651), .ZN(n4037) );
  NAND2_X1 U5012 ( .A1(n2975), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4035) );
  OAI211_X1 U5013 ( .C1(n2960), .C2(EBX_REG_11__SCAN_IN), .A(n4005), .B(n4035), 
        .ZN(n4036) );
  INV_X1 U5014 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4312) );
  NAND2_X1 U5015 ( .A1(n4005), .A2(n4312), .ZN(n4038) );
  OAI211_X1 U5016 ( .C1(n2959), .C2(EBX_REG_12__SCAN_IN), .A(n2975), .B(n4038), 
        .ZN(n4039) );
  OAI21_X1 U5017 ( .B1(n4085), .B2(EBX_REG_12__SCAN_IN), .A(n4039), .ZN(n4040)
         );
  INV_X1 U5018 ( .A(n4040), .ZN(n5333) );
  NAND2_X1 U5019 ( .A1(n2975), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4042) );
  OAI211_X1 U5020 ( .C1(n2960), .C2(EBX_REG_13__SCAN_IN), .A(n4005), .B(n4042), 
        .ZN(n4043) );
  OAI21_X1 U5021 ( .B1(n4081), .B2(EBX_REG_13__SCAN_IN), .A(n4043), .ZN(n5320)
         );
  NOR2_X2 U5022 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  INV_X1 U5023 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U5024 ( .A1(n4005), .A2(n5878), .ZN(n4044) );
  OAI211_X1 U5025 ( .C1(n2960), .C2(EBX_REG_14__SCAN_IN), .A(n2975), .B(n4044), 
        .ZN(n4045) );
  OAI21_X1 U5026 ( .B1(n4085), .B2(EBX_REG_14__SCAN_IN), .A(n4045), .ZN(n5308)
         );
  MUX2_X1 U5027 ( .A(n4081), .B(n2975), .S(EBX_REG_15__SCAN_IN), .Z(n4047) );
  INV_X1 U5028 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5864) );
  INV_X1 U5029 ( .A(n4629), .ZN(n4156) );
  NAND2_X1 U5030 ( .A1(n5864), .A2(n4156), .ZN(n4046) );
  INV_X2 U5031 ( .A(n5297), .ZN(n4054) );
  INV_X1 U5032 ( .A(n4085), .ZN(n4048) );
  INV_X1 U5033 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U5034 ( .A1(n4048), .A2(n5436), .ZN(n4051) );
  INV_X1 U5035 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U5036 ( .A1(n4005), .A2(n5852), .ZN(n4049) );
  OAI211_X1 U5037 ( .C1(n2959), .C2(EBX_REG_16__SCAN_IN), .A(n2975), .B(n4049), 
        .ZN(n4050) );
  NAND2_X1 U5038 ( .A1(n2975), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4052) );
  OAI211_X1 U5039 ( .C1(n2959), .C2(EBX_REG_17__SCAN_IN), .A(n4005), .B(n4052), 
        .ZN(n4053) );
  OAI21_X1 U5040 ( .B1(n4081), .B2(EBX_REG_17__SCAN_IN), .A(n4053), .ZN(n5431)
         );
  INV_X1 U5041 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U5042 ( .A1(n4005), .A2(n5833), .ZN(n4055) );
  OAI211_X1 U5043 ( .C1(n2960), .C2(EBX_REG_19__SCAN_IN), .A(n2975), .B(n4055), 
        .ZN(n4056) );
  OAI21_X1 U5044 ( .B1(n4085), .B2(EBX_REG_19__SCAN_IN), .A(n4056), .ZN(n4057)
         );
  INV_X1 U5045 ( .A(n4057), .ZN(n5421) );
  OR2_X1 U5046 ( .A1(n4629), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4059)
         );
  OR2_X1 U5047 ( .A1(n2959), .A2(EBX_REG_20__SCAN_IN), .ZN(n4058) );
  AND2_X1 U5048 ( .A1(n4059), .A2(n4058), .ZN(n5284) );
  OR2_X1 U5049 ( .A1(n2959), .A2(EBX_REG_18__SCAN_IN), .ZN(n5417) );
  OR2_X1 U5050 ( .A1(n4629), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4060)
         );
  NAND2_X1 U5051 ( .A1(n5417), .A2(n4060), .ZN(n5418) );
  NAND2_X1 U5052 ( .A1(n4001), .A2(EBX_REG_20__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U5053 ( .A1(n5418), .A2(n2975), .ZN(n4061) );
  OAI211_X1 U5054 ( .C1(n5284), .C2(n5418), .A(n4062), .B(n4061), .ZN(n4063)
         );
  INV_X1 U5055 ( .A(n4063), .ZN(n4064) );
  NAND2_X1 U5056 ( .A1(n2975), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4065) );
  OAI211_X1 U5057 ( .C1(n2959), .C2(EBX_REG_21__SCAN_IN), .A(n4005), .B(n4065), 
        .ZN(n4066) );
  OAI21_X1 U5058 ( .B1(n4081), .B2(EBX_REG_21__SCAN_IN), .A(n4066), .ZN(n5270)
         );
  MUX2_X1 U5059 ( .A(n4081), .B(n2975), .S(EBX_REG_23__SCAN_IN), .Z(n4067) );
  OAI21_X1 U5060 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n4629), .A(n4067), 
        .ZN(n5248) );
  INV_X1 U5061 ( .A(n5248), .ZN(n4070) );
  MUX2_X1 U5062 ( .A(n4085), .B(n4005), .S(EBX_REG_22__SCAN_IN), .Z(n4069) );
  NAND2_X1 U5063 ( .A1(n2960), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4068) );
  NAND2_X1 U5064 ( .A1(n4069), .A2(n4068), .ZN(n5260) );
  NAND2_X1 U5065 ( .A1(n4070), .A2(n5260), .ZN(n4071) );
  NOR2_X4 U5066 ( .A1(n5273), .A2(n4071), .ZN(n5247) );
  INV_X1 U5067 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U5068 ( .A1(n4005), .A2(n5774), .ZN(n4072) );
  OAI211_X1 U5069 ( .C1(n2960), .C2(EBX_REG_24__SCAN_IN), .A(n2975), .B(n4072), 
        .ZN(n4073) );
  OAI21_X1 U5070 ( .B1(n4085), .B2(EBX_REG_24__SCAN_IN), .A(n4073), .ZN(n5240)
         );
  INV_X1 U5071 ( .A(n5240), .ZN(n4075) );
  MUX2_X1 U5072 ( .A(n4081), .B(n2975), .S(EBX_REG_25__SCAN_IN), .Z(n4074) );
  OAI21_X1 U5073 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4629), .A(n4074), 
        .ZN(n5225) );
  NOR2_X1 U5074 ( .A1(n4075), .A2(n5225), .ZN(n4076) );
  AND2_X2 U5075 ( .A1(n5247), .A2(n4076), .ZN(n5228) );
  MUX2_X1 U5076 ( .A(n4085), .B(n4005), .S(EBX_REG_26__SCAN_IN), .Z(n4078) );
  NAND2_X1 U5077 ( .A1(n2960), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4077) );
  NAND2_X1 U5078 ( .A1(n4078), .A2(n4077), .ZN(n5213) );
  NAND2_X1 U5079 ( .A1(n2975), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4079) );
  OAI211_X1 U5080 ( .C1(n2959), .C2(EBX_REG_27__SCAN_IN), .A(n4005), .B(n4079), 
        .ZN(n4080) );
  OAI21_X1 U5081 ( .B1(n4081), .B2(EBX_REG_27__SCAN_IN), .A(n4080), .ZN(n5199)
         );
  INV_X1 U5082 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U5083 ( .A1(n4005), .A2(n5500), .ZN(n4083) );
  OAI211_X1 U5084 ( .C1(n2960), .C2(EBX_REG_28__SCAN_IN), .A(n2975), .B(n4083), 
        .ZN(n4084) );
  OAI21_X1 U5085 ( .B1(n4085), .B2(EBX_REG_28__SCAN_IN), .A(n4084), .ZN(n4087)
         );
  INV_X1 U5086 ( .A(n4087), .ZN(n4086) );
  INV_X1 U5087 ( .A(n5183), .ZN(n4193) );
  OAI21_X1 U5088 ( .B1(n3175), .B2(n4087), .A(n4193), .ZN(n5734) );
  INV_X1 U5089 ( .A(n5164), .ZN(n4672) );
  AOI22_X1 U5090 ( .A1(n2978), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5091 ( .A1(n2961), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5092 ( .A1(n2973), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5093 ( .A1(n4092), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4093) );
  NAND4_X1 U5094 ( .A1(n4096), .A2(n4095), .A3(n4094), .A4(n4093), .ZN(n4102)
         );
  AOI22_X1 U5095 ( .A1(n2971), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5096 ( .A1(n3489), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5097 ( .A1(n4120), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5098 ( .A1(n2979), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4097) );
  NAND4_X1 U5099 ( .A1(n4100), .A2(n4099), .A3(n4098), .A4(n4097), .ZN(n4101)
         );
  NOR2_X1 U5100 ( .A1(n4102), .A2(n4101), .ZN(n4114) );
  NAND2_X1 U5101 ( .A1(n4104), .A2(n4103), .ZN(n4113) );
  XNOR2_X1 U5102 ( .A(n4114), .B(n4113), .ZN(n4107) );
  AOI22_X1 U5103 ( .A1(n3721), .A2(EAX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5978), .ZN(n4105) );
  OAI21_X1 U5104 ( .B1(n4107), .B2(n4106), .A(n4105), .ZN(n4111) );
  INV_X1 U5105 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U5106 ( .A1(n4109), .A2(n5180), .ZN(n4110) );
  NAND2_X1 U5107 ( .A1(n4149), .A2(n4110), .ZN(n5494) );
  MUX2_X1 U5108 ( .A(n4111), .B(n5494), .S(n3438), .Z(n5179) );
  NOR2_X1 U5109 ( .A1(n4114), .A2(n4113), .ZN(n4129) );
  AOI22_X1 U5110 ( .A1(n2978), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3489), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5111 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n2971), .B1(n3407), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5112 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n3313), .B1(n2969), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5113 ( .A1(n2961), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4115) );
  NAND4_X1 U5114 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(n4127)
         );
  AOI22_X1 U5115 ( .A1(n2979), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5116 ( .A1(n2976), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5117 ( .A1(n2973), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5118 ( .A1(n4121), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4122) );
  NAND4_X1 U5119 ( .A1(n4125), .A2(n4124), .A3(n4123), .A4(n4122), .ZN(n4126)
         );
  NOR2_X1 U5120 ( .A1(n4127), .A2(n4126), .ZN(n4128) );
  XNOR2_X1 U5121 ( .A(n4129), .B(n4128), .ZN(n4133) );
  INV_X1 U5122 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4130) );
  INV_X1 U5123 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5159) );
  OAI22_X1 U5124 ( .A1(n3032), .A2(n4130), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5159), .ZN(n4131) );
  AOI21_X1 U5125 ( .B1(n4133), .B2(n4132), .A(n4131), .ZN(n4134) );
  XNOR2_X1 U5126 ( .A(n4149), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5161)
         );
  MUX2_X1 U5127 ( .A(n4134), .B(n5161), .S(n3859), .Z(n4191) );
  AOI22_X1 U5128 ( .A1(n3721), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4135), .ZN(n4136) );
  NAND3_X1 U5129 ( .A1(n4141), .A2(n4140), .A3(n4139), .ZN(n4142) );
  NAND2_X1 U5130 ( .A1(n4143), .A2(n4142), .ZN(n4145) );
  AND2_X1 U5131 ( .A1(n4145), .A2(n4144), .ZN(n4411) );
  INV_X1 U5132 ( .A(n4411), .ZN(n4146) );
  NAND2_X1 U5133 ( .A1(n5170), .A2(n5978), .ZN(n6568) );
  NOR3_X1 U5134 ( .A1(n6566), .A2(n6588), .A3(n6568), .ZN(n6564) );
  AND2_X1 U5135 ( .A1(n3438), .A2(n4222), .ZN(n6575) );
  INV_X1 U5136 ( .A(n6575), .ZN(n4147) );
  OR2_X2 U5137 ( .A1(n4225), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U5138 ( .A1(n4147), .A2(n6287), .ZN(n4148) );
  INV_X1 U5139 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4151) );
  NOR2_X1 U5140 ( .A1(n4230), .A2(n5170), .ZN(n4153) );
  NAND2_X1 U5141 ( .A1(n4232), .A2(n6152), .ZN(n4190) );
  NAND2_X1 U5142 ( .A1(n4629), .A2(EBX_REG_30__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U5143 ( .A1(n2960), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4154) );
  NAND2_X1 U5144 ( .A1(n4155), .A2(n4154), .ZN(n4195) );
  INV_X1 U5145 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6650) );
  INV_X1 U5146 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U5147 ( .A1(n4156), .A2(n5726), .ZN(n4160) );
  INV_X1 U5148 ( .A(n4160), .ZN(n4157) );
  MUX2_X1 U5149 ( .A(EBX_REG_29__SCAN_IN), .B(n4157), .S(n2975), .Z(n4158) );
  AOI21_X1 U5150 ( .B1(n4159), .B2(n6650), .A(n4158), .ZN(n5182) );
  NAND2_X1 U5151 ( .A1(n5183), .A2(n5182), .ZN(n5181) );
  OAI21_X1 U5152 ( .B1(EBX_REG_29__SCAN_IN), .B2(n2959), .A(n4160), .ZN(n4161)
         );
  NAND2_X1 U5153 ( .A1(n4197), .A2(n2975), .ZN(n4192) );
  OAI22_X1 U5154 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n4629), .B1(n2959), .B2(EBX_REG_31__SCAN_IN), .ZN(n4162) );
  INV_X1 U5155 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5406) );
  NOR2_X1 U5156 ( .A1(n4343), .A2(n5406), .ZN(n4167) );
  NOR2_X1 U5157 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n4200) );
  NOR2_X1 U5158 ( .A1(n2959), .A2(n4200), .ZN(n4165) );
  OR2_X1 U5159 ( .A1(n4166), .A2(STATE_REG_0__SCAN_IN), .ZN(n6018) );
  INV_X1 U5160 ( .A(n6018), .ZN(n4563) );
  NAND2_X1 U5161 ( .A1(n4563), .A2(n4200), .ZN(n6563) );
  AND2_X1 U5162 ( .A1(n4464), .A2(n6563), .ZN(n4203) );
  AOI22_X1 U5163 ( .A1(n4167), .A2(n4203), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n6142), .ZN(n4181) );
  NAND2_X1 U5164 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5327) );
  INV_X1 U5165 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6150) );
  INV_X1 U5166 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5372) );
  INV_X1 U5167 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4368) );
  INV_X1 U5168 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5390) );
  NOR3_X1 U5169 ( .A1(n5372), .A2(n4368), .A3(n5390), .ZN(n6157) );
  NAND3_X1 U5170 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .A3(
        n6157), .ZN(n6140) );
  NOR2_X1 U5171 ( .A1(n6150), .A2(n6140), .ZN(n6115) );
  NAND3_X1 U5172 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n6115), .ZN(n4182) );
  NOR2_X1 U5173 ( .A1(n6135), .A2(n4182), .ZN(n5360) );
  NAND4_X1 U5174 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n5360), .ZN(n5324) );
  NOR2_X1 U5175 ( .A1(n5327), .A2(n5324), .ZN(n4168) );
  NAND2_X1 U5176 ( .A1(n4168), .A2(REIP_REG_14__SCAN_IN), .ZN(n4170) );
  NAND2_X1 U5177 ( .A1(n4691), .A2(n6018), .ZN(n4535) );
  AND3_X1 U5178 ( .A1(n4535), .A2(n4200), .A3(n4537), .ZN(n4169) );
  NAND2_X1 U5179 ( .A1(n6159), .A2(n5371), .ZN(n6134) );
  AND2_X1 U5180 ( .A1(n4170), .A2(n6134), .ZN(n6098) );
  NAND3_X1 U5181 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4171) );
  AND2_X1 U5182 ( .A1(n6134), .A2(n4171), .ZN(n4172) );
  INV_X1 U5183 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U5184 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n6025) );
  OAI21_X1 U5185 ( .B1(n5588), .B2(n6025), .A(n6134), .ZN(n4173) );
  NAND2_X1 U5186 ( .A1(n6093), .A2(n4173), .ZN(n5287) );
  NAND3_X1 U5187 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4174) );
  AND2_X1 U5188 ( .A1(n6134), .A2(n4174), .ZN(n4175) );
  NAND2_X1 U5189 ( .A1(REIP_REG_25__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .ZN(
        n4184) );
  INV_X1 U5190 ( .A(n4184), .ZN(n4176) );
  NAND2_X1 U5191 ( .A1(n4176), .A2(REIP_REG_24__SCAN_IN), .ZN(n4177) );
  AND2_X1 U5192 ( .A1(n6134), .A2(n4177), .ZN(n4178) );
  NOR2_X2 U5193 ( .A1(n5254), .A2(n4178), .ZN(n5202) );
  NAND2_X1 U5194 ( .A1(n5202), .A2(n6159), .ZN(n4208) );
  AND2_X1 U5195 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4185) );
  NAND2_X1 U5196 ( .A1(n5202), .A2(n4185), .ZN(n4179) );
  NAND2_X1 U5197 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n4186) );
  OAI211_X1 U5198 ( .C1(n5186), .C2(n4186), .A(REIP_REG_31__SCAN_IN), .B(n4208), .ZN(n4180) );
  OAI211_X1 U5199 ( .C1(n5687), .C2(n6172), .A(n4181), .B(n4180), .ZN(n4188)
         );
  INV_X1 U5200 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5307) );
  INV_X1 U5201 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5354) );
  NAND3_X1 U5202 ( .A1(n5339), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n5306) );
  AND3_X1 U5203 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_17__SCAN_IN), .ZN(n4183) );
  INV_X1 U5204 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5572) );
  NAND3_X1 U5205 ( .A1(n5255), .A2(REIP_REG_24__SCAN_IN), .A3(
        REIP_REG_23__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U5206 ( .A1(n5208), .A2(n4185), .ZN(n5187) );
  NOR3_X1 U5207 ( .A1(n5187), .A2(REIP_REG_31__SCAN_IN), .A3(n4186), .ZN(n4187) );
  NAND2_X1 U5208 ( .A1(n4190), .A2(n4189), .ZN(U2796) );
  XNOR2_X2 U5209 ( .A(n5178), .B(n4191), .ZN(n5169) );
  INV_X1 U5210 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5493) );
  INV_X1 U5211 ( .A(n4197), .ZN(n4194) );
  OAI211_X1 U5212 ( .C1(n4194), .C2(n4193), .A(n4192), .B(n4195), .ZN(n4199)
         );
  INV_X1 U5213 ( .A(n4195), .ZN(n4196) );
  OAI211_X1 U5214 ( .C1(n5183), .C2(n3981), .A(n4197), .B(n4196), .ZN(n4198)
         );
  NAND2_X1 U5215 ( .A1(n4199), .A2(n4198), .ZN(n5716) );
  NOR2_X1 U5216 ( .A1(n4200), .A2(EBX_REG_31__SCAN_IN), .ZN(n4201) );
  AND2_X1 U5217 ( .A1(n4537), .A2(n4201), .ZN(n4202) );
  NOR2_X1 U5218 ( .A1(n4203), .A2(n4202), .ZN(n4204) );
  NOR2_X2 U5219 ( .A1(n4343), .A2(n4204), .ZN(n6143) );
  INV_X1 U5220 ( .A(n5161), .ZN(n4206) );
  OAI22_X1 U5221 ( .A1(n5159), .A2(n6186), .B1(n6155), .B2(n4206), .ZN(n4207)
         );
  AOI21_X1 U5222 ( .B1(EBX_REG_30__SCAN_IN), .B2(n6143), .A(n4207), .ZN(n4210)
         );
  OAI211_X1 U5223 ( .C1(n5186), .C2(n5493), .A(REIP_REG_30__SCAN_IN), .B(n4208), .ZN(n4209) );
  OAI211_X1 U5224 ( .C1(n5716), .C2(n6172), .A(n4210), .B(n4209), .ZN(n4211)
         );
  INV_X1 U5225 ( .A(n4211), .ZN(n4212) );
  OR2_X1 U5226 ( .A1(n4543), .A2(n2959), .ZN(n4557) );
  NOR2_X1 U5227 ( .A1(READY_N), .A2(n4411), .ZN(n4530) );
  INV_X1 U5228 ( .A(n4530), .ZN(n4214) );
  NOR2_X1 U5229 ( .A1(n6048), .A2(n4214), .ZN(n4428) );
  NOR2_X1 U5230 ( .A1(n4215), .A2(n3346), .ZN(n4216) );
  AOI21_X1 U5231 ( .B1(n4428), .B2(n6559), .A(n4216), .ZN(n4219) );
  NAND2_X1 U5232 ( .A1(n4421), .A2(n4406), .ZN(n4444) );
  NAND2_X1 U5233 ( .A1(n4232), .A2(n3214), .ZN(n4221) );
  AOI22_X1 U5234 ( .A1(n3031), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6779), .ZN(n4220) );
  NAND2_X1 U5235 ( .A1(n4221), .A2(n4220), .ZN(U2860) );
  NAND2_X1 U5236 ( .A1(n4222), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6579) );
  OR2_X2 U5237 ( .A1(n6579), .A2(n6476), .ZN(n6258) );
  INV_X1 U5238 ( .A(n4223), .ZN(n4224) );
  NAND2_X1 U5239 ( .A1(n4421), .A2(n4224), .ZN(n6552) );
  NAND2_X1 U5240 ( .A1(n6476), .A2(n4225), .ZN(n6610) );
  NAND2_X1 U5241 ( .A1(n6610), .A2(n6566), .ZN(n4226) );
  NAND2_X1 U5242 ( .A1(n6566), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4228) );
  NAND2_X1 U5243 ( .A1(n6059), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4227) );
  NAND2_X1 U5244 ( .A1(n4228), .A2(n4227), .ZN(n4484) );
  NAND2_X1 U5245 ( .A1(n6246), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4229)
         );
  INV_X1 U5246 ( .A(n6287), .ZN(n6247) );
  NAND2_X1 U5247 ( .A1(n6247), .A2(REIP_REG_31__SCAN_IN), .ZN(n5688) );
  OAI211_X1 U5248 ( .C1(n6254), .C2(n4230), .A(n4229), .B(n5688), .ZN(n4231)
         );
  AOI21_X1 U5249 ( .B1(n4232), .B2(n6265), .A(n4231), .ZN(n4331) );
  INV_X1 U5250 ( .A(n4280), .ZN(n4294) );
  NAND2_X1 U5251 ( .A1(n4259), .A2(n4260), .ZN(n4258) );
  INV_X1 U5252 ( .A(n4233), .ZN(n4249) );
  NAND2_X1 U5253 ( .A1(n4258), .A2(n4249), .ZN(n4248) );
  NAND2_X1 U5254 ( .A1(n4248), .A2(n4241), .ZN(n4235) );
  INV_X1 U5255 ( .A(n4235), .ZN(n4237) );
  INV_X1 U5256 ( .A(n4236), .ZN(n4234) );
  OR2_X1 U5257 ( .A1(n4235), .A2(n4234), .ZN(n4285) );
  OAI211_X1 U5258 ( .C1(n4237), .C2(n4236), .A(n4464), .B(n4285), .ZN(n4238)
         );
  INV_X1 U5259 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4240) );
  INV_X1 U5260 ( .A(n4241), .ZN(n4242) );
  XNOR2_X1 U5261 ( .A(n4248), .B(n4242), .ZN(n4243) );
  NAND2_X1 U5262 ( .A1(n4243), .A2(n4464), .ZN(n4244) );
  NAND2_X1 U5263 ( .A1(n4245), .A2(n4244), .ZN(n4270) );
  INV_X1 U5264 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4642) );
  XNOR2_X1 U5265 ( .A(n4270), .B(n4642), .ZN(n4634) );
  OAI21_X1 U5266 ( .B1(n4249), .B2(n4258), .A(n4248), .ZN(n4251) );
  AOI21_X1 U5267 ( .B1(n4251), .B2(n4464), .A(n4253), .ZN(n4252) );
  NAND2_X1 U5268 ( .A1(n4268), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4568)
         );
  INV_X1 U5269 ( .A(n4464), .ZN(n6614) );
  INV_X1 U5270 ( .A(n4253), .ZN(n4254) );
  OAI21_X1 U5271 ( .B1(n6614), .B2(n4260), .A(n4254), .ZN(n4255) );
  INV_X1 U5272 ( .A(n4255), .ZN(n4256) );
  NAND2_X1 U5273 ( .A1(n4257), .A2(n4256), .ZN(n4486) );
  NAND2_X2 U5274 ( .A1(n4486), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5911)
         );
  OR2_X1 U5275 ( .A1(n5041), .A2(n4294), .ZN(n4265) );
  OAI21_X1 U5276 ( .B1(n4260), .B2(n4259), .A(n4258), .ZN(n4262) );
  OAI211_X1 U5277 ( .C1(n4262), .C2(n6614), .A(n4261), .B(n3324), .ZN(n4263)
         );
  INV_X1 U5278 ( .A(n4263), .ZN(n4264) );
  NAND2_X1 U5279 ( .A1(n4265), .A2(n4264), .ZN(n4552) );
  INV_X1 U5280 ( .A(n5911), .ZN(n4266) );
  NAND2_X1 U5281 ( .A1(n4266), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4267)
         );
  NAND2_X1 U5282 ( .A1(n4568), .A2(n4570), .ZN(n4269) );
  AND2_X2 U5283 ( .A1(n4269), .A2(n4569), .ZN(n4633) );
  NAND2_X1 U5284 ( .A1(n4270), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4271)
         );
  NAND2_X1 U5285 ( .A1(n4273), .A2(n4280), .ZN(n4276) );
  XNOR2_X1 U5286 ( .A(n4285), .B(n4283), .ZN(n4274) );
  NAND2_X1 U5287 ( .A1(n4274), .A2(n4464), .ZN(n4275) );
  NAND2_X1 U5288 ( .A1(n4276), .A2(n4275), .ZN(n4277) );
  INV_X1 U5289 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5116) );
  XNOR2_X1 U5290 ( .A(n4277), .B(n5116), .ZN(n5103) );
  NAND2_X1 U5291 ( .A1(n5102), .A2(n5103), .ZN(n4279) );
  NAND2_X1 U5292 ( .A1(n4277), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4278)
         );
  NAND2_X1 U5293 ( .A1(n4279), .A2(n4278), .ZN(n5088) );
  NAND2_X1 U5294 ( .A1(n4302), .A2(n4282), .ZN(n4289) );
  INV_X1 U5295 ( .A(n4283), .ZN(n4284) );
  NOR2_X1 U5296 ( .A1(n4285), .A2(n4284), .ZN(n4287) );
  NAND2_X1 U5297 ( .A1(n4287), .A2(n4286), .ZN(n4303) );
  OAI211_X1 U5298 ( .C1(n4287), .C2(n4286), .A(n4303), .B(n4464), .ZN(n4288)
         );
  NAND2_X1 U5299 ( .A1(n4289), .A2(n4288), .ZN(n4290) );
  INV_X1 U5300 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5096) );
  XNOR2_X1 U5301 ( .A(n4290), .B(n5096), .ZN(n5087) );
  NAND2_X1 U5302 ( .A1(n5088), .A2(n5087), .ZN(n4292) );
  NAND2_X1 U5303 ( .A1(n4290), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4291)
         );
  INV_X1 U5304 ( .A(n4293), .ZN(n4295) );
  XNOR2_X1 U5305 ( .A(n4303), .B(n4304), .ZN(n4296) );
  NAND2_X1 U5306 ( .A1(n4296), .A2(n4464), .ZN(n4297) );
  NAND2_X1 U5307 ( .A1(n4298), .A2(n4297), .ZN(n4300) );
  INV_X1 U5308 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4299) );
  XNOR2_X1 U5309 ( .A(n4300), .B(n4299), .ZN(n5130) );
  NAND2_X1 U5310 ( .A1(n4300), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4301)
         );
  INV_X1 U5311 ( .A(n4303), .ZN(n4305) );
  NAND3_X1 U5312 ( .A1(n4305), .A2(n4464), .A3(n4304), .ZN(n4306) );
  NAND2_X1 U5313 ( .A1(n4309), .A2(n4306), .ZN(n4308) );
  INV_X1 U5314 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6307) );
  INV_X1 U5315 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4311) );
  NAND2_X1 U5316 ( .A1(n2989), .A2(n4311), .ZN(n5887) );
  NAND2_X1 U5317 ( .A1(n5674), .A2(n4312), .ZN(n5653) );
  NOR2_X1 U5318 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4313) );
  OR2_X1 U5319 ( .A1(n4309), .A2(n4313), .ZN(n4314) );
  NOR2_X1 U5320 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4316) );
  INV_X1 U5321 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U5322 ( .A1(n4309), .A2(n6045), .ZN(n5636) );
  NAND2_X1 U5323 ( .A1(n4309), .A2(n5878), .ZN(n4317) );
  AND2_X1 U5324 ( .A1(n5636), .A2(n4317), .ZN(n4318) );
  NAND2_X1 U5325 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U5326 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5693) );
  OAI21_X1 U5327 ( .B1(n5703), .B2(n5693), .A(n5609), .ZN(n4319) );
  INV_X1 U5328 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U5329 ( .A1(n5852), .A2(n5848), .ZN(n5603) );
  NOR2_X1 U5330 ( .A1(n5603), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4320)
         );
  AND2_X1 U5331 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5790) );
  AND2_X1 U5332 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U5333 ( .A1(n5790), .A2(n5704), .ZN(n5559) );
  NAND2_X1 U5334 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5708) );
  OAI21_X1 U5335 ( .B1(n5559), .B2(n5708), .A(n5609), .ZN(n4323) );
  INV_X1 U5336 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6736) );
  INV_X1 U5337 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5564) );
  NAND4_X1 U5338 ( .A1(n6736), .A2(n5833), .A3(n5564), .A4(n5774), .ZN(n4324)
         );
  INV_X1 U5339 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5545) );
  INV_X1 U5340 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U5341 ( .A1(n5545), .A2(n5795), .ZN(n5788) );
  NOR2_X1 U5342 ( .A1(n4324), .A2(n5788), .ZN(n4325) );
  INV_X1 U5343 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5764) );
  XNOR2_X1 U5344 ( .A(n5674), .B(n5764), .ZN(n5535) );
  NAND2_X1 U5345 ( .A1(n5609), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U5346 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5737) );
  NOR3_X2 U5347 ( .A1(n5516), .A2(n5737), .A3(n5726), .ZN(n5155) );
  INV_X1 U5348 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U5349 ( .A1(n5500), .A2(n5517), .ZN(n5738) );
  INV_X1 U5350 ( .A(n6256), .ZN(n4329) );
  NAND2_X1 U5351 ( .A1(n4331), .A2(n4330), .ZN(U2955) );
  INV_X1 U5352 ( .A(n4461), .ZN(n4337) );
  NAND2_X1 U5353 ( .A1(n4332), .A2(n4406), .ZN(n4333) );
  NAND2_X1 U5354 ( .A1(n4333), .A2(n6095), .ZN(n6182) );
  INV_X1 U5355 ( .A(n4334), .ZN(n4491) );
  OAI21_X1 U5356 ( .B1(n4336), .B2(n4335), .A(n4491), .ZN(n4590) );
  OAI22_X1 U5357 ( .A1(n6172), .A2(n4337), .B1(n5405), .B2(n4590), .ZN(n4346)
         );
  INV_X1 U5358 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U5359 ( .A1(n6174), .A2(n4585), .ZN(n4340) );
  NAND2_X1 U5360 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4339)
         );
  AOI22_X1 U5361 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6143), .B1(n6135), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n4338) );
  NAND3_X1 U5362 ( .A1(n4340), .A2(n4339), .A3(n4338), .ZN(n4345) );
  NOR2_X1 U5363 ( .A1(n4343), .A2(n4342), .ZN(n6177) );
  AND2_X1 U5364 ( .A1(n4341), .A2(n6177), .ZN(n4344) );
  NOR2_X1 U5365 ( .A1(n6159), .A2(REIP_REG_1__SCAN_IN), .ZN(n5391) );
  INV_X1 U5366 ( .A(READY_N), .ZN(n6611) );
  AOI221_X1 U5367 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6611), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4348) );
  INV_X1 U5368 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6014) );
  INV_X1 U5369 ( .A(HOLD), .ZN(n4381) );
  NAND2_X1 U5370 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6019) );
  INV_X1 U5371 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4353) );
  AOI21_X1 U5372 ( .B1(n4381), .B2(n6019), .A(n4353), .ZN(n4347) );
  AOI211_X1 U5373 ( .C1(n4348), .C2(HOLD), .A(n6014), .B(n4347), .ZN(n4352) );
  INV_X1 U5374 ( .A(NA_N), .ZN(n4349) );
  NAND2_X1 U5375 ( .A1(STATE_REG_2__SCAN_IN), .A2(n4349), .ZN(n4350) );
  AND3_X1 U5376 ( .A1(n4380), .A2(n6014), .A3(n4350), .ZN(n4378) );
  INV_X1 U5377 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6760) );
  OR3_X1 U5378 ( .A1(n6014), .A2(n6760), .A3(n6019), .ZN(n4351) );
  OAI22_X1 U5379 ( .A1(n4352), .A2(n4378), .B1(NA_N), .B2(n4351), .ZN(U3183)
         );
  NAND2_X1 U5380 ( .A1(n6021), .A2(n4353), .ZN(n4395) );
  INV_X1 U5381 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5537) );
  INV_X1 U5382 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6740) );
  INV_X1 U5383 ( .A(REIP_REG_24__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U5384 ( .A1(n6021), .A2(STATE_REG_2__SCAN_IN), .ZN(n4387) );
  OAI222_X1 U5385 ( .A1(n4395), .A2(n5537), .B1(n6021), .B2(n6740), .C1(n4363), 
        .C2(n4387), .ZN(U3207) );
  INV_X1 U5386 ( .A(REIP_REG_16__SCAN_IN), .ZN(n4355) );
  INV_X1 U5387 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n4354) );
  INV_X1 U5388 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5294) );
  OAI222_X1 U5389 ( .A1(n4395), .A2(n4355), .B1(n4354), .B2(n6021), .C1(n4387), 
        .C2(n5294), .ZN(U3198) );
  INV_X1 U5390 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5616) );
  INV_X1 U5391 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n4356) );
  OAI222_X1 U5392 ( .A1(n4395), .A2(n5616), .B1(n4356), .B2(n6021), .C1(n4387), 
        .C2(n4355), .ZN(U3199) );
  INV_X1 U5393 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n4357) );
  OAI222_X1 U5394 ( .A1(n4395), .A2(n5572), .B1(n4357), .B2(n6021), .C1(n4387), 
        .C2(n3059), .ZN(U3204) );
  INV_X1 U5395 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6761) );
  INV_X1 U5396 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5507) );
  OAI222_X1 U5397 ( .A1(n4395), .A2(n5493), .B1(n6021), .B2(n6761), .C1(n5507), 
        .C2(n4387), .ZN(U3211) );
  INV_X1 U5398 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n4358) );
  INV_X1 U5399 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6023) );
  OAI222_X1 U5400 ( .A1(n4395), .A2(n5588), .B1(n4358), .B2(n6021), .C1(n4387), 
        .C2(n6023), .ZN(U3202) );
  INV_X1 U5401 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5158) );
  INV_X1 U5402 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6724) );
  INV_X1 U5403 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4359) );
  OAI222_X1 U5404 ( .A1(n4387), .A2(n5158), .B1(n6021), .B2(n6724), .C1(n4359), 
        .C2(n4395), .ZN(U3213) );
  INV_X1 U5405 ( .A(REIP_REG_23__SCAN_IN), .ZN(n5554) );
  AOI22_X1 U5406 ( .A1(n4398), .A2(REIP_REG_22__SCAN_IN), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n4375), .ZN(n4360) );
  OAI21_X1 U5407 ( .B1(n5554), .B2(n4395), .A(n4360), .ZN(U3205) );
  INV_X1 U5408 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6168) );
  AOI22_X1 U5409 ( .A1(n4398), .A2(REIP_REG_3__SCAN_IN), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n4375), .ZN(n4361) );
  OAI21_X1 U5410 ( .B1(n6168), .B2(n4395), .A(n4361), .ZN(U3186) );
  AOI22_X1 U5411 ( .A1(n4398), .A2(REIP_REG_23__SCAN_IN), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n4375), .ZN(n4362) );
  OAI21_X1 U5412 ( .B1(n4363), .B2(n4395), .A(n4362), .ZN(U3206) );
  AOI22_X1 U5413 ( .A1(n4398), .A2(REIP_REG_27__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n4375), .ZN(n4364) );
  OAI21_X1 U5414 ( .B1(n5507), .B2(n4395), .A(n4364), .ZN(U3210) );
  AOI22_X1 U5415 ( .A1(n4398), .A2(REIP_REG_1__SCAN_IN), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n4375), .ZN(n4365) );
  OAI21_X1 U5416 ( .B1(n5390), .B2(n4395), .A(n4365), .ZN(U3184) );
  INV_X1 U5417 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5512) );
  AOI22_X1 U5418 ( .A1(n4398), .A2(REIP_REG_26__SCAN_IN), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n4375), .ZN(n4366) );
  OAI21_X1 U5419 ( .B1(n5512), .B2(n4395), .A(n4366), .ZN(U3209) );
  AOI22_X1 U5420 ( .A1(n4398), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n4375), .ZN(n4367) );
  OAI21_X1 U5421 ( .B1(n4368), .B2(n4395), .A(n4367), .ZN(U3185) );
  INV_X1 U5422 ( .A(n4395), .ZN(n4385) );
  AOI22_X1 U5423 ( .A1(n4398), .A2(REIP_REG_14__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n4375), .ZN(n4369) );
  OAI21_X1 U5424 ( .B1(n5294), .B2(n4400), .A(n4369), .ZN(U3197) );
  INV_X1 U5425 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5212) );
  AOI22_X1 U5426 ( .A1(n4398), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n4375), .ZN(n4370) );
  OAI21_X1 U5427 ( .B1(n5212), .B2(n4400), .A(n4370), .ZN(U3208) );
  AOI22_X1 U5428 ( .A1(n4398), .A2(REIP_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n4375), .ZN(n4371) );
  OAI21_X1 U5429 ( .B1(n3059), .B2(n4400), .A(n4371), .ZN(U3203) );
  AOI22_X1 U5430 ( .A1(n4398), .A2(REIP_REG_18__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n4375), .ZN(n4372) );
  OAI21_X1 U5431 ( .B1(n6023), .B2(n4400), .A(n4372), .ZN(U3201) );
  INV_X1 U5432 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6077) );
  AOI22_X1 U5433 ( .A1(n4398), .A2(REIP_REG_17__SCAN_IN), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n4375), .ZN(n4373) );
  OAI21_X1 U5434 ( .B1(n6077), .B2(n4400), .A(n4373), .ZN(U3200) );
  AOI22_X1 U5435 ( .A1(n4398), .A2(REIP_REG_13__SCAN_IN), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n4375), .ZN(n4374) );
  OAI21_X1 U5436 ( .B1(n5307), .B2(n4400), .A(n4374), .ZN(U3196) );
  INV_X1 U5437 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4377) );
  NAND2_X1 U5438 ( .A1(M_IO_N_REG_SCAN_IN), .A2(n4375), .ZN(n4376) );
  OAI21_X1 U5439 ( .B1(n4375), .B2(n4377), .A(n4376), .ZN(U3473) );
  NAND2_X1 U5440 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6015) );
  NAND2_X1 U5441 ( .A1(n6019), .A2(n6015), .ZN(n4379) );
  AOI21_X1 U5442 ( .B1(n4380), .B2(n4379), .A(n4378), .ZN(n4383) );
  INV_X1 U5443 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4401) );
  NOR2_X1 U5444 ( .A1(n4401), .A2(n4381), .ZN(n6017) );
  OAI21_X1 U5445 ( .B1(n6017), .B2(n6760), .A(n4375), .ZN(n4382) );
  NAND2_X1 U5446 ( .A1(n4383), .A2(n4382), .ZN(U3181) );
  NOR2_X1 U5447 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6058) );
  OAI21_X1 U5448 ( .B1(n6058), .B2(D_C_N_REG_SCAN_IN), .A(n4375), .ZN(n4384)
         );
  OAI21_X1 U5449 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n4375), .A(n4384), .ZN(
        U2791) );
  AOI22_X1 U5450 ( .A1(n4385), .A2(REIP_REG_5__SCAN_IN), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n4375), .ZN(n4386) );
  OAI21_X1 U5451 ( .B1(n6168), .B2(n4387), .A(n4386), .ZN(U3187) );
  INV_X1 U5452 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6132) );
  AOI22_X1 U5453 ( .A1(n4398), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n4375), .ZN(n4388) );
  OAI21_X1 U5454 ( .B1(n6132), .B2(n4395), .A(n4388), .ZN(U3189) );
  AOI22_X1 U5455 ( .A1(n4398), .A2(REIP_REG_29__SCAN_IN), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n4375), .ZN(n4389) );
  OAI21_X1 U5456 ( .B1(n5158), .B2(n4400), .A(n4389), .ZN(U3212) );
  AOI22_X1 U5457 ( .A1(n4398), .A2(REIP_REG_5__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n4375), .ZN(n4390) );
  OAI21_X1 U5458 ( .B1(n6150), .B2(n4395), .A(n4390), .ZN(U3188) );
  INV_X1 U5459 ( .A(REIP_REG_10__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U5460 ( .A1(n4398), .A2(REIP_REG_9__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n4375), .ZN(n4391) );
  OAI21_X1 U5461 ( .B1(n4392), .B2(n4400), .A(n4391), .ZN(U3192) );
  INV_X1 U5462 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5361) );
  AOI22_X1 U5463 ( .A1(n4398), .A2(REIP_REG_8__SCAN_IN), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n4375), .ZN(n4393) );
  OAI21_X1 U5464 ( .B1(n5361), .B2(n4400), .A(n4393), .ZN(U3191) );
  INV_X1 U5465 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5682) );
  AOI22_X1 U5466 ( .A1(n4398), .A2(REIP_REG_7__SCAN_IN), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n4375), .ZN(n4394) );
  OAI21_X1 U5467 ( .B1(n5682), .B2(n4395), .A(n4394), .ZN(U3190) );
  INV_X1 U5468 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5646) );
  AOI22_X1 U5469 ( .A1(n4398), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n4375), .ZN(n4396) );
  OAI21_X1 U5470 ( .B1(n5646), .B2(n4400), .A(n4396), .ZN(U3195) );
  INV_X1 U5471 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5338) );
  AOI22_X1 U5472 ( .A1(n4398), .A2(REIP_REG_11__SCAN_IN), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n4375), .ZN(n4397) );
  OAI21_X1 U5473 ( .B1(n5338), .B2(n4400), .A(n4397), .ZN(U3194) );
  AOI22_X1 U5474 ( .A1(n4398), .A2(REIP_REG_10__SCAN_IN), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n4375), .ZN(n4399) );
  OAI21_X1 U5475 ( .B1(n5354), .B2(n4400), .A(n4399), .ZN(U3193) );
  INV_X1 U5476 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4403) );
  OAI21_X1 U5477 ( .B1(n4401), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n4402) );
  OAI21_X1 U5478 ( .B1(n6021), .B2(n4403), .A(n6582), .ZN(U2789) );
  INV_X1 U5479 ( .A(n4408), .ZN(n4405) );
  OAI22_X1 U5480 ( .A1(n4431), .A2(n4406), .B1(n4405), .B2(n4404), .ZN(n6055)
         );
  NOR2_X1 U5481 ( .A1(n3003), .A2(n4406), .ZN(n5174) );
  NOR2_X1 U5482 ( .A1(n6018), .A2(READY_N), .ZN(n4416) );
  INV_X1 U5483 ( .A(n4416), .ZN(n4407) );
  OAI21_X1 U5484 ( .B1(n5174), .B2(READY_N), .A(n4407), .ZN(n6613) );
  NOR2_X1 U5485 ( .A1(n6055), .A2(n6613), .ZN(n6550) );
  NOR2_X1 U5486 ( .A1(n6550), .A2(n6573), .ZN(n6061) );
  INV_X1 U5487 ( .A(MORE_REG_SCAN_IN), .ZN(n4414) );
  INV_X1 U5488 ( .A(n4445), .ZN(n4546) );
  AND2_X1 U5489 ( .A1(n4444), .A2(n6552), .ZN(n4558) );
  NAND2_X1 U5490 ( .A1(n4558), .A2(n4408), .ZN(n4409) );
  MUX2_X1 U5491 ( .A(n4546), .B(n4409), .S(n4528), .Z(n4410) );
  AOI21_X1 U5492 ( .B1(n4411), .B2(n4419), .A(n4410), .ZN(n6553) );
  INV_X1 U5493 ( .A(n6553), .ZN(n4412) );
  NAND2_X1 U5494 ( .A1(n6061), .A2(n4412), .ZN(n4413) );
  OAI21_X1 U5495 ( .B1(n6061), .B2(n4414), .A(n4413), .ZN(U3471) );
  INV_X1 U5496 ( .A(n6567), .ZN(n5148) );
  INV_X1 U5497 ( .A(n4415), .ZN(n4452) );
  MUX2_X1 U5498 ( .A(n4444), .B(n4445), .S(n4528), .Z(n4433) );
  OAI21_X1 U5499 ( .B1(n5144), .B2(n4213), .A(n4416), .ZN(n4418) );
  NAND2_X1 U5500 ( .A1(n4418), .A2(n4417), .ZN(n4430) );
  INV_X1 U5501 ( .A(n4419), .ZN(n4424) );
  INV_X1 U5502 ( .A(n4420), .ZN(n4422) );
  NAND2_X1 U5503 ( .A1(n4422), .A2(n4421), .ZN(n4423) );
  NAND2_X1 U5504 ( .A1(n4424), .A2(n4423), .ZN(n4532) );
  INV_X1 U5505 ( .A(n4425), .ZN(n4426) );
  NAND2_X1 U5506 ( .A1(n4532), .A2(n4426), .ZN(n4427) );
  OR2_X1 U5507 ( .A1(n4428), .A2(n4427), .ZN(n4429) );
  AOI21_X1 U5508 ( .B1(n4431), .B2(n4430), .A(n4429), .ZN(n4432) );
  INV_X1 U5509 ( .A(n6540), .ZN(n4435) );
  INV_X1 U5510 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6060) );
  NAND2_X1 U5511 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4734) );
  NAND2_X1 U5512 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4651), .ZN(n6586) );
  NOR2_X1 U5513 ( .A1(n6060), .A2(n6586), .ZN(n4434) );
  AOI21_X1 U5514 ( .B1(n4435), .B2(n6559), .A(n4434), .ZN(n6047) );
  NOR2_X1 U5515 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6588), .ZN(n4652) );
  INV_X1 U5516 ( .A(n4652), .ZN(n6587) );
  NAND2_X1 U5517 ( .A1(n6047), .A2(n6587), .ZN(n6054) );
  INV_X1 U5518 ( .A(n6054), .ZN(n5151) );
  AOI21_X1 U5519 ( .B1(n5148), .B2(n4452), .A(n5151), .ZN(n4456) );
  INV_X1 U5520 ( .A(n4438), .ZN(n4439) );
  AND3_X1 U5521 ( .A1(n4440), .A2(n4543), .A3(n4439), .ZN(n4441) );
  NAND2_X1 U5522 ( .A1(n6048), .A2(n4441), .ZN(n4442) );
  NOR2_X1 U5523 ( .A1(n4443), .A2(n4442), .ZN(n5146) );
  NAND2_X1 U5524 ( .A1(n4445), .A2(n4444), .ZN(n4710) );
  XNOR2_X1 U5525 ( .A(n4415), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4449)
         );
  INV_X1 U5526 ( .A(n5144), .ZN(n4447) );
  XNOR2_X1 U5527 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4446) );
  OAI22_X1 U5528 ( .A1(n4447), .A2(n4446), .B1(n4712), .B2(n4449), .ZN(n4448)
         );
  AOI21_X1 U5529 ( .B1(n4710), .B2(n4449), .A(n4448), .ZN(n4450) );
  OAI21_X1 U5530 ( .B1(n4437), .B2(n5146), .A(n4450), .ZN(n4705) );
  INV_X1 U5531 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5905) );
  INV_X1 U5532 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4451) );
  INV_X1 U5533 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U5534 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4451), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4573), .ZN(n5150) );
  NOR3_X1 U5535 ( .A1(n5170), .A2(n5905), .A3(n5150), .ZN(n4454) );
  NOR3_X1 U5536 ( .A1(n6567), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4452), 
        .ZN(n4453) );
  AOI211_X1 U5537 ( .C1(n6049), .C2(n4705), .A(n4454), .B(n4453), .ZN(n4455)
         );
  OAI22_X1 U5538 ( .A1(n4456), .A2(n4436), .B1(n4455), .B2(n5151), .ZN(U3459)
         );
  NAND2_X1 U5539 ( .A1(n5144), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6538) );
  INV_X1 U5540 ( .A(n6049), .ZN(n5925) );
  OAI21_X1 U5541 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6567), .A(n6054), 
        .ZN(n5141) );
  INV_X1 U5542 ( .A(n5146), .ZN(n4720) );
  INV_X1 U5543 ( .A(n5142), .ZN(n4458) );
  AOI22_X1 U5544 ( .A1(n6421), .A2(n4720), .B1(n4458), .B2(n4457), .ZN(n6539)
         );
  OAI22_X1 U5545 ( .A1(n6539), .A2(n5925), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5170), .ZN(n4459) );
  OAI22_X1 U5546 ( .A1(n5141), .A2(n4459), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6054), .ZN(n4460) );
  OAI21_X1 U5547 ( .B1(n6538), .B2(n5925), .A(n4460), .ZN(U3461) );
  XNOR2_X1 U5548 ( .A(n4461), .B(n3003), .ZN(n4551) );
  INV_X1 U5549 ( .A(n4551), .ZN(n4463) );
  INV_X1 U5550 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4462) );
  OAI222_X1 U5551 ( .A1(n4463), .A2(n5428), .B1(n6195), .B2(n4462), .C1(n2970), 
        .C2(n4590), .ZN(U2858) );
  INV_X1 U5552 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U5553 ( .A1(n4495), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4465) );
  NAND2_X1 U5554 ( .A1(n6243), .A2(DATAI_11_), .ZN(n4504) );
  OAI211_X1 U5555 ( .C1(n4526), .C2(n4612), .A(n4465), .B(n4504), .ZN(U2935)
         );
  NAND2_X1 U5556 ( .A1(n4495), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4466) );
  NAND2_X1 U5557 ( .A1(n6243), .A2(DATAI_7_), .ZN(n4468) );
  OAI211_X1 U5558 ( .C1(n4526), .C2(n3571), .A(n4466), .B(n4468), .ZN(U2946)
         );
  NAND2_X1 U5559 ( .A1(n4495), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U5560 ( .A1(n6243), .A2(DATAI_5_), .ZN(n4520) );
  OAI211_X1 U5561 ( .C1(n4526), .C2(n3526), .A(n4467), .B(n4520), .ZN(U2944)
         );
  INV_X1 U5562 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4610) );
  NAND2_X1 U5563 ( .A1(n4495), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4469) );
  OAI211_X1 U5564 ( .C1(n4526), .C2(n4610), .A(n4469), .B(n4468), .ZN(U2931)
         );
  INV_X1 U5565 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6674) );
  NAND2_X1 U5566 ( .A1(n4495), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4470) );
  NAND2_X1 U5567 ( .A1(n6243), .A2(DATAI_13_), .ZN(n4508) );
  OAI211_X1 U5568 ( .C1(n4526), .C2(n6674), .A(n4470), .B(n4508), .ZN(U2937)
         );
  INV_X1 U5569 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U5570 ( .A1(n4495), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U5571 ( .A1(n6243), .A2(DATAI_3_), .ZN(n4506) );
  OAI211_X1 U5572 ( .C1(n4526), .C2(n6226), .A(n4471), .B(n4506), .ZN(U2942)
         );
  INV_X1 U5573 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U5574 ( .A1(n4495), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4472) );
  NAND2_X1 U5575 ( .A1(n6243), .A2(DATAI_2_), .ZN(n4510) );
  OAI211_X1 U5576 ( .C1(n4526), .C2(n6228), .A(n4472), .B(n4510), .ZN(U2941)
         );
  INV_X1 U5577 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U5578 ( .A1(n4495), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4473) );
  NAND2_X1 U5579 ( .A1(n6243), .A2(DATAI_1_), .ZN(n4518) );
  OAI211_X1 U5580 ( .C1(n4526), .C2(n6231), .A(n4473), .B(n4518), .ZN(U2940)
         );
  NAND2_X1 U5581 ( .A1(n4495), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4474) );
  NAND2_X1 U5582 ( .A1(n6243), .A2(DATAI_10_), .ZN(n4512) );
  OAI211_X1 U5583 ( .C1(n4526), .C2(n3896), .A(n4474), .B(n4512), .ZN(U2934)
         );
  INV_X1 U5584 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U5585 ( .A1(n4495), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U5586 ( .A1(n6243), .A2(DATAI_6_), .ZN(n4502) );
  OAI211_X1 U5587 ( .C1(n4526), .C2(n4598), .A(n4475), .B(n4502), .ZN(U2930)
         );
  INV_X1 U5588 ( .A(n4476), .ZN(n4480) );
  INV_X1 U5589 ( .A(n4477), .ZN(n4479) );
  OAI21_X1 U5590 ( .B1(n4480), .B2(n4479), .A(n4478), .ZN(n5404) );
  NOR2_X1 U5591 ( .A1(n4481), .A2(n4672), .ZN(n4482) );
  INV_X1 U5592 ( .A(n4482), .ZN(n4483) );
  INV_X1 U5593 ( .A(DATAI_0_), .ZN(n6713) );
  INV_X1 U5594 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6234) );
  OAI222_X1 U5595 ( .A1(n5404), .A2(n6776), .B1(n5491), .B2(n6713), .C1(n6234), 
        .C2(n5489), .ZN(U2891) );
  INV_X1 U5596 ( .A(DATAI_1_), .ZN(n4692) );
  OAI222_X1 U5597 ( .A1(n4590), .A2(n6776), .B1(n5491), .B2(n4692), .C1(n5489), 
        .C2(n6231), .ZN(U2890) );
  OR2_X1 U5598 ( .A1(n6246), .A2(n4484), .ZN(n4485) );
  INV_X1 U5599 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6752) );
  NOR2_X1 U5600 ( .A1(n6287), .A2(n6752), .ZN(n5908) );
  AOI21_X1 U5601 ( .B1(n4485), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5908), 
        .ZN(n4488) );
  OR2_X1 U5602 ( .A1(n4486), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5910)
         );
  NAND3_X1 U5603 ( .A1(n4329), .A2(n5910), .A3(n5911), .ZN(n4487) );
  OAI211_X1 U5604 ( .C1(n5404), .C2(n6258), .A(n4488), .B(n4487), .ZN(U2986)
         );
  INV_X1 U5605 ( .A(n4490), .ZN(n4493) );
  NAND3_X1 U5606 ( .A1(n4493), .A2(n4492), .A3(n4491), .ZN(n4494) );
  NAND2_X1 U5607 ( .A1(n4489), .A2(n4494), .ZN(n5398) );
  INV_X1 U5608 ( .A(DATAI_2_), .ZN(n4680) );
  OAI222_X1 U5609 ( .A1(n5398), .A2(n6776), .B1(n5491), .B2(n4680), .C1(n5489), 
        .C2(n6228), .ZN(U2889) );
  INV_X1 U5610 ( .A(DATAI_12_), .ZN(n4498) );
  INV_X1 U5611 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6643) );
  OAI222_X1 U5612 ( .A1(n4498), .A2(n4497), .B1(n4499), .B2(n6643), .C1(n4496), 
        .C2(n4526), .ZN(U2936) );
  NAND2_X1 U5613 ( .A1(n6243), .A2(DATAI_0_), .ZN(n4516) );
  NAND2_X1 U5614 ( .A1(n6242), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4500) );
  OAI211_X1 U5615 ( .C1(n4526), .C2(n6234), .A(n4516), .B(n4500), .ZN(U2939)
         );
  INV_X1 U5616 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U5617 ( .A1(n6243), .A2(DATAI_4_), .ZN(n4514) );
  NAND2_X1 U5618 ( .A1(n6242), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4501) );
  OAI211_X1 U5619 ( .C1(n4526), .C2(n6224), .A(n4514), .B(n4501), .ZN(U2943)
         );
  NAND2_X1 U5620 ( .A1(n6242), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4503) );
  OAI211_X1 U5621 ( .C1(n4526), .C2(n3545), .A(n4503), .B(n4502), .ZN(U2945)
         );
  INV_X1 U5622 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U5623 ( .A1(n6242), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4505) );
  OAI211_X1 U5624 ( .C1(n4526), .C2(n6679), .A(n4505), .B(n4504), .ZN(U2950)
         );
  NAND2_X1 U5625 ( .A1(n6242), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4507) );
  OAI211_X1 U5626 ( .C1(n4526), .C2(n3757), .A(n4507), .B(n4506), .ZN(U2927)
         );
  INV_X1 U5627 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U5628 ( .A1(n6242), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4509) );
  OAI211_X1 U5629 ( .C1(n4526), .C2(n6208), .A(n4509), .B(n4508), .ZN(U2952)
         );
  INV_X1 U5630 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U5631 ( .A1(n6242), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4511) );
  OAI211_X1 U5632 ( .C1(n4526), .C2(n4605), .A(n4511), .B(n4510), .ZN(U2926)
         );
  INV_X1 U5633 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U5634 ( .A1(n6242), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4513) );
  OAI211_X1 U5635 ( .C1(n4526), .C2(n6693), .A(n4513), .B(n4512), .ZN(U2949)
         );
  INV_X1 U5636 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6687) );
  NAND2_X1 U5637 ( .A1(n6242), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4515) );
  OAI211_X1 U5638 ( .C1(n4526), .C2(n6687), .A(n4515), .B(n4514), .ZN(U2928)
         );
  INV_X1 U5639 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U5640 ( .A1(n6242), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4517) );
  OAI211_X1 U5641 ( .C1(n4526), .C2(n4616), .A(n4517), .B(n4516), .ZN(U2924)
         );
  INV_X1 U5642 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U5643 ( .A1(n6242), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4519) );
  OAI211_X1 U5644 ( .C1(n4526), .C2(n4618), .A(n4519), .B(n4518), .ZN(U2925)
         );
  INV_X1 U5645 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4601) );
  NAND2_X1 U5646 ( .A1(n6242), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4521) );
  OAI211_X1 U5647 ( .C1(n4526), .C2(n4601), .A(n4521), .B(n4520), .ZN(U2929)
         );
  INV_X1 U5648 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5649 ( .A1(n6242), .A2(UWORD_REG_8__SCAN_IN), .B1(n6243), .B2(
        DATAI_8_), .ZN(n4522) );
  OAI21_X1 U5650 ( .B1(n4603), .B2(n4526), .A(n4522), .ZN(U2932) );
  INV_X1 U5651 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6204) );
  AOI22_X1 U5652 ( .A1(n6242), .A2(LWORD_REG_15__SCAN_IN), .B1(n6243), .B2(
        DATAI_15_), .ZN(n4523) );
  OAI21_X1 U5653 ( .B1(n6204), .B2(n4526), .A(n4523), .ZN(U2954) );
  AOI22_X1 U5654 ( .A1(n6242), .A2(UWORD_REG_14__SCAN_IN), .B1(n6243), .B2(
        DATAI_14_), .ZN(n4524) );
  OAI21_X1 U5655 ( .B1(n4130), .B2(n4526), .A(n4524), .ZN(U2938) );
  INV_X1 U5656 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4607) );
  AOI22_X1 U5657 ( .A1(n6242), .A2(UWORD_REG_9__SCAN_IN), .B1(n6243), .B2(
        DATAI_9_), .ZN(n4525) );
  OAI21_X1 U5658 ( .B1(n4607), .B2(n4526), .A(n4525), .ZN(U2933) );
  NAND2_X1 U5659 ( .A1(n4528), .A2(n4527), .ZN(n4533) );
  OAI211_X1 U5660 ( .C1(n4691), .C2(n4563), .A(n4530), .B(n4529), .ZN(n4531)
         );
  NAND3_X1 U5661 ( .A1(n4533), .A2(n4532), .A3(n4531), .ZN(n4534) );
  NAND2_X1 U5662 ( .A1(n4534), .A2(n6559), .ZN(n4542) );
  NAND2_X1 U5663 ( .A1(n4535), .A2(n6611), .ZN(n4538) );
  OAI211_X1 U5664 ( .C1(n4543), .C2(n4538), .A(n4537), .B(n4536), .ZN(n4539)
         );
  NAND2_X1 U5665 ( .A1(n4539), .A2(n4679), .ZN(n4540) );
  OR2_X1 U5666 ( .A1(n4543), .A2(n6614), .ZN(n6562) );
  OAI21_X1 U5667 ( .B1(n4555), .B2(n4544), .A(n6562), .ZN(n4545) );
  NOR2_X1 U5668 ( .A1(n6287), .A2(n5372), .ZN(n4584) );
  OR2_X1 U5669 ( .A1(n4560), .A2(n6247), .ZN(n5906) );
  INV_X1 U5670 ( .A(n4547), .ZN(n4548) );
  NAND2_X1 U5671 ( .A1(n4560), .A2(n4548), .ZN(n4572) );
  OAI21_X1 U5672 ( .B1(n5870), .B2(n5905), .A(n6039), .ZN(n4549) );
  MUX2_X1 U5673 ( .A(n5133), .B(n4549), .S(n4573), .Z(n4550) );
  AOI211_X1 U5674 ( .C1(n6300), .C2(n4551), .A(n4584), .B(n4550), .ZN(n4562)
         );
  OR2_X1 U5675 ( .A1(n4553), .A2(n4552), .ZN(n4587) );
  OR2_X1 U5676 ( .A1(n4555), .A2(n4554), .ZN(n4556) );
  NAND4_X1 U5677 ( .A1(n6048), .A2(n4558), .A3(n4557), .A4(n4556), .ZN(n4559)
         );
  NAND3_X1 U5678 ( .A1(n4587), .A2(n4586), .A3(n6304), .ZN(n4561) );
  NAND2_X1 U5679 ( .A1(n4562), .A2(n4561), .ZN(U3017) );
  INV_X1 U5680 ( .A(n6562), .ZN(n4564) );
  OAI21_X1 U5681 ( .B1(n5144), .B2(n4564), .A(n4563), .ZN(n4565) );
  NAND2_X1 U5682 ( .A1(n4651), .A2(n6566), .ZN(n6214) );
  NOR2_X4 U5683 ( .A1(n6212), .A2(n6612), .ZN(n6222) );
  AOI22_X1 U5684 ( .A1(DATAO_REG_20__SCAN_IN), .A2(n6222), .B1(n6229), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4567) );
  OAI21_X1 U5685 ( .B1(n6687), .B2(n6201), .A(n4567), .ZN(U2903) );
  NAND2_X1 U5686 ( .A1(n4569), .A2(n4568), .ZN(n4571) );
  XNOR2_X1 U5687 ( .A(n4571), .B(n4570), .ZN(n4596) );
  INV_X1 U5688 ( .A(n4572), .ZN(n4575) );
  OR2_X1 U5689 ( .A1(n5872), .A2(n4575), .ZN(n5700) );
  NAND2_X1 U5690 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5109) );
  AOI22_X1 U5691 ( .A1(n5700), .A2(n5109), .B1(n6277), .B2(n5133), .ZN(n4640)
         );
  INV_X1 U5692 ( .A(n4640), .ZN(n5093) );
  NOR3_X1 U5693 ( .A1(n6277), .A2(n5905), .A3(n4573), .ZN(n4574) );
  OAI21_X1 U5694 ( .B1(n5093), .B2(n4574), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4582) );
  NAND2_X1 U5695 ( .A1(n4575), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5874)
         );
  NAND2_X1 U5696 ( .A1(n5874), .A2(n6039), .ZN(n5699) );
  NAND3_X1 U5697 ( .A1(n5699), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n3180), 
        .ZN(n4580) );
  NOR2_X1 U5698 ( .A1(n4577), .A2(n4576), .ZN(n4578) );
  NOR2_X1 U5699 ( .A1(n4578), .A2(n4624), .ZN(n5396) );
  NOR2_X1 U5700 ( .A1(n6287), .A2(n5390), .ZN(n4591) );
  AOI21_X1 U5701 ( .B1(n6300), .B2(n5396), .A(n4591), .ZN(n4579) );
  AOI21_X1 U5702 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n5092) );
  NAND2_X1 U5703 ( .A1(n5114), .A2(n5092), .ZN(n4639) );
  AND3_X1 U5704 ( .A1(n4580), .A2(n4579), .A3(n4639), .ZN(n4581) );
  OAI211_X1 U5705 ( .C1(n4596), .C2(n5903), .A(n4582), .B(n4581), .ZN(U3016)
         );
  NOR2_X1 U5706 ( .A1(n6271), .A2(n4585), .ZN(n4583) );
  AOI211_X1 U5707 ( .C1(n6266), .C2(n4585), .A(n4584), .B(n4583), .ZN(n4589)
         );
  NAND3_X1 U5708 ( .A1(n4587), .A2(n4586), .A3(n4329), .ZN(n4588) );
  OAI211_X1 U5709 ( .C1(n6258), .C2(n4590), .A(n4589), .B(n4588), .ZN(U2985)
         );
  INV_X1 U5710 ( .A(n5398), .ZN(n4594) );
  AOI21_X1 U5711 ( .B1(n6246), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4591), 
        .ZN(n4592) );
  OAI21_X1 U5712 ( .B1(n5384), .B2(n6254), .A(n4592), .ZN(n4593) );
  AOI21_X1 U5713 ( .B1(n4594), .B2(n6265), .A(n4593), .ZN(n4595) );
  OAI21_X1 U5714 ( .B1(n4596), .B2(n6256), .A(n4595), .ZN(U2984) );
  AOI22_X1 U5715 ( .A1(n6229), .A2(UWORD_REG_6__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4597) );
  OAI21_X1 U5716 ( .B1(n4598), .B2(n6201), .A(n4597), .ZN(U2901) );
  AOI22_X1 U5717 ( .A1(n6229), .A2(UWORD_REG_3__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4599) );
  OAI21_X1 U5718 ( .B1(n3757), .B2(n6201), .A(n4599), .ZN(U2904) );
  AOI22_X1 U5719 ( .A1(n6229), .A2(UWORD_REG_5__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4600) );
  OAI21_X1 U5720 ( .B1(n4601), .B2(n6201), .A(n4600), .ZN(U2902) );
  AOI22_X1 U5721 ( .A1(n6229), .A2(UWORD_REG_8__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4602) );
  OAI21_X1 U5722 ( .B1(n4603), .B2(n6201), .A(n4602), .ZN(U2899) );
  AOI22_X1 U5723 ( .A1(n6229), .A2(UWORD_REG_2__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4604) );
  OAI21_X1 U5724 ( .B1(n4605), .B2(n6201), .A(n4604), .ZN(U2905) );
  AOI22_X1 U5725 ( .A1(n6229), .A2(UWORD_REG_9__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4606) );
  OAI21_X1 U5726 ( .B1(n4607), .B2(n6201), .A(n4606), .ZN(U2898) );
  AOI22_X1 U5727 ( .A1(n6229), .A2(UWORD_REG_13__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4608) );
  OAI21_X1 U5728 ( .B1(n6674), .B2(n6201), .A(n4608), .ZN(U2894) );
  AOI22_X1 U5729 ( .A1(n6229), .A2(UWORD_REG_7__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4609) );
  OAI21_X1 U5730 ( .B1(n4610), .B2(n6201), .A(n4609), .ZN(U2900) );
  AOI22_X1 U5731 ( .A1(n6229), .A2(UWORD_REG_11__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4611) );
  OAI21_X1 U5732 ( .B1(n4612), .B2(n6201), .A(n4611), .ZN(U2896) );
  AOI22_X1 U5733 ( .A1(n6229), .A2(UWORD_REG_10__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4613) );
  OAI21_X1 U5734 ( .B1(n3896), .B2(n6201), .A(n4613), .ZN(U2897) );
  AOI22_X1 U5735 ( .A1(n6612), .A2(UWORD_REG_14__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4614) );
  OAI21_X1 U5736 ( .B1(n4130), .B2(n6201), .A(n4614), .ZN(U2893) );
  AOI22_X1 U5737 ( .A1(n6612), .A2(UWORD_REG_0__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4615) );
  OAI21_X1 U5738 ( .B1(n4616), .B2(n6201), .A(n4615), .ZN(U2907) );
  AOI22_X1 U5739 ( .A1(n6612), .A2(UWORD_REG_1__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4617) );
  OAI21_X1 U5740 ( .B1(n4618), .B2(n6201), .A(n4617), .ZN(U2906) );
  OAI21_X1 U5741 ( .B1(n4619), .B2(n4621), .A(n4620), .ZN(n4740) );
  INV_X1 U5742 ( .A(DATAI_4_), .ZN(n4667) );
  OAI222_X1 U5743 ( .A1(n4740), .A2(n6776), .B1(n5491), .B2(n4667), .C1(n6224), 
        .C2(n5489), .ZN(U2887) );
  AOI21_X1 U5744 ( .B1(n4622), .B2(n4489), .A(n4619), .ZN(n4637) );
  INV_X1 U5745 ( .A(n4637), .ZN(n5383) );
  NOR2_X1 U5746 ( .A1(n4624), .A2(n4623), .ZN(n4625) );
  NOR2_X1 U5747 ( .A1(n3036), .A2(n4625), .ZN(n5376) );
  AOI22_X1 U5748 ( .A1(n6192), .A2(n5376), .B1(n5452), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4626) );
  OAI21_X1 U5749 ( .B1(n5383), .B2(n2970), .A(n4626), .ZN(U2856) );
  OAI21_X1 U5750 ( .B1(n3036), .B2(n4627), .A(n5105), .ZN(n6171) );
  INV_X1 U5751 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6737) );
  OAI222_X1 U5752 ( .A1(n6171), .A2(n5428), .B1(n6195), .B2(n6737), .C1(n2970), 
        .C2(n4740), .ZN(U2855) );
  INV_X1 U5753 ( .A(DATAI_3_), .ZN(n4686) );
  OAI222_X1 U5754 ( .A1(n5383), .A2(n6776), .B1(n5491), .B2(n4686), .C1(n5489), 
        .C2(n6226), .ZN(U2888) );
  INV_X1 U5755 ( .A(n5396), .ZN(n4628) );
  INV_X1 U5756 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6657) );
  OAI222_X1 U5757 ( .A1(n4628), .A2(n5428), .B1(n6195), .B2(n6657), .C1(n2970), 
        .C2(n5398), .ZN(U2857) );
  OR2_X1 U5758 ( .A1(n4629), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4631)
         );
  NAND2_X1 U5759 ( .A1(n4631), .A2(n4630), .ZN(n5904) );
  OAI222_X1 U5760 ( .A1(n5904), .A2(n5428), .B1(n6195), .B2(n4632), .C1(n5404), 
        .C2(n2970), .ZN(U2859) );
  XNOR2_X1 U5761 ( .A(n4634), .B(n4633), .ZN(n4646) );
  NOR2_X1 U5762 ( .A1(n6287), .A2(n4368), .ZN(n4643) );
  AOI21_X1 U5763 ( .B1(n6246), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4643), 
        .ZN(n4635) );
  OAI21_X1 U5764 ( .B1(n5374), .B2(n6254), .A(n4635), .ZN(n4636) );
  AOI21_X1 U5765 ( .B1(n4637), .B2(n6265), .A(n4636), .ZN(n4638) );
  OAI21_X1 U5766 ( .B1(n4646), .B2(n6256), .A(n4638), .ZN(U2983) );
  NAND2_X1 U5767 ( .A1(n4640), .A2(n4639), .ZN(n4747) );
  INV_X1 U5768 ( .A(n5109), .ZN(n4641) );
  AOI21_X1 U5769 ( .B1(n4641), .B2(n5699), .A(n5114), .ZN(n5095) );
  NOR2_X1 U5770 ( .A1(n5092), .A2(n5095), .ZN(n4744) );
  AOI22_X1 U5771 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4747), .B1(n4744), 
        .B2(n4642), .ZN(n4645) );
  AOI21_X1 U5772 ( .B1(n6300), .B2(n5376), .A(n4643), .ZN(n4644) );
  OAI211_X1 U5773 ( .C1(n4646), .C2(n5903), .A(n4645), .B(n4644), .ZN(U3015)
         );
  NAND2_X1 U5774 ( .A1(n4620), .A2(n4648), .ZN(n4649) );
  AND2_X1 U5775 ( .A1(n4647), .A2(n4649), .ZN(n6264) );
  INV_X1 U5776 ( .A(n6264), .ZN(n4650) );
  INV_X1 U5777 ( .A(DATAI_5_), .ZN(n6675) );
  OAI222_X1 U5778 ( .A1(n4650), .A2(n6776), .B1(n5491), .B2(n6675), .C1(n5489), 
        .C2(n3526), .ZN(U2886) );
  INV_X1 U5779 ( .A(n6516), .ZN(n5022) );
  NAND3_X1 U5780 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6547), .A3(n4916), .ZN(n6386) );
  NOR2_X1 U5781 ( .A1(n6309), .A2(n6386), .ZN(n4655) );
  INV_X1 U5782 ( .A(n4655), .ZN(n4704) );
  INV_X1 U5783 ( .A(n4751), .ZN(n4913) );
  OAI21_X1 U5784 ( .B1(n6428), .B2(n4913), .A(n6419), .ZN(n4660) );
  AND2_X1 U5785 ( .A1(n4654), .A2(n6421), .ZN(n4996) );
  INV_X1 U5786 ( .A(n4341), .ZN(n5917) );
  NAND2_X1 U5787 ( .A1(n5917), .A2(n4437), .ZN(n4752) );
  INV_X1 U5788 ( .A(n4752), .ZN(n6387) );
  AOI21_X1 U5789 ( .B1(n4996), .B2(n6387), .A(n4655), .ZN(n4659) );
  INV_X1 U5790 ( .A(n4659), .ZN(n4658) );
  AOI21_X1 U5791 ( .B1(n6476), .B2(n6386), .A(n4840), .ZN(n4657) );
  OAI21_X1 U5792 ( .B1(n4660), .B2(n4658), .A(n4657), .ZN(n4700) );
  OAI22_X1 U5793 ( .A1(n4660), .A2(n4659), .B1(n5978), .B2(n6386), .ZN(n4699)
         );
  AOI22_X1 U5794 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4700), .B1(n6515), 
        .B2(n4699), .ZN(n4666) );
  INV_X1 U5795 ( .A(DATAI_21_), .ZN(n4661) );
  NOR2_X1 U5796 ( .A1(n6258), .A2(n4661), .ZN(n6517) );
  INV_X1 U5797 ( .A(n4662), .ZN(n4663) );
  NAND2_X1 U5798 ( .A1(n4663), .A2(n5041), .ZN(n5929) );
  NAND2_X1 U5799 ( .A1(n4662), .A2(n5041), .ZN(n4920) );
  INV_X1 U5800 ( .A(DATAI_29_), .ZN(n4664) );
  NOR2_X1 U5801 ( .A1(n6258), .A2(n4664), .ZN(n6454) );
  AOI22_X1 U5802 ( .A1(n6517), .A2(n6007), .B1(n6414), .B2(n6454), .ZN(n4665)
         );
  OAI211_X1 U5803 ( .C1(n5022), .C2(n4704), .A(n4666), .B(n4665), .ZN(U3097)
         );
  INV_X1 U5804 ( .A(n6510), .ZN(n5038) );
  AOI22_X1 U5805 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4700), .B1(n6509), 
        .B2(n4699), .ZN(n4671) );
  INV_X1 U5806 ( .A(DATAI_20_), .ZN(n4668) );
  NOR2_X1 U5807 ( .A1(n6258), .A2(n4668), .ZN(n6511) );
  INV_X1 U5808 ( .A(DATAI_28_), .ZN(n4669) );
  NOR2_X1 U5809 ( .A1(n6258), .A2(n4669), .ZN(n6450) );
  AOI22_X1 U5810 ( .A1(n6511), .A2(n6007), .B1(n6414), .B2(n6450), .ZN(n4670)
         );
  OAI211_X1 U5811 ( .C1(n5038), .C2(n4704), .A(n4671), .B(n4670), .ZN(U3096)
         );
  INV_X1 U5812 ( .A(DATAI_7_), .ZN(n5040) );
  AOI22_X1 U5813 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4700), .B1(n6528), 
        .B2(n4699), .ZN(n4675) );
  NAND2_X1 U5814 ( .A1(n6265), .A2(DATAI_23_), .ZN(n6469) );
  INV_X1 U5815 ( .A(n6469), .ZN(n6532) );
  INV_X1 U5816 ( .A(DATAI_31_), .ZN(n4673) );
  NOR2_X1 U5817 ( .A1(n6258), .A2(n4673), .ZN(n6463) );
  AOI22_X1 U5818 ( .A1(n6532), .A2(n6007), .B1(n6414), .B2(n6463), .ZN(n4674)
         );
  OAI211_X1 U5819 ( .C1(n5018), .C2(n4704), .A(n4675), .B(n4674), .ZN(U3099)
         );
  INV_X1 U5820 ( .A(n6522), .ZN(n5014) );
  INV_X1 U5821 ( .A(DATAI_6_), .ZN(n4837) );
  AOI22_X1 U5822 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4700), .B1(n6521), 
        .B2(n4699), .ZN(n4678) );
  NAND2_X1 U5823 ( .A1(n6265), .A2(DATAI_22_), .ZN(n6461) );
  INV_X1 U5824 ( .A(n6461), .ZN(n6523) );
  INV_X1 U5825 ( .A(DATAI_30_), .ZN(n4676) );
  NOR2_X1 U5826 ( .A1(n6258), .A2(n4676), .ZN(n6457) );
  AOI22_X1 U5827 ( .A1(n6523), .A2(n6007), .B1(n6414), .B2(n6457), .ZN(n4677)
         );
  OAI211_X1 U5828 ( .C1(n5014), .C2(n4704), .A(n4678), .B(n4677), .ZN(U3098)
         );
  INV_X1 U5829 ( .A(n6498), .ZN(n5026) );
  AOI22_X1 U5830 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4700), .B1(n6497), 
        .B2(n4699), .ZN(n4684) );
  INV_X1 U5831 ( .A(DATAI_18_), .ZN(n4681) );
  NOR2_X1 U5832 ( .A1(n6258), .A2(n4681), .ZN(n6499) );
  INV_X1 U5833 ( .A(DATAI_26_), .ZN(n4682) );
  NOR2_X1 U5834 ( .A1(n6258), .A2(n4682), .ZN(n6442) );
  AOI22_X1 U5835 ( .A1(n6499), .A2(n6007), .B1(n6414), .B2(n6442), .ZN(n4683)
         );
  OAI211_X1 U5836 ( .C1(n5026), .C2(n4704), .A(n4684), .B(n4683), .ZN(U3094)
         );
  AOI22_X1 U5838 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4700), .B1(n6503), 
        .B2(n4699), .ZN(n4690) );
  INV_X1 U5839 ( .A(DATAI_19_), .ZN(n4687) );
  NOR2_X1 U5840 ( .A1(n6258), .A2(n4687), .ZN(n6505) );
  INV_X1 U5841 ( .A(DATAI_27_), .ZN(n4688) );
  NOR2_X1 U5842 ( .A1(n6258), .A2(n4688), .ZN(n6446) );
  AOI22_X1 U5843 ( .A1(n6505), .A2(n6007), .B1(n6414), .B2(n6446), .ZN(n4689)
         );
  OAI211_X1 U5844 ( .C1(n6504), .C2(n4704), .A(n4690), .B(n4689), .ZN(U3095)
         );
  AOI22_X1 U5845 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4700), .B1(n6491), 
        .B2(n4699), .ZN(n4696) );
  INV_X1 U5846 ( .A(DATAI_17_), .ZN(n4693) );
  NOR2_X1 U5847 ( .A1(n6258), .A2(n4693), .ZN(n6493) );
  INV_X1 U5848 ( .A(DATAI_25_), .ZN(n4694) );
  NOR2_X1 U5849 ( .A1(n6258), .A2(n4694), .ZN(n6438) );
  AOI22_X1 U5850 ( .A1(n6493), .A2(n6007), .B1(n6414), .B2(n6438), .ZN(n4695)
         );
  OAI211_X1 U5851 ( .C1(n5010), .C2(n4704), .A(n4696), .B(n4695), .ZN(U3093)
         );
  INV_X1 U5852 ( .A(n4697), .ZN(n4698) );
  NAND2_X1 U5853 ( .A1(n4698), .A2(n4537), .ZN(n5006) );
  AOI22_X1 U5854 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4700), .B1(n6474), 
        .B2(n4699), .ZN(n4703) );
  INV_X1 U5855 ( .A(DATAI_24_), .ZN(n6714) );
  NOR2_X1 U5856 ( .A1(n6258), .A2(n6714), .ZN(n6435) );
  INV_X1 U5857 ( .A(DATAI_16_), .ZN(n4701) );
  NOR2_X1 U5858 ( .A1(n6258), .A2(n4701), .ZN(n6487) );
  AOI22_X1 U5859 ( .A1(n6435), .A2(n6414), .B1(n6007), .B2(n6487), .ZN(n4702)
         );
  OAI211_X1 U5860 ( .C1(n4704), .C2(n5006), .A(n4703), .B(n4702), .ZN(U3092)
         );
  MUX2_X1 U5861 ( .A(n4705), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n6540), 
        .Z(n6546) );
  NAND2_X1 U5862 ( .A1(n6546), .A2(n5170), .ZN(n4722) );
  MUX2_X1 U5863 ( .A(n4706), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4415), 
        .Z(n4708) );
  NOR2_X1 U5864 ( .A1(n4708), .A2(n4707), .ZN(n4709) );
  NAND2_X1 U5865 ( .A1(n4710), .A2(n4709), .ZN(n4718) );
  XNOR2_X1 U5866 ( .A(n4711), .B(n3481), .ZN(n4716) );
  INV_X1 U5867 ( .A(n4712), .ZN(n4715) );
  AOI21_X1 U5868 ( .B1(n4415), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4714) );
  NOR2_X1 U5869 ( .A1(n3314), .A2(n4714), .ZN(n5923) );
  AOI22_X1 U5870 ( .A1(n5144), .A2(n4716), .B1(n4715), .B2(n5923), .ZN(n4717)
         );
  NAND2_X1 U5871 ( .A1(n4718), .A2(n4717), .ZN(n4719) );
  AOI21_X1 U5872 ( .B1(n4654), .B2(n4720), .A(n4719), .ZN(n5926) );
  MUX2_X1 U5873 ( .A(n5926), .B(n3481), .S(n6540), .Z(n6548) );
  NAND2_X1 U5874 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6060), .ZN(n4724) );
  INV_X1 U5875 ( .A(n4707), .ZN(n4721) );
  OAI22_X1 U5876 ( .A1(n4722), .A2(n6548), .B1(n4724), .B2(n4721), .ZN(n6556)
         );
  INV_X1 U5877 ( .A(n6556), .ZN(n4732) );
  NAND2_X1 U5878 ( .A1(n6540), .A2(n5170), .ZN(n4725) );
  NAND2_X1 U5879 ( .A1(n4725), .A2(n4724), .ZN(n4731) );
  INV_X1 U5880 ( .A(n4727), .ZN(n6479) );
  NOR2_X1 U5881 ( .A1(n3190), .A2(n6479), .ZN(n4728) );
  XNOR2_X1 U5882 ( .A(n4728), .B(n6053), .ZN(n6176) );
  NOR2_X1 U5883 ( .A1(n6048), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4729) );
  AND2_X1 U5884 ( .A1(n6176), .A2(n4729), .ZN(n4730) );
  AOI21_X1 U5885 ( .B1(n4731), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n4730), 
        .ZN(n6554) );
  OAI21_X1 U5886 ( .B1(n4732), .B2(n2981), .A(n6554), .ZN(n4735) );
  NOR2_X1 U5887 ( .A1(n4735), .A2(FLUSH_REG_SCAN_IN), .ZN(n4733) );
  NOR2_X1 U5888 ( .A1(n4735), .A2(n4734), .ZN(n6565) );
  INV_X1 U5889 ( .A(n6421), .ZN(n5046) );
  NOR2_X1 U5890 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5170), .ZN(n6591) );
  OAI22_X1 U5891 ( .A1(n4662), .A2(n6476), .B1(n5046), .B2(n6591), .ZN(n4736)
         );
  OAI21_X1 U5892 ( .B1(n6565), .B2(n4736), .A(n6599), .ZN(n4737) );
  OAI21_X1 U5893 ( .B1(n6599), .B2(n6309), .A(n4737), .ZN(U3465) );
  XNOR2_X1 U5894 ( .A(n4739), .B(n4738), .ZN(n4750) );
  INV_X1 U5895 ( .A(n4740), .ZN(n6183) );
  NOR2_X1 U5896 ( .A1(n6287), .A2(n6168), .ZN(n4746) );
  AOI21_X1 U5897 ( .B1(n6246), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4746), 
        .ZN(n4741) );
  OAI21_X1 U5898 ( .B1(n6173), .B2(n6254), .A(n4741), .ZN(n4742) );
  AOI21_X1 U5899 ( .B1(n6183), .B2(n6265), .A(n4742), .ZN(n4743) );
  OAI21_X1 U5900 ( .B1(n6256), .B2(n4750), .A(n4743), .ZN(U2982) );
  NAND2_X1 U5901 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5108) );
  OAI211_X1 U5902 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4744), .B(n5108), .ZN(n4749) );
  NOR2_X1 U5903 ( .A1(n6288), .A2(n6171), .ZN(n4745) );
  AOI211_X1 U5904 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n4747), .A(n4746), 
        .B(n4745), .ZN(n4748) );
  OAI211_X1 U5905 ( .C1(n5903), .C2(n4750), .A(n4749), .B(n4748), .ZN(U3014)
         );
  NOR2_X1 U5906 ( .A1(n4654), .A2(n4752), .ZN(n4794) );
  NAND3_X1 U5907 ( .A1(n6598), .A2(n6547), .A3(n4916), .ZN(n4787) );
  NOR2_X1 U5908 ( .A1(n6309), .A2(n4787), .ZN(n4781) );
  AOI21_X1 U5909 ( .B1(n4794), .B2(n6421), .A(n4781), .ZN(n4755) );
  INV_X1 U5910 ( .A(n4755), .ZN(n4754) );
  INV_X1 U5911 ( .A(n4787), .ZN(n4753) );
  AOI22_X1 U5912 ( .A1(n4790), .A2(n4754), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4753), .ZN(n4784) );
  AOI22_X1 U5913 ( .A1(n4790), .A2(n4755), .B1(n4787), .B2(n6476), .ZN(n4756)
         );
  NAND2_X1 U5914 ( .A1(n6426), .A2(n4756), .ZN(n4779) );
  NAND2_X1 U5915 ( .A1(n4779), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4760) );
  NOR2_X1 U5916 ( .A1(n4866), .A2(n5929), .ZN(n4867) );
  INV_X1 U5917 ( .A(n6463), .ZN(n6537) );
  INV_X1 U5918 ( .A(n4920), .ZN(n4757) );
  OAI22_X1 U5919 ( .A1(n4898), .A2(n6469), .B1(n6537), .B2(n4824), .ZN(n4758)
         );
  AOI21_X1 U5920 ( .B1(n6530), .B2(n4781), .A(n4758), .ZN(n4759) );
  OAI211_X1 U5921 ( .C1(n4784), .C2(n6384), .A(n4760), .B(n4759), .ZN(U3035)
         );
  NAND2_X1 U5922 ( .A1(n4779), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4763) );
  INV_X1 U5923 ( .A(n6457), .ZN(n6526) );
  OAI22_X1 U5924 ( .A1(n4898), .A2(n6461), .B1(n6526), .B2(n4824), .ZN(n4761)
         );
  AOI21_X1 U5925 ( .B1(n6522), .B2(n4781), .A(n4761), .ZN(n4762) );
  OAI211_X1 U5926 ( .C1(n4784), .C2(n6378), .A(n4763), .B(n4762), .ZN(U3034)
         );
  NAND2_X1 U5927 ( .A1(n4779), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4766) );
  INV_X1 U5928 ( .A(n6517), .ZN(n6000) );
  INV_X1 U5929 ( .A(n6454), .ZN(n6520) );
  OAI22_X1 U5930 ( .A1(n4898), .A2(n6000), .B1(n6520), .B2(n4824), .ZN(n4764)
         );
  AOI21_X1 U5931 ( .B1(n6516), .B2(n4781), .A(n4764), .ZN(n4765) );
  OAI211_X1 U5932 ( .C1(n4784), .C2(n6375), .A(n4766), .B(n4765), .ZN(U3033)
         );
  NAND2_X1 U5933 ( .A1(n4779), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4769) );
  INV_X1 U5934 ( .A(n6505), .ZN(n5992) );
  INV_X1 U5935 ( .A(n6446), .ZN(n6508) );
  OAI22_X1 U5936 ( .A1(n4898), .A2(n5992), .B1(n6508), .B2(n4824), .ZN(n4767)
         );
  AOI21_X1 U5937 ( .B1(n6782), .B2(n4781), .A(n4767), .ZN(n4768) );
  OAI211_X1 U5938 ( .C1(n4784), .C2(n6369), .A(n4769), .B(n4768), .ZN(U3031)
         );
  NAND2_X1 U5939 ( .A1(n4779), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4772) );
  INV_X1 U5940 ( .A(n6499), .ZN(n5988) );
  INV_X1 U5941 ( .A(n6442), .ZN(n6502) );
  OAI22_X1 U5942 ( .A1(n4898), .A2(n5988), .B1(n6502), .B2(n4824), .ZN(n4770)
         );
  AOI21_X1 U5943 ( .B1(n6498), .B2(n4781), .A(n4770), .ZN(n4771) );
  OAI211_X1 U5944 ( .C1(n4784), .C2(n6366), .A(n4772), .B(n4771), .ZN(U3030)
         );
  NAND2_X1 U5945 ( .A1(n4779), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4775) );
  INV_X1 U5946 ( .A(n6493), .ZN(n5984) );
  INV_X1 U5947 ( .A(n6438), .ZN(n6496) );
  OAI22_X1 U5948 ( .A1(n4898), .A2(n5984), .B1(n6496), .B2(n4824), .ZN(n4773)
         );
  AOI21_X1 U5949 ( .B1(n6492), .B2(n4781), .A(n4773), .ZN(n4774) );
  OAI211_X1 U5950 ( .C1(n4784), .C2(n6363), .A(n4775), .B(n4774), .ZN(U3029)
         );
  NAND2_X1 U5951 ( .A1(n4779), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4778) );
  INV_X1 U5952 ( .A(n6487), .ZN(n5980) );
  INV_X1 U5953 ( .A(n6435), .ZN(n6490) );
  OAI22_X1 U5954 ( .A1(n4898), .A2(n5980), .B1(n6490), .B2(n4824), .ZN(n4776)
         );
  AOI21_X1 U5955 ( .B1(n6475), .B2(n4781), .A(n4776), .ZN(n4777) );
  OAI211_X1 U5956 ( .C1(n4784), .C2(n6360), .A(n4778), .B(n4777), .ZN(U3028)
         );
  NAND2_X1 U5957 ( .A1(n4779), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4783) );
  INV_X1 U5958 ( .A(n6511), .ZN(n5996) );
  INV_X1 U5959 ( .A(n6450), .ZN(n6514) );
  OAI22_X1 U5960 ( .A1(n4898), .A2(n5996), .B1(n6514), .B2(n4824), .ZN(n4780)
         );
  AOI21_X1 U5961 ( .B1(n6510), .B2(n4781), .A(n4780), .ZN(n4782) );
  OAI211_X1 U5962 ( .C1(n4784), .C2(n6372), .A(n4783), .B(n4782), .ZN(U3032)
         );
  INV_X1 U5963 ( .A(n5032), .ZN(n4786) );
  NAND2_X1 U5964 ( .A1(n6419), .A2(n6059), .ZN(n6593) );
  AOI21_X1 U5965 ( .B1(n4786), .B2(n6593), .A(n4794), .ZN(n4789) );
  NOR2_X1 U5966 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4787), .ZN(n4827)
         );
  NOR2_X1 U5967 ( .A1(n4791), .A2(n5978), .ZN(n4870) );
  INV_X1 U5968 ( .A(n4870), .ZN(n6471) );
  OR2_X1 U5969 ( .A1(n6388), .A2(n6389), .ZN(n4922) );
  AOI21_X1 U5970 ( .B1(n4922), .B2(STATE2_REG_2__SCAN_IN), .A(n6394), .ZN(
        n4917) );
  OAI211_X1 U5971 ( .C1(n4827), .C2(n6588), .A(n6471), .B(n4917), .ZN(n4788)
         );
  INV_X1 U5972 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4798) );
  INV_X1 U5973 ( .A(n4791), .ZN(n4792) );
  NOR2_X1 U5974 ( .A1(n4792), .A2(n5978), .ZN(n5934) );
  INV_X1 U5975 ( .A(n4922), .ZN(n4793) );
  AOI22_X1 U5976 ( .A1(n4794), .A2(n6419), .B1(n5934), .B2(n4793), .ZN(n4823)
         );
  OAI22_X1 U5977 ( .A1(n5032), .A2(n6508), .B1(n4823), .B2(n6369), .ZN(n4796)
         );
  NOR2_X1 U5978 ( .A1(n4824), .A2(n5992), .ZN(n4795) );
  AOI211_X1 U5979 ( .C1(n6782), .C2(n4827), .A(n4796), .B(n4795), .ZN(n4797)
         );
  OAI21_X1 U5980 ( .B1(n4830), .B2(n4798), .A(n4797), .ZN(U3023) );
  INV_X1 U5981 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4802) );
  OAI22_X1 U5982 ( .A1(n5032), .A2(n6502), .B1(n4823), .B2(n6366), .ZN(n4800)
         );
  NOR2_X1 U5983 ( .A1(n4824), .A2(n5988), .ZN(n4799) );
  AOI211_X1 U5984 ( .C1(n6498), .C2(n4827), .A(n4800), .B(n4799), .ZN(n4801)
         );
  OAI21_X1 U5985 ( .B1(n4830), .B2(n4802), .A(n4801), .ZN(U3022) );
  OAI22_X1 U5986 ( .A1(n5032), .A2(n6496), .B1(n4823), .B2(n6363), .ZN(n4804)
         );
  NOR2_X1 U5987 ( .A1(n4824), .A2(n5984), .ZN(n4803) );
  AOI211_X1 U5988 ( .C1(n6492), .C2(n4827), .A(n4804), .B(n4803), .ZN(n4805)
         );
  OAI21_X1 U5989 ( .B1(n4830), .B2(n4806), .A(n4805), .ZN(U3021) );
  OAI22_X1 U5990 ( .A1(n5032), .A2(n6490), .B1(n4823), .B2(n6360), .ZN(n4808)
         );
  NOR2_X1 U5991 ( .A1(n4824), .A2(n5980), .ZN(n4807) );
  AOI211_X1 U5992 ( .C1(n6475), .C2(n4827), .A(n4808), .B(n4807), .ZN(n4809)
         );
  OAI21_X1 U5993 ( .B1(n4830), .B2(n4810), .A(n4809), .ZN(U3020) );
  INV_X1 U5994 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4814) );
  OAI22_X1 U5995 ( .A1(n5032), .A2(n6520), .B1(n4823), .B2(n6375), .ZN(n4812)
         );
  NOR2_X1 U5996 ( .A1(n4824), .A2(n6000), .ZN(n4811) );
  AOI211_X1 U5997 ( .C1(n6516), .C2(n4827), .A(n4812), .B(n4811), .ZN(n4813)
         );
  OAI21_X1 U5998 ( .B1(n4830), .B2(n4814), .A(n4813), .ZN(U3025) );
  INV_X1 U5999 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4818) );
  OAI22_X1 U6000 ( .A1(n5032), .A2(n6514), .B1(n4823), .B2(n6372), .ZN(n4816)
         );
  NOR2_X1 U6001 ( .A1(n4824), .A2(n5996), .ZN(n4815) );
  AOI211_X1 U6002 ( .C1(n6510), .C2(n4827), .A(n4816), .B(n4815), .ZN(n4817)
         );
  OAI21_X1 U6003 ( .B1(n4830), .B2(n4818), .A(n4817), .ZN(U3024) );
  INV_X1 U6004 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4822) );
  OAI22_X1 U6005 ( .A1(n5032), .A2(n6537), .B1(n4823), .B2(n6384), .ZN(n4820)
         );
  NOR2_X1 U6006 ( .A1(n4824), .A2(n6469), .ZN(n4819) );
  AOI211_X1 U6007 ( .C1(n6530), .C2(n4827), .A(n4820), .B(n4819), .ZN(n4821)
         );
  OAI21_X1 U6008 ( .B1(n4830), .B2(n4822), .A(n4821), .ZN(U3027) );
  INV_X1 U6009 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4829) );
  OAI22_X1 U6010 ( .A1(n5032), .A2(n6526), .B1(n4823), .B2(n6378), .ZN(n4826)
         );
  NOR2_X1 U6011 ( .A1(n4824), .A2(n6461), .ZN(n4825) );
  AOI211_X1 U6012 ( .C1(n6522), .C2(n4827), .A(n4826), .B(n4825), .ZN(n4828)
         );
  OAI21_X1 U6013 ( .B1(n4830), .B2(n4829), .A(n4828), .ZN(U3026) );
  NAND2_X1 U6014 ( .A1(n4647), .A2(n4832), .ZN(n4833) );
  AND2_X1 U6015 ( .A1(n4831), .A2(n4833), .ZN(n6153) );
  INV_X1 U6016 ( .A(n6153), .ZN(n4838) );
  XNOR2_X1 U6017 ( .A(n5107), .B(n4834), .ZN(n6148) );
  INV_X1 U6018 ( .A(n6148), .ZN(n4836) );
  INV_X1 U6019 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4835) );
  OAI222_X1 U6020 ( .A1(n4838), .A2(n2970), .B1(n5428), .B2(n4836), .C1(n6195), 
        .C2(n4835), .ZN(U2853) );
  OAI222_X1 U6021 ( .A1(n4838), .A2(n6776), .B1(n5491), .B2(n4837), .C1(n5489), 
        .C2(n3545), .ZN(U2885) );
  NAND3_X1 U6022 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n4916), .ZN(n6470) );
  NOR2_X1 U6023 ( .A1(n6309), .A2(n6470), .ZN(n4839) );
  INV_X1 U6024 ( .A(n4839), .ZN(n4865) );
  NAND2_X1 U6025 ( .A1(n6419), .A2(n5043), .ZN(n4843) );
  INV_X1 U6026 ( .A(n4437), .ZN(n5386) );
  NAND2_X1 U6027 ( .A1(n5386), .A2(n5917), .ZN(n6478) );
  INV_X1 U6028 ( .A(n6478), .ZN(n4921) );
  AOI21_X1 U6029 ( .B1(n4921), .B2(n4996), .A(n4839), .ZN(n4844) );
  INV_X1 U6030 ( .A(n4844), .ZN(n4842) );
  AOI21_X1 U6031 ( .B1(n6476), .B2(n6470), .A(n4840), .ZN(n4841) );
  OAI22_X1 U6032 ( .A1(n4844), .A2(n4843), .B1(n5978), .B2(n6470), .ZN(n4861)
         );
  AOI22_X1 U6033 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4862), .B1(n6515), 
        .B2(n4861), .ZN(n4848) );
  INV_X1 U6034 ( .A(n4845), .ZN(n4846) );
  AOI22_X1 U6035 ( .A1(n6517), .A2(n4990), .B1(n6531), .B2(n6454), .ZN(n4847)
         );
  OAI211_X1 U6036 ( .C1(n5022), .C2(n4865), .A(n4848), .B(n4847), .ZN(U3129)
         );
  AOI22_X1 U6037 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4862), .B1(n6503), 
        .B2(n4861), .ZN(n4850) );
  AOI22_X1 U6038 ( .A1(n6505), .A2(n4990), .B1(n6531), .B2(n6446), .ZN(n4849)
         );
  OAI211_X1 U6039 ( .C1(n6504), .C2(n4865), .A(n4850), .B(n4849), .ZN(U3127)
         );
  AOI22_X1 U6040 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4862), .B1(n6497), 
        .B2(n4861), .ZN(n4852) );
  AOI22_X1 U6041 ( .A1(n6499), .A2(n4990), .B1(n6531), .B2(n6442), .ZN(n4851)
         );
  OAI211_X1 U6042 ( .C1(n5026), .C2(n4865), .A(n4852), .B(n4851), .ZN(U3126)
         );
  AOI22_X1 U6043 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4862), .B1(n6528), 
        .B2(n4861), .ZN(n4854) );
  AOI22_X1 U6044 ( .A1(n6532), .A2(n4990), .B1(n6531), .B2(n6463), .ZN(n4853)
         );
  OAI211_X1 U6045 ( .C1(n5018), .C2(n4865), .A(n4854), .B(n4853), .ZN(U3131)
         );
  AOI22_X1 U6046 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4862), .B1(n6521), 
        .B2(n4861), .ZN(n4856) );
  AOI22_X1 U6047 ( .A1(n6523), .A2(n4990), .B1(n6531), .B2(n6457), .ZN(n4855)
         );
  OAI211_X1 U6048 ( .C1(n5014), .C2(n4865), .A(n4856), .B(n4855), .ZN(U3130)
         );
  AOI22_X1 U6049 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4862), .B1(n6509), 
        .B2(n4861), .ZN(n4858) );
  AOI22_X1 U6050 ( .A1(n6511), .A2(n4990), .B1(n6531), .B2(n6450), .ZN(n4857)
         );
  OAI211_X1 U6051 ( .C1(n5038), .C2(n4865), .A(n4858), .B(n4857), .ZN(U3128)
         );
  AOI22_X1 U6052 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4862), .B1(n6491), 
        .B2(n4861), .ZN(n4860) );
  AOI22_X1 U6053 ( .A1(n6493), .A2(n4990), .B1(n6531), .B2(n6438), .ZN(n4859)
         );
  OAI211_X1 U6054 ( .C1(n5010), .C2(n4865), .A(n4860), .B(n4859), .ZN(U3125)
         );
  AOI22_X1 U6055 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4862), .B1(n6474), 
        .B2(n4861), .ZN(n4864) );
  AOI22_X1 U6056 ( .A1(n6487), .A2(n4990), .B1(n6531), .B2(n6435), .ZN(n4863)
         );
  OAI211_X1 U6057 ( .C1(n5006), .C2(n4865), .A(n4864), .B(n4863), .ZN(U3124)
         );
  NAND2_X1 U6058 ( .A1(n5972), .A2(n6598), .ZN(n5052) );
  NOR2_X1 U6059 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5052), .ZN(n4872)
         );
  INV_X1 U6060 ( .A(n4872), .ZN(n4902) );
  INV_X1 U6061 ( .A(n5041), .ZN(n5915) );
  OAI21_X1 U6062 ( .B1(n5057), .B2(n4867), .A(n6593), .ZN(n4868) );
  AND2_X1 U6063 ( .A1(n4341), .A2(n4437), .ZN(n5970) );
  NAND2_X1 U6064 ( .A1(n6592), .A2(n5970), .ZN(n5047) );
  AOI21_X1 U6065 ( .B1(n4868), .B2(n5047), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4871) );
  NOR2_X1 U6066 ( .A1(n4870), .A2(n5933), .ZN(n5977) );
  NAND2_X1 U6067 ( .A1(n4896), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4877) );
  INV_X1 U6068 ( .A(n5047), .ZN(n4874) );
  INV_X1 U6069 ( .A(n5934), .ZN(n6484) );
  NOR2_X1 U6070 ( .A1(n6484), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4873)
         );
  AOI22_X1 U6071 ( .A1(n4874), .A2(n6419), .B1(n6389), .B2(n4873), .ZN(n4897)
         );
  OAI22_X1 U6072 ( .A1(n4898), .A2(n6514), .B1(n4897), .B2(n6372), .ZN(n4875)
         );
  AOI21_X1 U6073 ( .B1(n6511), .B2(n5057), .A(n4875), .ZN(n4876) );
  OAI211_X1 U6074 ( .C1(n4902), .C2(n5038), .A(n4877), .B(n4876), .ZN(U3040)
         );
  NAND2_X1 U6075 ( .A1(n4896), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4880) );
  OAI22_X1 U6076 ( .A1(n4898), .A2(n6520), .B1(n4897), .B2(n6375), .ZN(n4878)
         );
  AOI21_X1 U6077 ( .B1(n6517), .B2(n5057), .A(n4878), .ZN(n4879) );
  OAI211_X1 U6078 ( .C1(n4902), .C2(n5022), .A(n4880), .B(n4879), .ZN(U3041)
         );
  NAND2_X1 U6079 ( .A1(n4896), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4883) );
  OAI22_X1 U6080 ( .A1(n4898), .A2(n6526), .B1(n4897), .B2(n6378), .ZN(n4881)
         );
  AOI21_X1 U6081 ( .B1(n6523), .B2(n5057), .A(n4881), .ZN(n4882) );
  OAI211_X1 U6082 ( .C1(n4902), .C2(n5014), .A(n4883), .B(n4882), .ZN(U3042)
         );
  NAND2_X1 U6083 ( .A1(n4896), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4886) );
  OAI22_X1 U6084 ( .A1(n4898), .A2(n6537), .B1(n4897), .B2(n6384), .ZN(n4884)
         );
  AOI21_X1 U6085 ( .B1(n6532), .B2(n5057), .A(n4884), .ZN(n4885) );
  OAI211_X1 U6086 ( .C1(n4902), .C2(n5018), .A(n4886), .B(n4885), .ZN(U3043)
         );
  NAND2_X1 U6087 ( .A1(n4896), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4889) );
  OAI22_X1 U6088 ( .A1(n4898), .A2(n6496), .B1(n4897), .B2(n6363), .ZN(n4887)
         );
  AOI21_X1 U6089 ( .B1(n6493), .B2(n5057), .A(n4887), .ZN(n4888) );
  OAI211_X1 U6090 ( .C1(n4902), .C2(n5010), .A(n4889), .B(n4888), .ZN(U3037)
         );
  NAND2_X1 U6091 ( .A1(n4896), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4892) );
  OAI22_X1 U6092 ( .A1(n4898), .A2(n6502), .B1(n4897), .B2(n6366), .ZN(n4890)
         );
  AOI21_X1 U6093 ( .B1(n6499), .B2(n5057), .A(n4890), .ZN(n4891) );
  OAI211_X1 U6094 ( .C1(n4902), .C2(n5026), .A(n4892), .B(n4891), .ZN(U3038)
         );
  NAND2_X1 U6095 ( .A1(n4896), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4895) );
  OAI22_X1 U6096 ( .A1(n4898), .A2(n6490), .B1(n4897), .B2(n6360), .ZN(n4893)
         );
  AOI21_X1 U6097 ( .B1(n6487), .B2(n5057), .A(n4893), .ZN(n4894) );
  OAI211_X1 U6098 ( .C1(n5006), .C2(n4902), .A(n4895), .B(n4894), .ZN(U3036)
         );
  NAND2_X1 U6099 ( .A1(n4896), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4901) );
  OAI22_X1 U6100 ( .A1(n4898), .A2(n6508), .B1(n4897), .B2(n6369), .ZN(n4899)
         );
  AOI21_X1 U6101 ( .B1(n6505), .B2(n5057), .A(n4899), .ZN(n4900) );
  OAI211_X1 U6102 ( .C1(n4902), .C2(n6504), .A(n4901), .B(n4900), .ZN(U3039)
         );
  NAND2_X1 U6103 ( .A1(n4831), .A2(n4905), .ZN(n4906) );
  NAND2_X1 U6104 ( .A1(n4904), .A2(n4906), .ZN(n6259) );
  OR2_X1 U6105 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  NAND2_X1 U6106 ( .A1(n5126), .A2(n4909), .ZN(n6128) );
  INV_X1 U6107 ( .A(n6128), .ZN(n4910) );
  AOI22_X1 U6108 ( .A1(n4910), .A2(n6192), .B1(n5452), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4911) );
  OAI21_X1 U6109 ( .B1(n6259), .B2(n2970), .A(n4911), .ZN(U2852) );
  OAI21_X1 U6110 ( .B1(n6352), .B2(n4913), .A(n6419), .ZN(n6315) );
  INV_X1 U6111 ( .A(n6593), .ZN(n6480) );
  NOR2_X1 U6112 ( .A1(n5080), .A2(n6480), .ZN(n4915) );
  AOI211_X1 U6113 ( .C1(n4921), .C2(n6479), .A(n6315), .B(n4915), .ZN(n4919)
         );
  NAND3_X1 U6114 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6598), .A3(n4916), .ZN(n6312) );
  NOR2_X1 U6115 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6312), .ZN(n4954)
         );
  OAI211_X1 U6116 ( .C1(n4954), .C2(n6588), .A(n6484), .B(n4917), .ZN(n4918)
         );
  INV_X1 U6117 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4926) );
  NOR2_X2 U6118 ( .A1(n6352), .A2(n4920), .ZN(n6333) );
  NAND2_X1 U6119 ( .A1(n4921), .A2(n6419), .ZN(n6473) );
  OAI22_X1 U6120 ( .A1(n6473), .A2(n4654), .B1(n6471), .B2(n4922), .ZN(n4951)
         );
  AOI22_X1 U6121 ( .A1(n6333), .A2(n6505), .B1(n6503), .B2(n4951), .ZN(n4923)
         );
  OAI21_X1 U6122 ( .B1(n5080), .B2(n6508), .A(n4923), .ZN(n4924) );
  AOI21_X1 U6123 ( .B1(n6782), .B2(n4954), .A(n4924), .ZN(n4925) );
  OAI21_X1 U6124 ( .B1(n4957), .B2(n4926), .A(n4925), .ZN(U3055) );
  INV_X1 U6125 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4930) );
  AOI22_X1 U6126 ( .A1(n6333), .A2(n6523), .B1(n6521), .B2(n4951), .ZN(n4927)
         );
  OAI21_X1 U6127 ( .B1(n5080), .B2(n6526), .A(n4927), .ZN(n4928) );
  AOI21_X1 U6128 ( .B1(n6522), .B2(n4954), .A(n4928), .ZN(n4929) );
  OAI21_X1 U6129 ( .B1(n4957), .B2(n4930), .A(n4929), .ZN(U3058) );
  INV_X1 U6130 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4934) );
  AOI22_X1 U6131 ( .A1(n6333), .A2(n6517), .B1(n6515), .B2(n4951), .ZN(n4931)
         );
  OAI21_X1 U6132 ( .B1(n5080), .B2(n6520), .A(n4931), .ZN(n4932) );
  AOI21_X1 U6133 ( .B1(n6516), .B2(n4954), .A(n4932), .ZN(n4933) );
  OAI21_X1 U6134 ( .B1(n4957), .B2(n4934), .A(n4933), .ZN(U3057) );
  INV_X1 U6135 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4938) );
  AOI22_X1 U6136 ( .A1(n6333), .A2(n6499), .B1(n6497), .B2(n4951), .ZN(n4935)
         );
  OAI21_X1 U6137 ( .B1(n5080), .B2(n6502), .A(n4935), .ZN(n4936) );
  AOI21_X1 U6138 ( .B1(n6498), .B2(n4954), .A(n4936), .ZN(n4937) );
  OAI21_X1 U6139 ( .B1(n4957), .B2(n4938), .A(n4937), .ZN(U3054) );
  INV_X1 U6140 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4942) );
  AOI22_X1 U6141 ( .A1(n6333), .A2(n6493), .B1(n6491), .B2(n4951), .ZN(n4939)
         );
  OAI21_X1 U6142 ( .B1(n5080), .B2(n6496), .A(n4939), .ZN(n4940) );
  AOI21_X1 U6143 ( .B1(n6492), .B2(n4954), .A(n4940), .ZN(n4941) );
  OAI21_X1 U6144 ( .B1(n4957), .B2(n4942), .A(n4941), .ZN(U3053) );
  INV_X1 U6145 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4946) );
  AOI22_X1 U6146 ( .A1(n6333), .A2(n6487), .B1(n6474), .B2(n4951), .ZN(n4943)
         );
  OAI21_X1 U6147 ( .B1(n5080), .B2(n6490), .A(n4943), .ZN(n4944) );
  AOI21_X1 U6148 ( .B1(n6475), .B2(n4954), .A(n4944), .ZN(n4945) );
  OAI21_X1 U6149 ( .B1(n4957), .B2(n4946), .A(n4945), .ZN(U3052) );
  INV_X1 U6150 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4950) );
  AOI22_X1 U6151 ( .A1(n6333), .A2(n6511), .B1(n6509), .B2(n4951), .ZN(n4947)
         );
  OAI21_X1 U6152 ( .B1(n5080), .B2(n6514), .A(n4947), .ZN(n4948) );
  AOI21_X1 U6153 ( .B1(n6510), .B2(n4954), .A(n4948), .ZN(n4949) );
  OAI21_X1 U6154 ( .B1(n4957), .B2(n4950), .A(n4949), .ZN(U3056) );
  INV_X1 U6155 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4956) );
  AOI22_X1 U6156 ( .A1(n6333), .A2(n6532), .B1(n6528), .B2(n4951), .ZN(n4952)
         );
  OAI21_X1 U6157 ( .B1(n5080), .B2(n6537), .A(n4952), .ZN(n4953) );
  AOI21_X1 U6158 ( .B1(n6530), .B2(n4954), .A(n4953), .ZN(n4955) );
  OAI21_X1 U6159 ( .B1(n4957), .B2(n4956), .A(n4955), .ZN(U3059) );
  NOR2_X1 U6160 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4958), .ZN(n4963)
         );
  INV_X1 U6161 ( .A(n4963), .ZN(n4993) );
  NOR3_X1 U6162 ( .A1(n5933), .A2(n6598), .A3(n5934), .ZN(n4962) );
  NAND2_X1 U6163 ( .A1(n5386), .A2(n4341), .ZN(n6347) );
  INV_X1 U6164 ( .A(n5967), .ZN(n4959) );
  OAI21_X1 U6165 ( .B1(n4990), .B2(n4964), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4960) );
  NAND3_X1 U6166 ( .A1(n6347), .A2(n6419), .A3(n4960), .ZN(n4961) );
  NAND2_X1 U6167 ( .A1(n4987), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4968)
         );
  NOR2_X1 U6168 ( .A1(n6347), .A2(n6476), .ZN(n5936) );
  NOR2_X1 U6169 ( .A1(n6471), .A2(n6598), .ZN(n4965) );
  AOI22_X1 U6170 ( .A1(n5936), .A2(n4654), .B1(n6389), .B2(n4965), .ZN(n4988)
         );
  OAI22_X1 U6171 ( .A1(n5033), .A2(n5988), .B1(n4988), .B2(n6366), .ZN(n4966)
         );
  AOI21_X1 U6172 ( .B1(n6442), .B2(n4990), .A(n4966), .ZN(n4967) );
  OAI211_X1 U6173 ( .C1(n4993), .C2(n5026), .A(n4968), .B(n4967), .ZN(U3134)
         );
  NAND2_X1 U6174 ( .A1(n4987), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4971)
         );
  OAI22_X1 U6175 ( .A1(n5033), .A2(n6000), .B1(n4988), .B2(n6375), .ZN(n4969)
         );
  AOI21_X1 U6176 ( .B1(n6454), .B2(n4990), .A(n4969), .ZN(n4970) );
  OAI211_X1 U6177 ( .C1(n4993), .C2(n5022), .A(n4971), .B(n4970), .ZN(U3137)
         );
  NAND2_X1 U6178 ( .A1(n4987), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4974)
         );
  OAI22_X1 U6179 ( .A1(n5033), .A2(n5992), .B1(n4988), .B2(n6369), .ZN(n4972)
         );
  AOI21_X1 U6180 ( .B1(n6446), .B2(n4990), .A(n4972), .ZN(n4973) );
  OAI211_X1 U6181 ( .C1(n4993), .C2(n6504), .A(n4974), .B(n4973), .ZN(U3135)
         );
  NAND2_X1 U6182 ( .A1(n4987), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4977)
         );
  OAI22_X1 U6183 ( .A1(n5033), .A2(n6469), .B1(n4988), .B2(n6384), .ZN(n4975)
         );
  AOI21_X1 U6184 ( .B1(n6463), .B2(n4990), .A(n4975), .ZN(n4976) );
  OAI211_X1 U6185 ( .C1(n4993), .C2(n5018), .A(n4977), .B(n4976), .ZN(U3139)
         );
  NAND2_X1 U6186 ( .A1(n4987), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4980)
         );
  OAI22_X1 U6187 ( .A1(n5033), .A2(n5996), .B1(n4988), .B2(n6372), .ZN(n4978)
         );
  AOI21_X1 U6188 ( .B1(n6450), .B2(n4990), .A(n4978), .ZN(n4979) );
  OAI211_X1 U6189 ( .C1(n4993), .C2(n5038), .A(n4980), .B(n4979), .ZN(U3136)
         );
  NAND2_X1 U6190 ( .A1(n4987), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4983)
         );
  OAI22_X1 U6191 ( .A1(n5033), .A2(n5980), .B1(n4988), .B2(n6360), .ZN(n4981)
         );
  AOI21_X1 U6192 ( .B1(n4990), .B2(n6435), .A(n4981), .ZN(n4982) );
  OAI211_X1 U6193 ( .C1(n5006), .C2(n4993), .A(n4983), .B(n4982), .ZN(U3132)
         );
  NAND2_X1 U6194 ( .A1(n4987), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4986)
         );
  OAI22_X1 U6195 ( .A1(n5033), .A2(n5984), .B1(n4988), .B2(n6363), .ZN(n4984)
         );
  AOI21_X1 U6196 ( .B1(n6438), .B2(n4990), .A(n4984), .ZN(n4985) );
  OAI211_X1 U6197 ( .C1(n4993), .C2(n5010), .A(n4986), .B(n4985), .ZN(U3133)
         );
  NAND2_X1 U6198 ( .A1(n4987), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4992)
         );
  OAI22_X1 U6199 ( .A1(n5033), .A2(n6461), .B1(n4988), .B2(n6378), .ZN(n4989)
         );
  AOI21_X1 U6200 ( .B1(n6457), .B2(n4990), .A(n4989), .ZN(n4991) );
  OAI211_X1 U6201 ( .C1(n4993), .C2(n5014), .A(n4992), .B(n4991), .ZN(U3138)
         );
  AOI21_X1 U6202 ( .B1(n4994), .B2(n5915), .A(n6258), .ZN(n4998) );
  INV_X1 U6203 ( .A(n6347), .ZN(n4997) );
  INV_X1 U6204 ( .A(n5039), .ZN(n4995) );
  AOI21_X1 U6205 ( .B1(n4997), .B2(n4996), .A(n4995), .ZN(n5000) );
  OAI21_X1 U6206 ( .B1(n4998), .B2(n6480), .A(n5000), .ZN(n4999) );
  OAI211_X1 U6207 ( .C1(n6419), .C2(n5001), .A(n4999), .B(n6426), .ZN(n5036)
         );
  INV_X1 U6208 ( .A(n5000), .ZN(n5002) );
  AOI22_X1 U6209 ( .A1(n5002), .A2(n6419), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5001), .ZN(n5031) );
  OAI22_X1 U6210 ( .A1(n5980), .A2(n5032), .B1(n5031), .B2(n6360), .ZN(n5004)
         );
  NOR2_X1 U6211 ( .A1(n5033), .A2(n6490), .ZN(n5003) );
  AOI211_X1 U6212 ( .C1(INSTQUEUE_REG_15__0__SCAN_IN), .C2(n5036), .A(n5004), 
        .B(n5003), .ZN(n5005) );
  OAI21_X1 U6213 ( .B1(n5039), .B2(n5006), .A(n5005), .ZN(U3140) );
  OAI22_X1 U6214 ( .A1(n5984), .A2(n5032), .B1(n5031), .B2(n6363), .ZN(n5008)
         );
  NOR2_X1 U6215 ( .A1(n5033), .A2(n6496), .ZN(n5007) );
  AOI211_X1 U6216 ( .C1(INSTQUEUE_REG_15__1__SCAN_IN), .C2(n5036), .A(n5008), 
        .B(n5007), .ZN(n5009) );
  OAI21_X1 U6217 ( .B1(n5039), .B2(n5010), .A(n5009), .ZN(U3141) );
  OAI22_X1 U6218 ( .A1(n6461), .A2(n5032), .B1(n5031), .B2(n6378), .ZN(n5012)
         );
  NOR2_X1 U6219 ( .A1(n5033), .A2(n6526), .ZN(n5011) );
  AOI211_X1 U6220 ( .C1(INSTQUEUE_REG_15__6__SCAN_IN), .C2(n5036), .A(n5012), 
        .B(n5011), .ZN(n5013) );
  OAI21_X1 U6221 ( .B1(n5039), .B2(n5014), .A(n5013), .ZN(U3146) );
  OAI22_X1 U6222 ( .A1(n6469), .A2(n5032), .B1(n5031), .B2(n6384), .ZN(n5016)
         );
  NOR2_X1 U6223 ( .A1(n5033), .A2(n6537), .ZN(n5015) );
  AOI211_X1 U6224 ( .C1(INSTQUEUE_REG_15__7__SCAN_IN), .C2(n5036), .A(n5016), 
        .B(n5015), .ZN(n5017) );
  OAI21_X1 U6225 ( .B1(n5039), .B2(n5018), .A(n5017), .ZN(U3147) );
  OAI22_X1 U6226 ( .A1(n6000), .A2(n5032), .B1(n5031), .B2(n6375), .ZN(n5020)
         );
  NOR2_X1 U6227 ( .A1(n5033), .A2(n6520), .ZN(n5019) );
  AOI211_X1 U6228 ( .C1(INSTQUEUE_REG_15__5__SCAN_IN), .C2(n5036), .A(n5020), 
        .B(n5019), .ZN(n5021) );
  OAI21_X1 U6229 ( .B1(n5039), .B2(n5022), .A(n5021), .ZN(U3145) );
  OAI22_X1 U6230 ( .A1(n5988), .A2(n5032), .B1(n5031), .B2(n6366), .ZN(n5024)
         );
  NOR2_X1 U6231 ( .A1(n5033), .A2(n6502), .ZN(n5023) );
  AOI211_X1 U6232 ( .C1(INSTQUEUE_REG_15__2__SCAN_IN), .C2(n5036), .A(n5024), 
        .B(n5023), .ZN(n5025) );
  OAI21_X1 U6233 ( .B1(n5039), .B2(n5026), .A(n5025), .ZN(U3142) );
  OAI22_X1 U6234 ( .A1(n5992), .A2(n5032), .B1(n5031), .B2(n6369), .ZN(n5028)
         );
  NOR2_X1 U6235 ( .A1(n5033), .A2(n6508), .ZN(n5027) );
  AOI211_X1 U6236 ( .C1(INSTQUEUE_REG_15__3__SCAN_IN), .C2(n5036), .A(n5028), 
        .B(n5027), .ZN(n5029) );
  OAI21_X1 U6237 ( .B1(n5039), .B2(n6504), .A(n5029), .ZN(U3143) );
  OAI22_X1 U6238 ( .A1(n5996), .A2(n5032), .B1(n5031), .B2(n6372), .ZN(n5035)
         );
  NOR2_X1 U6239 ( .A1(n5033), .A2(n6514), .ZN(n5034) );
  AOI211_X1 U6240 ( .C1(INSTQUEUE_REG_15__4__SCAN_IN), .C2(n5036), .A(n5035), 
        .B(n5034), .ZN(n5037) );
  OAI21_X1 U6241 ( .B1(n5039), .B2(n5038), .A(n5037), .ZN(U3144) );
  OAI222_X1 U6242 ( .A1(n6259), .A2(n6776), .B1(n5491), .B2(n5040), .C1(n5489), 
        .C2(n3571), .ZN(U2884) );
  OR2_X1 U6243 ( .A1(n5041), .A2(n6059), .ZN(n6420) );
  OR2_X1 U6244 ( .A1(n6352), .A2(n6420), .ZN(n6345) );
  AND2_X1 U6245 ( .A1(n6428), .A2(n6345), .ZN(n5042) );
  AOI21_X1 U6246 ( .B1(n5043), .B2(n5042), .A(n6476), .ZN(n6596) );
  INV_X1 U6247 ( .A(n6420), .ZN(n5919) );
  AOI21_X1 U6248 ( .B1(n5044), .B2(n5919), .A(n6476), .ZN(n5045) );
  NOR2_X1 U6249 ( .A1(n6596), .A2(n5045), .ZN(n5055) );
  INV_X1 U6250 ( .A(n5055), .ZN(n5051) );
  OR2_X1 U6251 ( .A1(n5047), .A2(n5046), .ZN(n5049) );
  INV_X1 U6252 ( .A(n6423), .ZN(n5048) );
  NAND2_X1 U6253 ( .A1(n5048), .A2(n6598), .ZN(n5056) );
  NAND2_X1 U6254 ( .A1(n5049), .A2(n5056), .ZN(n5054) );
  INV_X1 U6255 ( .A(n5052), .ZN(n5050) );
  NAND2_X1 U6256 ( .A1(n6476), .A2(n5052), .ZN(n5053) );
  NAND2_X1 U6257 ( .A1(n5079), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5060) );
  INV_X1 U6258 ( .A(n5056), .ZN(n5083) );
  OAI22_X1 U6259 ( .A1(n5081), .A2(n6537), .B1(n6469), .B2(n5080), .ZN(n5058)
         );
  AOI21_X1 U6260 ( .B1(n6530), .B2(n5083), .A(n5058), .ZN(n5059) );
  OAI211_X1 U6261 ( .C1(n5086), .C2(n6384), .A(n5060), .B(n5059), .ZN(U3051)
         );
  NAND2_X1 U6262 ( .A1(n5079), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5063) );
  OAI22_X1 U6263 ( .A1(n5081), .A2(n6514), .B1(n5996), .B2(n5080), .ZN(n5061)
         );
  AOI21_X1 U6264 ( .B1(n6510), .B2(n5083), .A(n5061), .ZN(n5062) );
  OAI211_X1 U6265 ( .C1(n5086), .C2(n6372), .A(n5063), .B(n5062), .ZN(U3048)
         );
  NAND2_X1 U6266 ( .A1(n5079), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5066) );
  OAI22_X1 U6267 ( .A1(n5081), .A2(n6490), .B1(n5980), .B2(n5080), .ZN(n5064)
         );
  AOI21_X1 U6268 ( .B1(n6475), .B2(n5083), .A(n5064), .ZN(n5065) );
  OAI211_X1 U6269 ( .C1(n5086), .C2(n6360), .A(n5066), .B(n5065), .ZN(U3044)
         );
  NAND2_X1 U6270 ( .A1(n5079), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5069) );
  OAI22_X1 U6271 ( .A1(n5081), .A2(n6520), .B1(n6000), .B2(n5080), .ZN(n5067)
         );
  AOI21_X1 U6272 ( .B1(n6516), .B2(n5083), .A(n5067), .ZN(n5068) );
  OAI211_X1 U6273 ( .C1(n5086), .C2(n6375), .A(n5069), .B(n5068), .ZN(U3049)
         );
  NAND2_X1 U6274 ( .A1(n5079), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5072) );
  OAI22_X1 U6275 ( .A1(n5081), .A2(n6508), .B1(n5992), .B2(n5080), .ZN(n5070)
         );
  AOI21_X1 U6276 ( .B1(n6782), .B2(n5083), .A(n5070), .ZN(n5071) );
  OAI211_X1 U6277 ( .C1(n5086), .C2(n6369), .A(n5072), .B(n5071), .ZN(U3047)
         );
  NAND2_X1 U6278 ( .A1(n5079), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5075) );
  OAI22_X1 U6279 ( .A1(n5081), .A2(n6496), .B1(n5984), .B2(n5080), .ZN(n5073)
         );
  AOI21_X1 U6280 ( .B1(n6492), .B2(n5083), .A(n5073), .ZN(n5074) );
  OAI211_X1 U6281 ( .C1(n5086), .C2(n6363), .A(n5075), .B(n5074), .ZN(U3045)
         );
  NAND2_X1 U6282 ( .A1(n5079), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5078) );
  OAI22_X1 U6283 ( .A1(n5081), .A2(n6526), .B1(n6461), .B2(n5080), .ZN(n5076)
         );
  AOI21_X1 U6284 ( .B1(n6522), .B2(n5083), .A(n5076), .ZN(n5077) );
  OAI211_X1 U6285 ( .C1(n5086), .C2(n6378), .A(n5078), .B(n5077), .ZN(U3050)
         );
  NAND2_X1 U6286 ( .A1(n5079), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5085) );
  OAI22_X1 U6287 ( .A1(n5081), .A2(n6502), .B1(n5988), .B2(n5080), .ZN(n5082)
         );
  AOI21_X1 U6288 ( .B1(n6498), .B2(n5083), .A(n5082), .ZN(n5084) );
  OAI211_X1 U6289 ( .C1(n5086), .C2(n6366), .A(n5085), .B(n5084), .ZN(U3046)
         );
  XNOR2_X1 U6290 ( .A(n5088), .B(n5087), .ZN(n5101) );
  NOR2_X1 U6291 ( .A1(n6287), .A2(n6150), .ZN(n5098) );
  AOI21_X1 U6292 ( .B1(n6246), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5098), 
        .ZN(n5089) );
  OAI21_X1 U6293 ( .B1(n6156), .B2(n6254), .A(n5089), .ZN(n5090) );
  AOI21_X1 U6294 ( .B1(n6153), .B2(n6265), .A(n5090), .ZN(n5091) );
  OAI21_X1 U6295 ( .B1(n5101), .B2(n6256), .A(n5091), .ZN(U2980) );
  NAND2_X1 U6296 ( .A1(n5870), .A2(n6039), .ZN(n6286) );
  NOR2_X1 U6297 ( .A1(n5092), .A2(n5108), .ZN(n5113) );
  NAND2_X1 U6298 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5113), .ZN(n5094)
         );
  AOI21_X1 U6299 ( .B1(n6286), .B2(n5094), .A(n5093), .ZN(n5115) );
  INV_X1 U6300 ( .A(n5115), .ZN(n5097) );
  NOR2_X1 U6301 ( .A1(n5095), .A2(n5094), .ZN(n5137) );
  AOI22_X1 U6302 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5097), .B1(n5137), 
        .B2(n5096), .ZN(n5100) );
  AOI21_X1 U6303 ( .B1(n6300), .B2(n6148), .A(n5098), .ZN(n5099) );
  OAI211_X1 U6304 ( .C1(n5903), .C2(n5101), .A(n5100), .B(n5099), .ZN(U3012)
         );
  XOR2_X1 U6305 ( .A(n5103), .B(n5102), .Z(n6268) );
  NAND2_X1 U6306 ( .A1(n5105), .A2(n5104), .ZN(n5106) );
  AND2_X1 U6307 ( .A1(n5107), .A2(n5106), .ZN(n6191) );
  INV_X1 U6308 ( .A(n6191), .ZN(n5112) );
  NOR2_X1 U6309 ( .A1(n5109), .A2(n5108), .ZN(n5132) );
  NAND3_X1 U6310 ( .A1(n5699), .A2(n5132), .A3(n5116), .ZN(n5111) );
  INV_X1 U6311 ( .A(REIP_REG_5__SCAN_IN), .ZN(n5110) );
  OR2_X1 U6312 ( .A1(n6287), .A2(n5110), .ZN(n6269) );
  OAI211_X1 U6313 ( .C1(n6288), .C2(n5112), .A(n5111), .B(n6269), .ZN(n5118)
         );
  NAND2_X1 U6314 ( .A1(n5114), .A2(n5113), .ZN(n5135) );
  AOI21_X1 U6315 ( .B1(n5116), .B2(n5135), .A(n5115), .ZN(n5117) );
  AOI211_X1 U6316 ( .C1(n6304), .C2(n6268), .A(n5118), .B(n5117), .ZN(n5119)
         );
  INV_X1 U6317 ( .A(n5119), .ZN(U3013) );
  OAI21_X1 U6318 ( .B1(n3009), .B2(n5121), .A(n5120), .ZN(n6111) );
  AOI22_X1 U6319 ( .A1(n5486), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6779), .ZN(n5122) );
  OAI21_X1 U6320 ( .B1(n6111), .B2(n6776), .A(n5122), .ZN(U2882) );
  XOR2_X1 U6321 ( .A(n4904), .B(n5123), .Z(n6123) );
  INV_X1 U6322 ( .A(n6123), .ZN(n5125) );
  AOI22_X1 U6323 ( .A1(n5486), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6779), .ZN(n5124) );
  OAI21_X1 U6324 ( .B1(n5125), .B2(n6776), .A(n5124), .ZN(U2883) );
  NAND2_X1 U6325 ( .A1(n5126), .A2(n3164), .ZN(n5127) );
  NAND2_X1 U6326 ( .A1(n6106), .A2(n5127), .ZN(n6118) );
  INV_X1 U6327 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6119) );
  OAI22_X1 U6328 ( .A1(n6118), .A2(n5428), .B1(n6119), .B2(n6195), .ZN(n5128)
         );
  AOI21_X1 U6329 ( .B1(n6123), .B2(n6193), .A(n5128), .ZN(n5129) );
  INV_X1 U6330 ( .A(n5129), .ZN(U2851) );
  XNOR2_X1 U6331 ( .A(n5131), .B(n5130), .ZN(n6257) );
  INV_X1 U6332 ( .A(n5700), .ZN(n5815) );
  AND3_X1 U6333 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n5132), .ZN(n5691) );
  INV_X1 U6334 ( .A(n5133), .ZN(n5134) );
  AND2_X1 U6335 ( .A1(n6277), .A2(n5134), .ZN(n5814) );
  NAND2_X1 U6336 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5136) );
  NOR2_X1 U6337 ( .A1(n5136), .A2(n5135), .ZN(n5689) );
  OAI22_X1 U6338 ( .A1(n5815), .A2(n5691), .B1(n5814), .B2(n5689), .ZN(n6285)
         );
  OR2_X1 U6339 ( .A1(n6287), .A2(n6132), .ZN(n6261) );
  OAI21_X1 U6340 ( .B1(n6288), .B2(n6128), .A(n6261), .ZN(n5139) );
  NAND2_X1 U6341 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5137), .ZN(n6292)
         );
  NOR2_X1 U6342 ( .A1(n6292), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5138)
         );
  AOI211_X1 U6343 ( .C1(n6285), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5139), 
        .B(n5138), .ZN(n5140) );
  OAI21_X1 U6344 ( .B1(n5903), .B2(n6257), .A(n5140), .ZN(U3011) );
  INV_X1 U6345 ( .A(n5141), .ZN(n5154) );
  NOR3_X1 U6346 ( .A1(n5142), .A2(n2980), .A3(n4415), .ZN(n5143) );
  AOI21_X1 U6347 ( .B1(n5144), .B2(n5153), .A(n5143), .ZN(n5145) );
  OAI21_X1 U6348 ( .B1(n5917), .B2(n5146), .A(n5145), .ZN(n6542) );
  NOR2_X1 U6349 ( .A1(n5170), .A2(n5905), .ZN(n5149) );
  AOI222_X1 U6350 ( .A1(n6542), .A2(n6049), .B1(n5150), .B2(n5149), .C1(n5147), 
        .C2(n5148), .ZN(n5152) );
  OAI22_X1 U6351 ( .A1(n5154), .A2(n5153), .B1(n5152), .B2(n5151), .ZN(U3460)
         );
  XOR2_X1 U6352 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5156), .Z(n5723) );
  NAND2_X1 U6353 ( .A1(n5157), .A2(n6265), .ZN(n5163) );
  NOR2_X1 U6354 ( .A1(n6287), .A2(n5158), .ZN(n5720) );
  NOR2_X1 U6355 ( .A1(n6271), .A2(n5159), .ZN(n5160) );
  AOI211_X1 U6356 ( .C1(n6266), .C2(n5161), .A(n5720), .B(n5160), .ZN(n5162)
         );
  OAI211_X1 U6357 ( .C1(n5723), .C2(n6256), .A(n5163), .B(n5162), .ZN(U2956)
         );
  AOI22_X1 U6358 ( .A1(n3031), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6779), .ZN(n5167) );
  NAND2_X1 U6359 ( .A1(n3343), .A2(n5164), .ZN(n5165) );
  NAND2_X1 U6360 ( .A1(n6774), .A2(DATAI_14_), .ZN(n5166) );
  OAI211_X1 U6361 ( .C1(n5169), .C2(n6776), .A(n5167), .B(n5166), .ZN(U2861)
         );
  INV_X1 U6362 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5168) );
  OAI222_X1 U6363 ( .A1(n5428), .A2(n5716), .B1(n2970), .B2(n5169), .C1(n5168), 
        .C2(n6195), .ZN(U2829) );
  NAND2_X1 U6364 ( .A1(n6419), .A2(n5170), .ZN(n6057) );
  NAND2_X1 U6365 ( .A1(n5171), .A2(MEMORYFETCH_REG_SCAN_IN), .ZN(n5172) );
  NAND3_X1 U6366 ( .A1(n5173), .A2(n6057), .A3(n5172), .ZN(U2788) );
  INV_X1 U6367 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6368 ( .A1(n6057), .A2(n5177), .ZN(n5176) );
  INV_X1 U6369 ( .A(n5174), .ZN(n5175) );
  MUX2_X1 U6370 ( .A(n5176), .B(n5175), .S(n6609), .Z(U3474) );
  MUX2_X1 U6371 ( .A(W_R_N_REG_SCAN_IN), .B(n5177), .S(n6021), .Z(U3470) );
  OAI22_X1 U6372 ( .A1(n5180), .A2(n6186), .B1(n6155), .B2(n5494), .ZN(n5185)
         );
  OAI21_X1 U6373 ( .B1(n5183), .B2(n5182), .A(n5181), .ZN(n5725) );
  NOR2_X1 U6374 ( .A1(n5725), .A2(n6172), .ZN(n5184) );
  AOI211_X1 U6375 ( .C1(EBX_REG_29__SCAN_IN), .C2(n6143), .A(n5185), .B(n5184), 
        .ZN(n5189) );
  INV_X1 U6376 ( .A(n5186), .ZN(n5193) );
  MUX2_X1 U6377 ( .A(n5187), .B(n5193), .S(REIP_REG_29__SCAN_IN), .Z(n5188) );
  OAI211_X1 U6378 ( .C1(n5499), .C2(n6095), .A(n5189), .B(n5188), .ZN(U2798)
         );
  INV_X1 U6379 ( .A(n5509), .ZN(n5190) );
  OAI22_X1 U6380 ( .A1(n6678), .A2(n6186), .B1(n6155), .B2(n5190), .ZN(n5192)
         );
  NOR2_X1 U6381 ( .A1(n5734), .A2(n6172), .ZN(n5191) );
  AOI211_X1 U6382 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6143), .A(n5192), .B(n5191), 
        .ZN(n5196) );
  NAND2_X1 U6383 ( .A1(n5208), .A2(REIP_REG_27__SCAN_IN), .ZN(n5194) );
  MUX2_X1 U6384 ( .A(n5194), .B(n5193), .S(REIP_REG_28__SCAN_IN), .Z(n5195) );
  OAI211_X1 U6385 ( .C1(n5461), .C2(n6095), .A(n5196), .B(n5195), .ZN(U2799)
         );
  NAND2_X1 U6386 ( .A1(n5215), .A2(n5199), .ZN(n5200) );
  NAND2_X1 U6387 ( .A1(n5201), .A2(n5200), .ZN(n5744) );
  INV_X1 U6388 ( .A(n5202), .ZN(n5219) );
  NAND2_X1 U6389 ( .A1(n5219), .A2(REIP_REG_27__SCAN_IN), .ZN(n5206) );
  OAI22_X1 U6390 ( .A1(n5203), .A2(n6186), .B1(n6155), .B2(n5513), .ZN(n5204)
         );
  AOI21_X1 U6391 ( .B1(n6143), .B2(EBX_REG_27__SCAN_IN), .A(n5204), .ZN(n5205)
         );
  OAI211_X1 U6392 ( .C1(n5744), .C2(n6172), .A(n5206), .B(n5205), .ZN(n5207)
         );
  AOI21_X1 U6393 ( .B1(n5208), .B2(n5512), .A(n5207), .ZN(n5209) );
  OAI21_X1 U6394 ( .B1(n5521), .B2(n6095), .A(n5209), .ZN(U2800) );
  AOI21_X1 U6395 ( .B1(n5211), .B2(n5210), .A(n5197), .ZN(n5530) );
  INV_X1 U6396 ( .A(n5530), .ZN(n5466) );
  OAI21_X1 U6397 ( .B1(n5224), .B2(n5537), .A(n5212), .ZN(n5220) );
  OR2_X1 U6398 ( .A1(n5228), .A2(n5213), .ZN(n5214) );
  NAND2_X1 U6399 ( .A1(n5215), .A2(n5214), .ZN(n5752) );
  AOI22_X1 U6400 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6142), .B1(n6174), 
        .B2(n5526), .ZN(n5217) );
  NAND2_X1 U6401 ( .A1(n6143), .A2(EBX_REG_26__SCAN_IN), .ZN(n5216) );
  OAI211_X1 U6402 ( .C1(n5752), .C2(n6172), .A(n5217), .B(n5216), .ZN(n5218)
         );
  AOI21_X1 U6403 ( .B1(n5220), .B2(n5219), .A(n5218), .ZN(n5221) );
  OAI21_X1 U6404 ( .B1(n5466), .B2(n6095), .A(n5221), .ZN(U2801) );
  OAI21_X1 U6405 ( .B1(n5222), .B2(n5223), .A(n5210), .ZN(n5536) );
  INV_X1 U6406 ( .A(n5224), .ZN(n5233) );
  INV_X1 U6407 ( .A(n5225), .ZN(n5226) );
  AOI21_X1 U6408 ( .B1(n5247), .B2(n5240), .A(n5226), .ZN(n5227) );
  OR2_X1 U6409 ( .A1(n5228), .A2(n5227), .ZN(n5759) );
  INV_X1 U6410 ( .A(n5539), .ZN(n5229) );
  AOI22_X1 U6411 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6142), .B1(n6174), 
        .B2(n5229), .ZN(n5231) );
  NAND2_X1 U6412 ( .A1(n6143), .A2(EBX_REG_25__SCAN_IN), .ZN(n5230) );
  OAI211_X1 U6413 ( .C1(n5759), .C2(n6172), .A(n5231), .B(n5230), .ZN(n5232)
         );
  AOI21_X1 U6414 ( .B1(n5233), .B2(n5537), .A(n5232), .ZN(n5236) );
  INV_X1 U6415 ( .A(n5255), .ZN(n5234) );
  NOR3_X1 U6416 ( .A1(n5234), .A2(REIP_REG_24__SCAN_IN), .A3(n5554), .ZN(n5243) );
  OAI21_X1 U6417 ( .B1(n5243), .B2(n5254), .A(REIP_REG_25__SCAN_IN), .ZN(n5235) );
  OAI211_X1 U6418 ( .C1(n5536), .C2(n6095), .A(n5236), .B(n5235), .ZN(U2802)
         );
  AOI21_X1 U6419 ( .B1(n5239), .B2(n5238), .A(n5222), .ZN(n5552) );
  INV_X1 U6420 ( .A(n5552), .ZN(n5471) );
  XNOR2_X1 U6421 ( .A(n5247), .B(n5240), .ZN(n5769) );
  OAI22_X1 U6422 ( .A1(n5241), .A2(n6186), .B1(n6155), .B2(n5550), .ZN(n5242)
         );
  OAI21_X1 U6423 ( .B1(n5244), .B2(n5245), .A(n5238), .ZN(n5568) );
  OAI22_X1 U6424 ( .A1(n5246), .A2(n6186), .B1(n6155), .B2(n5555), .ZN(n5253)
         );
  INV_X1 U6425 ( .A(n5247), .ZN(n5251) );
  INV_X1 U6426 ( .A(n5260), .ZN(n5249) );
  OAI21_X1 U6427 ( .B1(n5273), .B2(n5249), .A(n5248), .ZN(n5250) );
  NAND2_X1 U6428 ( .A1(n5251), .A2(n5250), .ZN(n5781) );
  NOR2_X1 U6429 ( .A1(n5781), .A2(n6172), .ZN(n5252) );
  AOI211_X1 U6430 ( .C1(n6143), .C2(EBX_REG_23__SCAN_IN), .A(n5253), .B(n5252), 
        .ZN(n5257) );
  OAI21_X1 U6431 ( .B1(n5255), .B2(REIP_REG_23__SCAN_IN), .A(n5254), .ZN(n5256) );
  OAI211_X1 U6432 ( .C1(n5568), .C2(n6095), .A(n5257), .B(n5256), .ZN(U2804)
         );
  AOI21_X1 U6433 ( .B1(n5259), .B2(n5258), .A(n5244), .ZN(n5576) );
  INV_X1 U6434 ( .A(n5576), .ZN(n5476) );
  XNOR2_X1 U6435 ( .A(n5273), .B(n5260), .ZN(n5792) );
  INV_X1 U6436 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5409) );
  INV_X1 U6437 ( .A(n5574), .ZN(n5261) );
  AOI22_X1 U6438 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6142), .B1(n6174), 
        .B2(n5261), .ZN(n5262) );
  OAI21_X1 U6439 ( .B1(n6179), .B2(n5409), .A(n5262), .ZN(n5264) );
  NOR2_X1 U6440 ( .A1(n3030), .A2(REIP_REG_22__SCAN_IN), .ZN(n5263) );
  AOI211_X1 U6441 ( .C1(n6161), .C2(n5792), .A(n5264), .B(n5263), .ZN(n5267)
         );
  NOR2_X1 U6442 ( .A1(n5588), .A2(REIP_REG_21__SCAN_IN), .ZN(n5265) );
  AND2_X1 U6443 ( .A1(n3027), .A2(n5265), .ZN(n5276) );
  OAI21_X1 U6444 ( .B1(n5276), .B2(n5287), .A(REIP_REG_22__SCAN_IN), .ZN(n5266) );
  OAI211_X1 U6445 ( .C1(n5476), .C2(n6095), .A(n5267), .B(n5266), .ZN(U2805)
         );
  OAI21_X1 U6446 ( .B1(n5268), .B2(n5269), .A(n5258), .ZN(n5585) );
  NAND2_X1 U6447 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  NAND2_X1 U6448 ( .A1(n5273), .A2(n5272), .ZN(n5801) );
  OAI21_X1 U6449 ( .B1(n5801), .B2(n6172), .A(n5275), .ZN(n5277) );
  AOI211_X1 U6450 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5287), .A(n5277), .B(n5276), .ZN(n5278) );
  OAI21_X1 U6451 ( .B1(n5585), .B2(n6095), .A(n5278), .ZN(U2806) );
  AOI21_X1 U6452 ( .B1(n5280), .B2(n5279), .A(n5268), .ZN(n5592) );
  INV_X1 U6453 ( .A(n5592), .ZN(n5481) );
  OAI22_X1 U6454 ( .A1(n3106), .A2(n6186), .B1(n6155), .B2(n5590), .ZN(n5286)
         );
  MUX2_X1 U6455 ( .A(n2975), .B(n5418), .S(n5281), .Z(n5283) );
  XOR2_X1 U6456 ( .A(n5284), .B(n5283), .Z(n5808) );
  NOR2_X1 U6457 ( .A1(n5808), .A2(n6172), .ZN(n5285) );
  AOI211_X1 U6458 ( .C1(n6143), .C2(EBX_REG_20__SCAN_IN), .A(n5286), .B(n5285), 
        .ZN(n5289) );
  OAI21_X1 U6459 ( .B1(n3027), .B2(REIP_REG_20__SCAN_IN), .A(n5287), .ZN(n5288) );
  OAI211_X1 U6460 ( .C1(n5481), .C2(n6095), .A(n5289), .B(n5288), .ZN(U2807)
         );
  AND2_X1 U6461 ( .A1(n5290), .A2(n5291), .ZN(n5292) );
  OR2_X1 U6462 ( .A1(n5292), .A2(n3006), .ZN(n5626) );
  INV_X1 U6464 ( .A(n5293), .ZN(n5295) );
  NOR2_X1 U6465 ( .A1(n5295), .A2(n5294), .ZN(n6085) );
  NOR2_X1 U6466 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5295), .ZN(n6103) );
  OAI33_X1 U6467 ( .A1(1'b0), .A2(n6085), .A3(REIP_REG_16__SCAN_IN), .B1(n4355), .B2(n6098), .B3(n6103), .ZN(n5301) );
  XNOR2_X1 U6468 ( .A(n5297), .B(n5432), .ZN(n5855) );
  AOI22_X1 U6469 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6143), .B1(n5629), .B2(n6174), .ZN(n5298) );
  OAI21_X1 U6470 ( .B1(n6172), .B2(n5855), .A(n5298), .ZN(n5299) );
  AOI211_X1 U6471 ( .C1(n6142), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6167), 
        .B(n5299), .ZN(n5300) );
  OAI211_X1 U6472 ( .C1(n6095), .C2(n5626), .A(n5301), .B(n5300), .ZN(U2811)
         );
  OAI21_X1 U6473 ( .B1(n5302), .B2(n5305), .A(n5304), .ZN(n5643) );
  NAND2_X1 U6474 ( .A1(n5307), .A2(n5306), .ZN(n5313) );
  INV_X1 U6475 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5445) );
  NOR2_X1 U6476 ( .A1(n5322), .A2(n5308), .ZN(n5309) );
  OR2_X1 U6477 ( .A1(n5442), .A2(n5309), .ZN(n5879) );
  OAI22_X1 U6478 ( .A1(n5445), .A2(n6179), .B1(n6172), .B2(n5879), .ZN(n5310)
         );
  AOI211_X1 U6479 ( .C1(n6142), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6167), 
        .B(n5310), .ZN(n5311) );
  OAI21_X1 U6480 ( .B1(n5639), .B2(n6155), .A(n5311), .ZN(n5312) );
  AOI21_X1 U6481 ( .B1(n5313), .B2(n6098), .A(n5312), .ZN(n5314) );
  OAI21_X1 U6482 ( .B1(n5643), .B2(n6095), .A(n5314), .ZN(U2813) );
  INV_X1 U6483 ( .A(n5315), .ZN(n5316) );
  NOR2_X1 U6484 ( .A1(n5316), .A2(n5317), .ZN(n5318) );
  INV_X1 U6485 ( .A(n5648), .ZN(n5319) );
  OAI22_X1 U6486 ( .A1(n5651), .A2(n6095), .B1(n6155), .B2(n5319), .ZN(n5331)
         );
  AND2_X1 U6487 ( .A1(n5321), .A2(n5320), .ZN(n5323) );
  OR2_X1 U6488 ( .A1(n5323), .A2(n5322), .ZN(n6035) );
  NAND2_X1 U6489 ( .A1(n6134), .A2(n5324), .ZN(n5353) );
  OAI22_X1 U6490 ( .A1(n5325), .A2(n6186), .B1(n5646), .B2(n5353), .ZN(n5326)
         );
  AOI211_X1 U6491 ( .C1(n6143), .C2(EBX_REG_13__SCAN_IN), .A(n6167), .B(n5326), 
        .ZN(n5329) );
  OAI211_X1 U6492 ( .C1(REIP_REG_13__SCAN_IN), .C2(REIP_REG_12__SCAN_IN), .A(
        n5339), .B(n5327), .ZN(n5328) );
  OAI211_X1 U6493 ( .C1(n6035), .C2(n6172), .A(n5329), .B(n5328), .ZN(n5330)
         );
  OR2_X1 U6494 ( .A1(n5331), .A2(n5330), .ZN(U2814) );
  OAI21_X1 U6495 ( .B1(n3022), .B2(n5332), .A(n5315), .ZN(n5662) );
  INV_X1 U6496 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6690) );
  OAI22_X1 U6497 ( .A1(n6690), .A2(n6179), .B1(n5338), .B2(n5353), .ZN(n5337)
         );
  XNOR2_X1 U6498 ( .A(n5347), .B(n5333), .ZN(n5450) );
  NOR2_X1 U6499 ( .A1(n5450), .A2(n6172), .ZN(n5336) );
  INV_X1 U6500 ( .A(n6167), .ZN(n6144) );
  OAI21_X1 U6501 ( .B1(n6186), .B2(n3112), .A(n6144), .ZN(n5335) );
  NOR2_X1 U6502 ( .A1(n6155), .A2(n5658), .ZN(n5334) );
  NOR4_X1 U6503 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n5341)
         );
  NAND2_X1 U6504 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  OAI211_X1 U6505 ( .C1(n5662), .C2(n6095), .A(n5341), .B(n5340), .ZN(U2815)
         );
  AND2_X1 U6506 ( .A1(n5342), .A2(n5343), .ZN(n5344) );
  OR2_X1 U6507 ( .A1(n5344), .A2(n3022), .ZN(n6248) );
  OAI22_X1 U6508 ( .A1(n6248), .A2(n6095), .B1(n6155), .B2(n5345), .ZN(n5357)
         );
  OAI21_X1 U6509 ( .B1(n5346), .B2(n5348), .A(n5347), .ZN(n5349) );
  INV_X1 U6510 ( .A(n5349), .ZN(n5892) );
  OAI22_X1 U6511 ( .A1(n6651), .A2(n6179), .B1(n5350), .B2(n6186), .ZN(n5351)
         );
  AOI211_X1 U6512 ( .C1(n6161), .C2(n5892), .A(n6167), .B(n5351), .ZN(n5352)
         );
  OAI221_X1 U6513 ( .B1(REIP_REG_11__SCAN_IN), .B2(n5355), .C1(n5354), .C2(
        n5353), .A(n5352), .ZN(n5356) );
  OR2_X1 U6514 ( .A1(n5357), .A2(n5356), .ZN(U2816) );
  INV_X1 U6515 ( .A(n5342), .ZN(n5358) );
  AOI21_X1 U6516 ( .B1(n5359), .B2(n5120), .A(n5358), .ZN(n5671) );
  INV_X1 U6517 ( .A(n5671), .ZN(n5492) );
  INV_X1 U6518 ( .A(n6134), .ZN(n5399) );
  NOR2_X1 U6519 ( .A1(n5399), .A2(n5360), .ZN(n6117) );
  AND2_X1 U6520 ( .A1(n5361), .A2(n5364), .ZN(n6110) );
  OAI21_X1 U6521 ( .B1(n6117), .B2(n6110), .A(REIP_REG_10__SCAN_IN), .ZN(n5370) );
  INV_X1 U6522 ( .A(n5669), .ZN(n5368) );
  INV_X1 U6523 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5454) );
  NOR2_X1 U6524 ( .A1(n3043), .A2(n5362), .ZN(n5363) );
  OR2_X1 U6525 ( .A1(n5346), .A2(n5363), .ZN(n6289) );
  OAI22_X1 U6526 ( .A1(n5454), .A2(n6179), .B1(n6172), .B2(n6289), .ZN(n5367)
         );
  NAND3_X1 U6527 ( .A1(n5364), .A2(REIP_REG_9__SCAN_IN), .A3(n4392), .ZN(n5365) );
  OAI211_X1 U6528 ( .C1(n6186), .C2(n3604), .A(n6144), .B(n5365), .ZN(n5366)
         );
  AOI211_X1 U6529 ( .C1(n6174), .C2(n5368), .A(n5367), .B(n5366), .ZN(n5369)
         );
  OAI211_X1 U6530 ( .C1(n5492), .C2(n6095), .A(n5370), .B(n5369), .ZN(U2817)
         );
  OAI21_X1 U6531 ( .B1(n6159), .B2(n6157), .A(n5371), .ZN(n6170) );
  INV_X1 U6532 ( .A(n6159), .ZN(n6116) );
  NOR3_X1 U6533 ( .A1(n6157), .A2(n5390), .A3(n5372), .ZN(n5373) );
  AOI22_X1 U6534 ( .A1(n6116), .A2(n5373), .B1(n6143), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5380) );
  INV_X1 U6535 ( .A(n5374), .ZN(n5375) );
  AOI22_X1 U6536 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6142), .B1(n6174), 
        .B2(n5375), .ZN(n5379) );
  NAND2_X1 U6537 ( .A1(n6161), .A2(n5376), .ZN(n5378) );
  NAND2_X1 U6538 ( .A1(n6177), .A2(n4654), .ZN(n5377) );
  NAND4_X1 U6539 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), .ZN(n5381)
         );
  AOI21_X1 U6540 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6170), .A(n5381), .ZN(n5382)
         );
  OAI21_X1 U6541 ( .B1(n5383), .B2(n5405), .A(n5382), .ZN(U2824) );
  NAND2_X1 U6542 ( .A1(n6143), .A2(EBX_REG_2__SCAN_IN), .ZN(n5389) );
  INV_X1 U6543 ( .A(n5384), .ZN(n5385) );
  AOI22_X1 U6544 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6174), 
        .B2(n5385), .ZN(n5388) );
  NAND2_X1 U6545 ( .A1(n6177), .A2(n5386), .ZN(n5387) );
  NAND3_X1 U6546 ( .A1(n5389), .A2(n5388), .A3(n5387), .ZN(n5395) );
  NOR3_X1 U6547 ( .A1(n5391), .A2(n6135), .A3(n5390), .ZN(n5393) );
  AOI21_X1 U6548 ( .B1(n6116), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5392) );
  NOR2_X1 U6549 ( .A1(n5393), .A2(n5392), .ZN(n5394) );
  AOI211_X1 U6550 ( .C1(n5396), .C2(n6161), .A(n5395), .B(n5394), .ZN(n5397)
         );
  OAI21_X1 U6551 ( .B1(n5405), .B2(n5398), .A(n5397), .ZN(U2825) );
  AOI22_X1 U6552 ( .A1(EBX_REG_0__SCAN_IN), .A2(n6143), .B1(n6177), .B2(n6421), 
        .ZN(n5403) );
  NAND2_X1 U6553 ( .A1(n6186), .A2(n6155), .ZN(n5401) );
  OAI22_X1 U6554 ( .A1(n5399), .A2(n6752), .B1(n6172), .B2(n5904), .ZN(n5400)
         );
  AOI21_X1 U6555 ( .B1(n5401), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5400), 
        .ZN(n5402) );
  OAI211_X1 U6556 ( .C1(n5405), .C2(n5404), .A(n5403), .B(n5402), .ZN(U2827)
         );
  OAI22_X1 U6557 ( .A1(n5687), .A2(n5428), .B1(n5406), .B2(n6195), .ZN(U2828)
         );
  OAI222_X1 U6558 ( .A1(n6650), .A2(n6195), .B1(n5428), .B2(n5725), .C1(n5499), 
        .C2(n2970), .ZN(U2830) );
  INV_X1 U6559 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5407) );
  OAI222_X1 U6560 ( .A1(n5744), .A2(n5428), .B1(n5407), .B2(n6195), .C1(n5521), 
        .C2(n2970), .ZN(U2832) );
  INV_X1 U6561 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6648) );
  OAI222_X1 U6562 ( .A1(n5752), .A2(n5428), .B1(n6648), .B2(n6195), .C1(n5466), 
        .C2(n2970), .ZN(U2833) );
  INV_X1 U6563 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6742) );
  OAI222_X1 U6564 ( .A1(n5759), .A2(n5428), .B1(n6742), .B2(n6195), .C1(n5536), 
        .C2(n2970), .ZN(U2834) );
  INV_X1 U6565 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6677) );
  OAI222_X1 U6566 ( .A1(n6677), .A2(n6195), .B1(n5428), .B2(n5769), .C1(n2970), 
        .C2(n5471), .ZN(U2835) );
  INV_X1 U6567 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5408) );
  OAI222_X1 U6568 ( .A1(n5408), .A2(n6195), .B1(n5428), .B2(n5781), .C1(n5568), 
        .C2(n2970), .ZN(U2836) );
  INV_X1 U6569 ( .A(n5792), .ZN(n5410) );
  OAI222_X1 U6570 ( .A1(n5476), .A2(n2970), .B1(n5428), .B2(n5410), .C1(n6195), 
        .C2(n5409), .ZN(U2837) );
  INV_X1 U6571 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5411) );
  OAI222_X1 U6572 ( .A1(n5801), .A2(n5428), .B1(n5411), .B2(n6195), .C1(n5585), 
        .C2(n2970), .ZN(U2838) );
  INV_X1 U6573 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5412) );
  OAI222_X1 U6574 ( .A1(n5808), .A2(n5428), .B1(n6195), .B2(n5412), .C1(n2970), 
        .C2(n5481), .ZN(U2839) );
  NAND2_X1 U6575 ( .A1(n5413), .A2(n5414), .ZN(n5415) );
  AND2_X1 U6576 ( .A1(n5279), .A2(n5415), .ZN(n6032) );
  INV_X1 U6577 ( .A(n6032), .ZN(n5601) );
  INV_X1 U6578 ( .A(n5416), .ZN(n5420) );
  MUX2_X1 U6579 ( .A(n5418), .B(n5417), .S(n4001), .Z(n5423) );
  INV_X1 U6580 ( .A(n5423), .ZN(n5419) );
  NAND2_X1 U6581 ( .A1(n5420), .A2(n5419), .ZN(n5425) );
  XNOR2_X1 U6582 ( .A(n5425), .B(n5421), .ZN(n6026) );
  INV_X1 U6583 ( .A(n6026), .ZN(n5830) );
  AOI22_X1 U6584 ( .A1(n5830), .A2(n6192), .B1(n5452), .B2(EBX_REG_19__SCAN_IN), .ZN(n5422) );
  OAI21_X1 U6585 ( .B1(n5601), .B2(n2970), .A(n5422), .ZN(U2840) );
  NAND2_X1 U6586 ( .A1(n5416), .A2(n5423), .ZN(n5424) );
  NAND2_X1 U6587 ( .A1(n5425), .A2(n5424), .ZN(n6079) );
  INV_X1 U6588 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6706) );
  OAI21_X1 U6589 ( .B1(n5426), .B2(n5427), .A(n5413), .ZN(n6777) );
  OAI222_X1 U6590 ( .A1(n6079), .A2(n5428), .B1(n6195), .B2(n6706), .C1(n2970), 
        .C2(n6777), .ZN(U2841) );
  INV_X1 U6591 ( .A(n5426), .ZN(n5429) );
  OAI21_X1 U6592 ( .B1(n3006), .B2(n5430), .A(n5429), .ZN(n6088) );
  OAI21_X1 U6593 ( .B1(n5297), .B2(n5432), .A(n5431), .ZN(n5433) );
  AND2_X1 U6594 ( .A1(n5433), .A2(n5416), .ZN(n6089) );
  INV_X1 U6595 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6661) );
  NOR2_X1 U6596 ( .A1(n6195), .A2(n6661), .ZN(n5434) );
  AOI21_X1 U6597 ( .B1(n6089), .B2(n6192), .A(n5434), .ZN(n5435) );
  OAI21_X1 U6598 ( .B1(n6088), .B2(n2970), .A(n5435), .ZN(U2842) );
  OAI22_X1 U6599 ( .A1(n5855), .A2(n5428), .B1(n5436), .B2(n6195), .ZN(n5437)
         );
  INV_X1 U6600 ( .A(n5437), .ZN(n5438) );
  OAI21_X1 U6601 ( .B1(n5626), .B2(n2970), .A(n5438), .ZN(U2843) );
  NAND2_X1 U6602 ( .A1(n5304), .A2(n5439), .ZN(n5440) );
  NAND2_X1 U6603 ( .A1(n5290), .A2(n5440), .ZN(n6096) );
  OR2_X1 U6604 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  AND2_X1 U6605 ( .A1(n5297), .A2(n5443), .ZN(n6099) );
  AOI22_X1 U6606 ( .A1(n6099), .A2(n6192), .B1(EBX_REG_15__SCAN_IN), .B2(n5452), .ZN(n5444) );
  OAI21_X1 U6607 ( .B1(n6096), .B2(n2970), .A(n5444), .ZN(U2844) );
  OAI22_X1 U6608 ( .A1(n5879), .A2(n5428), .B1(n5445), .B2(n6195), .ZN(n5446)
         );
  INV_X1 U6609 ( .A(n5446), .ZN(n5447) );
  OAI21_X1 U6610 ( .B1(n5643), .B2(n2970), .A(n5447), .ZN(U2845) );
  INV_X1 U6611 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6755) );
  OAI22_X1 U6612 ( .A1(n6035), .A2(n5428), .B1(n6755), .B2(n6195), .ZN(n5448)
         );
  INV_X1 U6613 ( .A(n5448), .ZN(n5449) );
  OAI21_X1 U6614 ( .B1(n5651), .B2(n2970), .A(n5449), .ZN(U2846) );
  INV_X1 U6615 ( .A(n5450), .ZN(n6275) );
  AOI22_X1 U6616 ( .A1(n6275), .A2(n6192), .B1(n5452), .B2(EBX_REG_12__SCAN_IN), .ZN(n5451) );
  OAI21_X1 U6617 ( .B1(n5662), .B2(n2970), .A(n5451), .ZN(U2847) );
  AOI22_X1 U6618 ( .A1(n5892), .A2(n6192), .B1(n5452), .B2(EBX_REG_11__SCAN_IN), .ZN(n5453) );
  OAI21_X1 U6619 ( .B1(n6248), .B2(n2970), .A(n5453), .ZN(U2848) );
  OAI22_X1 U6620 ( .A1(n6289), .A2(n5428), .B1(n5454), .B2(n6195), .ZN(n5455)
         );
  INV_X1 U6621 ( .A(n5455), .ZN(n5456) );
  OAI21_X1 U6622 ( .B1(n5492), .B2(n2970), .A(n5456), .ZN(U2849) );
  AOI22_X1 U6623 ( .A1(n3031), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6779), .ZN(n5458) );
  NAND2_X1 U6624 ( .A1(n6774), .A2(DATAI_13_), .ZN(n5457) );
  OAI211_X1 U6625 ( .C1(n5499), .C2(n6776), .A(n5458), .B(n5457), .ZN(U2862)
         );
  AOI22_X1 U6626 ( .A1(n3031), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6779), .ZN(n5460) );
  NAND2_X1 U6627 ( .A1(n6774), .A2(DATAI_12_), .ZN(n5459) );
  OAI211_X1 U6628 ( .C1(n5461), .C2(n6776), .A(n5460), .B(n5459), .ZN(U2863)
         );
  AOI22_X1 U6629 ( .A1(n3031), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6779), .ZN(n5463) );
  NAND2_X1 U6630 ( .A1(n6774), .A2(DATAI_11_), .ZN(n5462) );
  OAI211_X1 U6631 ( .C1(n5521), .C2(n6776), .A(n5463), .B(n5462), .ZN(U2864)
         );
  AOI22_X1 U6632 ( .A1(n3031), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6779), .ZN(n5465) );
  NAND2_X1 U6633 ( .A1(n6774), .A2(DATAI_10_), .ZN(n5464) );
  OAI211_X1 U6634 ( .C1(n5466), .C2(n6776), .A(n5465), .B(n5464), .ZN(U2865)
         );
  AOI22_X1 U6635 ( .A1(n3031), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6779), .ZN(n5468) );
  NAND2_X1 U6636 ( .A1(n6774), .A2(DATAI_9_), .ZN(n5467) );
  OAI211_X1 U6637 ( .C1(n5536), .C2(n6776), .A(n5468), .B(n5467), .ZN(U2866)
         );
  AOI22_X1 U6638 ( .A1(n3031), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6779), .ZN(n5470) );
  NAND2_X1 U6639 ( .A1(n6774), .A2(DATAI_8_), .ZN(n5469) );
  OAI211_X1 U6640 ( .C1(n5471), .C2(n6776), .A(n5470), .B(n5469), .ZN(U2867)
         );
  AOI22_X1 U6641 ( .A1(n3031), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6779), .ZN(n5473) );
  NAND2_X1 U6642 ( .A1(n6774), .A2(DATAI_7_), .ZN(n5472) );
  OAI211_X1 U6643 ( .C1(n5568), .C2(n6776), .A(n5473), .B(n5472), .ZN(U2868)
         );
  AOI22_X1 U6644 ( .A1(n3031), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6779), .ZN(n5475) );
  NAND2_X1 U6645 ( .A1(n6774), .A2(DATAI_6_), .ZN(n5474) );
  OAI211_X1 U6646 ( .C1(n5476), .C2(n6776), .A(n5475), .B(n5474), .ZN(U2869)
         );
  AOI22_X1 U6647 ( .A1(n3031), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6779), .ZN(n5478) );
  NAND2_X1 U6648 ( .A1(n6774), .A2(DATAI_5_), .ZN(n5477) );
  OAI211_X1 U6649 ( .C1(n5585), .C2(n6776), .A(n5478), .B(n5477), .ZN(U2870)
         );
  AOI22_X1 U6650 ( .A1(n3031), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6779), .ZN(n5480) );
  NAND2_X1 U6651 ( .A1(n6774), .A2(DATAI_4_), .ZN(n5479) );
  OAI211_X1 U6652 ( .C1(n5481), .C2(n6776), .A(n5480), .B(n5479), .ZN(U2871)
         );
  AOI22_X1 U6653 ( .A1(n3031), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6779), .ZN(n5483) );
  NAND2_X1 U6654 ( .A1(n6774), .A2(DATAI_0_), .ZN(n5482) );
  OAI211_X1 U6655 ( .C1(n5626), .C2(n6776), .A(n5483), .B(n5482), .ZN(U2875)
         );
  AOI22_X1 U6656 ( .A1(n5486), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6779), .ZN(n5484) );
  OAI21_X1 U6657 ( .B1(n6096), .B2(n6776), .A(n5484), .ZN(U2876) );
  AOI22_X1 U6658 ( .A1(n5486), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6779), .ZN(n5485) );
  OAI21_X1 U6659 ( .B1(n5643), .B2(n6776), .A(n5485), .ZN(U2877) );
  INV_X1 U6660 ( .A(DATAI_13_), .ZN(n6723) );
  OAI222_X1 U6661 ( .A1(n5651), .A2(n6776), .B1(n5491), .B2(n6723), .C1(n5489), 
        .C2(n6208), .ZN(U2878) );
  AOI22_X1 U6662 ( .A1(n5486), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n6779), .ZN(n5487) );
  OAI21_X1 U6663 ( .B1(n5662), .B2(n6776), .A(n5487), .ZN(U2879) );
  INV_X1 U6664 ( .A(DATAI_11_), .ZN(n5488) );
  OAI222_X1 U6665 ( .A1(n6248), .A2(n6776), .B1(n5491), .B2(n5488), .C1(n5489), 
        .C2(n6679), .ZN(U2880) );
  INV_X1 U6666 ( .A(DATAI_10_), .ZN(n5490) );
  OAI222_X1 U6667 ( .A1(n5492), .A2(n6776), .B1(n5491), .B2(n5490), .C1(n5489), 
        .C2(n6693), .ZN(U2881) );
  NOR2_X1 U6668 ( .A1(n6287), .A2(n5493), .ZN(n5729) );
  NOR2_X1 U6669 ( .A1(n6254), .A2(n5494), .ZN(n5495) );
  AOI211_X1 U6670 ( .C1(n6246), .C2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5729), 
        .B(n5495), .ZN(n5498) );
  INV_X1 U6671 ( .A(n5737), .ZN(n5697) );
  INV_X1 U6672 ( .A(n5516), .ZN(n5501) );
  AOI21_X1 U6673 ( .B1(n5697), .B2(n5501), .A(n2992), .ZN(n5496) );
  XNOR2_X1 U6674 ( .A(n5496), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5724)
         );
  NAND2_X1 U6675 ( .A1(n5724), .A2(n4329), .ZN(n5497) );
  OAI211_X1 U6676 ( .C1(n5499), .C2(n6258), .A(n5498), .B(n5497), .ZN(U2957)
         );
  INV_X1 U6677 ( .A(n2992), .ZN(n5504) );
  NAND3_X1 U6678 ( .A1(n5501), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5500), .ZN(n5503) );
  NAND3_X1 U6679 ( .A1(n5515), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n5517), .ZN(n5502) );
  NAND3_X1 U6680 ( .A1(n5504), .A2(n5503), .A3(n5502), .ZN(n5505) );
  NAND2_X1 U6681 ( .A1(n5506), .A2(n6265), .ZN(n5511) );
  NOR2_X1 U6682 ( .A1(n6287), .A2(n5507), .ZN(n5736) );
  NOR2_X1 U6683 ( .A1(n6271), .A2(n6678), .ZN(n5508) );
  AOI211_X1 U6684 ( .C1(n6266), .C2(n5509), .A(n5736), .B(n5508), .ZN(n5510)
         );
  OAI211_X1 U6685 ( .C1(n5741), .C2(n6256), .A(n5511), .B(n5510), .ZN(U2958)
         );
  NOR2_X1 U6686 ( .A1(n6287), .A2(n5512), .ZN(n5746) );
  NOR2_X1 U6687 ( .A1(n6254), .A2(n5513), .ZN(n5514) );
  AOI211_X1 U6688 ( .C1(n6246), .C2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5746), 
        .B(n5514), .ZN(n5520) );
  NAND2_X1 U6689 ( .A1(n5516), .A2(n5515), .ZN(n5518) );
  XNOR2_X1 U6690 ( .A(n5518), .B(n5517), .ZN(n5743) );
  NAND2_X1 U6691 ( .A1(n5743), .A2(n4329), .ZN(n5519) );
  OAI211_X1 U6692 ( .C1(n5521), .C2(n6258), .A(n5520), .B(n5519), .ZN(U2959)
         );
  NAND2_X1 U6693 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  XNOR2_X1 U6694 ( .A(n5525), .B(n5524), .ZN(n5758) );
  NAND2_X1 U6695 ( .A1(n6266), .A2(n5526), .ZN(n5527) );
  NAND2_X1 U6696 ( .A1(n6247), .A2(REIP_REG_26__SCAN_IN), .ZN(n5751) );
  OAI211_X1 U6697 ( .C1(n6271), .C2(n5528), .A(n5527), .B(n5751), .ZN(n5529)
         );
  AOI21_X1 U6698 ( .B1(n5530), .B2(n6265), .A(n5529), .ZN(n5531) );
  OAI21_X1 U6699 ( .B1(n5758), .B2(n6256), .A(n5531), .ZN(U2960) );
  INV_X1 U6700 ( .A(n5532), .ZN(n5533) );
  AOI21_X1 U6701 ( .B1(n5535), .B2(n5534), .A(n5533), .ZN(n5768) );
  INV_X1 U6702 ( .A(n5536), .ZN(n5541) );
  NOR2_X1 U6703 ( .A1(n6287), .A2(n5537), .ZN(n5761) );
  AOI21_X1 U6704 ( .B1(n6246), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5761), 
        .ZN(n5538) );
  OAI21_X1 U6705 ( .B1(n5539), .B2(n6254), .A(n5538), .ZN(n5540) );
  AOI21_X1 U6706 ( .B1(n5541), .B2(n6265), .A(n5540), .ZN(n5542) );
  OAI21_X1 U6707 ( .B1(n5768), .B2(n6256), .A(n5542), .ZN(U2961) );
  XNOR2_X1 U6708 ( .A(n5609), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5597)
         );
  OR2_X1 U6709 ( .A1(n5609), .A2(n5833), .ZN(n5543) );
  NAND2_X1 U6710 ( .A1(n5609), .A2(n6736), .ZN(n5544) );
  XNOR2_X1 U6711 ( .A(n5674), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5580)
         );
  AOI21_X1 U6712 ( .B1(n2989), .B2(n5545), .A(n5546), .ZN(n5571) );
  NOR3_X1 U6713 ( .A1(n5655), .A2(n5795), .A3(n5564), .ZN(n5547) );
  INV_X1 U6714 ( .A(n5546), .ZN(n5578) );
  OR2_X1 U6715 ( .A1(n2989), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5569)
         );
  AOI22_X1 U6716 ( .A1(n5571), .A2(n5547), .B1(n5563), .B2(n5564), .ZN(n5548)
         );
  XNOR2_X1 U6717 ( .A(n5548), .B(n5774), .ZN(n5779) );
  NAND2_X1 U6718 ( .A1(n6246), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5549)
         );
  NAND2_X1 U6719 ( .A1(n6247), .A2(REIP_REG_24__SCAN_IN), .ZN(n5770) );
  OAI211_X1 U6720 ( .C1(n6254), .C2(n5550), .A(n5549), .B(n5770), .ZN(n5551)
         );
  AOI21_X1 U6721 ( .B1(n5552), .B2(n6265), .A(n5551), .ZN(n5553) );
  OAI21_X1 U6722 ( .B1(n5779), .B2(n6256), .A(n5553), .ZN(U2962) );
  NOR2_X1 U6723 ( .A1(n6287), .A2(n5554), .ZN(n5783) );
  NOR2_X1 U6724 ( .A1(n6254), .A2(n5555), .ZN(n5556) );
  AOI211_X1 U6725 ( .C1(n6246), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5783), 
        .B(n5556), .ZN(n5567) );
  NAND2_X1 U6726 ( .A1(n5609), .A2(n5864), .ZN(n5557) );
  NAND2_X1 U6727 ( .A1(n5558), .A2(n5557), .ZN(n5624) );
  AND2_X1 U6728 ( .A1(n5674), .A2(n5852), .ZN(n5620) );
  NOR2_X1 U6729 ( .A1(n5559), .A2(n5703), .ZN(n5560) );
  NAND2_X1 U6730 ( .A1(n2989), .A2(n5560), .ZN(n5561) );
  NOR2_X1 U6731 ( .A1(n5610), .A2(n5561), .ZN(n5562) );
  NAND2_X1 U6732 ( .A1(n5780), .A2(n4329), .ZN(n5566) );
  OAI211_X1 U6733 ( .C1(n5568), .C2(n6258), .A(n5567), .B(n5566), .ZN(U2963)
         );
  OAI21_X1 U6734 ( .B1(n5655), .B2(n5795), .A(n5569), .ZN(n5570) );
  XNOR2_X1 U6735 ( .A(n5571), .B(n5570), .ZN(n5798) );
  NOR2_X1 U6736 ( .A1(n6287), .A2(n5572), .ZN(n5791) );
  AOI21_X1 U6737 ( .B1(n6246), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5791), 
        .ZN(n5573) );
  OAI21_X1 U6738 ( .B1(n5574), .B2(n6254), .A(n5573), .ZN(n5575) );
  AOI21_X1 U6739 ( .B1(n5576), .B2(n6265), .A(n5575), .ZN(n5577) );
  OAI21_X1 U6740 ( .B1(n5798), .B2(n6256), .A(n5577), .ZN(U2964) );
  OAI21_X1 U6741 ( .B1(n5580), .B2(n5579), .A(n5578), .ZN(n5799) );
  NAND2_X1 U6742 ( .A1(n5799), .A2(n4329), .ZN(n5584) );
  NOR2_X1 U6743 ( .A1(n6287), .A2(n3059), .ZN(n5803) );
  NOR2_X1 U6744 ( .A1(n6254), .A2(n5581), .ZN(n5582) );
  AOI211_X1 U6745 ( .C1(n6246), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5803), 
        .B(n5582), .ZN(n5583) );
  OAI211_X1 U6746 ( .C1(n6258), .C2(n5585), .A(n5584), .B(n5583), .ZN(U2965)
         );
  XNOR2_X1 U6747 ( .A(n2989), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5586)
         );
  XNOR2_X1 U6748 ( .A(n5587), .B(n5586), .ZN(n5824) );
  NOR2_X1 U6749 ( .A1(n6287), .A2(n5588), .ZN(n5811) );
  AOI21_X1 U6750 ( .B1(n6246), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5811), 
        .ZN(n5589) );
  OAI21_X1 U6751 ( .B1(n5590), .B2(n6254), .A(n5589), .ZN(n5591) );
  AOI21_X1 U6752 ( .B1(n5592), .B2(n6265), .A(n5591), .ZN(n5593) );
  OAI21_X1 U6753 ( .B1(n5824), .B2(n6256), .A(n5593), .ZN(U2966) );
  NOR2_X1 U6754 ( .A1(n6287), .A2(n6023), .ZN(n5829) );
  NOR2_X1 U6755 ( .A1(n6271), .A2(n5594), .ZN(n5595) );
  AOI211_X1 U6756 ( .C1(n6266), .C2(n5596), .A(n5829), .B(n5595), .ZN(n5600)
         );
  OR2_X1 U6757 ( .A1(n5598), .A2(n5597), .ZN(n5827) );
  NAND3_X1 U6758 ( .A1(n5827), .A2(n5826), .A3(n4329), .ZN(n5599) );
  OAI211_X1 U6759 ( .C1(n5601), .C2(n6258), .A(n5600), .B(n5599), .ZN(U2967)
         );
  NAND2_X1 U6760 ( .A1(n5674), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5614) );
  INV_X1 U6761 ( .A(n5603), .ZN(n5604) );
  NAND4_X1 U6762 ( .A1(n5602), .A2(n5604), .A3(n5655), .A4(n5864), .ZN(n5612)
         );
  OAI21_X1 U6763 ( .B1(n5610), .B2(n5614), .A(n5612), .ZN(n5605) );
  XNOR2_X1 U6764 ( .A(n5605), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5841)
         );
  NAND2_X1 U6765 ( .A1(n6247), .A2(REIP_REG_18__SCAN_IN), .ZN(n5836) );
  OAI21_X1 U6766 ( .B1(n6271), .B2(n3108), .A(n5836), .ZN(n5607) );
  NOR2_X1 U6767 ( .A1(n6777), .A2(n6258), .ZN(n5606) );
  AOI211_X1 U6768 ( .C1(n6266), .C2(n6075), .A(n5607), .B(n5606), .ZN(n5608)
         );
  OAI21_X1 U6769 ( .B1(n5841), .B2(n6256), .A(n5608), .ZN(U2968) );
  INV_X1 U6770 ( .A(n5610), .ZN(n5615) );
  OR2_X1 U6771 ( .A1(n5674), .A2(n5852), .ZN(n5621) );
  NAND2_X1 U6772 ( .A1(n5610), .A2(n5621), .ZN(n5611) );
  OAI211_X1 U6773 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5674), .A(n5611), .B(n5614), .ZN(n5613) );
  OAI211_X1 U6774 ( .C1(n5615), .C2(n5614), .A(n5613), .B(n5612), .ZN(n5842)
         );
  NAND2_X1 U6775 ( .A1(n5842), .A2(n4329), .ZN(n5619) );
  NOR2_X1 U6776 ( .A1(n6287), .A2(n5616), .ZN(n5845) );
  NOR2_X1 U6777 ( .A1(n6254), .A2(n6086), .ZN(n5617) );
  AOI211_X1 U6778 ( .C1(n6246), .C2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n5845), 
        .B(n5617), .ZN(n5618) );
  OAI211_X1 U6779 ( .C1(n6258), .C2(n6088), .A(n5619), .B(n5618), .ZN(U2969)
         );
  INV_X1 U6780 ( .A(n5620), .ZN(n5622) );
  NAND2_X1 U6781 ( .A1(n5622), .A2(n5621), .ZN(n5623) );
  XNOR2_X1 U6782 ( .A(n5624), .B(n5623), .ZN(n5860) );
  NAND2_X1 U6783 ( .A1(n6247), .A2(REIP_REG_16__SCAN_IN), .ZN(n5854) );
  OAI21_X1 U6784 ( .B1(n6271), .B2(n5625), .A(n5854), .ZN(n5628) );
  NOR2_X1 U6785 ( .A1(n5626), .A2(n6258), .ZN(n5627) );
  AOI211_X1 U6786 ( .C1(n6266), .C2(n5629), .A(n5628), .B(n5627), .ZN(n5630)
         );
  OAI21_X1 U6787 ( .B1(n6256), .B2(n5860), .A(n5630), .ZN(U2970) );
  XNOR2_X1 U6788 ( .A(n5609), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5631)
         );
  XNOR2_X1 U6789 ( .A(n5602), .B(n5631), .ZN(n5867) );
  NAND2_X1 U6790 ( .A1(n5867), .A2(n4329), .ZN(n5635) );
  NOR2_X1 U6791 ( .A1(n6287), .A2(n5294), .ZN(n5861) );
  INV_X1 U6792 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6101) );
  NOR2_X1 U6793 ( .A1(n6271), .A2(n6101), .ZN(n5632) );
  AOI211_X1 U6794 ( .C1(n5633), .C2(n6266), .A(n5861), .B(n5632), .ZN(n5634)
         );
  OAI211_X1 U6795 ( .C1(n6258), .C2(n6096), .A(n5635), .B(n5634), .ZN(U2971)
         );
  XNOR2_X1 U6796 ( .A(n5609), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5645)
         );
  NAND2_X1 U6797 ( .A1(n3004), .A2(n5645), .ZN(n5644) );
  NAND2_X1 U6798 ( .A1(n5644), .A2(n5636), .ZN(n5638) );
  XNOR2_X1 U6799 ( .A(n5674), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5637)
         );
  XNOR2_X1 U6800 ( .A(n5638), .B(n5637), .ZN(n5869) );
  NAND2_X1 U6801 ( .A1(n5869), .A2(n4329), .ZN(n5642) );
  AND2_X1 U6802 ( .A1(n6247), .A2(REIP_REG_14__SCAN_IN), .ZN(n5883) );
  NOR2_X1 U6803 ( .A1(n6254), .A2(n5639), .ZN(n5640) );
  AOI211_X1 U6804 ( .C1(n6246), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5883), 
        .B(n5640), .ZN(n5641) );
  OAI211_X1 U6805 ( .C1(n6258), .C2(n5643), .A(n5642), .B(n5641), .ZN(U2972)
         );
  OAI21_X1 U6806 ( .B1(n3004), .B2(n5645), .A(n5644), .ZN(n6042) );
  NAND2_X1 U6807 ( .A1(n6042), .A2(n4329), .ZN(n5650) );
  OAI22_X1 U6808 ( .A1(n6271), .A2(n5325), .B1(n6287), .B2(n5646), .ZN(n5647)
         );
  AOI21_X1 U6809 ( .B1(n6266), .B2(n5648), .A(n5647), .ZN(n5649) );
  OAI211_X1 U6810 ( .C1(n6258), .C2(n5651), .A(n5650), .B(n5649), .ZN(U2973)
         );
  NAND2_X1 U6811 ( .A1(n5652), .A2(n5663), .ZN(n5891) );
  AND2_X1 U6812 ( .A1(n5655), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5889)
         );
  AOI21_X1 U6813 ( .B1(n5891), .B2(n5887), .A(n5889), .ZN(n5657) );
  INV_X1 U6814 ( .A(n5653), .ZN(n5654) );
  AOI21_X1 U6815 ( .B1(n5655), .B2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5654), 
        .ZN(n5656) );
  XNOR2_X1 U6816 ( .A(n5657), .B(n5656), .ZN(n6281) );
  NAND2_X1 U6817 ( .A1(n6281), .A2(n4329), .ZN(n5661) );
  NOR2_X1 U6818 ( .A1(n6287), .A2(n5338), .ZN(n6274) );
  NOR2_X1 U6819 ( .A1(n6254), .A2(n5658), .ZN(n5659) );
  AOI211_X1 U6820 ( .C1(n6246), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6274), 
        .B(n5659), .ZN(n5660) );
  OAI211_X1 U6821 ( .C1(n6258), .C2(n5662), .A(n5661), .B(n5660), .ZN(U2974)
         );
  INV_X1 U6822 ( .A(n5663), .ZN(n5665) );
  NOR2_X1 U6823 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  XNOR2_X1 U6824 ( .A(n5667), .B(n5666), .ZN(n6291) );
  INV_X1 U6825 ( .A(n6291), .ZN(n5673) );
  AOI22_X1 U6826 ( .A1(n6246), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6247), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5668) );
  OAI21_X1 U6827 ( .B1(n5669), .B2(n6254), .A(n5668), .ZN(n5670) );
  AOI21_X1 U6828 ( .B1(n5671), .B2(n6265), .A(n5670), .ZN(n5672) );
  OAI21_X1 U6829 ( .B1(n5673), .B2(n6256), .A(n5672), .ZN(U2976) );
  XNOR2_X1 U6830 ( .A(n5674), .B(n6307), .ZN(n5675) );
  XNOR2_X1 U6831 ( .A(n5676), .B(n5675), .ZN(n6303) );
  NAND2_X1 U6832 ( .A1(n6303), .A2(n4329), .ZN(n5679) );
  NAND2_X1 U6833 ( .A1(n6247), .A2(REIP_REG_9__SCAN_IN), .ZN(n6298) );
  OAI21_X1 U6834 ( .B1(n6271), .B2(n3111), .A(n6298), .ZN(n5677) );
  AOI21_X1 U6835 ( .B1(n6266), .B2(n6112), .A(n5677), .ZN(n5678) );
  OAI211_X1 U6836 ( .C1(n6258), .C2(n6111), .A(n5679), .B(n5678), .ZN(U2977)
         );
  XNOR2_X1 U6837 ( .A(n5681), .B(n5680), .ZN(n5902) );
  NAND2_X1 U6838 ( .A1(n6246), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5683)
         );
  OR2_X1 U6839 ( .A1(n6287), .A2(n5682), .ZN(n5897) );
  OAI211_X1 U6840 ( .C1(n6254), .C2(n6121), .A(n5683), .B(n5897), .ZN(n5684)
         );
  AOI21_X1 U6841 ( .B1(n6123), .B2(n6265), .A(n5684), .ZN(n5685) );
  OAI21_X1 U6842 ( .B1(n5902), .B2(n6256), .A(n5685), .ZN(U2978) );
  INV_X1 U6843 ( .A(n5687), .ZN(n5713) );
  INV_X1 U6844 ( .A(n5688), .ZN(n5712) );
  NAND2_X1 U6845 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U6846 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6294) );
  NOR2_X1 U6847 ( .A1(n6293), .A2(n6294), .ZN(n5690) );
  NAND2_X1 U6848 ( .A1(n5689), .A2(n5690), .ZN(n5873) );
  NAND2_X1 U6849 ( .A1(n5691), .A2(n5690), .ZN(n5875) );
  INV_X1 U6850 ( .A(n5875), .ZN(n6037) );
  NAND2_X1 U6851 ( .A1(n6037), .A2(n5699), .ZN(n6276) );
  NAND2_X1 U6852 ( .A1(n5873), .A2(n6276), .ZN(n6273) );
  NAND3_X1 U6853 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5880) );
  INV_X1 U6854 ( .A(n5880), .ZN(n5692) );
  NAND2_X1 U6855 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5692), .ZN(n5853) );
  NOR2_X1 U6856 ( .A1(n5693), .A2(n5853), .ZN(n5813) );
  INV_X1 U6857 ( .A(n5813), .ZN(n5843) );
  NOR2_X1 U6858 ( .A1(n5843), .A2(n5848), .ZN(n5694) );
  NAND2_X1 U6859 ( .A1(n6273), .A2(n5694), .ZN(n5835) );
  INV_X1 U6860 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5809) );
  NOR2_X1 U6861 ( .A1(n5835), .A2(n5809), .ZN(n5821) );
  NAND2_X1 U6862 ( .A1(n5821), .A2(n5704), .ZN(n5807) );
  INV_X1 U6863 ( .A(n5790), .ZN(n5695) );
  AND2_X1 U6864 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5753) );
  INV_X1 U6865 ( .A(n5753), .ZN(n5696) );
  NOR2_X1 U6866 ( .A1(n5763), .A2(n5696), .ZN(n5742) );
  NAND2_X1 U6867 ( .A1(n5742), .A2(n5697), .ZN(n5733) );
  AND2_X1 U6868 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5709) );
  INV_X1 U6869 ( .A(n5709), .ZN(n5698) );
  NOR2_X1 U6870 ( .A1(n5733), .A2(n5698), .ZN(n5710) );
  INV_X1 U6871 ( .A(n6286), .ZN(n5820) );
  INV_X1 U6872 ( .A(n5699), .ZN(n5818) );
  NAND2_X1 U6873 ( .A1(n5818), .A2(n6277), .ZN(n5707) );
  INV_X1 U6874 ( .A(n5814), .ZN(n5817) );
  NAND2_X1 U6875 ( .A1(n5873), .A2(n5817), .ZN(n5702) );
  NAND2_X1 U6876 ( .A1(n5700), .A2(n5875), .ZN(n5701) );
  NAND2_X1 U6877 ( .A1(n5702), .A2(n5701), .ZN(n6279) );
  INV_X1 U6878 ( .A(n5703), .ZN(n5705) );
  NAND3_X1 U6879 ( .A1(n5813), .A2(n5705), .A3(n5704), .ZN(n5706) );
  NOR2_X1 U6880 ( .A1(n6279), .A2(n3215), .ZN(n5800) );
  OAI21_X1 U6881 ( .B1(n5709), .B2(n5820), .A(n5727), .ZN(n5717) );
  MUX2_X1 U6882 ( .A(n5710), .B(n5717), .S(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .Z(n5711) );
  AOI211_X2 U6883 ( .C1(n5713), .C2(n6300), .A(n5712), .B(n5711), .ZN(n5714)
         );
  OAI21_X1 U6884 ( .B1(n5715), .B2(n5903), .A(n5714), .ZN(U2987) );
  INV_X1 U6885 ( .A(n5716), .ZN(n5721) );
  NOR2_X1 U6886 ( .A1(n5733), .A2(n5726), .ZN(n5718) );
  MUX2_X1 U6887 ( .A(n5718), .B(n5717), .S(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .Z(n5719) );
  AOI211_X1 U6888 ( .C1(n6300), .C2(n5721), .A(n5720), .B(n5719), .ZN(n5722)
         );
  OAI21_X1 U6889 ( .B1(n5723), .B2(n5903), .A(n5722), .ZN(U2988) );
  NAND2_X1 U6890 ( .A1(n5724), .A2(n6304), .ZN(n5732) );
  INV_X1 U6891 ( .A(n5725), .ZN(n5730) );
  NOR2_X1 U6892 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  AOI211_X1 U6893 ( .C1(n6300), .C2(n5730), .A(n5729), .B(n5728), .ZN(n5731)
         );
  OAI211_X1 U6894 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n5733), .A(n5732), .B(n5731), .ZN(U2989) );
  NOR2_X1 U6895 ( .A1(n5734), .A2(n6288), .ZN(n5735) );
  AOI211_X1 U6896 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5747), .A(n5736), .B(n5735), .ZN(n5740) );
  NAND3_X1 U6897 ( .A1(n5742), .A2(n5738), .A3(n5737), .ZN(n5739) );
  OAI211_X1 U6898 ( .C1(n5741), .C2(n5903), .A(n5740), .B(n5739), .ZN(U2990)
         );
  INV_X1 U6899 ( .A(n5742), .ZN(n5750) );
  NAND2_X1 U6900 ( .A1(n5743), .A2(n6304), .ZN(n5749) );
  NOR2_X1 U6901 ( .A1(n5744), .A2(n6288), .ZN(n5745) );
  AOI211_X1 U6902 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5747), .A(n5746), .B(n5745), .ZN(n5748) );
  OAI211_X1 U6903 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5750), .A(n5749), .B(n5748), .ZN(U2991) );
  INV_X1 U6904 ( .A(n5772), .ZN(n5762) );
  OAI21_X1 U6905 ( .B1(n5752), .B2(n6288), .A(n5751), .ZN(n5756) );
  INV_X1 U6906 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5754) );
  AOI211_X1 U6907 ( .C1(n5754), .C2(n5764), .A(n5753), .B(n5763), .ZN(n5755)
         );
  AOI211_X1 U6908 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5762), .A(n5756), .B(n5755), .ZN(n5757) );
  OAI21_X1 U6909 ( .B1(n5758), .B2(n5903), .A(n5757), .ZN(U2992) );
  NOR2_X1 U6910 ( .A1(n5759), .A2(n6288), .ZN(n5760) );
  AOI211_X1 U6911 ( .C1(n5762), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5761), .B(n5760), .ZN(n5767) );
  INV_X1 U6912 ( .A(n5763), .ZN(n5765) );
  NAND2_X1 U6913 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  OAI211_X1 U6914 ( .C1(n5768), .C2(n5903), .A(n5767), .B(n5766), .ZN(U2993)
         );
  INV_X1 U6915 ( .A(n5769), .ZN(n5777) );
  INV_X1 U6916 ( .A(n5770), .ZN(n5776) );
  INV_X1 U6917 ( .A(n5807), .ZN(n5771) );
  NAND3_X1 U6918 ( .A1(n5771), .A2(n5790), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5773) );
  AOI21_X1 U6919 ( .B1(n5774), .B2(n5773), .A(n5772), .ZN(n5775) );
  AOI211_X1 U6920 ( .C1(n6300), .C2(n5777), .A(n5776), .B(n5775), .ZN(n5778)
         );
  OAI21_X1 U6921 ( .B1(n5779), .B2(n5903), .A(n5778), .ZN(U2994) );
  NAND2_X1 U6922 ( .A1(n5780), .A2(n6304), .ZN(n5786) );
  NOR2_X1 U6923 ( .A1(n5781), .A2(n6288), .ZN(n5782) );
  AOI211_X1 U6924 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5784), .A(n5783), .B(n5782), .ZN(n5785) );
  OAI211_X1 U6925 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5787), .A(n5786), .B(n5785), .ZN(U2995) );
  INV_X1 U6926 ( .A(n5788), .ZN(n5789) );
  OR3_X1 U6927 ( .A1(n5807), .A2(n5790), .A3(n5789), .ZN(n5794) );
  AOI21_X1 U6928 ( .B1(n5792), .B2(n6300), .A(n5791), .ZN(n5793) );
  OAI211_X1 U6929 ( .C1(n5800), .C2(n5795), .A(n5794), .B(n5793), .ZN(n5796)
         );
  INV_X1 U6930 ( .A(n5796), .ZN(n5797) );
  OAI21_X1 U6931 ( .B1(n5798), .B2(n5903), .A(n5797), .ZN(U2996) );
  NAND2_X1 U6932 ( .A1(n5799), .A2(n6304), .ZN(n5806) );
  INV_X1 U6933 ( .A(n5800), .ZN(n5804) );
  NOR2_X1 U6934 ( .A1(n5801), .A2(n6288), .ZN(n5802) );
  AOI211_X1 U6935 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5804), .A(n5803), .B(n5802), .ZN(n5805) );
  OAI211_X1 U6936 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5807), .A(n5806), .B(n5805), .ZN(U2997) );
  INV_X1 U6937 ( .A(n5808), .ZN(n5812) );
  NOR4_X1 U6938 ( .A1(n5835), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5809), 
        .A4(n5833), .ZN(n5810) );
  AOI211_X1 U6939 ( .C1(n5812), .C2(n6300), .A(n5811), .B(n5810), .ZN(n5823)
         );
  AOI21_X1 U6940 ( .B1(n5815), .B2(n5814), .A(n5813), .ZN(n5816) );
  AOI211_X1 U6941 ( .C1(n5848), .C2(n5817), .A(n5816), .B(n6279), .ZN(n5849)
         );
  OAI21_X1 U6942 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5818), .A(n5849), 
        .ZN(n5839) );
  INV_X1 U6943 ( .A(n5839), .ZN(n5819) );
  OAI21_X1 U6944 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5820), .A(n5819), 
        .ZN(n5825) );
  AND2_X1 U6945 ( .A1(n5821), .A2(n5833), .ZN(n5828) );
  OAI21_X1 U6946 ( .B1(n5825), .B2(n5828), .A(INSTADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n5822) );
  OAI211_X1 U6947 ( .C1(n5824), .C2(n5903), .A(n5823), .B(n5822), .ZN(U2998)
         );
  INV_X1 U6948 ( .A(n5825), .ZN(n5834) );
  NAND3_X1 U6949 ( .A1(n5827), .A2(n5826), .A3(n6304), .ZN(n5832) );
  AOI211_X1 U6950 ( .C1(n6300), .C2(n5830), .A(n5829), .B(n5828), .ZN(n5831)
         );
  OAI211_X1 U6951 ( .C1(n5834), .C2(n5833), .A(n5832), .B(n5831), .ZN(U2999)
         );
  NOR2_X1 U6952 ( .A1(n5835), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5838)
         );
  OAI21_X1 U6953 ( .B1(n6079), .B2(n6288), .A(n5836), .ZN(n5837) );
  AOI211_X1 U6954 ( .C1(n5839), .C2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5838), .B(n5837), .ZN(n5840) );
  OAI21_X1 U6955 ( .B1(n5841), .B2(n5903), .A(n5840), .ZN(U3000) );
  NAND2_X1 U6956 ( .A1(n5842), .A2(n6304), .ZN(n5847) );
  INV_X1 U6957 ( .A(n6273), .ZN(n5894) );
  NOR3_X1 U6958 ( .A1(n5894), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5843), 
        .ZN(n5844) );
  AOI211_X1 U6959 ( .C1(n6300), .C2(n6089), .A(n5845), .B(n5844), .ZN(n5846)
         );
  OAI211_X1 U6960 ( .C1(n5849), .C2(n5848), .A(n5847), .B(n5846), .ZN(U3001)
         );
  AND2_X1 U6961 ( .A1(n6286), .A2(n5853), .ZN(n5850) );
  NOR2_X1 U6962 ( .A1(n6279), .A2(n5850), .ZN(n5865) );
  NOR2_X1 U6963 ( .A1(n5853), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5851)
         );
  NAND2_X1 U6964 ( .A1(n6273), .A2(n5851), .ZN(n5862) );
  AOI21_X1 U6965 ( .B1(n5865), .B2(n5862), .A(n5852), .ZN(n5858) );
  NOR4_X1 U6966 ( .A1(n5894), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5864), 
        .A4(n5853), .ZN(n5857) );
  OAI21_X1 U6967 ( .B1(n5855), .B2(n6288), .A(n5854), .ZN(n5856) );
  NOR3_X1 U6968 ( .A1(n5858), .A2(n5857), .A3(n5856), .ZN(n5859) );
  OAI21_X1 U6969 ( .B1(n5860), .B2(n5903), .A(n5859), .ZN(U3002) );
  AOI21_X1 U6970 ( .B1(n6099), .B2(n6300), .A(n5861), .ZN(n5863) );
  OAI211_X1 U6971 ( .C1(n5865), .C2(n5864), .A(n5863), .B(n5862), .ZN(n5866)
         );
  AOI21_X1 U6972 ( .B1(n5867), .B2(n6304), .A(n5866), .ZN(n5868) );
  INV_X1 U6973 ( .A(n5868), .ZN(U3003) );
  INV_X1 U6974 ( .A(n5869), .ZN(n5886) );
  AOI21_X1 U6975 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5870), .ZN(n5871) );
  AOI211_X1 U6976 ( .C1(n5872), .C2(n5880), .A(n5871), .B(n6279), .ZN(n6046)
         );
  OAI21_X1 U6977 ( .B1(n5875), .B2(n5874), .A(n5873), .ZN(n5877) );
  NAND2_X1 U6978 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5876) );
  NOR2_X1 U6979 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5876), .ZN(n6036)
         );
  NAND2_X1 U6980 ( .A1(n5877), .A2(n6036), .ZN(n6044) );
  AOI21_X1 U6981 ( .B1(n6046), .B2(n6044), .A(n5878), .ZN(n5884) );
  NOR2_X1 U6982 ( .A1(n5879), .A2(n6288), .ZN(n5882) );
  NOR3_X1 U6983 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5894), .A3(n5880), 
        .ZN(n5881) );
  NOR4_X1 U6984 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n5885)
         );
  OAI21_X1 U6985 ( .B1(n5886), .B2(n5903), .A(n5885), .ZN(U3004) );
  INV_X1 U6986 ( .A(n5887), .ZN(n5888) );
  NOR2_X1 U6987 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  XNOR2_X1 U6988 ( .A(n5891), .B(n5890), .ZN(n6253) );
  AOI22_X1 U6989 ( .A1(n5892), .A2(n6300), .B1(n6247), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5893) );
  OAI21_X1 U6990 ( .B1(n5894), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5893), 
        .ZN(n5895) );
  AOI21_X1 U6991 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6279), .A(n5895), 
        .ZN(n5896) );
  OAI21_X1 U6992 ( .B1(n6253), .B2(n5903), .A(n5896), .ZN(U3007) );
  OAI21_X1 U6993 ( .B1(n6118), .B2(n6288), .A(n5897), .ZN(n5900) );
  OAI21_X1 U6994 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6293), .ZN(n5898) );
  NOR2_X1 U6995 ( .A1(n6292), .A2(n5898), .ZN(n5899) );
  AOI211_X1 U6996 ( .C1(n6285), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5900), 
        .B(n5899), .ZN(n5901) );
  OAI21_X1 U6997 ( .B1(n5903), .B2(n5902), .A(n5901), .ZN(U3010) );
  INV_X1 U6998 ( .A(n5904), .ZN(n5909) );
  AOI21_X1 U6999 ( .B1(n6039), .B2(n5906), .A(n5905), .ZN(n5907) );
  AOI211_X1 U7000 ( .C1(n6300), .C2(n5909), .A(n5908), .B(n5907), .ZN(n5914)
         );
  NAND3_X1 U7001 ( .A1(n6304), .A2(n5911), .A3(n5910), .ZN(n5912) );
  NAND3_X1 U7002 ( .A1(n5914), .A2(n5913), .A3(n5912), .ZN(U3018) );
  OAI211_X1 U7003 ( .C1(n5915), .C2(STATEBS16_REG_SCAN_IN), .A(n6419), .B(
        n6420), .ZN(n5916) );
  OAI21_X1 U7004 ( .B1(n5917), .B2(n6591), .A(n5916), .ZN(n5918) );
  MUX2_X1 U7005 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5918), .S(n6599), 
        .Z(U3464) );
  XNOR2_X1 U7006 ( .A(n5920), .B(n5919), .ZN(n5921) );
  OAI22_X1 U7007 ( .A1(n5921), .A2(n6476), .B1(n4437), .B2(n6591), .ZN(n5922)
         );
  MUX2_X1 U7008 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5922), .S(n6599), 
        .Z(U3463) );
  INV_X1 U7009 ( .A(n5923), .ZN(n5924) );
  OAI22_X1 U7010 ( .A1(n5926), .A2(n5925), .B1(n5924), .B2(n6567), .ZN(n5927)
         );
  MUX2_X1 U7011 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5927), .S(n6054), 
        .Z(U3456) );
  INV_X1 U7012 ( .A(n6353), .ZN(n5928) );
  NOR2_X1 U7013 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5928), .ZN(n6340)
         );
  OAI21_X1 U7014 ( .B1(n6380), .B2(n6341), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5930) );
  NAND3_X1 U7015 ( .A1(n6347), .A2(n6419), .A3(n5930), .ZN(n5931) );
  OAI21_X1 U7016 ( .B1(n6340), .B2(n6588), .A(n5931), .ZN(n5932) );
  NOR4_X2 U7017 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5934), .A3(n5933), 
        .A4(n5932), .ZN(n6344) );
  INV_X1 U7018 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5940) );
  NOR2_X1 U7019 ( .A1(n6471), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5935)
         );
  AOI22_X1 U7020 ( .A1(n5936), .A2(n6592), .B1(n6389), .B2(n5935), .ZN(n6338)
         );
  OAI22_X1 U7021 ( .A1(n5961), .A2(n6496), .B1(n6338), .B2(n6363), .ZN(n5937)
         );
  AOI21_X1 U7022 ( .B1(n6493), .B2(n6380), .A(n5937), .ZN(n5939) );
  NAND2_X1 U7023 ( .A1(n6492), .A2(n6340), .ZN(n5938) );
  OAI211_X1 U7024 ( .C1(n6344), .C2(n5940), .A(n5939), .B(n5938), .ZN(U3069)
         );
  INV_X1 U7025 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5944) );
  OAI22_X1 U7026 ( .A1(n5961), .A2(n6502), .B1(n6338), .B2(n6366), .ZN(n5941)
         );
  AOI21_X1 U7027 ( .B1(n6380), .B2(n6499), .A(n5941), .ZN(n5943) );
  NAND2_X1 U7028 ( .A1(n6498), .A2(n6340), .ZN(n5942) );
  OAI211_X1 U7029 ( .C1(n6344), .C2(n5944), .A(n5943), .B(n5942), .ZN(U3070)
         );
  INV_X1 U7030 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5948) );
  OAI22_X1 U7031 ( .A1(n5961), .A2(n6508), .B1(n6338), .B2(n6369), .ZN(n5945)
         );
  AOI21_X1 U7032 ( .B1(n6380), .B2(n6505), .A(n5945), .ZN(n5947) );
  NAND2_X1 U7033 ( .A1(n6782), .A2(n6340), .ZN(n5946) );
  OAI211_X1 U7034 ( .C1(n6344), .C2(n5948), .A(n5947), .B(n5946), .ZN(U3071)
         );
  OAI22_X1 U7035 ( .A1(n5961), .A2(n6514), .B1(n6338), .B2(n6372), .ZN(n5949)
         );
  AOI21_X1 U7036 ( .B1(n6380), .B2(n6511), .A(n5949), .ZN(n5951) );
  NAND2_X1 U7037 ( .A1(n6510), .A2(n6340), .ZN(n5950) );
  OAI211_X1 U7038 ( .C1(n6344), .C2(n5952), .A(n5951), .B(n5950), .ZN(U3072)
         );
  INV_X1 U7039 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5956) );
  OAI22_X1 U7040 ( .A1(n5961), .A2(n6520), .B1(n6338), .B2(n6375), .ZN(n5953)
         );
  AOI21_X1 U7041 ( .B1(n6380), .B2(n6517), .A(n5953), .ZN(n5955) );
  NAND2_X1 U7042 ( .A1(n6516), .A2(n6340), .ZN(n5954) );
  OAI211_X1 U7043 ( .C1(n6344), .C2(n5956), .A(n5955), .B(n5954), .ZN(U3073)
         );
  OAI22_X1 U7044 ( .A1(n5961), .A2(n6526), .B1(n6338), .B2(n6378), .ZN(n5958)
         );
  INV_X1 U7045 ( .A(n6380), .ZN(n5962) );
  NOR2_X1 U7046 ( .A1(n5962), .A2(n6461), .ZN(n5957) );
  AOI211_X1 U7047 ( .C1(n6522), .C2(n6340), .A(n5958), .B(n5957), .ZN(n5959)
         );
  OAI21_X1 U7048 ( .B1(n6344), .B2(n5960), .A(n5959), .ZN(U3074) );
  INV_X1 U7049 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5966) );
  OAI22_X1 U7050 ( .A1(n5961), .A2(n6537), .B1(n6338), .B2(n6384), .ZN(n5964)
         );
  NOR2_X1 U7051 ( .A1(n5962), .A2(n6469), .ZN(n5963) );
  AOI211_X1 U7052 ( .C1(n6530), .C2(n6340), .A(n5964), .B(n5963), .ZN(n5965)
         );
  OAI21_X1 U7053 ( .B1(n6344), .B2(n5966), .A(n5965), .ZN(U3075) );
  INV_X1 U7054 ( .A(n6007), .ZN(n5968) );
  AOI21_X1 U7055 ( .B1(n6009), .B2(n5968), .A(n6059), .ZN(n5969) );
  NOR2_X1 U7056 ( .A1(n5969), .A2(n6476), .ZN(n5974) );
  NOR2_X1 U7057 ( .A1(n6484), .A2(n6598), .ZN(n5971) );
  AOI22_X1 U7058 ( .A1(n5974), .A2(n6422), .B1(n6389), .B2(n5971), .ZN(n6013)
         );
  NAND2_X1 U7059 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5972), .ZN(n6432) );
  NOR2_X1 U7060 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6432), .ZN(n6011)
         );
  INV_X1 U7061 ( .A(n6011), .ZN(n5975) );
  INV_X1 U7062 ( .A(n6422), .ZN(n5973) );
  AOI22_X1 U7063 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5975), .B1(n5974), .B2(
        n5973), .ZN(n5976) );
  OAI211_X1 U7064 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n5978), .A(n5977), .B(n5976), .ZN(n6006) );
  AOI22_X1 U7065 ( .A1(n6007), .A2(n6435), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n6006), .ZN(n5979) );
  OAI21_X1 U7066 ( .B1(n6009), .B2(n5980), .A(n5979), .ZN(n5981) );
  AOI21_X1 U7067 ( .B1(n6475), .B2(n6011), .A(n5981), .ZN(n5982) );
  OAI21_X1 U7068 ( .B1(n6013), .B2(n6360), .A(n5982), .ZN(U3100) );
  AOI22_X1 U7069 ( .A1(n6007), .A2(n6438), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n6006), .ZN(n5983) );
  OAI21_X1 U7070 ( .B1(n6009), .B2(n5984), .A(n5983), .ZN(n5985) );
  AOI21_X1 U7071 ( .B1(n6492), .B2(n6011), .A(n5985), .ZN(n5986) );
  OAI21_X1 U7072 ( .B1(n6013), .B2(n6363), .A(n5986), .ZN(U3101) );
  AOI22_X1 U7073 ( .A1(n6007), .A2(n6442), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n6006), .ZN(n5987) );
  OAI21_X1 U7074 ( .B1(n6009), .B2(n5988), .A(n5987), .ZN(n5989) );
  AOI21_X1 U7075 ( .B1(n6498), .B2(n6011), .A(n5989), .ZN(n5990) );
  OAI21_X1 U7076 ( .B1(n6013), .B2(n6366), .A(n5990), .ZN(U3102) );
  AOI22_X1 U7077 ( .A1(n6007), .A2(n6446), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n6006), .ZN(n5991) );
  OAI21_X1 U7078 ( .B1(n6009), .B2(n5992), .A(n5991), .ZN(n5993) );
  AOI21_X1 U7079 ( .B1(n6782), .B2(n6011), .A(n5993), .ZN(n5994) );
  OAI21_X1 U7080 ( .B1(n6013), .B2(n6369), .A(n5994), .ZN(U3103) );
  AOI22_X1 U7081 ( .A1(n6007), .A2(n6450), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n6006), .ZN(n5995) );
  OAI21_X1 U7082 ( .B1(n6009), .B2(n5996), .A(n5995), .ZN(n5997) );
  AOI21_X1 U7083 ( .B1(n6510), .B2(n6011), .A(n5997), .ZN(n5998) );
  OAI21_X1 U7084 ( .B1(n6013), .B2(n6372), .A(n5998), .ZN(U3104) );
  AOI22_X1 U7085 ( .A1(n6007), .A2(n6454), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n6006), .ZN(n5999) );
  OAI21_X1 U7086 ( .B1(n6009), .B2(n6000), .A(n5999), .ZN(n6001) );
  AOI21_X1 U7087 ( .B1(n6516), .B2(n6011), .A(n6001), .ZN(n6002) );
  OAI21_X1 U7088 ( .B1(n6013), .B2(n6375), .A(n6002), .ZN(U3105) );
  AOI22_X1 U7089 ( .A1(n6007), .A2(n6457), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n6006), .ZN(n6003) );
  OAI21_X1 U7090 ( .B1(n6009), .B2(n6461), .A(n6003), .ZN(n6004) );
  AOI21_X1 U7091 ( .B1(n6522), .B2(n6011), .A(n6004), .ZN(n6005) );
  OAI21_X1 U7092 ( .B1(n6013), .B2(n6378), .A(n6005), .ZN(U3106) );
  AOI22_X1 U7093 ( .A1(n6007), .A2(n6463), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n6006), .ZN(n6008) );
  OAI21_X1 U7094 ( .B1(n6009), .B2(n6469), .A(n6008), .ZN(n6010) );
  AOI21_X1 U7095 ( .B1(n6530), .B2(n6011), .A(n6010), .ZN(n6012) );
  OAI21_X1 U7096 ( .B1(n6013), .B2(n6384), .A(n6012), .ZN(U3107) );
  NOR2_X1 U7097 ( .A1(n6014), .A2(n6760), .ZN(n6016) );
  OAI21_X1 U7098 ( .B1(n6017), .B2(n6016), .A(n6015), .ZN(n6020) );
  NAND3_X1 U7099 ( .A1(n6020), .A2(n6019), .A3(n6018), .ZN(U3182) );
  MUX2_X1 U7100 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6021), .Z(U3448) );
  MUX2_X1 U7101 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6021), .Z(U3447) );
  MUX2_X1 U7102 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6021), .Z(U3446) );
  MUX2_X1 U7103 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6021), .Z(U3445) );
  AND2_X1 U7104 ( .A1(n6222), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7105 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6031) );
  OAI22_X1 U7106 ( .A1(n6093), .A2(n6023), .B1(n6022), .B2(n6155), .ZN(n6024)
         );
  AOI211_X1 U7107 ( .C1(n6142), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6167), 
        .B(n6024), .ZN(n6030) );
  OAI21_X1 U7108 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n6025), .ZN(n6027) );
  OAI22_X1 U7109 ( .A1(n6084), .A2(n6027), .B1(n6026), .B2(n6172), .ZN(n6028)
         );
  AOI21_X1 U7110 ( .B1(n6032), .B2(n6152), .A(n6028), .ZN(n6029) );
  OAI211_X1 U7111 ( .C1(n6031), .C2(n6179), .A(n6030), .B(n6029), .ZN(U2808)
         );
  AOI22_X1 U7112 ( .A1(n6032), .A2(n6197), .B1(n3031), .B2(DATAI_19_), .ZN(
        n6034) );
  AOI22_X1 U7113 ( .A1(n6774), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6779), .ZN(n6033) );
  NAND2_X1 U7114 ( .A1(n6034), .A2(n6033), .ZN(U2872) );
  NOR2_X1 U7115 ( .A1(n6035), .A2(n6288), .ZN(n6041) );
  NAND2_X1 U7116 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  OAI22_X1 U7117 ( .A1(n6039), .A2(n6038), .B1(n5646), .B2(n6287), .ZN(n6040)
         );
  AOI211_X1 U7118 ( .C1(n6042), .C2(n6304), .A(n6041), .B(n6040), .ZN(n6043)
         );
  OAI211_X1 U7119 ( .C1(n6046), .C2(n6045), .A(n6044), .B(n6043), .ZN(U3005)
         );
  INV_X1 U7120 ( .A(n6047), .ZN(n6051) );
  INV_X1 U7121 ( .A(n6048), .ZN(n6050) );
  NAND4_X1 U7122 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6176), .ZN(n6052)
         );
  OAI21_X1 U7123 ( .B1(n6054), .B2(n6053), .A(n6052), .ZN(U3455) );
  OAI21_X1 U7124 ( .B1(n6055), .B2(n6573), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6056) );
  OAI21_X1 U7125 ( .B1(n6057), .B2(n6566), .A(n6056), .ZN(U2790) );
  INV_X1 U7126 ( .A(n6582), .ZN(n6585) );
  OAI21_X1 U7127 ( .B1(BS16_N), .B2(n6058), .A(n6585), .ZN(n6583) );
  OAI21_X1 U7128 ( .B1(n6585), .B2(n6059), .A(n6583), .ZN(U2792) );
  OAI21_X1 U7129 ( .B1(n6061), .B2(n6060), .A(n6256), .ZN(U2793) );
  NOR4_X1 U7130 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6065) );
  NOR4_X1 U7131 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6064) );
  NOR4_X1 U7132 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6063) );
  NOR4_X1 U7133 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6062) );
  NAND4_X1 U7134 ( .A1(n6065), .A2(n6064), .A3(n6063), .A4(n6062), .ZN(n6071)
         );
  NOR4_X1 U7135 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6069) );
  AOI211_X1 U7136 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_7__SCAN_IN), .B(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n6068) );
  NOR4_X1 U7137 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n6067) );
  NOR4_X1 U7138 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n6066) );
  NAND4_X1 U7139 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n6070)
         );
  NOR2_X1 U7140 ( .A1(n6071), .A2(n6070), .ZN(n6608) );
  INV_X1 U7141 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6665) );
  NOR3_X1 U7142 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6073) );
  OAI21_X1 U7143 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6073), .A(n6608), .ZN(n6072)
         );
  OAI21_X1 U7144 ( .B1(n6608), .B2(n6665), .A(n6072), .ZN(U2794) );
  INV_X1 U7145 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6758) );
  NOR2_X1 U7146 ( .A1(REIP_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n6602) );
  OAI21_X1 U7147 ( .B1(n6073), .B2(n6602), .A(n6608), .ZN(n6074) );
  OAI21_X1 U7148 ( .B1(n6608), .B2(n6758), .A(n6074), .ZN(U2795) );
  AOI22_X1 U7149 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6143), .B1(n6075), .B2(n6174), .ZN(n6076) );
  OAI21_X1 U7150 ( .B1(n6093), .B2(n6077), .A(n6076), .ZN(n6078) );
  AOI211_X1 U7151 ( .C1(n6142), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6167), 
        .B(n6078), .ZN(n6083) );
  INV_X1 U7152 ( .A(n6777), .ZN(n6081) );
  INV_X1 U7153 ( .A(n6079), .ZN(n6080) );
  AOI22_X1 U7154 ( .A1(n6081), .A2(n6152), .B1(n6161), .B2(n6080), .ZN(n6082)
         );
  OAI211_X1 U7155 ( .C1(REIP_REG_18__SCAN_IN), .C2(n6084), .A(n6083), .B(n6082), .ZN(U2809) );
  AOI21_X1 U7156 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6085), .A(
        REIP_REG_17__SCAN_IN), .ZN(n6092) );
  OAI22_X1 U7157 ( .A1(n3725), .A2(n6186), .B1(n6086), .B2(n6155), .ZN(n6087)
         );
  AOI211_X1 U7158 ( .C1(n6143), .C2(EBX_REG_17__SCAN_IN), .A(n6167), .B(n6087), 
        .ZN(n6091) );
  INV_X1 U7159 ( .A(n6088), .ZN(n6198) );
  AOI22_X1 U7160 ( .A1(n6198), .A2(n6152), .B1(n6161), .B2(n6089), .ZN(n6090)
         );
  OAI211_X1 U7161 ( .C1(n6093), .C2(n6092), .A(n6091), .B(n6090), .ZN(U2810)
         );
  OAI22_X1 U7162 ( .A1(n6096), .A2(n6095), .B1(n6155), .B2(n6094), .ZN(n6097)
         );
  INV_X1 U7163 ( .A(n6097), .ZN(n6105) );
  AOI22_X1 U7164 ( .A1(n6161), .A2(n6099), .B1(REIP_REG_15__SCAN_IN), .B2(
        n6098), .ZN(n6100) );
  OAI211_X1 U7165 ( .C1(n6186), .C2(n6101), .A(n6100), .B(n6144), .ZN(n6102)
         );
  AOI211_X1 U7166 ( .C1(n6143), .C2(EBX_REG_15__SCAN_IN), .A(n6103), .B(n6102), 
        .ZN(n6104) );
  NAND2_X1 U7167 ( .A1(n6105), .A2(n6104), .ZN(U2812) );
  AOI21_X1 U7168 ( .B1(n6107), .B2(n6106), .A(n3043), .ZN(n6301) );
  INV_X1 U7169 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6190) );
  AOI22_X1 U7170 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6142), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6117), .ZN(n6108) );
  OAI211_X1 U7171 ( .C1(n6179), .C2(n6190), .A(n6108), .B(n6144), .ZN(n6109)
         );
  AOI211_X1 U7172 ( .C1(n6301), .C2(n6161), .A(n6110), .B(n6109), .ZN(n6114)
         );
  INV_X1 U7173 ( .A(n6111), .ZN(n6188) );
  AOI22_X1 U7174 ( .A1(n6188), .A2(n6152), .B1(n6174), .B2(n6112), .ZN(n6113)
         );
  NAND2_X1 U7175 ( .A1(n6114), .A2(n6113), .ZN(U2818) );
  AND2_X1 U7176 ( .A1(n6116), .A2(n6115), .ZN(n6133) );
  AOI21_X1 U7177 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6133), .A(
        REIP_REG_8__SCAN_IN), .ZN(n6127) );
  INV_X1 U7178 ( .A(n6117), .ZN(n6126) );
  OAI22_X1 U7179 ( .A1(n6119), .A2(n6179), .B1(n6172), .B2(n6118), .ZN(n6120)
         );
  AOI211_X1 U7180 ( .C1(n6142), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6167), 
        .B(n6120), .ZN(n6125) );
  INV_X1 U7181 ( .A(n6121), .ZN(n6122) );
  AOI22_X1 U7182 ( .A1(n6123), .A2(n6152), .B1(n6122), .B2(n6174), .ZN(n6124)
         );
  OAI211_X1 U7183 ( .C1(n6127), .C2(n6126), .A(n6125), .B(n6124), .ZN(U2819)
         );
  OAI21_X1 U7184 ( .B1(n6186), .B2(n6263), .A(n6144), .ZN(n6131) );
  OAI22_X1 U7185 ( .A1(n6129), .A2(n6179), .B1(n6172), .B2(n6128), .ZN(n6130)
         );
  AOI211_X1 U7186 ( .C1(n6133), .C2(n6132), .A(n6131), .B(n6130), .ZN(n6139)
         );
  INV_X1 U7187 ( .A(n6259), .ZN(n6137) );
  OAI21_X1 U7188 ( .B1(n6135), .B2(n6140), .A(n6134), .ZN(n6165) );
  OAI21_X1 U7189 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6159), .A(n6165), .ZN(n6136)
         );
  AOI22_X1 U7190 ( .A1(n6137), .A2(n6152), .B1(REIP_REG_7__SCAN_IN), .B2(n6136), .ZN(n6138) );
  OAI211_X1 U7191 ( .C1(n6255), .C2(n6155), .A(n6139), .B(n6138), .ZN(U2820)
         );
  INV_X1 U7192 ( .A(n6140), .ZN(n6141) );
  NAND2_X1 U7193 ( .A1(n6141), .A2(n6150), .ZN(n6146) );
  AOI22_X1 U7194 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6143), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6142), .ZN(n6145) );
  OAI211_X1 U7195 ( .C1(n6159), .C2(n6146), .A(n6145), .B(n6144), .ZN(n6147)
         );
  AOI21_X1 U7196 ( .B1(n6161), .B2(n6148), .A(n6147), .ZN(n6149) );
  OAI21_X1 U7197 ( .B1(n6150), .B2(n6165), .A(n6149), .ZN(n6151) );
  AOI21_X1 U7198 ( .B1(n6153), .B2(n6152), .A(n6151), .ZN(n6154) );
  OAI21_X1 U7199 ( .B1(n6156), .B2(n6155), .A(n6154), .ZN(U2821) );
  INV_X1 U7200 ( .A(n6157), .ZN(n6158) );
  NOR2_X1 U7201 ( .A1(n6159), .A2(n6158), .ZN(n6169) );
  AOI21_X1 U7202 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6169), .A(
        REIP_REG_5__SCAN_IN), .ZN(n6166) );
  INV_X1 U7203 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6196) );
  OAI22_X1 U7204 ( .A1(n6196), .A2(n6179), .B1(n6272), .B2(n6186), .ZN(n6160)
         );
  AOI211_X1 U7205 ( .C1(n6161), .C2(n6191), .A(n6167), .B(n6160), .ZN(n6164)
         );
  INV_X1 U7206 ( .A(n6162), .ZN(n6267) );
  AOI22_X1 U7207 ( .A1(n6264), .A2(n6182), .B1(n6267), .B2(n6174), .ZN(n6163)
         );
  OAI211_X1 U7208 ( .C1(n6166), .C2(n6165), .A(n6164), .B(n6163), .ZN(U2822)
         );
  INV_X1 U7209 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6187) );
  AOI221_X1 U7210 ( .B1(n6170), .B2(REIP_REG_4__SCAN_IN), .C1(n6169), .C2(
        n6168), .A(n6167), .ZN(n6185) );
  NOR2_X1 U7211 ( .A1(n6172), .A2(n6171), .ZN(n6181) );
  INV_X1 U7212 ( .A(n6173), .ZN(n6175) );
  AOI22_X1 U7213 ( .A1(n6177), .A2(n6176), .B1(n6175), .B2(n6174), .ZN(n6178)
         );
  OAI21_X1 U7214 ( .B1(n6179), .B2(n6737), .A(n6178), .ZN(n6180) );
  AOI211_X1 U7215 ( .C1(n6183), .C2(n6182), .A(n6181), .B(n6180), .ZN(n6184)
         );
  OAI211_X1 U7216 ( .C1(n6187), .C2(n6186), .A(n6185), .B(n6184), .ZN(U2823)
         );
  AOI22_X1 U7217 ( .A1(n6188), .A2(n6193), .B1(n6192), .B2(n6301), .ZN(n6189)
         );
  OAI21_X1 U7218 ( .B1(n6190), .B2(n6195), .A(n6189), .ZN(U2850) );
  AOI22_X1 U7219 ( .A1(n6264), .A2(n6193), .B1(n6192), .B2(n6191), .ZN(n6194)
         );
  OAI21_X1 U7220 ( .B1(n6196), .B2(n6195), .A(n6194), .ZN(U2854) );
  AOI22_X1 U7221 ( .A1(n6198), .A2(n6197), .B1(n3031), .B2(DATAI_17_), .ZN(
        n6200) );
  AOI22_X1 U7222 ( .A1(n6774), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6779), .ZN(n6199) );
  NAND2_X1 U7223 ( .A1(n6200), .A2(n6199), .ZN(U2874) );
  AOI22_X1 U7224 ( .A1(n6222), .A2(DATAO_REG_28__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n3090), .ZN(n6202) );
  OAI21_X1 U7225 ( .B1(n6643), .B2(n6214), .A(n6202), .ZN(U2895) );
  AOI22_X1 U7226 ( .A1(n6612), .A2(LWORD_REG_15__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6203) );
  OAI21_X1 U7227 ( .B1(n6204), .B2(n6233), .A(n6203), .ZN(U2908) );
  INV_X1 U7228 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6206) );
  AOI22_X1 U7229 ( .A1(n6612), .A2(LWORD_REG_14__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6205) );
  OAI21_X1 U7230 ( .B1(n6206), .B2(n6233), .A(n6205), .ZN(U2909) );
  AOI22_X1 U7231 ( .A1(n6612), .A2(LWORD_REG_13__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6207) );
  OAI21_X1 U7232 ( .B1(n6208), .B2(n6233), .A(n6207), .ZN(U2910) );
  INV_X1 U7233 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6210) );
  AOI22_X1 U7234 ( .A1(n6612), .A2(LWORD_REG_12__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6209) );
  OAI21_X1 U7235 ( .B1(n6210), .B2(n6233), .A(n6209), .ZN(U2911) );
  AOI22_X1 U7236 ( .A1(n6612), .A2(LWORD_REG_11__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6211) );
  OAI21_X1 U7237 ( .B1(n6679), .B2(n6233), .A(n6211), .ZN(U2912) );
  INV_X1 U7238 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7239 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6212), .B1(n6222), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6213) );
  OAI21_X1 U7240 ( .B1(n6721), .B2(n6214), .A(n6213), .ZN(U2913) );
  INV_X1 U7241 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6216) );
  AOI22_X1 U7242 ( .A1(n6612), .A2(LWORD_REG_9__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6215) );
  OAI21_X1 U7243 ( .B1(n6216), .B2(n6233), .A(n6215), .ZN(U2914) );
  INV_X1 U7244 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6218) );
  AOI22_X1 U7245 ( .A1(n6612), .A2(LWORD_REG_8__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6217) );
  OAI21_X1 U7246 ( .B1(n6218), .B2(n6233), .A(n6217), .ZN(U2915) );
  AOI22_X1 U7247 ( .A1(n6612), .A2(LWORD_REG_7__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6219) );
  OAI21_X1 U7248 ( .B1(n3571), .B2(n6233), .A(n6219), .ZN(U2916) );
  AOI22_X1 U7249 ( .A1(n6612), .A2(LWORD_REG_6__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6220) );
  OAI21_X1 U7250 ( .B1(n3545), .B2(n6233), .A(n6220), .ZN(U2917) );
  AOI22_X1 U7251 ( .A1(n6612), .A2(LWORD_REG_5__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6221) );
  OAI21_X1 U7252 ( .B1(n3526), .B2(n6233), .A(n6221), .ZN(U2918) );
  AOI22_X1 U7253 ( .A1(n6612), .A2(LWORD_REG_4__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6223) );
  OAI21_X1 U7254 ( .B1(n6224), .B2(n6233), .A(n6223), .ZN(U2919) );
  AOI22_X1 U7255 ( .A1(n6612), .A2(LWORD_REG_3__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6225) );
  OAI21_X1 U7256 ( .B1(n6226), .B2(n6233), .A(n6225), .ZN(U2920) );
  AOI22_X1 U7257 ( .A1(n6612), .A2(LWORD_REG_2__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6227) );
  OAI21_X1 U7258 ( .B1(n6228), .B2(n6233), .A(n6227), .ZN(U2921) );
  AOI22_X1 U7259 ( .A1(DATAO_REG_1__SCAN_IN), .A2(n6222), .B1(n6229), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n6230) );
  OAI21_X1 U7260 ( .B1(n6231), .B2(n6233), .A(n6230), .ZN(U2922) );
  AOI22_X1 U7261 ( .A1(n6612), .A2(LWORD_REG_0__SCAN_IN), .B1(n6222), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6232) );
  OAI21_X1 U7262 ( .B1(n6234), .B2(n6233), .A(n6232), .ZN(U2923) );
  AOI22_X1 U7263 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6242), .B1(n6241), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7264 ( .A1(n6243), .A2(DATAI_8_), .ZN(n6235) );
  NAND2_X1 U7265 ( .A1(n6236), .A2(n6235), .ZN(U2947) );
  AOI22_X1 U7266 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6242), .B1(n6241), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7267 ( .A1(n6243), .A2(DATAI_9_), .ZN(n6237) );
  NAND2_X1 U7268 ( .A1(n6238), .A2(n6237), .ZN(U2948) );
  AOI22_X1 U7269 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6242), .B1(n6241), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7270 ( .A1(n6243), .A2(DATAI_12_), .ZN(n6239) );
  NAND2_X1 U7271 ( .A1(n6240), .A2(n6239), .ZN(U2951) );
  AOI22_X1 U7272 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6242), .B1(n6241), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7273 ( .A1(n6243), .A2(DATAI_14_), .ZN(n6244) );
  NAND2_X1 U7274 ( .A1(n6245), .A2(n6244), .ZN(U2953) );
  AOI22_X1 U7275 ( .A1(n6247), .A2(REIP_REG_11__SCAN_IN), .B1(n6246), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6252) );
  INV_X1 U7276 ( .A(n6248), .ZN(n6250) );
  AOI22_X1 U7277 ( .A1(n6250), .A2(n6265), .B1(n6266), .B2(n6249), .ZN(n6251)
         );
  OAI211_X1 U7278 ( .C1(n6253), .C2(n6256), .A(n6252), .B(n6251), .ZN(U2975)
         );
  OAI222_X1 U7279 ( .A1(n6259), .A2(n6258), .B1(n6257), .B2(n6256), .C1(n6255), 
        .C2(n6254), .ZN(n6260) );
  INV_X1 U7280 ( .A(n6260), .ZN(n6262) );
  OAI211_X1 U7281 ( .C1(n6263), .C2(n6271), .A(n6262), .B(n6261), .ZN(U2979)
         );
  AOI222_X1 U7282 ( .A1(n6268), .A2(n4329), .B1(n6267), .B2(n6266), .C1(n6265), 
        .C2(n6264), .ZN(n6270) );
  OAI211_X1 U7283 ( .C1(n6272), .C2(n6271), .A(n6270), .B(n6269), .ZN(U2981)
         );
  NAND2_X1 U7284 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6273), .ZN(n6284) );
  AOI21_X1 U7285 ( .B1(n6275), .B2(n6300), .A(n6274), .ZN(n6283) );
  AOI21_X1 U7286 ( .B1(n6277), .B2(n6276), .A(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n6278) );
  OR2_X1 U7287 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  AOI22_X1 U7288 ( .A1(n6281), .A2(n6304), .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6280), .ZN(n6282) );
  OAI211_X1 U7289 ( .C1(INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n6284), .A(n6283), .B(n6282), .ZN(U3006) );
  AOI21_X1 U7290 ( .B1(n6293), .B2(n6286), .A(n6285), .ZN(n6308) );
  OAI22_X1 U7291 ( .A1(n6289), .A2(n6288), .B1(n4392), .B2(n6287), .ZN(n6290)
         );
  AOI21_X1 U7292 ( .B1(n6291), .B2(n6304), .A(n6290), .ZN(n6296) );
  NOR2_X1 U7293 ( .A1(n6293), .A2(n6292), .ZN(n6302) );
  OAI211_X1 U7294 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6302), .B(n6294), .ZN(n6295) );
  OAI211_X1 U7295 ( .C1(n6308), .C2(n6297), .A(n6296), .B(n6295), .ZN(U3008)
         );
  INV_X1 U7296 ( .A(n6298), .ZN(n6299) );
  AOI21_X1 U7297 ( .B1(n6301), .B2(n6300), .A(n6299), .ZN(n6306) );
  AOI22_X1 U7298 ( .A1(n6304), .A2(n6303), .B1(n6302), .B2(n6307), .ZN(n6305)
         );
  OAI211_X1 U7299 ( .C1(n6308), .C2(n6307), .A(n6306), .B(n6305), .ZN(U3009)
         );
  NOR2_X1 U7300 ( .A1(n6662), .A2(n6599), .ZN(U3019) );
  INV_X1 U7301 ( .A(n6315), .ZN(n6313) );
  NAND2_X1 U7302 ( .A1(n6421), .A2(n6479), .ZN(n6346) );
  OR2_X1 U7303 ( .A1(n6478), .A2(n6346), .ZN(n6311) );
  NOR2_X1 U7304 ( .A1(n6309), .A2(n6312), .ZN(n6332) );
  INV_X1 U7305 ( .A(n6332), .ZN(n6310) );
  NAND2_X1 U7306 ( .A1(n6311), .A2(n6310), .ZN(n6314) );
  INV_X1 U7307 ( .A(n6312), .ZN(n6317) );
  AOI22_X1 U7308 ( .A1(n6475), .A2(n6332), .B1(n6341), .B2(n6487), .ZN(n6319)
         );
  OR2_X1 U7309 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  OAI211_X1 U7310 ( .C1(n6419), .C2(n6317), .A(n6316), .B(n6426), .ZN(n6334)
         );
  AOI22_X1 U7311 ( .A1(n6334), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n6435), 
        .B2(n6333), .ZN(n6318) );
  OAI211_X1 U7312 ( .C1(n6337), .C2(n6360), .A(n6319), .B(n6318), .ZN(U3060)
         );
  AOI22_X1 U7313 ( .A1(n6492), .A2(n6332), .B1(n6493), .B2(n6341), .ZN(n6321)
         );
  AOI22_X1 U7314 ( .A1(n6334), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n6438), 
        .B2(n6333), .ZN(n6320) );
  OAI211_X1 U7315 ( .C1(n6337), .C2(n6363), .A(n6321), .B(n6320), .ZN(U3061)
         );
  AOI22_X1 U7316 ( .A1(n6498), .A2(n6332), .B1(n6341), .B2(n6499), .ZN(n6323)
         );
  AOI22_X1 U7317 ( .A1(n6334), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n6442), 
        .B2(n6333), .ZN(n6322) );
  OAI211_X1 U7318 ( .C1(n6337), .C2(n6366), .A(n6323), .B(n6322), .ZN(U3062)
         );
  AOI22_X1 U7319 ( .A1(n6782), .A2(n6332), .B1(n6341), .B2(n6505), .ZN(n6325)
         );
  AOI22_X1 U7320 ( .A1(n6334), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n6446), 
        .B2(n6333), .ZN(n6324) );
  OAI211_X1 U7321 ( .C1(n6337), .C2(n6369), .A(n6325), .B(n6324), .ZN(U3063)
         );
  AOI22_X1 U7322 ( .A1(n6510), .A2(n6332), .B1(n6341), .B2(n6511), .ZN(n6327)
         );
  AOI22_X1 U7323 ( .A1(n6334), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n6450), 
        .B2(n6333), .ZN(n6326) );
  OAI211_X1 U7324 ( .C1(n6337), .C2(n6372), .A(n6327), .B(n6326), .ZN(U3064)
         );
  AOI22_X1 U7325 ( .A1(n6516), .A2(n6332), .B1(n6341), .B2(n6517), .ZN(n6329)
         );
  AOI22_X1 U7326 ( .A1(n6334), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n6454), 
        .B2(n6333), .ZN(n6328) );
  OAI211_X1 U7327 ( .C1(n6337), .C2(n6375), .A(n6329), .B(n6328), .ZN(U3065)
         );
  AOI22_X1 U7328 ( .A1(n6522), .A2(n6332), .B1(n6341), .B2(n6523), .ZN(n6331)
         );
  AOI22_X1 U7329 ( .A1(n6334), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n6457), 
        .B2(n6333), .ZN(n6330) );
  OAI211_X1 U7330 ( .C1(n6337), .C2(n6378), .A(n6331), .B(n6330), .ZN(U3066)
         );
  AOI22_X1 U7331 ( .A1(n6530), .A2(n6332), .B1(n6341), .B2(n6532), .ZN(n6336)
         );
  AOI22_X1 U7332 ( .A1(n6334), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n6463), 
        .B2(n6333), .ZN(n6335) );
  OAI211_X1 U7333 ( .C1(n6337), .C2(n6384), .A(n6336), .B(n6335), .ZN(U3067)
         );
  INV_X1 U7334 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6727) );
  INV_X1 U7335 ( .A(n6338), .ZN(n6339) );
  AOI22_X1 U7336 ( .A1(n6475), .A2(n6340), .B1(n6474), .B2(n6339), .ZN(n6343)
         );
  AOI22_X1 U7337 ( .A1(n6380), .A2(n6487), .B1(n6341), .B2(n6435), .ZN(n6342)
         );
  OAI211_X1 U7338 ( .C1(n6344), .C2(n6727), .A(n6343), .B(n6342), .ZN(U3068)
         );
  NAND2_X1 U7339 ( .A1(n6345), .A2(n6419), .ZN(n6355) );
  INV_X1 U7340 ( .A(n6355), .ZN(n6349) );
  OR2_X1 U7341 ( .A1(n6347), .A2(n6346), .ZN(n6348) );
  NAND2_X1 U7342 ( .A1(n6348), .A2(n6350), .ZN(n6354) );
  AOI22_X1 U7343 ( .A1(n6349), .A2(n6354), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6353), .ZN(n6385) );
  INV_X1 U7344 ( .A(n6350), .ZN(n6379) );
  AOI22_X1 U7345 ( .A1(n6475), .A2(n6379), .B1(n6487), .B2(n6391), .ZN(n6359)
         );
  OAI22_X1 U7346 ( .A1(n6355), .A2(n6354), .B1(n6353), .B2(n6419), .ZN(n6356)
         );
  INV_X1 U7347 ( .A(n6356), .ZN(n6357) );
  NAND2_X1 U7348 ( .A1(n6426), .A2(n6357), .ZN(n6381) );
  AOI22_X1 U7349 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6381), .B1(n6435), 
        .B2(n6380), .ZN(n6358) );
  OAI211_X1 U7350 ( .C1(n6385), .C2(n6360), .A(n6359), .B(n6358), .ZN(U3076)
         );
  AOI22_X1 U7351 ( .A1(n6492), .A2(n6379), .B1(n6380), .B2(n6438), .ZN(n6362)
         );
  AOI22_X1 U7352 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6381), .B1(n6493), 
        .B2(n6391), .ZN(n6361) );
  OAI211_X1 U7353 ( .C1(n6385), .C2(n6363), .A(n6362), .B(n6361), .ZN(U3077)
         );
  AOI22_X1 U7354 ( .A1(n6498), .A2(n6379), .B1(n6380), .B2(n6442), .ZN(n6365)
         );
  AOI22_X1 U7355 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6381), .B1(n6499), 
        .B2(n6391), .ZN(n6364) );
  OAI211_X1 U7356 ( .C1(n6385), .C2(n6366), .A(n6365), .B(n6364), .ZN(U3078)
         );
  AOI22_X1 U7357 ( .A1(n6782), .A2(n6379), .B1(n6505), .B2(n6391), .ZN(n6368)
         );
  AOI22_X1 U7358 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6381), .B1(n6446), 
        .B2(n6380), .ZN(n6367) );
  OAI211_X1 U7359 ( .C1(n6385), .C2(n6369), .A(n6368), .B(n6367), .ZN(U3079)
         );
  AOI22_X1 U7360 ( .A1(n6510), .A2(n6379), .B1(n6380), .B2(n6450), .ZN(n6371)
         );
  AOI22_X1 U7361 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6381), .B1(n6511), 
        .B2(n6391), .ZN(n6370) );
  OAI211_X1 U7362 ( .C1(n6385), .C2(n6372), .A(n6371), .B(n6370), .ZN(U3080)
         );
  AOI22_X1 U7363 ( .A1(n6516), .A2(n6379), .B1(n6380), .B2(n6454), .ZN(n6374)
         );
  AOI22_X1 U7364 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6381), .B1(n6517), 
        .B2(n6391), .ZN(n6373) );
  OAI211_X1 U7365 ( .C1(n6385), .C2(n6375), .A(n6374), .B(n6373), .ZN(U3081)
         );
  AOI22_X1 U7366 ( .A1(n6522), .A2(n6379), .B1(n6523), .B2(n6391), .ZN(n6377)
         );
  AOI22_X1 U7367 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6381), .B1(n6457), 
        .B2(n6380), .ZN(n6376) );
  OAI211_X1 U7368 ( .C1(n6385), .C2(n6378), .A(n6377), .B(n6376), .ZN(U3082)
         );
  AOI22_X1 U7369 ( .A1(n6530), .A2(n6379), .B1(n6532), .B2(n6391), .ZN(n6383)
         );
  AOI22_X1 U7370 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6381), .B1(n6463), 
        .B2(n6380), .ZN(n6382) );
  OAI211_X1 U7371 ( .C1(n6385), .C2(n6384), .A(n6383), .B(n6382), .ZN(U3083)
         );
  NOR2_X1 U7372 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6386), .ZN(n6413)
         );
  NAND2_X1 U7373 ( .A1(n6387), .A2(n4654), .ZN(n6392) );
  INV_X1 U7374 ( .A(n6388), .ZN(n6390) );
  OR2_X1 U7375 ( .A1(n6390), .A2(n6389), .ZN(n6472) );
  OAI22_X1 U7376 ( .A1(n6392), .A2(n6476), .B1(n6484), .B2(n6472), .ZN(n6412)
         );
  AOI22_X1 U7377 ( .A1(n6475), .A2(n6413), .B1(n6474), .B2(n6412), .ZN(n6399)
         );
  NOR3_X1 U7378 ( .A1(n6414), .A2(n6391), .A3(n6476), .ZN(n6393) );
  OAI21_X1 U7379 ( .B1(n6393), .B2(n6480), .A(n6392), .ZN(n6397) );
  AOI21_X1 U7380 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6472), .A(n6394), .ZN(
        n6485) );
  INV_X1 U7381 ( .A(n6413), .ZN(n6395) );
  NAND2_X1 U7382 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6395), .ZN(n6396) );
  NAND4_X1 U7383 ( .A1(n6397), .A2(n6485), .A3(n6471), .A4(n6396), .ZN(n6415)
         );
  AOI22_X1 U7384 ( .A1(n6415), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6414), 
        .B2(n6487), .ZN(n6398) );
  OAI211_X1 U7385 ( .C1(n6490), .C2(n6418), .A(n6399), .B(n6398), .ZN(U3084)
         );
  AOI22_X1 U7386 ( .A1(n6492), .A2(n6413), .B1(n6491), .B2(n6412), .ZN(n6401)
         );
  AOI22_X1 U7387 ( .A1(n6415), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6493), 
        .B2(n6414), .ZN(n6400) );
  OAI211_X1 U7388 ( .C1(n6496), .C2(n6418), .A(n6401), .B(n6400), .ZN(U3085)
         );
  AOI22_X1 U7389 ( .A1(n6498), .A2(n6413), .B1(n6497), .B2(n6412), .ZN(n6403)
         );
  AOI22_X1 U7390 ( .A1(n6415), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6499), 
        .B2(n6414), .ZN(n6402) );
  OAI211_X1 U7391 ( .C1(n6502), .C2(n6418), .A(n6403), .B(n6402), .ZN(U3086)
         );
  AOI22_X1 U7392 ( .A1(n6782), .A2(n6413), .B1(n6503), .B2(n6412), .ZN(n6405)
         );
  AOI22_X1 U7393 ( .A1(n6415), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6505), 
        .B2(n6414), .ZN(n6404) );
  OAI211_X1 U7394 ( .C1(n6508), .C2(n6418), .A(n6405), .B(n6404), .ZN(U3087)
         );
  AOI22_X1 U7395 ( .A1(n6510), .A2(n6413), .B1(n6509), .B2(n6412), .ZN(n6407)
         );
  AOI22_X1 U7396 ( .A1(n6415), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6511), 
        .B2(n6414), .ZN(n6406) );
  OAI211_X1 U7397 ( .C1(n6514), .C2(n6418), .A(n6407), .B(n6406), .ZN(U3088)
         );
  AOI22_X1 U7398 ( .A1(n6516), .A2(n6413), .B1(n6515), .B2(n6412), .ZN(n6409)
         );
  AOI22_X1 U7399 ( .A1(n6415), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6517), 
        .B2(n6414), .ZN(n6408) );
  OAI211_X1 U7400 ( .C1(n6520), .C2(n6418), .A(n6409), .B(n6408), .ZN(U3089)
         );
  AOI22_X1 U7401 ( .A1(n6522), .A2(n6413), .B1(n6521), .B2(n6412), .ZN(n6411)
         );
  AOI22_X1 U7402 ( .A1(n6415), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6523), 
        .B2(n6414), .ZN(n6410) );
  OAI211_X1 U7403 ( .C1(n6526), .C2(n6418), .A(n6411), .B(n6410), .ZN(U3090)
         );
  AOI22_X1 U7404 ( .A1(n6530), .A2(n6413), .B1(n6528), .B2(n6412), .ZN(n6417)
         );
  AOI22_X1 U7405 ( .A1(n6415), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6532), 
        .B2(n6414), .ZN(n6416) );
  OAI211_X1 U7406 ( .C1(n6537), .C2(n6418), .A(n6417), .B(n6416), .ZN(U3091)
         );
  OAI21_X1 U7407 ( .B1(n6428), .B2(n6420), .A(n6419), .ZN(n6434) );
  NAND2_X1 U7408 ( .A1(n6422), .A2(n6421), .ZN(n6425) );
  NOR2_X1 U7409 ( .A1(n6598), .A2(n6423), .ZN(n6464) );
  INV_X1 U7410 ( .A(n6464), .ZN(n6424) );
  NAND2_X1 U7411 ( .A1(n6425), .A2(n6424), .ZN(n6431) );
  OAI21_X1 U7412 ( .B1(n6434), .B2(n6431), .A(n6426), .ZN(n6427) );
  INV_X1 U7413 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n6708) );
  INV_X1 U7414 ( .A(n6428), .ZN(n6430) );
  AOI22_X1 U7415 ( .A1(n6475), .A2(n6464), .B1(n6487), .B2(n6477), .ZN(n6437)
         );
  INV_X1 U7416 ( .A(n6431), .ZN(n6433) );
  OAI22_X1 U7417 ( .A1(n6434), .A2(n6433), .B1(n6432), .B2(n5978), .ZN(n6465)
         );
  AOI22_X1 U7418 ( .A1(n6435), .A2(n6462), .B1(n6474), .B2(n6465), .ZN(n6436)
         );
  OAI211_X1 U7419 ( .C1(n6458), .C2(n6708), .A(n6437), .B(n6436), .ZN(U3108)
         );
  INV_X1 U7420 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n6441) );
  AOI22_X1 U7421 ( .A1(n6492), .A2(n6464), .B1(n6493), .B2(n6477), .ZN(n6440)
         );
  AOI22_X1 U7422 ( .A1(n6438), .A2(n6462), .B1(n6491), .B2(n6465), .ZN(n6439)
         );
  OAI211_X1 U7423 ( .C1(n6458), .C2(n6441), .A(n6440), .B(n6439), .ZN(U3109)
         );
  INV_X1 U7424 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6445) );
  AOI22_X1 U7425 ( .A1(n6498), .A2(n6464), .B1(n6499), .B2(n6477), .ZN(n6444)
         );
  AOI22_X1 U7426 ( .A1(n6442), .A2(n6462), .B1(n6497), .B2(n6465), .ZN(n6443)
         );
  OAI211_X1 U7427 ( .C1(n6458), .C2(n6445), .A(n6444), .B(n6443), .ZN(U3110)
         );
  INV_X1 U7428 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6449) );
  AOI22_X1 U7429 ( .A1(n6782), .A2(n6464), .B1(n6505), .B2(n6477), .ZN(n6448)
         );
  AOI22_X1 U7430 ( .A1(n6446), .A2(n6462), .B1(n6503), .B2(n6465), .ZN(n6447)
         );
  OAI211_X1 U7431 ( .C1(n6458), .C2(n6449), .A(n6448), .B(n6447), .ZN(U3111)
         );
  INV_X1 U7432 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6453) );
  AOI22_X1 U7433 ( .A1(n6510), .A2(n6464), .B1(n6511), .B2(n6477), .ZN(n6452)
         );
  AOI22_X1 U7434 ( .A1(n6450), .A2(n6462), .B1(n6509), .B2(n6465), .ZN(n6451)
         );
  OAI211_X1 U7435 ( .C1(n6458), .C2(n6453), .A(n6452), .B(n6451), .ZN(U3112)
         );
  INV_X1 U7436 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6705) );
  AOI22_X1 U7437 ( .A1(n6516), .A2(n6464), .B1(n6517), .B2(n6477), .ZN(n6456)
         );
  AOI22_X1 U7438 ( .A1(n6454), .A2(n6462), .B1(n6515), .B2(n6465), .ZN(n6455)
         );
  OAI211_X1 U7439 ( .C1(n6458), .C2(n6705), .A(n6456), .B(n6455), .ZN(U3113)
         );
  AOI22_X1 U7440 ( .A1(n6522), .A2(n6464), .B1(n6457), .B2(n6462), .ZN(n6460)
         );
  INV_X1 U7441 ( .A(n6458), .ZN(n6466) );
  AOI22_X1 U7442 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6466), .B1(n6521), 
        .B2(n6465), .ZN(n6459) );
  OAI211_X1 U7443 ( .C1(n6461), .C2(n6536), .A(n6460), .B(n6459), .ZN(U3114)
         );
  AOI22_X1 U7444 ( .A1(n6530), .A2(n6464), .B1(n6463), .B2(n6462), .ZN(n6468)
         );
  AOI22_X1 U7445 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6466), .B1(n6528), 
        .B2(n6465), .ZN(n6467) );
  OAI211_X1 U7446 ( .C1(n6469), .C2(n6536), .A(n6468), .B(n6467), .ZN(U3115)
         );
  NOR2_X1 U7447 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6470), .ZN(n6529)
         );
  OAI22_X1 U7448 ( .A1(n6473), .A2(n6592), .B1(n6472), .B2(n6471), .ZN(n6527)
         );
  AOI22_X1 U7449 ( .A1(n6475), .A2(n6529), .B1(n6474), .B2(n6527), .ZN(n6489)
         );
  NOR3_X1 U7450 ( .A1(n6477), .A2(n6531), .A3(n6476), .ZN(n6481) );
  OAI22_X1 U7451 ( .A1(n6481), .A2(n6480), .B1(n6479), .B2(n6478), .ZN(n6486)
         );
  INV_X1 U7452 ( .A(n6529), .ZN(n6482) );
  NAND2_X1 U7453 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6482), .ZN(n6483) );
  NAND4_X1 U7454 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(n6533)
         );
  AOI22_X1 U7455 ( .A1(n6533), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6487), 
        .B2(n6531), .ZN(n6488) );
  OAI211_X1 U7456 ( .C1(n6490), .C2(n6536), .A(n6489), .B(n6488), .ZN(U3116)
         );
  AOI22_X1 U7457 ( .A1(n6492), .A2(n6529), .B1(n6491), .B2(n6527), .ZN(n6495)
         );
  AOI22_X1 U7458 ( .A1(n6533), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6493), 
        .B2(n6531), .ZN(n6494) );
  OAI211_X1 U7459 ( .C1(n6496), .C2(n6536), .A(n6495), .B(n6494), .ZN(U3117)
         );
  AOI22_X1 U7460 ( .A1(n6498), .A2(n6529), .B1(n6497), .B2(n6527), .ZN(n6501)
         );
  AOI22_X1 U7461 ( .A1(n6533), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6499), 
        .B2(n6531), .ZN(n6500) );
  OAI211_X1 U7462 ( .C1(n6502), .C2(n6536), .A(n6501), .B(n6500), .ZN(U3118)
         );
  AOI22_X1 U7463 ( .A1(n6782), .A2(n6529), .B1(n6503), .B2(n6527), .ZN(n6507)
         );
  AOI22_X1 U7464 ( .A1(n6533), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6505), 
        .B2(n6531), .ZN(n6506) );
  OAI211_X1 U7465 ( .C1(n6508), .C2(n6536), .A(n6507), .B(n6506), .ZN(U3119)
         );
  AOI22_X1 U7466 ( .A1(n6510), .A2(n6529), .B1(n6509), .B2(n6527), .ZN(n6513)
         );
  AOI22_X1 U7467 ( .A1(n6533), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6511), 
        .B2(n6531), .ZN(n6512) );
  OAI211_X1 U7468 ( .C1(n6514), .C2(n6536), .A(n6513), .B(n6512), .ZN(U3120)
         );
  AOI22_X1 U7469 ( .A1(n6516), .A2(n6529), .B1(n6515), .B2(n6527), .ZN(n6519)
         );
  AOI22_X1 U7470 ( .A1(n6533), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6517), 
        .B2(n6531), .ZN(n6518) );
  OAI211_X1 U7471 ( .C1(n6520), .C2(n6536), .A(n6519), .B(n6518), .ZN(U3121)
         );
  AOI22_X1 U7472 ( .A1(n6522), .A2(n6529), .B1(n6521), .B2(n6527), .ZN(n6525)
         );
  AOI22_X1 U7473 ( .A1(n6533), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6523), 
        .B2(n6531), .ZN(n6524) );
  OAI211_X1 U7474 ( .C1(n6526), .C2(n6536), .A(n6525), .B(n6524), .ZN(U3122)
         );
  AOI22_X1 U7475 ( .A1(n6530), .A2(n6529), .B1(n6528), .B2(n6527), .ZN(n6535)
         );
  AOI22_X1 U7476 ( .A1(n6533), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6532), 
        .B2(n6531), .ZN(n6534) );
  OAI211_X1 U7477 ( .C1(n6537), .C2(n6536), .A(n6535), .B(n6534), .ZN(U3123)
         );
  AND3_X1 U7478 ( .A1(n6539), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6538), 
        .ZN(n6544) );
  AOI21_X1 U7479 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6544), .A(n6540), 
        .ZN(n6541) );
  NAND2_X1 U7480 ( .A1(n6542), .A2(n6541), .ZN(n6543) );
  OAI21_X1 U7481 ( .B1(n6544), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6543), 
        .ZN(n6545) );
  AOI222_X1 U7482 ( .A1(n6547), .A2(n6546), .B1(n6547), .B2(n6545), .C1(n6546), 
        .C2(n6545), .ZN(n6549) );
  OAI21_X1 U7483 ( .B1(n6549), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6548), 
        .ZN(n6558) );
  AOI21_X1 U7484 ( .B1(n6549), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6557) );
  OAI21_X1 U7485 ( .B1(MORE_REG_SCAN_IN), .B2(FLUSH_REG_SCAN_IN), .A(n6550), 
        .ZN(n6551) );
  NAND4_X1 U7486 ( .A1(n6554), .A2(n6553), .A3(n6552), .A4(n6551), .ZN(n6555)
         );
  AOI211_X1 U7487 ( .C1(n6558), .C2(n6557), .A(n6556), .B(n6555), .ZN(n6571)
         );
  AOI22_X1 U7488 ( .A1(n6571), .A2(n6559), .B1(READY_N), .B2(n6612), .ZN(n6560) );
  INV_X1 U7489 ( .A(n6560), .ZN(n6561) );
  OAI21_X1 U7490 ( .B1(n6563), .B2(n6562), .A(n6561), .ZN(n6589) );
  OAI21_X1 U7491 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6611), .A(n6589), .ZN(
        n6572) );
  AOI221_X1 U7492 ( .B1(n6565), .B2(STATE2_REG_0__SCAN_IN), .C1(n6572), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6564), .ZN(n6570) );
  OAI211_X1 U7493 ( .C1(n6568), .C2(n6567), .A(n6566), .B(n6589), .ZN(n6569)
         );
  OAI211_X1 U7494 ( .C1(n6571), .C2(n6573), .A(n6570), .B(n6569), .ZN(U3148)
         );
  OAI211_X1 U7495 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6572), .ZN(n6578) );
  OAI21_X1 U7496 ( .B1(READY_N), .B2(n6574), .A(n6573), .ZN(n6576) );
  AOI21_X1 U7497 ( .B1(n6576), .B2(n6589), .A(n6575), .ZN(n6577) );
  NAND2_X1 U7498 ( .A1(n6578), .A2(n6577), .ZN(U3149) );
  OAI221_X1 U7499 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6611), .A(n6586), .ZN(n6580) );
  OAI21_X1 U7500 ( .B1(n6615), .B2(n6580), .A(n6579), .ZN(U3150) );
  AND2_X1 U7501 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6582), .ZN(U3151) );
  AND2_X1 U7502 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6582), .ZN(U3152) );
  AND2_X1 U7503 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6582), .ZN(U3153) );
  AND2_X1 U7504 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6582), .ZN(U3154) );
  AND2_X1 U7505 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6582), .ZN(U3155) );
  AND2_X1 U7506 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6582), .ZN(U3156) );
  AND2_X1 U7507 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6582), .ZN(U3157) );
  INV_X1 U7508 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6671) );
  NOR2_X1 U7509 ( .A1(n6585), .A2(n6671), .ZN(U3158) );
  AND2_X1 U7510 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6582), .ZN(U3159) );
  AND2_X1 U7511 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6582), .ZN(U3160) );
  AND2_X1 U7512 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6582), .ZN(U3161) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6582), .ZN(U3162) );
  INV_X1 U7514 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6688) );
  NOR2_X1 U7515 ( .A1(n6585), .A2(n6688), .ZN(U3163) );
  AND2_X1 U7516 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6582), .ZN(U3164) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6582), .ZN(U3165) );
  AND2_X1 U7518 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6582), .ZN(U3166) );
  AND2_X1 U7519 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6582), .ZN(U3167) );
  AND2_X1 U7520 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6582), .ZN(U3168) );
  AND2_X1 U7521 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6582), .ZN(U3169) );
  AND2_X1 U7522 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6582), .ZN(U3170) );
  AND2_X1 U7523 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6582), .ZN(U3171) );
  AND2_X1 U7524 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6582), .ZN(U3172) );
  AND2_X1 U7525 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6582), .ZN(U3173) );
  AND2_X1 U7526 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6582), .ZN(U3174) );
  INV_X1 U7527 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6645) );
  NOR2_X1 U7528 ( .A1(n6585), .A2(n6645), .ZN(U3175) );
  AND2_X1 U7529 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6582), .ZN(U3176) );
  AND2_X1 U7530 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6582), .ZN(U3177) );
  AND2_X1 U7531 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6582), .ZN(U3178) );
  AND2_X1 U7532 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6582), .ZN(U3179) );
  AND2_X1 U7533 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6582), .ZN(U3180) );
  INV_X1 U7534 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6601) );
  INV_X1 U7535 ( .A(n6583), .ZN(n6581) );
  AOI21_X1 U7536 ( .B1(n6601), .B2(n6582), .A(n6581), .ZN(U3451) );
  INV_X1 U7537 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6584) );
  OAI21_X1 U7538 ( .B1(n6585), .B2(n6584), .A(n6583), .ZN(U3452) );
  OAI211_X1 U7539 ( .C1(n6589), .C2(n6588), .A(n6587), .B(n6586), .ZN(U3453)
         );
  INV_X1 U7540 ( .A(n6590), .ZN(n6594) );
  OAI22_X1 U7541 ( .A1(n6594), .A2(n6593), .B1(n6592), .B2(n6591), .ZN(n6595)
         );
  OAI21_X1 U7542 ( .B1(n6596), .B2(n6595), .A(n6599), .ZN(n6597) );
  OAI21_X1 U7543 ( .B1(n6599), .B2(n6598), .A(n6597), .ZN(U3462) );
  NOR3_X1 U7544 ( .A1(n6601), .A2(REIP_REG_0__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6600) );
  AOI221_X1 U7545 ( .B1(n6602), .B2(n6601), .C1(REIP_REG_1__SCAN_IN), .C2(
        REIP_REG_0__SCAN_IN), .A(n6600), .ZN(n6604) );
  INV_X1 U7546 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6603) );
  INV_X1 U7547 ( .A(n6608), .ZN(n6605) );
  AOI22_X1 U7548 ( .A1(n6608), .A2(n6604), .B1(n6603), .B2(n6605), .ZN(U3468)
         );
  NOR2_X1 U7549 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6607) );
  INV_X1 U7550 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U7551 ( .A1(n6608), .A2(n6607), .B1(n6606), .B2(n6605), .ZN(U3469)
         );
  AOI211_X1 U7552 ( .C1(n6612), .C2(n6611), .A(n6610), .B(n6609), .ZN(n6619)
         );
  OAI211_X1 U7553 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6614), .A(n6613), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6616) );
  AOI21_X1 U7554 ( .B1(n6616), .B2(STATE2_REG_0__SCAN_IN), .A(n6615), .ZN(
        n6618) );
  NAND2_X1 U7555 ( .A1(n6619), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6617) );
  OAI21_X1 U7556 ( .B1(n6619), .B2(n6618), .A(n6617), .ZN(U3472) );
  INV_X1 U7557 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6642) );
  NAND4_X1 U7558 ( .A1(UWORD_REG_12__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(n6642), .A4(n3453), .ZN(n6623) );
  INV_X1 U7559 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6647) );
  NAND4_X1 U7560 ( .A1(EBX_REG_26__SCAN_IN), .A2(EBX_REG_11__SCAN_IN), .A3(
        n6647), .A4(n6650), .ZN(n6622) );
  NAND4_X1 U7561 ( .A1(EBX_REG_2__SCAN_IN), .A2(EAX_REG_7__SCAN_IN), .A3(n3771), .A4(n6659), .ZN(n6621) );
  INV_X1 U7562 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6664) );
  NAND4_X1 U7563 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        BYTEENABLE_REG_1__SCAN_IN), .A3(n6661), .A4(n6664), .ZN(n6620) );
  NOR4_X1 U7564 ( .A1(n6623), .A2(n6622), .A3(n6621), .A4(n6620), .ZN(n6773)
         );
  NAND4_X1 U7565 ( .A1(EAX_REG_29__SCAN_IN), .A2(DATAI_5_), .A3(n6677), .A4(
        n6678), .ZN(n6640) );
  NAND4_X1 U7566 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(n6679), .A4(n6672), .ZN(n6639) );
  NOR3_X1 U7567 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(EBX_REG_12__SCAN_IN), 
        .A3(EAX_REG_30__SCAN_IN), .ZN(n6626) );
  NOR3_X1 U7568 ( .A1(EAX_REG_20__SCAN_IN), .A2(DATAWIDTH_REG_19__SCAN_IN), 
        .A3(n6624), .ZN(n6625) );
  NAND4_X1 U7569 ( .A1(STATE_REG_1__SCAN_IN), .A2(EAX_REG_10__SCAN_IN), .A3(
        n6626), .A4(n6625), .ZN(n6638) );
  INV_X1 U7570 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6754) );
  NAND4_X1 U7571 ( .A1(EBX_REG_13__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_0__SCAN_IN), .A4(n6754), .ZN(n6629) );
  NAND3_X1 U7572 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(M_IO_N_REG_SCAN_IN), 
        .A3(n6760), .ZN(n6628) );
  INV_X1 U7573 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6739) );
  NAND4_X1 U7574 ( .A1(EBX_REG_4__SCAN_IN), .A2(ADDRESS_REG_23__SCAN_IN), .A3(
        n6736), .A4(n6739), .ZN(n6627) );
  NOR4_X1 U7575 ( .A1(ADDRESS_REG_27__SCAN_IN), .A2(n6629), .A3(n6628), .A4(
        n6627), .ZN(n6636) );
  NAND3_X1 U7576 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUE_REG_9__0__SCAN_IN), .A3(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n6632) );
  NAND4_X1 U7577 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(
        INSTQUEUE_REG_11__0__SCAN_IN), .A3(INSTQUEUE_REG_11__5__SCAN_IN), .A4(
        n6706), .ZN(n6631) );
  NAND4_X1 U7578 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(
        INSTQUEUE_REG_3__2__SCAN_IN), .A3(DATAI_24_), .A4(DATAI_0_), .ZN(n6630) );
  NOR4_X1 U7579 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6632), .A3(n6631), .A4(
        n6630), .ZN(n6635) );
  NOR4_X1 U7580 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(
        INSTQUEUE_REG_6__0__SCAN_IN), .A3(ADDRESS_REG_29__SCAN_IN), .A4(n6723), 
        .ZN(n6634) );
  AND4_X1 U7581 ( .A1(n6743), .A2(n6744), .A3(INSTQUEUE_REG_0__6__SCAN_IN), 
        .A4(EBX_REG_25__SCAN_IN), .ZN(n6633) );
  NAND4_X1 U7582 ( .A1(n6636), .A2(n6635), .A3(n6634), .A4(n6633), .ZN(n6637)
         );
  NOR4_X1 U7583 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n6772)
         );
  AOI22_X1 U7584 ( .A1(n6643), .A2(keyinput13), .B1(n6642), .B2(keyinput17), 
        .ZN(n6641) );
  OAI221_X1 U7585 ( .B1(n6643), .B2(keyinput13), .C1(n6642), .C2(keyinput17), 
        .A(n6641), .ZN(n6655) );
  AOI22_X1 U7586 ( .A1(n6645), .A2(keyinput8), .B1(n3453), .B2(keyinput7), 
        .ZN(n6644) );
  OAI221_X1 U7587 ( .B1(n6645), .B2(keyinput8), .C1(n3453), .C2(keyinput7), 
        .A(n6644), .ZN(n6654) );
  AOI22_X1 U7588 ( .A1(n6648), .A2(keyinput43), .B1(n6647), .B2(keyinput23), 
        .ZN(n6646) );
  OAI221_X1 U7589 ( .B1(n6648), .B2(keyinput43), .C1(n6647), .C2(keyinput23), 
        .A(n6646), .ZN(n6653) );
  AOI22_X1 U7590 ( .A1(n6651), .A2(keyinput5), .B1(n6650), .B2(keyinput59), 
        .ZN(n6649) );
  OAI221_X1 U7591 ( .B1(n6651), .B2(keyinput5), .C1(n6650), .C2(keyinput59), 
        .A(n6649), .ZN(n6652) );
  NOR4_X1 U7592 ( .A1(n6655), .A2(n6654), .A3(n6653), .A4(n6652), .ZN(n6703)
         );
  AOI22_X1 U7593 ( .A1(n3571), .A2(keyinput50), .B1(n6657), .B2(keyinput16), 
        .ZN(n6656) );
  OAI221_X1 U7594 ( .B1(n3571), .B2(keyinput50), .C1(n6657), .C2(keyinput16), 
        .A(n6656), .ZN(n6669) );
  AOI22_X1 U7595 ( .A1(n3771), .A2(keyinput0), .B1(keyinput40), .B2(n6659), 
        .ZN(n6658) );
  OAI221_X1 U7596 ( .B1(n3771), .B2(keyinput0), .C1(n6659), .C2(keyinput40), 
        .A(n6658), .ZN(n6668) );
  AOI22_X1 U7597 ( .A1(n6662), .A2(keyinput44), .B1(keyinput48), .B2(n6661), 
        .ZN(n6660) );
  OAI221_X1 U7598 ( .B1(n6662), .B2(keyinput44), .C1(n6661), .C2(keyinput48), 
        .A(n6660), .ZN(n6667) );
  AOI22_X1 U7599 ( .A1(n6665), .A2(keyinput11), .B1(n6664), .B2(keyinput34), 
        .ZN(n6663) );
  OAI221_X1 U7600 ( .B1(n6665), .B2(keyinput11), .C1(n6664), .C2(keyinput34), 
        .A(n6663), .ZN(n6666) );
  NOR4_X1 U7601 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6702)
         );
  AOI22_X1 U7602 ( .A1(n6672), .A2(keyinput61), .B1(keyinput51), .B2(n6671), 
        .ZN(n6670) );
  OAI221_X1 U7603 ( .B1(n6672), .B2(keyinput61), .C1(n6671), .C2(keyinput51), 
        .A(n6670), .ZN(n6685) );
  AOI22_X1 U7604 ( .A1(n6675), .A2(keyinput33), .B1(n6674), .B2(keyinput9), 
        .ZN(n6673) );
  OAI221_X1 U7605 ( .B1(n6675), .B2(keyinput33), .C1(n6674), .C2(keyinput9), 
        .A(n6673), .ZN(n6684) );
  AOI22_X1 U7606 ( .A1(n6678), .A2(keyinput47), .B1(n6677), .B2(keyinput36), 
        .ZN(n6676) );
  OAI221_X1 U7607 ( .B1(n6678), .B2(keyinput47), .C1(n6677), .C2(keyinput36), 
        .A(n6676), .ZN(n6683) );
  XOR2_X1 U7608 ( .A(n6679), .B(keyinput29), .Z(n6681) );
  XNOR2_X1 U7609 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .B(keyinput60), .ZN(n6680)
         );
  NAND2_X1 U7610 ( .A1(n6681), .A2(n6680), .ZN(n6682) );
  NOR4_X1 U7611 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .ZN(n6701)
         );
  AOI22_X1 U7612 ( .A1(n6688), .A2(keyinput28), .B1(n6687), .B2(keyinput31), 
        .ZN(n6686) );
  OAI221_X1 U7613 ( .B1(n6688), .B2(keyinput28), .C1(n6687), .C2(keyinput31), 
        .A(n6686), .ZN(n6699) );
  AOI22_X1 U7614 ( .A1(n4130), .A2(keyinput4), .B1(n6690), .B2(keyinput22), 
        .ZN(n6689) );
  OAI221_X1 U7615 ( .B1(n4130), .B2(keyinput4), .C1(n6690), .C2(keyinput22), 
        .A(n6689), .ZN(n6698) );
  INV_X1 U7616 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6692) );
  AOI22_X1 U7617 ( .A1(n6693), .A2(keyinput14), .B1(n6692), .B2(keyinput46), 
        .ZN(n6691) );
  OAI221_X1 U7618 ( .B1(n6693), .B2(keyinput14), .C1(n6692), .C2(keyinput46), 
        .A(n6691), .ZN(n6697) );
  XNOR2_X1 U7619 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput39), .ZN(n6695) );
  XNOR2_X1 U7620 ( .A(keyinput37), .B(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6694) );
  NAND2_X1 U7621 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  NOR4_X1 U7622 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n6700)
         );
  NAND4_X1 U7623 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6771)
         );
  AOI22_X1 U7624 ( .A1(n6706), .A2(keyinput12), .B1(n6705), .B2(keyinput53), 
        .ZN(n6704) );
  OAI221_X1 U7625 ( .B1(n6706), .B2(keyinput12), .C1(n6705), .C2(keyinput53), 
        .A(n6704), .ZN(n6718) );
  AOI22_X1 U7626 ( .A1(n4934), .A2(keyinput57), .B1(n6708), .B2(keyinput20), 
        .ZN(n6707) );
  OAI221_X1 U7627 ( .B1(n4934), .B2(keyinput57), .C1(n6708), .C2(keyinput20), 
        .A(n6707), .ZN(n6717) );
  INV_X1 U7628 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6711) );
  INV_X1 U7629 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6710) );
  AOI22_X1 U7630 ( .A1(n6711), .A2(keyinput52), .B1(keyinput21), .B2(n6710), 
        .ZN(n6709) );
  OAI221_X1 U7631 ( .B1(n6711), .B2(keyinput52), .C1(n6710), .C2(keyinput21), 
        .A(n6709), .ZN(n6716) );
  AOI22_X1 U7632 ( .A1(n6714), .A2(keyinput26), .B1(keyinput45), .B2(n6713), 
        .ZN(n6712) );
  OAI221_X1 U7633 ( .B1(n6714), .B2(keyinput26), .C1(n6713), .C2(keyinput45), 
        .A(n6712), .ZN(n6715) );
  NOR4_X1 U7634 ( .A1(n6718), .A2(n6717), .A3(n6716), .A4(n6715), .ZN(n6769)
         );
  INV_X1 U7635 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6720) );
  AOI22_X1 U7636 ( .A1(n6721), .A2(keyinput35), .B1(n6720), .B2(keyinput6), 
        .ZN(n6719) );
  OAI221_X1 U7637 ( .B1(n6721), .B2(keyinput35), .C1(n6720), .C2(keyinput6), 
        .A(n6719), .ZN(n6734) );
  AOI22_X1 U7638 ( .A1(n6724), .A2(keyinput10), .B1(n6723), .B2(keyinput3), 
        .ZN(n6722) );
  OAI221_X1 U7639 ( .B1(n6724), .B2(keyinput10), .C1(n6723), .C2(keyinput3), 
        .A(n6722), .ZN(n6733) );
  INV_X1 U7640 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6726) );
  AOI22_X1 U7641 ( .A1(n6727), .A2(keyinput25), .B1(n6726), .B2(keyinput41), 
        .ZN(n6725) );
  OAI221_X1 U7642 ( .B1(n6727), .B2(keyinput25), .C1(n6726), .C2(keyinput41), 
        .A(n6725), .ZN(n6732) );
  INV_X1 U7643 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6728) );
  XOR2_X1 U7644 ( .A(n6728), .B(keyinput56), .Z(n6730) );
  XNOR2_X1 U7645 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput49), .ZN(
        n6729) );
  NAND2_X1 U7646 ( .A1(n6730), .A2(n6729), .ZN(n6731) );
  NOR4_X1 U7647 ( .A1(n6734), .A2(n6733), .A3(n6732), .A4(n6731), .ZN(n6768)
         );
  AOI22_X1 U7648 ( .A1(n6737), .A2(keyinput38), .B1(keyinput18), .B2(n6736), 
        .ZN(n6735) );
  OAI221_X1 U7649 ( .B1(n6737), .B2(keyinput38), .C1(n6736), .C2(keyinput18), 
        .A(n6735), .ZN(n6750) );
  AOI22_X1 U7650 ( .A1(n6740), .A2(keyinput62), .B1(keyinput19), .B2(n6739), 
        .ZN(n6738) );
  OAI221_X1 U7651 ( .B1(n6740), .B2(keyinput62), .C1(n6739), .C2(keyinput19), 
        .A(n6738), .ZN(n6749) );
  AOI22_X1 U7652 ( .A1(n6743), .A2(keyinput32), .B1(keyinput42), .B2(n6742), 
        .ZN(n6741) );
  OAI221_X1 U7653 ( .B1(n6743), .B2(keyinput32), .C1(n6742), .C2(keyinput42), 
        .A(n6741), .ZN(n6748) );
  INV_X1 U7654 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6744) );
  XOR2_X1 U7655 ( .A(n6744), .B(keyinput63), .Z(n6746) );
  XNOR2_X1 U7656 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput58), .ZN(n6745)
         );
  NAND2_X1 U7657 ( .A1(n6746), .A2(n6745), .ZN(n6747) );
  NOR4_X1 U7658 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n6767)
         );
  AOI22_X1 U7659 ( .A1(n6752), .A2(keyinput15), .B1(n5212), .B2(keyinput2), 
        .ZN(n6751) );
  OAI221_X1 U7660 ( .B1(n6752), .B2(keyinput15), .C1(n5212), .C2(keyinput2), 
        .A(n6751), .ZN(n6765) );
  AOI22_X1 U7661 ( .A1(n6755), .A2(keyinput30), .B1(n6754), .B2(keyinput55), 
        .ZN(n6753) );
  OAI221_X1 U7662 ( .B1(n6755), .B2(keyinput30), .C1(n6754), .C2(keyinput55), 
        .A(n6753), .ZN(n6764) );
  INV_X1 U7663 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6757) );
  AOI22_X1 U7664 ( .A1(n6758), .A2(keyinput54), .B1(keyinput1), .B2(n6757), 
        .ZN(n6756) );
  OAI221_X1 U7665 ( .B1(n6758), .B2(keyinput54), .C1(n6757), .C2(keyinput1), 
        .A(n6756), .ZN(n6763) );
  AOI22_X1 U7666 ( .A1(n6761), .A2(keyinput27), .B1(keyinput24), .B2(n6760), 
        .ZN(n6759) );
  OAI221_X1 U7667 ( .B1(n6761), .B2(keyinput27), .C1(n6760), .C2(keyinput24), 
        .A(n6759), .ZN(n6762) );
  NOR4_X1 U7668 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n6766)
         );
  NAND4_X1 U7669 ( .A1(n6769), .A2(n6768), .A3(n6767), .A4(n6766), .ZN(n6770)
         );
  AOI211_X1 U7670 ( .C1(n6773), .C2(n6772), .A(n6771), .B(n6770), .ZN(n6781)
         );
  AOI22_X1 U7671 ( .A1(n3031), .A2(DATAI_18_), .B1(n6774), .B2(DATAI_2_), .ZN(
        n6775) );
  OAI21_X1 U7672 ( .B1(n6777), .B2(n6776), .A(n6775), .ZN(n6778) );
  AOI21_X1 U7673 ( .B1(EAX_REG_18__SCAN_IN), .B2(n6779), .A(n6778), .ZN(n6780)
         );
  XNOR2_X1 U7674 ( .A(n6781), .B(n6780), .ZN(U2873) );
  AND2_X1 U3575 ( .A1(n3226), .A2(n3225), .ZN(n3372) );
  AND2_X1 U3440 ( .A1(n3225), .A2(n4723), .ZN(n3470) );
  NAND2_X1 U4094 ( .A1(n3131), .A2(n3132), .ZN(n3530) );
  AND2_X2 U3458 ( .A1(n2980), .A2(n4707), .ZN(n2963) );
  XNOR2_X1 U4065 ( .A(n3440), .B(n3371), .ZN(n4341) );
  NAND2_X1 U4409 ( .A1(n3448), .A2(n3447), .ZN(n5041) );
  CLKBUF_X1 U3409 ( .A(n3407), .Z(n4092) );
  AND2_X1 U3424 ( .A1(n5147), .A2(n3220), .ZN(n3303) );
  CLKBUF_X1 U3428 ( .A(n3347), .Z(n3996) );
  INV_X2 U3441 ( .A(n5655), .ZN(n5609) );
  CLKBUF_X2 U3442 ( .A(n4723), .Z(n2981) );
  CLKBUF_X1 U34450 ( .A(n3359), .Z(n5164) );
  CLKBUF_X1 U3450 ( .A(n6229), .Z(n6612) );
  NAND2_X1 U34550 ( .A1(n5525), .A2(n4327), .ZN(n5516) );
  OR2_X1 U34600 ( .A1(n4697), .A2(n4685), .ZN(n6504) );
  INV_X1 U3479 ( .A(n6504), .ZN(n6782) );
endmodule

