

module b21_C_AntiSAT_k_256_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416;

  INV_X2 U4977 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X4 U4978 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4979 ( .A1(n6432), .A2(n6433), .ZN(n6431) );
  BUF_X1 U4980 ( .A(n5228), .Z(n5702) );
  BUF_X2 U4981 ( .A(n6318), .Z(n7893) );
  CLKBUF_X2 U4982 ( .A(n6322), .Z(n8005) );
  AND2_X1 U4983 ( .A1(n7643), .A2(n5084), .ZN(n5309) );
  CLKBUF_X1 U4984 ( .A(n5986), .Z(n4659) );
  OR3_X1 U4985 ( .A1(n8912), .A2(n8911), .A3(n8910), .ZN(n8916) );
  BUF_X1 U4986 ( .A(n6261), .Z(n7985) );
  INV_X2 U4987 ( .A(n8001), .ZN(n7996) );
  INV_X1 U4988 ( .A(n7690), .ZN(n6170) );
  NOR2_X1 U4989 ( .A1(n6835), .A2(n9961), .ZN(n6951) );
  NAND2_X1 U4990 ( .A1(n5081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U4992 ( .A1(n6149), .A2(n9457), .ZN(n6151) );
  OAI211_X1 U4993 ( .C1(P1_IR_REG_31__SCAN_IN), .C2(n5847), .A(n5846), .B(
        n6146), .ZN(n6249) );
  INV_X1 U4994 ( .A(n7069), .ZN(n7549) );
  AND4_X1 U4995 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .ZN(n6895)
         );
  INV_X1 U4996 ( .A(n6151), .ZN(n9466) );
  INV_X2 U4997 ( .A(n4659), .ZN(n7677) );
  INV_X1 U4998 ( .A(n9573), .ZN(n7687) );
  CLKBUF_X2 U4999 ( .A(n6256), .Z(n4473) );
  OAI21_X2 U5000 ( .B1(n5013), .B2(n5012), .A(n5010), .ZN(n6432) );
  OAI21_X2 U5001 ( .B1(n9189), .B2(n8928), .A(n8929), .ZN(n9177) );
  XNOR2_X2 U5002 ( .A(n5367), .B(n5365), .ZN(n7053) );
  NAND2_X2 U5003 ( .A1(n5333), .A2(n5332), .ZN(n6825) );
  OAI21_X2 U5004 ( .B1(n6431), .B2(n5036), .A(n5033), .ZN(n6718) );
  OR2_X1 U5005 ( .A1(n9961), .A2(n6828), .ZN(n7756) );
  NAND2_X2 U5006 ( .A1(n5355), .A2(n5354), .ZN(n9961) );
  XNOR2_X2 U5007 ( .A(n5094), .B(n5076), .ZN(n7878) );
  NAND2_X1 U5008 ( .A1(n7442), .A2(n7858), .ZN(n7648) );
  NOR2_X2 U5009 ( .A1(n7846), .A2(n5039), .ZN(n5038) );
  NAND2_X2 U5010 ( .A1(n7737), .A2(n7736), .ZN(n7846) );
  INV_X1 U5011 ( .A(n6249), .ZN(n6754) );
  NAND2_X2 U5012 ( .A1(n7878), .A2(n5794), .ZN(n6077) );
  NAND2_X1 U5013 ( .A1(n8021), .A2(n5718), .ZN(n5786) );
  NAND2_X1 U5014 ( .A1(n4677), .A2(n4676), .ZN(n4910) );
  AND2_X1 U5015 ( .A1(n4677), .A2(n4682), .ZN(n8046) );
  NAND2_X1 U5016 ( .A1(n8055), .A2(n8054), .ZN(n4677) );
  NAND2_X1 U5017 ( .A1(n4681), .A2(n4679), .ZN(n8055) );
  AND2_X1 U5018 ( .A1(n4682), .A2(n4911), .ZN(n4676) );
  NAND2_X1 U5019 ( .A1(n4683), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U5020 ( .A1(n8028), .A2(n8027), .ZN(n4683) );
  AND2_X1 U5021 ( .A1(n4494), .A2(n5654), .ZN(n4680) );
  NAND2_X1 U5022 ( .A1(n9229), .A2(n8932), .ZN(n4644) );
  CLKBUF_X1 U5023 ( .A(n7467), .Z(n4566) );
  NAND2_X1 U5024 ( .A1(n8430), .A2(n7782), .ZN(n8416) );
  AOI21_X1 U5025 ( .B1(n7906), .B2(n4858), .A(n4856), .ZN(n4855) );
  NAND2_X1 U5026 ( .A1(n7887), .A2(n7886), .ZN(n7906) );
  XNOR2_X1 U5027 ( .A(n8488), .B(n8111), .ZN(n8326) );
  NAND2_X1 U5028 ( .A1(n5666), .A2(n5665), .ZN(n8488) );
  NAND2_X1 U5029 ( .A1(n5680), .A2(n5679), .ZN(n8482) );
  NAND2_X1 U5030 ( .A1(n4870), .A2(n5444), .ZN(n7083) );
  NAND2_X1 U5031 ( .A1(n5582), .A2(n5581), .ZN(n8508) );
  NAND2_X1 U5032 ( .A1(n5545), .A2(n5544), .ZN(n8519) );
  OR2_X1 U5033 ( .A1(n7079), .A2(n8812), .ZN(n9501) );
  AND2_X1 U5034 ( .A1(n7747), .A2(n7746), .ZN(n7851) );
  AND2_X1 U5035 ( .A1(n7050), .A2(n7049), .ZN(n9526) );
  OAI21_X1 U5036 ( .B1(n5349), .B2(n4689), .A(n4685), .ZN(n5423) );
  NAND2_X1 U5037 ( .A1(n5284), .A2(n5283), .ZN(n6681) );
  XNOR2_X1 U5038 ( .A(n5298), .B(n5297), .ZN(n6750) );
  CLKBUF_X1 U5039 ( .A(n8692), .Z(n8717) );
  INV_X1 U5040 ( .A(n6612), .ZN(n6903) );
  INV_X2 U5041 ( .A(n9836), .ZN(n4474) );
  OAI211_X1 U5042 ( .C1(n6458), .C2(n6749), .A(n6457), .B(n6456), .ZN(n6612)
         );
  INV_X1 U5043 ( .A(n9914), .ZN(n5853) );
  NAND4_X1 U5044 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n6158)
         );
  CLKBUF_X1 U5045 ( .A(n5309), .Z(n5787) );
  INV_X2 U5046 ( .A(n5309), .ZN(n7668) );
  OR2_X1 U5047 ( .A1(n6224), .A2(n8795), .ZN(n6196) );
  NAND2_X1 U5048 ( .A1(n7869), .A2(n7689), .ZN(n9868) );
  OR2_X1 U5049 ( .A1(n5310), .A2(n5085), .ZN(n5086) );
  AND3_X1 U5050 ( .A1(n5143), .A2(n5142), .A3(n5141), .ZN(n9908) );
  INV_X2 U5051 ( .A(n5279), .ZN(n7680) );
  XNOR2_X1 U5052 ( .A(n6145), .B(n6144), .ZN(n6150) );
  AND2_X1 U5053 ( .A1(n4620), .A2(n4546), .ZN(n4589) );
  NAND2_X1 U5054 ( .A1(n8964), .A2(n6733), .ZN(n6572) );
  OR2_X1 U5055 ( .A1(n6148), .A2(n9456), .ZN(n6145) );
  XNOR2_X1 U5056 ( .A(n5837), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8964) );
  AND2_X1 U5057 ( .A1(n5823), .A2(n4537), .ZN(n6148) );
  XNOR2_X1 U5058 ( .A(n6194), .B(n6193), .ZN(n6733) );
  OR2_X1 U5059 ( .A1(n5080), .A2(n5077), .ZN(n4620) );
  AOI21_X1 U5060 ( .B1(n6187), .B2(P1_IR_REG_31__SCAN_IN), .A(n4851), .ZN(
        n4850) );
  NAND2_X1 U5061 ( .A1(n5738), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5748) );
  XNOR2_X1 U5062 ( .A(n5112), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U5063 ( .A1(n5095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5097) );
  XNOR2_X1 U5064 ( .A(n5105), .B(n5104), .ZN(n7669) );
  NAND2_X2 U5065 ( .A1(n7677), .A2(P1_U3084), .ZN(n9463) );
  NOR2_X1 U5066 ( .A1(n5904), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U5067 ( .A1(n4852), .A2(n6189), .ZN(n4851) );
  NOR2_X1 U5068 ( .A1(n5106), .A2(n5102), .ZN(n5103) );
  NAND2_X1 U5069 ( .A1(n5071), .A2(n5070), .ZN(n5501) );
  INV_X1 U5070 ( .A(n5164), .ZN(n5986) );
  NOR2_X1 U5071 ( .A1(n6188), .A2(n5004), .ZN(n4631) );
  AND2_X1 U5072 ( .A1(n5929), .A2(n5814), .ZN(n4824) );
  AND2_X1 U5073 ( .A1(n5813), .A2(n5002), .ZN(n5001) );
  NAND2_X1 U5074 ( .A1(n5907), .A2(n5005), .ZN(n5004) );
  AND2_X1 U5075 ( .A1(n5118), .A2(n5067), .ZN(n5184) );
  INV_X1 U5076 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5100) );
  INV_X1 U5077 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5747) );
  NOR2_X1 U5078 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5101) );
  INV_X1 U5079 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5104) );
  NOR2_X1 U5080 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5064) );
  NOR2_X1 U5081 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5063) );
  INV_X1 U5082 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5456) );
  INV_X1 U5083 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5183) );
  CLKBUF_X1 U5084 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9861) );
  INV_X1 U5085 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4709) );
  INV_X1 U5086 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8234) );
  NOR2_X2 U5087 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5118) );
  OR2_X2 U5088 ( .A1(n9518), .A2(n9431), .ZN(n7151) );
  XNOR2_X1 U5089 ( .A(n6190), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6256) );
  NOR2_X2 U5090 ( .A1(n8074), .A2(n5618), .ZN(n5639) );
  AOI22_X1 U5091 ( .A1(n5543), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6010), .B2(
        n8143), .ZN(n5187) );
  INV_X1 U5092 ( .A(n6749), .ZN(n4475) );
  XNOR2_X2 U5093 ( .A(n5097), .B(n5096), .ZN(n5794) );
  NAND2_X1 U5094 ( .A1(n5722), .A2(n5721), .ZN(n7637) );
  NAND2_X1 U5095 ( .A1(n5720), .A2(n5719), .ZN(n5722) );
  OR2_X1 U5096 ( .A1(n8476), .A2(n8262), .ZN(n7811) );
  NAND2_X1 U5097 ( .A1(n6555), .A2(n8064), .ZN(n7706) );
  OR2_X1 U5098 ( .A1(n9404), .A2(n9312), .ZN(n8860) );
  AND2_X1 U5099 ( .A1(n5845), .A2(n4783), .ZN(n4782) );
  INV_X1 U5100 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4783) );
  NAND2_X1 U5101 ( .A1(n5695), .A2(n5694), .ZN(n5720) );
  NOR3_X1 U5102 ( .A1(n8319), .A2(n8476), .A3(n4787), .ZN(n8266) );
  NAND2_X1 U5103 ( .A1(n6430), .A2(n4520), .ZN(n4573) );
  NAND2_X1 U5104 ( .A1(n4738), .A2(n4603), .ZN(n7745) );
  NOR2_X1 U5105 ( .A1(n7740), .A2(n7739), .ZN(n4738) );
  NAND2_X1 U5106 ( .A1(n4563), .A2(n4562), .ZN(n4561) );
  NOR2_X1 U5107 ( .A1(n8817), .A2(n8901), .ZN(n4562) );
  NAND2_X1 U5108 ( .A1(n8819), .A2(n8818), .ZN(n4563) );
  NAND2_X1 U5109 ( .A1(n4531), .A2(n7806), .ZN(n4623) );
  NOR2_X1 U5110 ( .A1(n9933), .A2(n8095), .ZN(n5039) );
  NAND2_X1 U5111 ( .A1(n5373), .A2(n5372), .ZN(n5398) );
  AND2_X1 U5112 ( .A1(n7714), .A2(n7871), .ZN(n7834) );
  OR2_X1 U5113 ( .A1(n8459), .A2(n7685), .ZN(n7835) );
  NAND2_X1 U5114 ( .A1(n8301), .A2(n8262), .ZN(n4816) );
  INV_X1 U5115 ( .A(n4795), .ZN(n4793) );
  OR2_X1 U5116 ( .A1(n8523), .A2(n9580), .ZN(n7784) );
  OR2_X1 U5117 ( .A1(n9568), .A2(n7649), .ZN(n7695) );
  OR2_X1 U5118 ( .A1(n7435), .A2(n7443), .ZN(n7766) );
  NOR2_X1 U5119 ( .A1(n7731), .A2(n5042), .ZN(n5041) );
  INV_X1 U5120 ( .A(n7729), .ZN(n5042) );
  NAND2_X1 U5121 ( .A1(n5103), .A2(n5104), .ZN(n5738) );
  NAND2_X1 U5122 ( .A1(n5071), .A2(n4900), .ZN(n5106) );
  AND2_X1 U5123 ( .A1(n4545), .A2(n5070), .ZN(n4900) );
  NOR2_X1 U5124 ( .A1(n9344), .A2(n9350), .ZN(n4708) );
  OR2_X1 U5125 ( .A1(n9356), .A2(n9166), .ZN(n8895) );
  AND2_X1 U5126 ( .A1(n9372), .A2(n9216), .ZN(n8928) );
  OR2_X1 U5127 ( .A1(n9372), .A2(n9216), .ZN(n8929) );
  AND2_X1 U5128 ( .A1(n9255), .A2(n9277), .ZN(n8934) );
  INV_X1 U5129 ( .A(n4992), .ZN(n4991) );
  NAND2_X1 U5130 ( .A1(n9628), .A2(n8761), .ZN(n4995) );
  NAND2_X1 U5131 ( .A1(n4473), .A2(n6733), .ZN(n6224) );
  XNOR2_X1 U5132 ( .A(n7675), .B(n7674), .ZN(n7673) );
  AND2_X1 U5133 ( .A1(n5580), .A2(n5566), .ZN(n5578) );
  XNOR2_X1 U5134 ( .A(n5537), .B(SI_18_), .ZN(n5534) );
  NAND2_X1 U5135 ( .A1(n4930), .A2(n5470), .ZN(n5497) );
  NAND2_X1 U5136 ( .A1(n4927), .A2(n4925), .ZN(n4930) );
  NOR2_X1 U5137 ( .A1(n5471), .A2(n4926), .ZN(n4925) );
  INV_X1 U5138 ( .A(n5451), .ZN(n4926) );
  AND2_X1 U5139 ( .A1(n5498), .A2(n5476), .ZN(n5496) );
  XNOR2_X1 U5140 ( .A(n5449), .B(SI_14_), .ZN(n5446) );
  NAND2_X1 U5141 ( .A1(n4931), .A2(n4935), .ZN(n5349) );
  INV_X1 U5142 ( .A(n4936), .ZN(n4935) );
  OAI21_X1 U5143 ( .B1(n5061), .B2(n4937), .A(n5058), .ZN(n4936) );
  NAND2_X1 U5144 ( .A1(n4710), .A2(n5115), .ZN(n5135) );
  INV_X1 U5145 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4914) );
  AND2_X1 U5146 ( .A1(n5558), .A2(n5559), .ZN(n7459) );
  NOR2_X1 U5147 ( .A1(n5796), .A2(n9886), .ZN(n5793) );
  NAND2_X2 U5148 ( .A1(n4890), .A2(n4889), .ZN(n7690) );
  INV_X1 U5149 ( .A(n5189), .ZN(n7665) );
  AND2_X1 U5150 ( .A1(n5689), .A2(n5688), .ZN(n8018) );
  AND3_X1 U5151 ( .A1(n5212), .A2(n5213), .A3(n4606), .ZN(n8064) );
  INV_X1 U5152 ( .A(n4607), .ZN(n4606) );
  AND2_X1 U5153 ( .A1(n5770), .A2(n5769), .ZN(n6074) );
  NAND2_X1 U5154 ( .A1(n8355), .A2(n8259), .ZN(n8327) );
  OR2_X1 U5155 ( .A1(n8513), .A2(n8254), .ZN(n7780) );
  NAND2_X1 U5156 ( .A1(n5508), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5549) );
  INV_X1 U5157 ( .A(n5509), .ZN(n5508) );
  NAND2_X1 U5158 ( .A1(n6713), .A2(n4822), .ZN(n6827) );
  AND2_X1 U5159 ( .A1(n6715), .A2(n6712), .ZN(n4822) );
  INV_X1 U5160 ( .A(n7851), .ZN(n6715) );
  NAND2_X1 U5161 ( .A1(n4567), .A2(n5858), .ZN(n6359) );
  INV_X1 U5162 ( .A(n9886), .ZN(n6008) );
  NAND2_X1 U5163 ( .A1(n5725), .A2(n5724), .ZN(n8471) );
  NAND2_X1 U5164 ( .A1(n5701), .A2(n5700), .ZN(n8476) );
  INV_X1 U5165 ( .A(n9973), .ZN(n9963) );
  INV_X1 U5166 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5076) );
  OR3_X1 U5167 ( .A1(n5951), .A2(n5844), .A3(n5843), .ZN(n5846) );
  NAND2_X1 U5168 ( .A1(n7029), .A2(n4521), .ZN(n7036) );
  NAND2_X1 U5169 ( .A1(n4840), .A2(n4838), .ZN(n8578) );
  AOI21_X1 U5170 ( .B1(n4841), .B2(n4477), .A(n4839), .ZN(n4838) );
  INV_X1 U5171 ( .A(n8580), .ZN(n4839) );
  OR2_X1 U5172 ( .A1(n7555), .A2(n8647), .ZN(n7579) );
  INV_X1 U5173 ( .A(n8721), .ZN(n7628) );
  INV_X1 U5174 ( .A(n6273), .ZN(n7624) );
  AND2_X1 U5175 ( .A1(n7585), .A2(n7584), .ZN(n9149) );
  NAND2_X1 U5176 ( .A1(n9162), .A2(n8779), .ZN(n4647) );
  OR2_X1 U5177 ( .A1(n9375), .A2(n9194), .ZN(n9190) );
  OAI22_X1 U5178 ( .A1(n9252), .A2(n7527), .B1(n9394), .B2(n9277), .ZN(n9247)
         );
  NOR2_X1 U5179 ( .A1(n9255), .A2(n8591), .ZN(n7527) );
  OAI21_X1 U5180 ( .B1(n9282), .B2(n7615), .A(n8849), .ZN(n9274) );
  OR2_X1 U5181 ( .A1(n9416), .A2(n9311), .ZN(n8845) );
  OR2_X1 U5182 ( .A1(n9322), .A2(n8630), .ZN(n5060) );
  OR2_X1 U5183 ( .A1(n9419), .A2(n9014), .ZN(n7401) );
  NAND2_X1 U5184 ( .A1(n7133), .A2(n7132), .ZN(n7212) );
  NAND2_X2 U5185 ( .A1(n6754), .A2(n7677), .ZN(n6749) );
  AND2_X1 U5186 ( .A1(n5642), .A2(n5626), .ZN(n5640) );
  INV_X1 U5187 ( .A(n8018), .ZN(n8305) );
  NAND2_X1 U5188 ( .A1(n8997), .A2(n4473), .ZN(n4973) );
  AOI21_X1 U5189 ( .B1(n8999), .B2(n9000), .A(n6733), .ZN(n4972) );
  AOI21_X1 U5190 ( .B1(n9002), .B2(n6733), .A(n9009), .ZN(n4969) );
  AND2_X1 U5191 ( .A1(n7755), .A2(n7756), .ZN(n4728) );
  NAND2_X1 U5192 ( .A1(n4612), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U5193 ( .A1(n7750), .A2(n7834), .ZN(n4737) );
  NAND2_X1 U5194 ( .A1(n4613), .A2(n7831), .ZN(n4612) );
  NAND2_X1 U5195 ( .A1(n4561), .A2(n4560), .ZN(n8823) );
  NAND2_X1 U5196 ( .A1(n8820), .A2(n8901), .ZN(n4560) );
  NOR3_X1 U5197 ( .A1(n4718), .A2(n7788), .A3(n7787), .ZN(n4717) );
  AOI21_X1 U5198 ( .B1(n7785), .B2(n7784), .A(n7783), .ZN(n4718) );
  AOI21_X1 U5199 ( .B1(n7779), .B2(n7786), .A(n7778), .ZN(n4619) );
  NOR2_X1 U5200 ( .A1(n4618), .A2(n4617), .ZN(n4616) );
  NAND2_X1 U5201 ( .A1(n7781), .A2(n7831), .ZN(n4617) );
  AND2_X1 U5202 ( .A1(n4622), .A2(n4621), .ZN(n4723) );
  AOI21_X1 U5203 ( .B1(n4484), .B2(n7806), .A(n7807), .ZN(n4621) );
  INV_X1 U5204 ( .A(n7636), .ZN(n4964) );
  OR2_X1 U5205 ( .A1(n7111), .A2(n7115), .ZN(n7755) );
  NAND2_X1 U5206 ( .A1(n6431), .A2(n5041), .ZN(n5040) );
  INV_X1 U5207 ( .A(n5039), .ZN(n5037) );
  INV_X1 U5208 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U5209 ( .A1(n4652), .A2(n4650), .ZN(n4649) );
  INV_X1 U5210 ( .A(n8818), .ZN(n4650) );
  INV_X1 U5211 ( .A(n5370), .ZN(n4688) );
  INV_X1 U5212 ( .A(n5399), .ZN(n4690) );
  INV_X1 U5213 ( .A(n5398), .ZN(n4686) );
  NAND2_X1 U5214 ( .A1(n5303), .A2(n5302), .ZN(n5325) );
  OR2_X1 U5215 ( .A1(n5298), .A2(n5297), .ZN(n5300) );
  NAND2_X1 U5216 ( .A1(n5276), .A2(n5275), .ZN(n5299) );
  OAI21_X1 U5217 ( .B1(n8284), .B2(n5019), .A(n7822), .ZN(n5018) );
  AOI21_X1 U5218 ( .B1(n7821), .B2(n7820), .A(n8273), .ZN(n4611) );
  INV_X1 U5219 ( .A(n7826), .ZN(n4609) );
  OR2_X1 U5220 ( .A1(n5306), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5380) );
  OR2_X1 U5221 ( .A1(n8482), .A2(n8305), .ZN(n4817) );
  INV_X1 U5222 ( .A(n5053), .ZN(n5050) );
  INV_X1 U5223 ( .A(n8335), .ZN(n5049) );
  AND2_X1 U5224 ( .A1(n5054), .A2(n7795), .ZN(n5052) );
  INV_X1 U5225 ( .A(n8356), .ZN(n5054) );
  NOR2_X1 U5226 ( .A1(n8362), .A2(n7794), .ZN(n5053) );
  NAND2_X1 U5227 ( .A1(n5583), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5607) );
  NOR2_X1 U5228 ( .A1(n4601), .A2(n8519), .ZN(n4599) );
  NAND2_X1 U5229 ( .A1(n8447), .A2(n4602), .ZN(n4601) );
  OR2_X1 U5230 ( .A1(n9609), .A2(n7163), .ZN(n7760) );
  NOR2_X1 U5231 ( .A1(n7111), .A2(n9615), .ZN(n4595) );
  AOI21_X1 U5232 ( .B1(n6832), .B2(n5029), .A(n5028), .ZN(n5027) );
  INV_X1 U5233 ( .A(n7756), .ZN(n5028) );
  INV_X1 U5234 ( .A(n7747), .ZN(n5029) );
  AND2_X1 U5235 ( .A1(n7755), .A2(n7757), .ZN(n6949) );
  OR2_X1 U5236 ( .A1(n6825), .A2(n6714), .ZN(n7747) );
  AND2_X1 U5237 ( .A1(n4576), .A2(n7846), .ZN(n4570) );
  NAND2_X1 U5238 ( .A1(n7731), .A2(n4575), .ZN(n4572) );
  NAND2_X1 U5239 ( .A1(n5861), .A2(n5862), .ZN(n4575) );
  NOR2_X1 U5240 ( .A1(n9926), .A2(n6555), .ZN(n4593) );
  INV_X1 U5241 ( .A(n7669), .ZN(n7871) );
  OR2_X1 U5242 ( .A1(n8491), .A2(n8031), .ZN(n8335) );
  NAND2_X1 U5243 ( .A1(n8235), .A2(n9599), .ZN(n9569) );
  NOR2_X1 U5244 ( .A1(n5074), .A2(n5073), .ZN(n5075) );
  INV_X1 U5245 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5739) );
  AND4_X1 U5246 ( .A1(n5066), .A2(n5065), .A3(n5064), .A4(n5063), .ZN(n5069)
         );
  AND4_X1 U5247 ( .A1(n5426), .A2(n5378), .A3(n5456), .A4(n5183), .ZN(n5068)
         );
  NOR2_X1 U5248 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5065) );
  INV_X1 U5249 ( .A(n8562), .ZN(n4861) );
  AOI21_X1 U5250 ( .B1(n4960), .B2(n8962), .A(n8964), .ZN(n8996) );
  NOR2_X1 U5251 ( .A1(n4961), .A2(n8991), .ZN(n4960) );
  OR2_X1 U5252 ( .A1(n8963), .A2(n4962), .ZN(n4961) );
  NAND2_X1 U5253 ( .A1(n4767), .A2(n4769), .ZN(n4766) );
  NAND2_X1 U5254 ( .A1(n6151), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4767) );
  NAND2_X1 U5255 ( .A1(n9466), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4769) );
  OR2_X1 U5256 ( .A1(n9362), .A2(n9149), .ZN(n8894) );
  AND2_X1 U5257 ( .A1(n9372), .A2(n8618), .ZN(n8893) );
  NOR2_X1 U5258 ( .A1(n4698), .A2(n9372), .ZN(n4697) );
  INV_X1 U5259 ( .A(n4699), .ZN(n4698) );
  NOR2_X1 U5260 ( .A1(n9375), .A2(n9380), .ZN(n4699) );
  OR2_X1 U5261 ( .A1(n9387), .A2(n9264), .ZN(n8886) );
  INV_X1 U5262 ( .A(n4639), .ZN(n4638) );
  OAI21_X1 U5263 ( .B1(n4641), .B2(n4640), .A(n8848), .ZN(n4639) );
  INV_X1 U5264 ( .A(n8845), .ZN(n4640) );
  INV_X1 U5265 ( .A(n4990), .ZN(n4989) );
  OAI21_X1 U5266 ( .B1(n4498), .B2(n4991), .A(n7394), .ZN(n4990) );
  NOR2_X1 U5267 ( .A1(n8762), .A2(n9634), .ZN(n4705) );
  AND2_X1 U5268 ( .A1(n4478), .A2(n8815), .ZN(n4652) );
  INV_X1 U5269 ( .A(n9130), .ZN(n4777) );
  NAND2_X1 U5270 ( .A1(n4774), .A2(n4773), .ZN(n4772) );
  NAND2_X1 U5271 ( .A1(n9130), .A2(n9128), .ZN(n4773) );
  OAI21_X1 U5272 ( .B1(n4778), .B2(n4775), .A(n4777), .ZN(n4774) );
  INV_X1 U5273 ( .A(n9128), .ZN(n4775) );
  INV_X1 U5274 ( .A(n5842), .ZN(n4780) );
  NAND2_X1 U5275 ( .A1(n4940), .A2(n4938), .ZN(n5693) );
  AOI21_X1 U5276 ( .B1(n4942), .B2(n4944), .A(n4939), .ZN(n4938) );
  INV_X1 U5277 ( .A(n4943), .ZN(n4942) );
  AND2_X1 U5278 ( .A1(n5694), .A2(n5678), .ZN(n5692) );
  NAND2_X1 U5279 ( .A1(n4941), .A2(n5642), .ZN(n5660) );
  NAND2_X1 U5280 ( .A1(n5540), .A2(n10158), .ZN(n5560) );
  NAND2_X1 U5281 ( .A1(n5539), .A2(n5538), .ZN(n5562) );
  INV_X1 U5282 ( .A(n5534), .ZN(n5535) );
  XNOR2_X1 U5283 ( .A(n5520), .B(SI_17_), .ZN(n5519) );
  NAND2_X1 U5284 ( .A1(n5425), .A2(n4928), .ZN(n4927) );
  NOR2_X1 U5285 ( .A1(n5447), .A2(n4929), .ZN(n4928) );
  INV_X1 U5286 ( .A(n5424), .ZN(n4929) );
  INV_X1 U5287 ( .A(n5446), .ZN(n5447) );
  INV_X1 U5288 ( .A(n5325), .ZN(n4937) );
  INV_X1 U5289 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U5290 ( .A1(n4671), .A2(n4670), .ZN(n4896) );
  AND2_X1 U5291 ( .A1(n4673), .A2(n4476), .ZN(n4897) );
  NAND2_X1 U5292 ( .A1(n7277), .A2(n4899), .ZN(n4895) );
  OAI21_X1 U5293 ( .B1(n5174), .B2(n4875), .A(n4873), .ZN(n6140) );
  AOI21_X1 U5294 ( .B1(n5195), .B2(n4874), .A(n4485), .ZN(n4873) );
  AND2_X1 U5295 ( .A1(n8068), .A2(n5194), .ZN(n5195) );
  NAND2_X1 U5296 ( .A1(n5267), .A2(n5266), .ZN(n5889) );
  AND2_X1 U5297 ( .A1(n5320), .A2(n4880), .ZN(n4879) );
  NAND2_X1 U5298 ( .A1(n6592), .A2(n4881), .ZN(n4880) );
  INV_X1 U5299 ( .A(n5268), .ZN(n4881) );
  INV_X1 U5300 ( .A(n6592), .ZN(n4882) );
  INV_X1 U5301 ( .A(n4887), .ZN(n4886) );
  OAI21_X1 U5302 ( .B1(n6699), .B2(n4888), .A(n6844), .ZN(n4887) );
  INV_X1 U5303 ( .A(n5364), .ZN(n4888) );
  AOI21_X1 U5304 ( .B1(n8036), .B2(n4669), .A(n5594), .ZN(n4668) );
  OR2_X1 U5305 ( .A1(n7466), .A2(n4666), .ZN(n4665) );
  NAND2_X1 U5306 ( .A1(n5345), .A2(n5344), .ZN(n6701) );
  AND2_X1 U5307 ( .A1(n5152), .A2(n5151), .ZN(n8085) );
  AND2_X1 U5308 ( .A1(n7835), .A2(n7826), .ZN(n7691) );
  AND2_X1 U5309 ( .A1(n8459), .A2(n7685), .ZN(n7692) );
  AND2_X1 U5310 ( .A1(n5712), .A2(n5711), .ZN(n8262) );
  AND4_X1 U5311 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n7114)
         );
  AND2_X1 U5312 ( .A1(n4814), .A2(n4813), .ZN(n4812) );
  NAND2_X1 U5313 ( .A1(n4815), .A2(n8261), .ZN(n4813) );
  NAND2_X1 U5314 ( .A1(n8302), .A2(n4816), .ZN(n4814) );
  AND2_X1 U5315 ( .A1(n4816), .A2(n4817), .ZN(n4815) );
  NAND2_X1 U5316 ( .A1(n8327), .A2(n8336), .ZN(n4803) );
  NOR2_X1 U5317 ( .A1(n8350), .A2(n8491), .ZN(n8349) );
  NAND2_X1 U5318 ( .A1(n5055), .A2(n5052), .ZN(n8334) );
  AND2_X1 U5319 ( .A1(n5637), .A2(n5636), .ZN(n8345) );
  NAND2_X1 U5320 ( .A1(n8379), .A2(n5053), .ZN(n5055) );
  AOI21_X1 U5321 ( .B1(n5022), .B2(n8415), .A(n4618), .ZN(n5021) );
  AOI21_X1 U5322 ( .B1(n9885), .B2(n10293), .A(n9891), .ZN(n8386) );
  AND2_X1 U5323 ( .A1(n8508), .A2(n8255), .ZN(n4800) );
  INV_X1 U5324 ( .A(n8416), .ZN(n5024) );
  OR2_X1 U5325 ( .A1(n4798), .A2(n4503), .ZN(n4795) );
  AND2_X1 U5326 ( .A1(n8253), .A2(n4511), .ZN(n4798) );
  NOR2_X1 U5327 ( .A1(n4503), .A2(n4797), .ZN(n4796) );
  INV_X1 U5328 ( .A(n8251), .ZN(n4797) );
  NOR2_X1 U5329 ( .A1(n9574), .A2(n5032), .ZN(n5031) );
  INV_X1 U5330 ( .A(n7771), .ZN(n5032) );
  AND2_X1 U5331 ( .A1(n9574), .A2(n8247), .ZN(n4591) );
  AND2_X1 U5332 ( .A1(n7772), .A2(n7771), .ZN(n7858) );
  INV_X1 U5333 ( .A(n7856), .ZN(n7433) );
  NAND2_X1 U5334 ( .A1(n5386), .A2(n5385), .ZN(n5412) );
  INV_X1 U5335 ( .A(n5388), .ZN(n5386) );
  NAND2_X1 U5336 ( .A1(n7113), .A2(n4509), .ZN(n7168) );
  OR2_X1 U5337 ( .A1(n5313), .A2(n5312), .ZN(n5334) );
  OR2_X1 U5338 ( .A1(n5334), .A2(n10102), .ZN(n5388) );
  NAND2_X1 U5339 ( .A1(n6685), .A2(n6684), .ZN(n6713) );
  INV_X1 U5340 ( .A(n7849), .ZN(n6684) );
  AOI21_X1 U5341 ( .B1(n5038), .B2(n5035), .A(n5034), .ZN(n5033) );
  INV_X1 U5342 ( .A(n5041), .ZN(n5035) );
  NAND2_X1 U5343 ( .A1(n4572), .A2(n4576), .ZN(n4574) );
  OAI21_X1 U5344 ( .B1(n6359), .B2(n5860), .A(n5859), .ZN(n6430) );
  OR2_X1 U5345 ( .A1(n7844), .A2(n5880), .ZN(n5859) );
  NOR2_X1 U5346 ( .A1(n9876), .A2(n5014), .ZN(n5013) );
  INV_X1 U5347 ( .A(n7696), .ZN(n5014) );
  NAND2_X1 U5348 ( .A1(n5854), .A2(n5853), .ZN(n7696) );
  INV_X1 U5349 ( .A(n5855), .ZN(n5854) );
  NAND2_X1 U5350 ( .A1(n6525), .A2(n7842), .ZN(n6524) );
  AND2_X1 U5351 ( .A1(n7696), .A2(n7719), .ZN(n7842) );
  OR2_X1 U5352 ( .A1(n6007), .A2(n6116), .ZN(n9581) );
  NAND2_X1 U5353 ( .A1(n6157), .A2(n6516), .ZN(n6533) );
  INV_X1 U5354 ( .A(n9581), .ZN(n9865) );
  AND2_X1 U5355 ( .A1(n4803), .A2(n4818), .ZN(n8310) );
  AND2_X1 U5356 ( .A1(n5075), .A2(n5043), .ZN(n5044) );
  AND2_X1 U5357 ( .A1(n5047), .A2(n5076), .ZN(n5043) );
  INV_X1 U5358 ( .A(n5501), .ZN(n5046) );
  OR2_X1 U5359 ( .A1(n5738), .A2(n5737), .ZN(n5743) );
  INV_X1 U5360 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5771) );
  INV_X1 U5361 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U5362 ( .A1(n5986), .A2(n5091), .ZN(n5115) );
  NOR2_X1 U5363 ( .A1(n4844), .A2(n4842), .ZN(n4841) );
  INV_X1 U5364 ( .A(n4493), .ZN(n4842) );
  OR2_X1 U5365 ( .A1(n6757), .A2(n6756), .ZN(n6987) );
  NAND2_X1 U5366 ( .A1(n7100), .A2(n7099), .ZN(n7101) );
  NAND2_X1 U5367 ( .A1(n7101), .A2(n7102), .ZN(n7310) );
  INV_X1 U5368 ( .A(n4866), .ZN(n6207) );
  AOI21_X1 U5369 ( .B1(n6318), .B2(n6583), .A(n6202), .ZN(n6203) );
  OAI21_X1 U5370 ( .B1(n7102), .B2(n4849), .A(n7346), .ZN(n4848) );
  AND2_X1 U5371 ( .A1(n8792), .A2(n8917), .ZN(n8991) );
  OR2_X1 U5372 ( .A1(n9703), .A2(n9702), .ZN(n4747) );
  AND2_X1 U5373 ( .A1(n4747), .A2(n4746), .ZN(n9716) );
  NAND2_X1 U5374 ( .A1(n9707), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4746) );
  OR2_X1 U5375 ( .A1(n9716), .A2(n9715), .ZN(n4745) );
  OR2_X1 U5376 ( .A1(n9072), .A2(n9071), .ZN(n4743) );
  INV_X1 U5377 ( .A(n4708), .ZN(n4706) );
  AND2_X1 U5378 ( .A1(n8914), .A2(n8987), .ZN(n9130) );
  NAND2_X1 U5379 ( .A1(n7610), .A2(n7621), .ZN(n9126) );
  OR2_X1 U5380 ( .A1(n9167), .A2(n9356), .ZN(n9154) );
  NAND2_X1 U5381 ( .A1(n4647), .A2(n4646), .ZN(n9152) );
  AND2_X1 U5382 ( .A1(n7620), .A2(n8880), .ZN(n4646) );
  NAND2_X1 U5383 ( .A1(n8895), .A2(n8881), .ZN(n9147) );
  OR2_X1 U5384 ( .A1(n9365), .A2(n9195), .ZN(n9161) );
  AND2_X1 U5385 ( .A1(n7597), .A2(n7596), .ZN(n9166) );
  NAND2_X1 U5386 ( .A1(n9161), .A2(n8877), .ZN(n9182) );
  NAND2_X1 U5387 ( .A1(n4644), .A2(n4518), .ZN(n9210) );
  NAND2_X1 U5388 ( .A1(n7551), .A2(n5059), .ZN(n9189) );
  OR2_X1 U5389 ( .A1(n9209), .A2(n9194), .ZN(n5059) );
  NAND2_X1 U5390 ( .A1(n9203), .A2(n7550), .ZN(n7551) );
  OR2_X1 U5391 ( .A1(n9375), .A2(n9230), .ZN(n7550) );
  AND2_X1 U5392 ( .A1(n8886), .A2(n8736), .ZN(n9246) );
  NAND2_X1 U5393 ( .A1(n4643), .A2(n7616), .ZN(n9237) );
  INV_X1 U5394 ( .A(n9260), .ZN(n4643) );
  AND2_X1 U5395 ( .A1(n7519), .A2(n7518), .ZN(n9255) );
  AND4_X1 U5396 ( .A1(n7414), .A2(n7413), .A3(n7412), .A4(n7411), .ZN(n9311)
         );
  NOR2_X1 U5397 ( .A1(n4784), .A2(n4642), .ZN(n4641) );
  INV_X1 U5398 ( .A(n8844), .ZN(n4784) );
  NOR2_X1 U5399 ( .A1(n9301), .A2(n9411), .ZN(n9300) );
  INV_X1 U5400 ( .A(n9283), .ZN(n8689) );
  OR2_X1 U5401 ( .A1(n7141), .A2(n7140), .ZN(n7223) );
  NAND2_X1 U5402 ( .A1(n4534), .A2(n4995), .ZN(n4992) );
  NAND2_X1 U5403 ( .A1(n7212), .A2(n8947), .ZN(n4994) );
  NOR2_X1 U5404 ( .A1(n7151), .A2(n9634), .ZN(n7232) );
  NAND2_X1 U5405 ( .A1(n9501), .A2(n8818), .ZN(n4653) );
  AND4_X1 U5406 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(n7357)
         );
  INV_X1 U5407 ( .A(n9017), .ZN(n8675) );
  NAND2_X1 U5408 ( .A1(n6889), .A2(n4497), .ZN(n6986) );
  NAND2_X1 U5409 ( .A1(n9769), .A2(n8972), .ZN(n6766) );
  AND4_X1 U5410 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(n7104)
         );
  NAND2_X1 U5411 ( .A1(n8800), .A2(n8801), .ZN(n8939) );
  AND4_X1 U5412 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(n7040)
         );
  NOR2_X1 U5413 ( .A1(n9781), .A2(n6798), .ZN(n6797) );
  NAND2_X1 U5414 ( .A1(n9770), .A2(n4513), .ZN(n9769) );
  NAND2_X1 U5415 ( .A1(n6658), .A2(n8971), .ZN(n9770) );
  NAND2_X1 U5416 ( .A1(n8732), .A2(n8731), .ZN(n9344) );
  NOR2_X1 U5417 ( .A1(n9247), .A2(n9246), .ZN(n9391) );
  INV_X1 U5418 ( .A(n9272), .ZN(n9398) );
  INV_X1 U5419 ( .A(n6882), .ZN(n9813) );
  AND2_X1 U5420 ( .A1(n6224), .A2(n6566), .ZN(n9524) );
  XNOR2_X1 U5421 ( .A(n4920), .B(n7679), .ZN(n8789) );
  OAI21_X1 U5422 ( .B1(n7673), .B2(n4921), .A(n7676), .ZN(n4920) );
  XNOR2_X1 U5423 ( .A(n5720), .B(n5719), .ZN(n7587) );
  XNOR2_X1 U5424 ( .A(n5835), .B(n5834), .ZN(n6017) );
  OAI21_X1 U5425 ( .B1(n5836), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5835) );
  XNOR2_X1 U5426 ( .A(n5840), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8795) );
  XNOR2_X1 U5427 ( .A(n5599), .B(n5595), .ZN(n7472) );
  NAND2_X1 U5428 ( .A1(n4949), .A2(n4953), .ZN(n5599) );
  OR2_X1 U5429 ( .A1(n5562), .A2(n4956), .ZN(n4949) );
  XNOR2_X1 U5430 ( .A(n4661), .B(n5519), .ZN(n7497) );
  NAND2_X1 U5431 ( .A1(n5499), .A2(n5498), .ZN(n4661) );
  NAND2_X1 U5432 ( .A1(n5425), .A2(n5424), .ZN(n5448) );
  NAND2_X1 U5433 ( .A1(n5003), .A2(n4869), .ZN(n5904) );
  NOR2_X1 U5434 ( .A1(n5913), .A2(n5004), .ZN(n5003) );
  NAND2_X1 U5435 ( .A1(n4684), .A2(n5370), .ZN(n5400) );
  NAND2_X1 U5436 ( .A1(n5349), .A2(n4691), .ZN(n4684) );
  NAND2_X1 U5437 ( .A1(n4922), .A2(n4924), .ZN(n5243) );
  AOI21_X1 U5438 ( .B1(n5220), .B2(n4483), .A(n4532), .ZN(n4924) );
  NAND2_X1 U5439 ( .A1(n4902), .A2(n4901), .ZN(n8021) );
  AOI21_X1 U5440 ( .B1(n4903), .B2(n4906), .A(n4550), .ZN(n4901) );
  NAND2_X1 U5441 ( .A1(n8046), .A2(n4903), .ZN(n4902) );
  INV_X1 U5442 ( .A(n4907), .ZN(n4906) );
  NAND2_X1 U5443 ( .A1(n4663), .A2(n8020), .ZN(n4662) );
  NAND2_X1 U5444 ( .A1(n4664), .A2(n8101), .ZN(n4663) );
  NAND2_X1 U5445 ( .A1(n4912), .A2(n4550), .ZN(n4664) );
  NAND2_X1 U5446 ( .A1(n5628), .A2(n5627), .ZN(n8497) );
  NAND2_X1 U5447 ( .A1(n5174), .A2(n6173), .ZN(n6174) );
  AND2_X1 U5448 ( .A1(n6349), .A2(n5114), .ZN(n6161) );
  AND3_X1 U5449 ( .A1(n5574), .A2(n5573), .A3(n5572), .ZN(n8254) );
  AND2_X1 U5450 ( .A1(n5614), .A2(n5613), .ZN(n8038) );
  AND2_X1 U5451 ( .A1(n5530), .A2(n5529), .ZN(n9580) );
  NAND2_X1 U5452 ( .A1(n5605), .A2(n5604), .ZN(n8504) );
  INV_X1 U5453 ( .A(n8051), .ZN(n8094) );
  NAND2_X1 U5454 ( .A1(n5525), .A2(n5524), .ZN(n8523) );
  AND2_X1 U5455 ( .A1(n8075), .A2(n9864), .ZN(n8106) );
  NAND2_X1 U5456 ( .A1(n5461), .A2(n5460), .ZN(n7435) );
  NAND2_X1 U5457 ( .A1(n4740), .A2(n4739), .ZN(n4565) );
  OR2_X1 U5458 ( .A1(n7873), .A2(n4741), .ZN(n4740) );
  OR2_X1 U5459 ( .A1(n6074), .A2(n5773), .ZN(n9886) );
  INV_X1 U5460 ( .A(n8064), .ZN(n9866) );
  NAND4_X1 U5461 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n8122)
         );
  OR2_X1 U5462 ( .A1(n5189), .A2(n6109), .ZN(n5191) );
  AOI21_X1 U5463 ( .B1(n8267), .B2(n8466), .A(n8266), .ZN(n8467) );
  AOI21_X1 U5464 ( .B1(n8278), .B2(n9868), .A(n8277), .ZN(n8469) );
  INV_X1 U5465 ( .A(n8276), .ZN(n8277) );
  INV_X1 U5466 ( .A(n4805), .ZN(n4804) );
  OAI211_X1 U5467 ( .C1(n8310), .C2(n4585), .A(n4582), .B(n4581), .ZN(n8480)
         );
  NAND2_X1 U5468 ( .A1(n8312), .A2(n8302), .ZN(n4585) );
  AOI21_X1 U5469 ( .B1(n4583), .B2(n8261), .A(n4528), .ZN(n4582) );
  NAND2_X1 U5470 ( .A1(n8310), .A2(n4583), .ZN(n4581) );
  AND2_X1 U5471 ( .A1(n8479), .A2(n8478), .ZN(n4587) );
  NAND2_X1 U5472 ( .A1(n5046), .A2(n5044), .ZN(n5095) );
  XNOR2_X1 U5473 ( .A(n5111), .B(n5110), .ZN(n7840) );
  AND4_X1 U5474 ( .A1(n7491), .A2(n7490), .A3(n7489), .A4(n7488), .ZN(n9312)
         );
  NAND2_X1 U5475 ( .A1(n7600), .A2(n7599), .ZN(n9350) );
  INV_X1 U5476 ( .A(n9014), .ZN(n8630) );
  NAND2_X1 U5477 ( .A1(n7405), .A2(n7404), .ZN(n9416) );
  NAND2_X1 U5478 ( .A1(n4857), .A2(n7911), .ZN(n4856) );
  NAND2_X1 U5479 ( .A1(n7055), .A2(n7054), .ZN(n9431) );
  INV_X1 U5480 ( .A(n9174), .ZN(n9362) );
  NAND2_X1 U5481 ( .A1(n7400), .A2(n7399), .ZN(n9419) );
  NAND2_X1 U5482 ( .A1(n7562), .A2(n7561), .ZN(n9216) );
  INV_X1 U5483 ( .A(n9264), .ZN(n9231) );
  INV_X1 U5484 ( .A(n7357), .ZN(n9016) );
  INV_X1 U5485 ( .A(n7104), .ZN(n9018) );
  OAI21_X1 U5486 ( .B1(n9109), .B2(n9108), .A(n4753), .ZN(n4752) );
  AOI21_X1 U5487 ( .B1(n9110), .B2(n9750), .A(n9742), .ZN(n4753) );
  AND2_X1 U5488 ( .A1(n5972), .A2(n6381), .ZN(n9750) );
  OR2_X1 U5489 ( .A1(n9354), .A2(n9335), .ZN(n4656) );
  INV_X1 U5490 ( .A(n9516), .ZN(n9321) );
  NAND2_X1 U5491 ( .A1(n9835), .A2(n6222), .ZN(n9790) );
  INV_X1 U5492 ( .A(n9139), .ZN(n9333) );
  NAND2_X1 U5493 ( .A1(n6242), .A2(n6241), .ZN(n9836) );
  INV_X1 U5494 ( .A(n8795), .ZN(n9003) );
  INV_X1 U5495 ( .A(n6191), .ZN(n6192) );
  NAND2_X1 U5496 ( .A1(n7705), .A2(n7706), .ZN(n4714) );
  NAND2_X1 U5497 ( .A1(n4713), .A2(n4711), .ZN(n7724) );
  NAND2_X1 U5498 ( .A1(n4712), .A2(n7831), .ZN(n4711) );
  NAND2_X1 U5499 ( .A1(n4714), .A2(n7834), .ZN(n4713) );
  NAND2_X1 U5500 ( .A1(n7720), .A2(n7722), .ZN(n4712) );
  NAND2_X1 U5501 ( .A1(n4605), .A2(n7735), .ZN(n4604) );
  OAI21_X1 U5502 ( .B1(n7749), .B2(n7748), .A(n4614), .ZN(n4613) );
  AND2_X1 U5503 ( .A1(n7747), .A2(n7756), .ZN(n4614) );
  AOI21_X1 U5504 ( .B1(n7745), .B2(n7744), .A(n7743), .ZN(n7749) );
  NAND2_X1 U5505 ( .A1(n4736), .A2(n4733), .ZN(n4732) );
  NOR2_X1 U5506 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  INV_X1 U5507 ( .A(n7751), .ZN(n4734) );
  OR2_X1 U5508 ( .A1(n7161), .A2(n7834), .ZN(n4731) );
  AOI21_X1 U5509 ( .B1(n4727), .B2(n7759), .A(n4726), .ZN(n4725) );
  NAND2_X1 U5510 ( .A1(n7758), .A2(n7834), .ZN(n4726) );
  NAND2_X1 U5511 ( .A1(n4736), .A2(n4728), .ZN(n4727) );
  NAND2_X1 U5512 ( .A1(n4729), .A2(n4724), .ZN(n7764) );
  INV_X1 U5513 ( .A(n4730), .ZN(n4729) );
  INV_X1 U5514 ( .A(n4725), .ZN(n4724) );
  AOI21_X1 U5515 ( .B1(n4732), .B2(n7754), .A(n4731), .ZN(n4730) );
  OAI21_X1 U5516 ( .B1(n4716), .B2(n4502), .A(n4715), .ZN(n7797) );
  NAND2_X1 U5517 ( .A1(n7794), .A2(n7831), .ZN(n4715) );
  NOR2_X1 U5518 ( .A1(n4717), .A2(n4524), .ZN(n4716) );
  NAND2_X1 U5519 ( .A1(n4615), .A2(n4517), .ZN(n7798) );
  OAI21_X1 U5520 ( .B1(n4619), .B2(n7788), .A(n4616), .ZN(n4615) );
  NOR2_X1 U5521 ( .A1(n5673), .A2(n4948), .ZN(n4947) );
  INV_X1 U5522 ( .A(n5658), .ZN(n4948) );
  INV_X1 U5523 ( .A(n4723), .ZN(n7816) );
  NAND2_X1 U5524 ( .A1(n4722), .A2(n4721), .ZN(n7818) );
  NAND2_X1 U5525 ( .A1(n7811), .A2(n7834), .ZN(n4721) );
  OAI21_X1 U5526 ( .B1(n4723), .B2(n8263), .A(n4525), .ZN(n4722) );
  NAND2_X1 U5527 ( .A1(n6195), .A2(n6572), .ZN(n6261) );
  OR2_X1 U5528 ( .A1(n9350), .A2(n9150), .ZN(n8896) );
  OAI21_X1 U5529 ( .B1(n7637), .B2(n4966), .A(n4963), .ZN(n7675) );
  AOI21_X1 U5530 ( .B1(n4965), .B2(n4964), .A(n4555), .ZN(n4963) );
  INV_X1 U5531 ( .A(n5642), .ZN(n4944) );
  OAI21_X1 U5532 ( .B1(n5640), .B2(n4944), .A(n4947), .ZN(n4943) );
  INV_X1 U5533 ( .A(n4945), .ZN(n4939) );
  AOI21_X1 U5534 ( .B1(n4947), .B2(n5659), .A(n4946), .ZN(n4945) );
  INV_X1 U5535 ( .A(n5672), .ZN(n4946) );
  AND2_X1 U5536 ( .A1(n4959), .A2(n5578), .ZN(n4958) );
  NAND2_X1 U5537 ( .A1(n5561), .A2(n5560), .ZN(n4959) );
  NOR2_X1 U5538 ( .A1(n4919), .A2(n4918), .ZN(n4917) );
  INV_X1 U5539 ( .A(n5498), .ZN(n4918) );
  INV_X1 U5540 ( .A(n5519), .ZN(n4919) );
  NOR2_X1 U5541 ( .A1(n4933), .A2(n4937), .ZN(n4932) );
  INV_X1 U5542 ( .A(n5299), .ZN(n4933) );
  INV_X1 U5543 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4658) );
  INV_X1 U5544 ( .A(n5735), .ZN(n5228) );
  NOR2_X1 U5545 ( .A1(n4507), .A2(n4872), .ZN(n4871) );
  INV_X1 U5546 ( .A(n5445), .ZN(n4872) );
  INV_X1 U5547 ( .A(n8036), .ZN(n4666) );
  INV_X1 U5548 ( .A(n5577), .ZN(n4669) );
  OR2_X1 U5549 ( .A1(n8044), .A2(n8043), .ZN(n4911) );
  OAI21_X1 U5550 ( .B1(n5189), .B2(n6552), .A(n5211), .ZN(n4607) );
  NAND2_X1 U5551 ( .A1(n4812), .A2(n8281), .ZN(n4811) );
  INV_X1 U5552 ( .A(n7780), .ZN(n5023) );
  OR2_X1 U5553 ( .A1(n8122), .A2(n9919), .ZN(n7705) );
  NAND2_X1 U5554 ( .A1(n7711), .A2(n7701), .ZN(n7839) );
  INV_X1 U5555 ( .A(n4817), .ZN(n4584) );
  NAND2_X1 U5556 ( .A1(n8349), .A2(n8260), .ZN(n8331) );
  NAND2_X1 U5557 ( .A1(n8426), .A2(n7652), .ZN(n8430) );
  NAND2_X1 U5558 ( .A1(n5040), .A2(n5038), .ZN(n6687) );
  NAND2_X1 U5559 ( .A1(n5040), .A2(n5037), .ZN(n5867) );
  OR2_X1 U5560 ( .A1(n5224), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U5561 ( .A1(n8560), .A2(n8562), .ZN(n8623) );
  NOR2_X1 U5562 ( .A1(n9058), .A2(n4749), .ZN(n5944) );
  AND2_X1 U5563 ( .A1(n9062), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4749) );
  OR2_X1 U5564 ( .A1(n9344), .A2(n7632), .ZN(n8914) );
  AND2_X1 U5565 ( .A1(n8871), .A2(n9190), .ZN(n8892) );
  NAND2_X1 U5566 ( .A1(n4705), .A2(n7396), .ZN(n4704) );
  OAI21_X1 U5567 ( .B1(n9501), .B2(n4651), .A(n4648), .ZN(n7219) );
  INV_X1 U5568 ( .A(n4652), .ZN(n4651) );
  AND2_X1 U5569 ( .A1(n4649), .A2(n8760), .ZN(n4648) );
  NAND2_X1 U5570 ( .A1(n8753), .A2(n8810), .ZN(n4760) );
  AND2_X1 U5571 ( .A1(n4504), .A2(n9820), .ZN(n4693) );
  NAND2_X1 U5572 ( .A1(n9022), .A2(n9808), .ZN(n8969) );
  NAND2_X1 U5573 ( .A1(n6808), .A2(n6607), .ZN(n8979) );
  OAI21_X1 U5574 ( .B1(n9177), .B2(n4979), .A(n4978), .ZN(n7610) );
  NAND2_X1 U5575 ( .A1(n4983), .A2(n4985), .ZN(n4979) );
  NAND2_X1 U5576 ( .A1(n4981), .A2(n4985), .ZN(n4978) );
  NAND2_X1 U5577 ( .A1(n9146), .A2(n9166), .ZN(n4985) );
  INV_X1 U5578 ( .A(SI_30_), .ZN(n4921) );
  AND2_X1 U5579 ( .A1(n5721), .A2(n5699), .ZN(n5719) );
  NAND2_X1 U5580 ( .A1(n4952), .A2(n4950), .ZN(n5621) );
  AND2_X1 U5581 ( .A1(n4951), .A2(n5598), .ZN(n4950) );
  AOI21_X1 U5582 ( .B1(n4958), .B2(n4955), .A(n4954), .ZN(n4953) );
  INV_X1 U5583 ( .A(n5580), .ZN(n4954) );
  INV_X1 U5584 ( .A(n5560), .ZN(n4955) );
  INV_X1 U5585 ( .A(n4958), .ZN(n4956) );
  INV_X1 U5586 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5817) );
  INV_X1 U5587 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5819) );
  INV_X1 U5588 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5818) );
  INV_X1 U5589 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5816) );
  INV_X1 U5590 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5942) );
  INV_X1 U5591 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U5592 ( .A1(n4854), .A2(n5817), .ZN(n4853) );
  INV_X1 U5593 ( .A(n6186), .ZN(n4854) );
  NAND2_X1 U5594 ( .A1(n5497), .A2(n5496), .ZN(n5499) );
  NAND2_X1 U5595 ( .A1(n5949), .A2(n5946), .ZN(n6186) );
  NAND2_X1 U5596 ( .A1(n5403), .A2(n5402), .ZN(n5424) );
  AOI21_X1 U5597 ( .B1(n4690), .B2(n4687), .A(n4686), .ZN(n4685) );
  NAND2_X1 U5598 ( .A1(n4690), .A2(n5370), .ZN(n4689) );
  NOR2_X1 U5599 ( .A1(n4691), .A2(n4688), .ZN(n4687) );
  INV_X1 U5600 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5005) );
  NOR2_X1 U5601 ( .A1(n5366), .A2(n4692), .ZN(n4691) );
  INV_X1 U5602 ( .A(n5348), .ZN(n4692) );
  INV_X1 U5603 ( .A(n5365), .ZN(n5366) );
  XNOR2_X1 U5604 ( .A(n5368), .B(SI_11_), .ZN(n5365) );
  NAND2_X1 U5605 ( .A1(n5274), .A2(n5273), .ZN(n5298) );
  AND2_X1 U5606 ( .A1(n5220), .A2(n5199), .ZN(n4923) );
  NOR2_X1 U5607 ( .A1(n4908), .A2(n5805), .ZN(n4907) );
  INV_X1 U5608 ( .A(n4909), .ZN(n4908) );
  AOI21_X1 U5609 ( .B1(n4905), .B2(n4907), .A(n4904), .ZN(n4903) );
  INV_X1 U5610 ( .A(n5691), .ZN(n4904) );
  INV_X1 U5611 ( .A(n4911), .ZN(n4905) );
  INV_X1 U5612 ( .A(n7085), .ZN(n4870) );
  NAND2_X1 U5613 ( .A1(n4877), .A2(n4876), .ZN(n5897) );
  AOI21_X1 U5614 ( .B1(n4879), .B2(n4882), .A(n4514), .ZN(n4876) );
  NAND2_X1 U5615 ( .A1(n5463), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5481) );
  INV_X1 U5616 ( .A(n5464), .ZN(n5463) );
  NAND2_X1 U5617 ( .A1(n4683), .A2(n4494), .ZN(n4675) );
  INV_X1 U5618 ( .A(n5654), .ZN(n4674) );
  NAND2_X1 U5619 ( .A1(n4894), .A2(n4892), .ZN(n7467) );
  AOI21_X1 U5620 ( .B1(n4896), .B2(n4897), .A(n4893), .ZN(n4892) );
  INV_X1 U5621 ( .A(n5559), .ZN(n4893) );
  NAND2_X1 U5622 ( .A1(n4910), .A2(n4907), .ZN(n4912) );
  NAND2_X1 U5623 ( .A1(n8044), .A2(n8043), .ZN(n4909) );
  AND2_X1 U5624 ( .A1(n7083), .A2(n5445), .ZN(n7288) );
  NAND2_X1 U5625 ( .A1(n5016), .A2(n5015), .ZN(n7670) );
  AOI21_X1 U5626 ( .B1(n5017), .B2(n5019), .A(n7824), .ZN(n5015) );
  INV_X1 U5627 ( .A(n5018), .ZN(n5017) );
  OAI21_X1 U5628 ( .B1(n4610), .B2(n4608), .A(n4529), .ZN(n7837) );
  OR2_X1 U5629 ( .A1(n7866), .A2(n4609), .ZN(n4608) );
  NOR2_X1 U5630 ( .A1(n4611), .A2(n7827), .ZN(n4610) );
  OR2_X1 U5631 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  INV_X1 U5632 ( .A(n7874), .ZN(n4741) );
  NOR4_X1 U5633 ( .A1(n7867), .A2(n7866), .A3(n8281), .A4(n7865), .ZN(n7868)
         );
  OR2_X1 U5634 ( .A1(n5380), .A2(n5379), .ZN(n5406) );
  NOR2_X1 U5635 ( .A1(n8462), .A2(n4787), .ZN(n4786) );
  NOR2_X1 U5636 ( .A1(n4811), .A2(n8326), .ZN(n4806) );
  OAI21_X1 U5637 ( .B1(n4811), .B2(n4818), .A(n4808), .ZN(n4805) );
  AOI21_X1 U5638 ( .B1(n4810), .B2(n4812), .A(n4809), .ZN(n4808) );
  NOR2_X1 U5639 ( .A1(n8471), .A2(n8304), .ZN(n4809) );
  NOR2_X1 U5640 ( .A1(n8284), .A2(n4815), .ZN(n4810) );
  OR2_X1 U5641 ( .A1(n8331), .A2(n8482), .ZN(n8319) );
  NOR2_X1 U5642 ( .A1(n8319), .A2(n8476), .ZN(n8297) );
  OR3_X1 U5643 ( .A1(n5682), .A2(n8047), .A3(n5681), .ZN(n5704) );
  OAI21_X1 U5644 ( .B1(n8379), .B2(n5051), .A(n5048), .ZN(n7654) );
  INV_X1 U5645 ( .A(n5052), .ZN(n5051) );
  AOI21_X1 U5646 ( .B1(n5052), .B2(n5050), .A(n5049), .ZN(n5048) );
  NOR2_X1 U5647 ( .A1(n8502), .A2(n4588), .ZN(n8357) );
  AND2_X1 U5648 ( .A1(n8497), .A2(n8258), .ZN(n4588) );
  NAND2_X1 U5649 ( .A1(n8357), .A2(n8356), .ZN(n8355) );
  OR2_X1 U5650 ( .A1(n8381), .A2(n8497), .ZN(n8350) );
  NAND2_X1 U5651 ( .A1(n8399), .A2(n8391), .ZN(n8381) );
  AOI21_X1 U5652 ( .B1(n4792), .B2(n4791), .A(n4535), .ZN(n4790) );
  INV_X1 U5653 ( .A(n4796), .ZN(n4791) );
  NOR2_X1 U5654 ( .A1(n8410), .A2(n8508), .ZN(n8399) );
  NAND2_X1 U5655 ( .A1(n8414), .A2(n4599), .ZN(n4598) );
  INV_X1 U5656 ( .A(n4599), .ZN(n4597) );
  AND2_X1 U5657 ( .A1(n7784), .A2(n7777), .ZN(n8449) );
  OR2_X1 U5658 ( .A1(n5481), .A2(n6973), .ZN(n5509) );
  AND2_X1 U5659 ( .A1(n7766), .A2(n7765), .ZN(n7856) );
  NAND2_X1 U5660 ( .A1(n6951), .A2(n4481), .ZN(n7267) );
  AND2_X1 U5661 ( .A1(n7168), .A2(n7167), .ZN(n7170) );
  NAND2_X1 U5662 ( .A1(n7170), .A2(n7169), .ZN(n7262) );
  INV_X1 U5663 ( .A(n5412), .ZN(n5410) );
  NAND2_X1 U5664 ( .A1(n6951), .A2(n4595), .ZN(n7171) );
  AND4_X1 U5665 ( .A1(n5438), .A2(n5437), .A3(n5436), .A4(n5435), .ZN(n7163)
         );
  AND2_X1 U5666 ( .A1(n6951), .A2(n9972), .ZN(n7121) );
  NAND2_X1 U5667 ( .A1(n5027), .A2(n5030), .ZN(n5026) );
  NAND2_X1 U5668 ( .A1(n6948), .A2(n4516), .ZN(n7113) );
  NAND2_X1 U5669 ( .A1(n6829), .A2(n5030), .ZN(n6948) );
  OR2_X1 U5670 ( .A1(n6726), .A2(n6825), .ZN(n6835) );
  NAND2_X1 U5671 ( .A1(n6830), .A2(n7747), .ZN(n6831) );
  NAND2_X1 U5672 ( .A1(n6831), .A2(n6832), .ZN(n6943) );
  INV_X1 U5673 ( .A(n7846), .ZN(n4571) );
  AOI21_X1 U5674 ( .B1(n4570), .B2(n4572), .A(n4527), .ZN(n4569) );
  NAND2_X1 U5675 ( .A1(n6693), .A2(n9948), .ZN(n6726) );
  AND2_X1 U5676 ( .A1(n7742), .A2(n7744), .ZN(n7849) );
  AND2_X1 U5677 ( .A1(n6360), .A2(n4490), .ZN(n5881) );
  NAND2_X1 U5678 ( .A1(n6360), .A2(n4593), .ZN(n6440) );
  INV_X1 U5679 ( .A(n5011), .ZN(n5010) );
  NAND2_X1 U5680 ( .A1(n7722), .A2(n7720), .ZN(n5012) );
  AND4_X1 U5681 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n8095)
         );
  NOR2_X1 U5682 ( .A1(n9870), .A2(n9869), .ZN(n6360) );
  NAND2_X1 U5683 ( .A1(n6360), .A2(n5880), .ZN(n6438) );
  NAND2_X1 U5684 ( .A1(n4568), .A2(n5857), .ZN(n9877) );
  NOR2_X1 U5685 ( .A1(n9618), .A2(n7871), .ZN(n6354) );
  NOR2_X1 U5686 ( .A1(n8302), .A2(n4584), .ZN(n4583) );
  NAND2_X1 U5687 ( .A1(n5644), .A2(n5643), .ZN(n8491) );
  NOR2_X1 U5688 ( .A1(n8367), .A2(n8366), .ZN(n8502) );
  OR2_X1 U5689 ( .A1(n4890), .A2(n9895), .ZN(n9971) );
  AND2_X1 U5690 ( .A1(n6535), .A2(n9894), .ZN(n9899) );
  OR2_X1 U5691 ( .A1(n9895), .A2(n7870), .ZN(n9973) );
  NAND2_X1 U5692 ( .A1(n4487), .A2(n5046), .ZN(n5079) );
  NAND2_X1 U5693 ( .A1(n4819), .A2(n5045), .ZN(n5093) );
  AND2_X1 U5694 ( .A1(n5075), .A2(n5047), .ZN(n5045) );
  INV_X1 U5695 ( .A(n5743), .ZN(n5740) );
  OR2_X1 U5696 ( .A1(n5107), .A2(n8542), .ZN(n5112) );
  NOR2_X1 U5697 ( .A1(n5501), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5099) );
  NOR2_X1 U5698 ( .A1(n5249), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5281) );
  INV_X1 U5699 ( .A(n6195), .ZN(n6204) );
  OR2_X1 U5700 ( .A1(n7590), .A2(n10138), .ZN(n7603) );
  NAND2_X1 U5701 ( .A1(n7906), .A2(n7905), .ZN(n8560) );
  NOR2_X1 U5702 ( .A1(n4862), .A2(n4859), .ZN(n4858) );
  NOR2_X1 U5703 ( .A1(n7905), .A2(n4861), .ZN(n4859) );
  INV_X1 U5704 ( .A(n7904), .ZN(n4862) );
  NAND2_X1 U5705 ( .A1(n4858), .A2(n4860), .ZN(n4857) );
  AND2_X1 U5706 ( .A1(n7905), .A2(n4861), .ZN(n4860) );
  INV_X1 U5707 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U5708 ( .A1(n6742), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U5709 ( .A1(n7531), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7544) );
  INV_X1 U5710 ( .A(n7532), .ZN(n7531) );
  OR2_X1 U5711 ( .A1(n7522), .A2(n8590), .ZN(n7532) );
  NAND2_X1 U5712 ( .A1(n7957), .A2(n7956), .ZN(n8666) );
  CLKBUF_X1 U5713 ( .A(n7893), .Z(n8011) );
  NAND2_X1 U5714 ( .A1(n9336), .A2(n9115), .ZN(n8962) );
  AND3_X1 U5715 ( .A1(n6447), .A2(n6446), .A3(n6449), .ZN(n4977) );
  OR2_X1 U5716 ( .A1(n6273), .A2(n9812), .ZN(n6447) );
  OR2_X1 U5717 ( .A1(n6273), .A2(n6272), .ZN(n6278) );
  NAND2_X1 U5718 ( .A1(n4766), .A2(n9461), .ZN(n4768) );
  OR2_X1 U5719 ( .A1(n6273), .A2(n6182), .ZN(n6185) );
  OR2_X1 U5720 ( .A1(n6069), .A2(n6068), .ZN(n4757) );
  AND2_X1 U5721 ( .A1(n4757), .A2(n4756), .ZN(n9645) );
  NAND2_X1 U5722 ( .A1(n6455), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4756) );
  AND2_X1 U5723 ( .A1(n4745), .A2(n4744), .ZN(n9730) );
  NAND2_X1 U5724 ( .A1(n9720), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4744) );
  NOR2_X1 U5725 ( .A1(n9045), .A2(n4750), .ZN(n9060) );
  AND2_X1 U5726 ( .A1(n9049), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4750) );
  NOR2_X1 U5727 ( .A1(n9060), .A2(n9059), .ZN(n9058) );
  XNOR2_X1 U5728 ( .A(n5944), .B(n6061), .ZN(n7010) );
  AND2_X1 U5729 ( .A1(n4743), .A2(n4742), .ZN(n9089) );
  NAND2_X1 U5730 ( .A1(n9091), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4742) );
  NOR2_X1 U5731 ( .A1(n9089), .A2(n9088), .ZN(n9099) );
  AND2_X1 U5732 ( .A1(n8791), .A2(n8790), .ZN(n8792) );
  NAND2_X1 U5733 ( .A1(n9119), .A2(n4708), .ZN(n4707) );
  NOR2_X1 U5734 ( .A1(n7621), .A2(n4779), .ZN(n4778) );
  INV_X1 U5735 ( .A(n8895), .ZN(n4779) );
  AOI21_X1 U5736 ( .B1(n9210), .B2(n8892), .A(n8893), .ZN(n9183) );
  AND2_X1 U5737 ( .A1(n9242), .A2(n4695), .ZN(n9178) );
  NOR2_X1 U5738 ( .A1(n9365), .A2(n4696), .ZN(n4695) );
  INV_X1 U5739 ( .A(n4697), .ZN(n4696) );
  AND2_X1 U5740 ( .A1(n7571), .A2(n7570), .ZN(n9195) );
  AND2_X1 U5741 ( .A1(n8930), .A2(n8929), .ZN(n9192) );
  NAND2_X1 U5742 ( .A1(n9242), .A2(n4699), .ZN(n9204) );
  OAI21_X1 U5743 ( .B1(n9247), .B2(n4997), .A(n4996), .ZN(n9203) );
  INV_X1 U5744 ( .A(n4998), .ZN(n4997) );
  AOI21_X1 U5745 ( .B1(n4998), .B2(n5000), .A(n4488), .ZN(n4996) );
  AOI21_X1 U5746 ( .B1(n9246), .B2(n4999), .A(n7538), .ZN(n4998) );
  AND2_X1 U5747 ( .A1(n9254), .A2(n8597), .ZN(n9242) );
  NAND2_X1 U5748 ( .A1(n9242), .A2(n9227), .ZN(n9221) );
  NAND2_X1 U5749 ( .A1(n9237), .A2(n7618), .ZN(n9238) );
  AND4_X1 U5750 ( .A1(n7513), .A2(n7512), .A3(n7511), .A4(n7510), .ZN(n9263)
         );
  NAND2_X1 U5751 ( .A1(n9273), .A2(n8863), .ZN(n9260) );
  NOR2_X1 U5752 ( .A1(n9268), .A2(n9394), .ZN(n9254) );
  NAND2_X1 U5753 ( .A1(n9274), .A2(n9275), .ZN(n9273) );
  OR2_X1 U5754 ( .A1(n9289), .A2(n9398), .ZN(n9268) );
  AND2_X1 U5755 ( .A1(n8861), .A2(n8863), .ZN(n9275) );
  NAND2_X1 U5756 ( .A1(n7476), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7508) );
  INV_X1 U5757 ( .A(n7486), .ZN(n7476) );
  NAND2_X1 U5758 ( .A1(n4636), .A2(n4634), .ZN(n9282) );
  AOI21_X1 U5759 ( .B1(n4638), .B2(n4640), .A(n4635), .ZN(n4634) );
  INV_X1 U5760 ( .A(n8843), .ZN(n4635) );
  AOI21_X1 U5761 ( .B1(n7496), .B2(n8956), .A(n7495), .ZN(n9299) );
  AND2_X1 U5762 ( .A1(n9416), .A2(n9329), .ZN(n7495) );
  NAND2_X1 U5763 ( .A1(n7407), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7421) );
  INV_X1 U5764 ( .A(n7409), .ZN(n7407) );
  OR2_X1 U5765 ( .A1(n9316), .A2(n9416), .ZN(n9301) );
  AOI21_X1 U5766 ( .B1(n4989), .B2(n4991), .A(n4526), .ZN(n4986) );
  NAND2_X1 U5767 ( .A1(n7221), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7251) );
  AOI21_X1 U5768 ( .B1(n7248), .B2(n8950), .A(n8743), .ZN(n7249) );
  NOR2_X1 U5769 ( .A1(n7151), .A2(n4703), .ZN(n7243) );
  INV_X1 U5770 ( .A(n4705), .ZN(n4703) );
  NAND2_X1 U5771 ( .A1(n4653), .A2(n4652), .ZN(n7218) );
  INV_X1 U5772 ( .A(n7058), .ZN(n7056) );
  OR2_X1 U5773 ( .A1(n6987), .A2(n7302), .ZN(n7058) );
  OAI21_X1 U5774 ( .B1(n6889), .B2(n5008), .A(n5006), .ZN(n9499) );
  INV_X1 U5775 ( .A(n5007), .ZN(n5006) );
  OAI22_X1 U5776 ( .A1(n4497), .A2(n5008), .B1(n7096), .B2(n9506), .ZN(n5007)
         );
  NAND2_X1 U5777 ( .A1(n4533), .A2(n6985), .ZN(n5008) );
  AND3_X1 U5778 ( .A1(n6797), .A2(n4693), .A3(n9829), .ZN(n9519) );
  NAND2_X1 U5779 ( .A1(n4627), .A2(n4761), .ZN(n7079) );
  AOI21_X1 U5780 ( .B1(n4764), .B2(n8810), .A(n4762), .ZN(n4761) );
  NAND2_X1 U5781 ( .A1(n6766), .A2(n4628), .ZN(n4627) );
  NOR2_X1 U5782 ( .A1(n4760), .A2(n8939), .ZN(n4628) );
  NAND2_X1 U5783 ( .A1(n4763), .A2(n8801), .ZN(n8804) );
  NAND2_X1 U5784 ( .A1(n6766), .A2(n4765), .ZN(n4763) );
  NOR2_X1 U5785 ( .A1(n8939), .A2(n4759), .ZN(n4765) );
  INV_X1 U5786 ( .A(n8753), .ZN(n4759) );
  NAND2_X1 U5787 ( .A1(n6797), .A2(n9813), .ZN(n6892) );
  AND2_X1 U5788 ( .A1(n8941), .A2(n6644), .ZN(n4974) );
  NAND2_X1 U5789 ( .A1(n9783), .A2(n9808), .ZN(n9781) );
  AND4_X1 U5790 ( .A1(n6485), .A2(n6484), .A3(n6483), .A4(n6482), .ZN(n9772)
         );
  AND2_X1 U5791 ( .A1(n6611), .A2(n6903), .ZN(n9783) );
  INV_X1 U5792 ( .A(n9022), .ZN(n6633) );
  NAND2_X1 U5793 ( .A1(n8979), .A2(n8937), .ZN(n6658) );
  AND4_X1 U5794 ( .A1(n6342), .A2(n6341), .A3(n6340), .A4(n6339), .ZN(n9774)
         );
  INV_X1 U5795 ( .A(n6235), .ZN(n4867) );
  INV_X1 U5796 ( .A(n9112), .ZN(n9137) );
  AOI21_X1 U5797 ( .B1(n9134), .B2(n9776), .A(n9133), .ZN(n9347) );
  NAND2_X1 U5798 ( .A1(n4777), .A2(n9128), .ZN(n4776) );
  OAI211_X1 U5799 ( .C1(n6642), .C2(n6749), .A(n6641), .B(n6640), .ZN(n6798)
         );
  INV_X1 U5800 ( .A(n9782), .ZN(n9830) );
  OR2_X1 U5801 ( .A1(n9792), .A2(n6221), .ZN(n6559) );
  INV_X1 U5802 ( .A(n6787), .ZN(n9835) );
  AND2_X1 U5803 ( .A1(n9003), .A2(n8992), .ZN(n6566) );
  INV_X1 U5804 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4781) );
  XNOR2_X1 U5805 ( .A(n7658), .B(n7657), .ZN(n8729) );
  NAND2_X1 U5806 ( .A1(n4967), .A2(n7640), .ZN(n7658) );
  XNOR2_X1 U5807 ( .A(n7637), .B(n7636), .ZN(n7598) );
  INV_X1 U5808 ( .A(n5826), .ZN(n5830) );
  OAI21_X1 U5809 ( .B1(n5660), .B2(n5659), .A(n5658), .ZN(n5674) );
  INV_X1 U5810 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U5811 ( .A1(n4957), .A2(n5560), .ZN(n5579) );
  NAND2_X1 U5812 ( .A1(n4853), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U5813 ( .A1(n4927), .A2(n5451), .ZN(n5472) );
  INV_X1 U5814 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5907) );
  NOR2_X1 U5815 ( .A1(n5913), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U5816 ( .A1(n5349), .A2(n5348), .ZN(n5367) );
  INV_X1 U5817 ( .A(n4934), .ZN(n5347) );
  AOI21_X1 U5818 ( .B1(n5324), .B2(n5061), .A(n4937), .ZN(n4934) );
  INV_X1 U5819 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5002) );
  NAND2_X1 U5820 ( .A1(n5180), .A2(n5179), .ZN(n5200) );
  XNOR2_X1 U5821 ( .A(n5135), .B(n5116), .ZN(n5134) );
  XNOR2_X1 U5822 ( .A(n4748), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U5823 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4748) );
  AND2_X1 U5824 ( .A1(n5164), .A2(SI_0_), .ZN(n6198) );
  AND4_X1 U5825 ( .A1(n5292), .A2(n5291), .A3(n5290), .A4(n5289), .ZN(n6620)
         );
  AND4_X1 U5826 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .ZN(n6828)
         );
  AND4_X1 U5827 ( .A1(n5318), .A2(n5317), .A3(n5316), .A4(n5315), .ZN(n6680)
         );
  OAI21_X1 U5828 ( .B1(n7277), .B2(n4897), .A(n4896), .ZN(n7458) );
  NAND2_X1 U5829 ( .A1(n4895), .A2(n4898), .ZN(n7460) );
  INV_X1 U5830 ( .A(n4897), .ZN(n4898) );
  AND2_X1 U5831 ( .A1(n5793), .A2(n4890), .ZN(n8075) );
  AND2_X1 U5832 ( .A1(n8268), .A2(n5728), .ZN(n8290) );
  OAI21_X1 U5833 ( .B1(n4566), .B2(n7466), .A(n5577), .ZN(n8037) );
  NAND2_X1 U5834 ( .A1(n6703), .A2(n5364), .ZN(n6845) );
  AND2_X1 U5835 ( .A1(n5480), .A2(n5479), .ZN(n9599) );
  AND3_X1 U5836 ( .A1(n5513), .A2(n5512), .A3(n5511), .ZN(n7649) );
  AND4_X1 U5837 ( .A1(n5469), .A2(n5468), .A3(n5467), .A4(n5466), .ZN(n7443)
         );
  NAND2_X1 U5838 ( .A1(n5219), .A2(n5218), .ZN(n8100) );
  NAND2_X1 U5839 ( .A1(n6174), .A2(n5195), .ZN(n8066) );
  NAND2_X1 U5840 ( .A1(n5889), .A2(n5268), .ZN(n4878) );
  OAI21_X1 U5841 ( .B1(n5889), .B2(n4882), .A(n4879), .ZN(n6626) );
  INV_X1 U5842 ( .A(n6533), .ZN(n4891) );
  AND2_X1 U5843 ( .A1(n5590), .A2(n5589), .ZN(n8419) );
  AOI21_X1 U5844 ( .B1(n4886), .B2(n4888), .A(n4884), .ZN(n4883) );
  INV_X1 U5845 ( .A(n6843), .ZN(n4884) );
  AND4_X1 U5846 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n6714)
         );
  AND4_X1 U5847 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n7115)
         );
  INV_X1 U5848 ( .A(n8084), .ZN(n8096) );
  NAND2_X1 U5849 ( .A1(n5360), .A2(n6699), .ZN(n6703) );
  AND2_X1 U5850 ( .A1(n8075), .A2(n9865), .ZN(n8084) );
  OAI21_X1 U5851 ( .B1(n7277), .B2(n7276), .A(n5518), .ZN(n7336) );
  INV_X1 U5852 ( .A(n4912), .ZN(n8017) );
  NAND2_X1 U5853 ( .A1(n4910), .A2(n4909), .ZN(n5804) );
  NAND2_X1 U5854 ( .A1(n5775), .A2(n9871), .ZN(n8098) );
  NAND2_X1 U5855 ( .A1(n7690), .A2(n7689), .ZN(n7875) );
  OR2_X1 U5856 ( .A1(n5310), .A2(n5144), .ZN(n5147) );
  CLKBUF_X1 U5857 ( .A(n6495), .Z(n8124) );
  INV_X1 U5858 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10102) );
  AND2_X1 U5859 ( .A1(n9851), .A2(n6116), .ZN(n9850) );
  NAND2_X1 U5860 ( .A1(n7683), .A2(n7682), .ZN(n8459) );
  XNOR2_X1 U5861 ( .A(n8240), .B(n8459), .ZN(n8461) );
  OR2_X1 U5862 ( .A1(n5727), .A2(n5726), .ZN(n8268) );
  AND2_X1 U5863 ( .A1(n8289), .A2(n8288), .ZN(n8474) );
  NAND2_X1 U5864 ( .A1(n4807), .A2(n4812), .ZN(n8282) );
  NAND2_X1 U5865 ( .A1(n4803), .A2(n4802), .ZN(n4807) );
  AND2_X1 U5866 ( .A1(n4815), .A2(n4818), .ZN(n4802) );
  NAND2_X1 U5867 ( .A1(n5055), .A2(n7795), .ZN(n8344) );
  NAND2_X1 U5868 ( .A1(n8379), .A2(n7793), .ZN(n8363) );
  INV_X1 U5869 ( .A(n8504), .ZN(n8391) );
  NAND2_X1 U5870 ( .A1(n8417), .A2(n7780), .ZN(n8395) );
  NAND2_X1 U5871 ( .A1(n4794), .A2(n4795), .ZN(n8409) );
  NAND2_X1 U5872 ( .A1(n8443), .A2(n4796), .ZN(n4794) );
  AND2_X1 U5873 ( .A1(n4799), .A2(n4511), .ZN(n8425) );
  NAND2_X1 U5874 ( .A1(n8443), .A2(n8251), .ZN(n4799) );
  NAND2_X1 U5875 ( .A1(n7648), .A2(n7771), .ZN(n9575) );
  AND2_X1 U5876 ( .A1(n8248), .A2(n8247), .ZN(n9566) );
  NAND2_X1 U5877 ( .A1(n7437), .A2(n7436), .ZN(n7439) );
  INV_X1 U5878 ( .A(n9599), .ZN(n8246) );
  NAND2_X1 U5879 ( .A1(n6713), .A2(n6712), .ZN(n6716) );
  NAND2_X1 U5880 ( .A1(n5863), .A2(n7846), .ZN(n6682) );
  NAND2_X1 U5881 ( .A1(n4573), .A2(n4574), .ZN(n5863) );
  OAI21_X1 U5882 ( .B1(n6430), .B2(n5862), .A(n5861), .ZN(n6420) );
  NAND2_X1 U5883 ( .A1(n5009), .A2(n7720), .ZN(n6363) );
  NAND2_X1 U5884 ( .A1(n5013), .A2(n6524), .ZN(n5009) );
  NAND2_X1 U5885 ( .A1(n6524), .A2(n7696), .ZN(n9863) );
  NAND2_X1 U5886 ( .A1(n9591), .A2(n9571), .ZN(n9881) );
  OR2_X1 U5887 ( .A1(n5884), .A2(n5883), .ZN(n9873) );
  NAND2_X1 U5888 ( .A1(n6008), .A2(n6354), .ZN(n9871) );
  INV_X1 U5889 ( .A(n9881), .ZN(n8440) );
  INV_X1 U5890 ( .A(n9873), .ZN(n8456) );
  AND2_X2 U5891 ( .A1(n6370), .A2(n6369), .ZN(n9995) );
  AOI22_X1 U5892 ( .A1(n8467), .A2(n9963), .B1(n8466), .B2(n9962), .ZN(n8468)
         );
  AND2_X1 U5893 ( .A1(n6009), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9892) );
  AND2_X1 U5894 ( .A1(n5044), .A2(n4821), .ZN(n4820) );
  AND2_X1 U5895 ( .A1(n5096), .A2(n5077), .ZN(n4821) );
  INV_X1 U5896 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8542) );
  XNOR2_X1 U5897 ( .A(n5752), .B(n5751), .ZN(n7092) );
  INV_X1 U5898 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10101) );
  INV_X1 U5899 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6399) );
  INV_X1 U5900 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6181) );
  INV_X1 U5901 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10243) );
  INV_X1 U5902 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6058) );
  INV_X1 U5903 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6035) );
  INV_X1 U5904 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6027) );
  INV_X1 U5905 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6015) );
  INV_X1 U5906 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5998) );
  INV_X1 U5907 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5994) );
  INV_X1 U5908 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10179) );
  NAND2_X1 U5909 ( .A1(n4660), .A2(n5090), .ZN(n5092) );
  NAND2_X1 U5910 ( .A1(n4659), .A2(SI_0_), .ZN(n4660) );
  NAND2_X1 U5911 ( .A1(n7589), .A2(n7588), .ZN(n9356) );
  NAND2_X1 U5912 ( .A1(n7587), .A2(n4475), .ZN(n7589) );
  NAND2_X1 U5913 ( .A1(n7242), .A2(n7241), .ZN(n9426) );
  NAND2_X1 U5914 ( .A1(n7963), .A2(n7966), .ZN(n8642) );
  NAND2_X1 U5915 ( .A1(n7541), .A2(n7540), .ZN(n9375) );
  NAND2_X1 U5916 ( .A1(n7310), .A2(n7309), .ZN(n7347) );
  NAND2_X1 U5917 ( .A1(n4837), .A2(n4477), .ZN(n8579) );
  OR2_X1 U5918 ( .A1(n7920), .A2(n4841), .ZN(n4837) );
  INV_X1 U5919 ( .A(n4834), .ZN(n4828) );
  NAND2_X1 U5920 ( .A1(n4833), .A2(n4832), .ZN(n4831) );
  INV_X1 U5921 ( .A(n8552), .ZN(n4832) );
  INV_X1 U5922 ( .A(n8554), .ZN(n4833) );
  NAND2_X1 U5923 ( .A1(n4836), .A2(n4835), .ZN(n4834) );
  INV_X1 U5924 ( .A(n8551), .ZN(n4835) );
  NAND2_X1 U5925 ( .A1(n8554), .A2(n8552), .ZN(n4836) );
  AND2_X1 U5926 ( .A1(n8009), .A2(n8645), .ZN(n4830) );
  NAND2_X1 U5927 ( .A1(n4826), .A2(n4500), .ZN(n4825) );
  INV_X1 U5928 ( .A(n4831), .ZN(n4826) );
  NAND2_X1 U5929 ( .A1(n4865), .A2(n6331), .ZN(n6268) );
  AND4_X1 U5930 ( .A1(n7526), .A2(n7525), .A3(n7524), .A4(n7523), .ZN(n8591)
         );
  NAND2_X1 U5931 ( .A1(n7499), .A2(n7498), .ZN(n9411) );
  INV_X1 U5932 ( .A(n9255), .ZN(n9394) );
  INV_X1 U5933 ( .A(n9328), .ZN(n8709) );
  INV_X1 U5934 ( .A(n4848), .ZN(n4847) );
  AND2_X1 U5935 ( .A1(n7920), .A2(n7919), .ZN(n4845) );
  NAND2_X1 U5936 ( .A1(n7494), .A2(n7493), .ZN(n9404) );
  OAI21_X1 U5937 ( .B1(n6223), .B2(n9784), .A(n9790), .ZN(n8692) );
  INV_X1 U5938 ( .A(n9149), .ZN(n9184) );
  INV_X1 U5939 ( .A(n9263), .ZN(n9284) );
  INV_X1 U5940 ( .A(n9311), .ZN(n9329) );
  INV_X1 U5941 ( .A(n9772), .ZN(n9021) );
  NAND2_X1 U5942 ( .A1(n4977), .A2(n6448), .ZN(n9022) );
  CLKBUF_X1 U5943 ( .A(n6235), .Z(n9026) );
  NAND2_X1 U5944 ( .A1(n6052), .A2(n6051), .ZN(n6050) );
  AND2_X1 U5945 ( .A1(n6388), .A2(n4758), .ZN(n6069) );
  NAND2_X1 U5946 ( .A1(n6391), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4758) );
  INV_X1 U5947 ( .A(n4757), .ZN(n6067) );
  INV_X1 U5948 ( .A(n4747), .ZN(n9701) );
  INV_X1 U5949 ( .A(n4745), .ZN(n9714) );
  NOR2_X1 U5950 ( .A1(n9068), .A2(n9069), .ZN(n9072) );
  INV_X1 U5951 ( .A(n4743), .ZN(n9086) );
  AND2_X1 U5952 ( .A1(n5977), .A2(n6374), .ZN(n9742) );
  INV_X1 U5953 ( .A(n8792), .ZN(n9336) );
  NAND2_X1 U5954 ( .A1(n8728), .A2(n8727), .ZN(n9340) );
  NAND2_X1 U5955 ( .A1(n4647), .A2(n8880), .ZN(n9148) );
  NAND2_X1 U5956 ( .A1(n4980), .A2(n4983), .ZN(n9145) );
  AND2_X1 U5957 ( .A1(n7574), .A2(n7573), .ZN(n9174) );
  NAND2_X1 U5958 ( .A1(n9177), .A2(n9182), .ZN(n4984) );
  NAND2_X1 U5959 ( .A1(n7554), .A2(n7553), .ZN(n9372) );
  NAND2_X1 U5960 ( .A1(n4644), .A2(n8931), .ZN(n9212) );
  NOR2_X1 U5961 ( .A1(n9391), .A2(n5000), .ZN(n9220) );
  NAND2_X1 U5962 ( .A1(n7475), .A2(n7474), .ZN(n9387) );
  AND2_X1 U5963 ( .A1(n7504), .A2(n7503), .ZN(n9272) );
  NAND2_X1 U5964 ( .A1(n4637), .A2(n8845), .ZN(n9309) );
  NAND2_X1 U5965 ( .A1(n9326), .A2(n4641), .ZN(n4637) );
  NAND2_X1 U5966 ( .A1(n9326), .A2(n8838), .ZN(n7614) );
  NAND2_X1 U5967 ( .A1(n4988), .A2(n4992), .ZN(n7395) );
  NAND2_X1 U5968 ( .A1(n7212), .A2(n4498), .ZN(n4988) );
  INV_X1 U5969 ( .A(n7211), .ZN(n4993) );
  NAND2_X1 U5970 ( .A1(n7136), .A2(n7135), .ZN(n9634) );
  NAND2_X1 U5971 ( .A1(n4653), .A2(n8815), .ZN(n7137) );
  NAND2_X1 U5972 ( .A1(n6986), .A2(n6985), .ZN(n7047) );
  OR2_X1 U5973 ( .A1(n7157), .A2(n9830), .ZN(n9139) );
  AND2_X1 U5974 ( .A1(n6889), .A2(n6740), .ZN(n6755) );
  NAND2_X1 U5975 ( .A1(n6766), .A2(n8753), .ZN(n6893) );
  OAI211_X1 U5976 ( .C1(n6656), .C2(n6749), .A(n6655), .B(n6654), .ZN(n6882)
         );
  BUF_X1 U5977 ( .A(n6279), .Z(n6599) );
  AND2_X1 U5978 ( .A1(n9786), .A2(n6567), .ZN(n9516) );
  INV_X1 U5979 ( .A(n7634), .ZN(n9353) );
  AND2_X1 U5980 ( .A1(n6195), .A2(n6016), .ZN(n9793) );
  AND2_X1 U5981 ( .A1(n6210), .A2(n6209), .ZN(n9455) );
  INV_X1 U5982 ( .A(n6150), .ZN(n9461) );
  INV_X1 U5983 ( .A(n6374), .ZN(n7456) );
  INV_X1 U5984 ( .A(n8964), .ZN(n8992) );
  INV_X1 U5985 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6397) );
  INV_X1 U5986 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6179) );
  INV_X1 U5987 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6059) );
  INV_X1 U5988 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5999) );
  INV_X1 U5989 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U5990 ( .A(n4720), .B(n4719), .ZN(n6642) );
  INV_X1 U5991 ( .A(n5220), .ZN(n4719) );
  AOI21_X1 U5992 ( .B1(n5200), .B2(n5199), .A(n4483), .ZN(n4720) );
  NOR2_X1 U5993 ( .A1(n9558), .A2(n10406), .ZN(n10023) );
  AOI21_X1 U5994 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10021), .ZN(n10020) );
  NOR2_X1 U5995 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  NAND2_X1 U5996 ( .A1(n4683), .A2(n4494), .ZN(n4678) );
  NAND2_X1 U5997 ( .A1(n4662), .A2(n8021), .ZN(n8026) );
  AOI21_X1 U5998 ( .B1(n7876), .B2(n7875), .A(n4565), .ZN(n7883) );
  NAND2_X1 U5999 ( .A1(n4578), .A2(n4587), .ZN(n8532) );
  NAND2_X1 U6000 ( .A1(n4580), .A2(n9978), .ZN(n4578) );
  INV_X1 U6001 ( .A(n8480), .ZN(n4580) );
  OAI211_X1 U6002 ( .C1(n8480), .C2(n4558), .A(n4586), .B(n4577), .ZN(P2_U3515) );
  NAND2_X1 U6003 ( .A1(n4579), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n4586) );
  OR2_X1 U6004 ( .A1(n4587), .A2(n4579), .ZN(n4577) );
  NOR2_X1 U6005 ( .A1(n5975), .A2(P1_U3084), .ZN(P1_U4006) );
  NAND2_X1 U6006 ( .A1(n4970), .A2(n4969), .ZN(n4968) );
  OAI211_X1 U6007 ( .C1(n9111), .C2(n9785), .A(n4754), .B(n4751), .ZN(P1_U3260) );
  NOR2_X1 U6008 ( .A1(n4755), .A2(n4559), .ZN(n4754) );
  NAND2_X1 U6009 ( .A1(n4752), .A2(n9785), .ZN(n4751) );
  AND2_X1 U6010 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  AOI21_X1 U6011 ( .B1(n9351), .B2(n9333), .A(n7635), .ZN(n4655) );
  OR2_X1 U6012 ( .A1(n8482), .A2(n8018), .ZN(n7806) );
  NAND2_X1 U6013 ( .A1(n7806), .A2(n7812), .ZN(n8312) );
  NAND2_X1 U6014 ( .A1(n6604), .A2(n8747), .ZN(n6576) );
  NAND2_X1 U6015 ( .A1(n5533), .A2(n5532), .ZN(n4476) );
  OR2_X1 U6016 ( .A1(n4843), .A2(n4505), .ZN(n4477) );
  NAND2_X1 U6017 ( .A1(n9431), .A2(n8599), .ZN(n4478) );
  OR2_X2 U6018 ( .A1(n6249), .A2(n7677), .ZN(n4479) );
  INV_X1 U6019 ( .A(n8981), .ZN(n4762) );
  NAND2_X1 U6020 ( .A1(n4788), .A2(n8293), .ZN(n4787) );
  AND4_X1 U6021 ( .A1(n5949), .A2(n5819), .A3(n4869), .A4(n5818), .ZN(n4480)
         );
  INV_X1 U6022 ( .A(n7814), .ZN(n5019) );
  OR2_X1 U6023 ( .A1(n5922), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U6024 ( .A1(n5383), .A2(n5382), .ZN(n7111) );
  AND2_X1 U6025 ( .A1(n4595), .A2(n4594), .ZN(n4481) );
  AND2_X1 U6026 ( .A1(n5026), .A2(n6949), .ZN(n4482) );
  AND2_X1 U6027 ( .A1(n5202), .A2(SI_4_), .ZN(n4483) );
  AND2_X1 U6028 ( .A1(n4624), .A2(n4626), .ZN(n4484) );
  NAND2_X1 U6029 ( .A1(n7811), .A2(n7808), .ZN(n8263) );
  INV_X1 U6030 ( .A(n8263), .ZN(n8302) );
  AND2_X1 U6031 ( .A1(n5198), .A2(n5197), .ZN(n4485) );
  OR2_X1 U6032 ( .A1(n9174), .A2(n9149), .ZN(n4486) );
  AND2_X1 U6033 ( .A1(n5044), .A2(n5096), .ZN(n4487) );
  NOR2_X1 U6034 ( .A1(n8592), .A2(n9227), .ZN(n4488) );
  AND2_X1 U6035 ( .A1(n4953), .A2(n5595), .ZN(n4489) );
  AND2_X1 U6036 ( .A1(n4593), .A2(n4592), .ZN(n4490) );
  OR2_X1 U6037 ( .A1(n9569), .A2(n9568), .ZN(n4491) );
  AND2_X1 U6038 ( .A1(n6797), .A2(n4504), .ZN(n4492) );
  CLKBUF_X3 U6039 ( .A(n6444), .Z(n8721) );
  XOR2_X1 U6040 ( .A(n7923), .B(n7996), .Z(n4493) );
  NAND2_X1 U6041 ( .A1(n5639), .A2(n5638), .ZN(n4494) );
  OR2_X1 U6042 ( .A1(n9154), .A2(n4707), .ZN(n4495) );
  AND2_X1 U6043 ( .A1(n8571), .A2(n8570), .ZN(n4496) );
  XNOR2_X1 U6044 ( .A(n8471), .B(n8304), .ZN(n8284) );
  AND2_X1 U6045 ( .A1(n8943), .A2(n6740), .ZN(n4497) );
  NAND2_X1 U6046 ( .A1(n7695), .A2(n7693), .ZN(n9574) );
  AND2_X1 U6047 ( .A1(n4995), .A2(n8947), .ZN(n4498) );
  OR2_X1 U6048 ( .A1(n9365), .A2(n9013), .ZN(n4499) );
  OAI211_X1 U6049 ( .C1(n6739), .C2(n6749), .A(n6738), .B(n6737), .ZN(n6896)
         );
  AND2_X1 U6050 ( .A1(n8008), .A2(n8645), .ZN(n4500) );
  OR2_X1 U6051 ( .A1(n7781), .A2(n7831), .ZN(n4501) );
  OR2_X1 U6052 ( .A1(n7794), .A2(n7831), .ZN(n4502) );
  INV_X1 U6053 ( .A(n8801), .ZN(n4764) );
  AND4_X1 U6054 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(n6262)
         );
  XNOR2_X1 U6055 ( .A(n5748), .B(n5747), .ZN(n5774) );
  AND2_X1 U6056 ( .A1(n8519), .A2(n8451), .ZN(n4503) );
  AND2_X1 U6057 ( .A1(n6912), .A2(n9813), .ZN(n4504) );
  AND2_X1 U6058 ( .A1(n4493), .A2(n7919), .ZN(n4505) );
  INV_X1 U6059 ( .A(n7733), .ZN(n4576) );
  AND2_X1 U6060 ( .A1(n4486), .A2(n9182), .ZN(n4506) );
  NAND2_X1 U6061 ( .A1(n5826), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5837) );
  INV_X1 U6062 ( .A(n7790), .ZN(n4618) );
  AND2_X1 U6063 ( .A1(n7289), .A2(n5488), .ZN(n4507) );
  INV_X1 U6064 ( .A(n7757), .ZN(n4735) );
  OR3_X1 U6065 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        n9861), .ZN(n4508) );
  AND2_X1 U6066 ( .A1(n7854), .A2(n7112), .ZN(n4509) );
  AND2_X1 U6067 ( .A1(n8326), .A2(n7804), .ZN(n4510) );
  NAND2_X1 U6068 ( .A1(n5024), .A2(n7653), .ZN(n8417) );
  OR2_X1 U6069 ( .A1(n8523), .A2(n8250), .ZN(n4511) );
  AND2_X1 U6070 ( .A1(n8762), .A2(n9015), .ZN(n4512) );
  OAI21_X1 U6071 ( .B1(n7467), .B2(n4665), .A(n4668), .ZN(n4667) );
  NAND2_X1 U6072 ( .A1(n5568), .A2(n5567), .ZN(n8513) );
  AND2_X1 U6073 ( .A1(n6764), .A2(n8969), .ZN(n4513) );
  NAND2_X1 U6074 ( .A1(n6599), .A2(n6262), .ZN(n6604) );
  AND2_X1 U6075 ( .A1(n5323), .A2(n5322), .ZN(n4514) );
  NAND2_X1 U6076 ( .A1(n7565), .A2(n7564), .ZN(n9365) );
  INV_X1 U6077 ( .A(n8762), .ZN(n9628) );
  NAND2_X1 U6078 ( .A1(n7215), .A2(n7214), .ZN(n8762) );
  OR2_X1 U6079 ( .A1(n8504), .A2(n8038), .ZN(n7793) );
  AND2_X1 U6080 ( .A1(n9152), .A2(n8895), .ZN(n4515) );
  AND2_X1 U6081 ( .A1(n7853), .A2(n6947), .ZN(n4516) );
  INV_X1 U6082 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9456) );
  AND2_X1 U6083 ( .A1(n8366), .A2(n4501), .ZN(n4517) );
  INV_X1 U6084 ( .A(n9380), .ZN(n9227) );
  NAND2_X1 U6085 ( .A1(n7530), .A2(n7529), .ZN(n9380) );
  INV_X1 U6086 ( .A(n4844), .ZN(n4843) );
  AND2_X1 U6087 ( .A1(n5207), .A2(n5206), .ZN(n5880) );
  INV_X1 U6088 ( .A(n5880), .ZN(n6555) );
  AND2_X1 U6089 ( .A1(n7619), .A2(n8931), .ZN(n4518) );
  AND2_X1 U6090 ( .A1(n6019), .A2(n6020), .ZN(n4519) );
  AND2_X1 U6091 ( .A1(n7663), .A2(n7662), .ZN(n8241) );
  INV_X1 U6092 ( .A(n8241), .ZN(n8462) );
  AND2_X1 U6093 ( .A1(n4576), .A2(n5861), .ZN(n4520) );
  AND2_X1 U6094 ( .A1(n7028), .A2(n7030), .ZN(n4521) );
  AND2_X1 U6095 ( .A1(n7756), .A2(n7751), .ZN(n6832) );
  INV_X1 U6096 ( .A(n6832), .ZN(n5030) );
  NAND2_X1 U6097 ( .A1(n5408), .A2(n5407), .ZN(n9615) );
  AND3_X1 U6098 ( .A1(n5946), .A2(n5942), .A3(n5817), .ZN(n4522) );
  AND2_X1 U6099 ( .A1(n4782), .A2(n4781), .ZN(n4523) );
  INV_X1 U6100 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5047) );
  INV_X1 U6101 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5946) );
  AND2_X1 U6102 ( .A1(n7792), .A2(n7791), .ZN(n4524) );
  NOR2_X1 U6103 ( .A1(n7810), .A2(n7834), .ZN(n4525) );
  NOR2_X1 U6104 ( .A1(n7396), .A2(n8709), .ZN(n4526) );
  INV_X1 U6105 ( .A(n4626), .ZN(n4625) );
  NAND2_X1 U6106 ( .A1(n8261), .A2(n7802), .ZN(n4626) );
  INV_X1 U6107 ( .A(n8933), .ZN(n7616) );
  AND2_X1 U6108 ( .A1(n9394), .A2(n8591), .ZN(n8933) );
  AND2_X1 U6109 ( .A1(n6681), .A2(n8119), .ZN(n4527) );
  AND2_X1 U6110 ( .A1(n8302), .A2(n4584), .ZN(n4528) );
  AND2_X1 U6111 ( .A1(n7833), .A2(n7832), .ZN(n4529) );
  INV_X1 U6112 ( .A(n7736), .ZN(n5034) );
  NAND2_X1 U6113 ( .A1(n4863), .A2(n4864), .ZN(n4530) );
  OR2_X1 U6114 ( .A1(n4624), .A2(n4510), .ZN(n4531) );
  AND2_X1 U6115 ( .A1(n5222), .A2(SI_5_), .ZN(n4532) );
  NAND2_X1 U6116 ( .A1(n9506), .A2(n7096), .ZN(n4533) );
  NAND2_X1 U6117 ( .A1(n9461), .A2(n9466), .ZN(n6338) );
  INV_X2 U6118 ( .A(n6646), .ZN(n7623) );
  OR2_X1 U6119 ( .A1(n7211), .A2(n4512), .ZN(n4534) );
  NOR2_X1 U6120 ( .A1(n8414), .A2(n8254), .ZN(n4535) );
  OAI21_X1 U6121 ( .B1(n4982), .B2(n4506), .A(n9147), .ZN(n4981) );
  NAND2_X1 U6122 ( .A1(n5880), .A2(n9866), .ZN(n7722) );
  INV_X1 U6123 ( .A(n4983), .ZN(n4982) );
  NAND2_X1 U6124 ( .A1(n4536), .A2(n4486), .ZN(n4983) );
  INV_X1 U6125 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U6126 ( .A1(n4499), .A2(n7586), .ZN(n4536) );
  AND2_X1 U6127 ( .A1(n5829), .A2(n4523), .ZN(n4537) );
  AND2_X1 U6128 ( .A1(n6448), .A2(n6673), .ZN(n4538) );
  OR2_X1 U6129 ( .A1(n8466), .A2(n7661), .ZN(n7823) );
  NAND2_X1 U6130 ( .A1(n5830), .A2(n5829), .ZN(n5842) );
  AND2_X1 U6131 ( .A1(n8643), .A2(n8570), .ZN(n4539) );
  AND2_X1 U6132 ( .A1(n4984), .A2(n4499), .ZN(n4540) );
  AND2_X1 U6133 ( .A1(n4778), .A2(n9130), .ZN(n4541) );
  NAND3_X1 U6134 ( .A1(n4632), .A2(n4824), .A3(n5001), .ZN(n4542) );
  NOR2_X1 U6135 ( .A1(n7734), .A2(n7846), .ZN(n4543) );
  NOR2_X1 U6136 ( .A1(n8404), .A2(n5023), .ZN(n5022) );
  INV_X1 U6137 ( .A(n7309), .ZN(n4849) );
  NOR2_X1 U6138 ( .A1(n7653), .A2(n4793), .ZN(n4792) );
  AND2_X1 U6139 ( .A1(n7438), .A2(n7436), .ZN(n4544) );
  AND2_X1 U6140 ( .A1(n5100), .A2(n5047), .ZN(n4545) );
  OR2_X1 U6141 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4546) );
  INV_X1 U6142 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5813) );
  AND2_X1 U6143 ( .A1(n4476), .A2(n5518), .ZN(n4899) );
  INV_X1 U6144 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4869) );
  INV_X1 U6145 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5815) );
  INV_X1 U6146 ( .A(n8838), .ZN(n4642) );
  OR2_X1 U6147 ( .A1(n7906), .A2(n7905), .ZN(n4547) );
  NAND2_X1 U6148 ( .A1(n9785), .A2(n9003), .ZN(n8921) );
  NAND2_X1 U6149 ( .A1(n9567), .A2(n8249), .ZN(n8443) );
  NAND2_X1 U6150 ( .A1(n4987), .A2(n4986), .ZN(n9315) );
  OAI21_X1 U6151 ( .B1(n6187), .B2(n4853), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6400) );
  INV_X1 U6152 ( .A(n8326), .ZN(n8336) );
  NAND2_X1 U6153 ( .A1(n7660), .A2(n7659), .ZN(n8466) );
  INV_X1 U6154 ( .A(n8466), .ZN(n4788) );
  NAND3_X1 U6155 ( .A1(n4824), .A2(n5001), .A3(n4823), .ZN(n5913) );
  NAND2_X1 U6156 ( .A1(n9242), .A2(n4697), .ZN(n4700) );
  INV_X1 U6157 ( .A(n4789), .ZN(n8434) );
  NOR2_X1 U6158 ( .A1(n9569), .A2(n4597), .ZN(n4789) );
  INV_X1 U6159 ( .A(n5000), .ZN(n4999) );
  AND2_X1 U6160 ( .A1(n9387), .A2(n9231), .ZN(n5000) );
  NOR2_X1 U6161 ( .A1(n9569), .A2(n4598), .ZN(n4596) );
  OR2_X1 U6162 ( .A1(n9380), .A2(n8592), .ZN(n8932) );
  INV_X1 U6163 ( .A(n4600), .ZN(n8444) );
  NOR2_X1 U6164 ( .A1(n9569), .A2(n4601), .ZN(n4600) );
  OR2_X1 U6165 ( .A1(n6187), .A2(n6186), .ZN(n4548) );
  NAND2_X1 U6166 ( .A1(n7920), .A2(n4505), .ZN(n4549) );
  NAND2_X1 U6167 ( .A1(n8260), .A2(n8346), .ZN(n4818) );
  NAND2_X1 U6168 ( .A1(n5718), .A2(n5717), .ZN(n4550) );
  AND4_X1 U6169 ( .A1(n5001), .A2(n5925), .A3(n5812), .A4(n5929), .ZN(n4551)
         );
  AND2_X1 U6170 ( .A1(n4994), .A2(n4993), .ZN(n4552) );
  AND2_X1 U6171 ( .A1(n7113), .A2(n7112), .ZN(n4553) );
  NAND2_X1 U6172 ( .A1(n5504), .A2(n5503), .ZN(n9568) );
  INV_X1 U6173 ( .A(n9568), .ZN(n4602) );
  NAND2_X1 U6174 ( .A1(n7840), .A2(n7687), .ZN(n7877) );
  INV_X1 U6175 ( .A(n7877), .ZN(n4890) );
  OAI21_X1 U6176 ( .B1(n5842), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U6177 ( .A1(n5793), .A2(n5782), .ZN(n8082) );
  AND2_X1 U6178 ( .A1(n4878), .A2(n6592), .ZN(n4554) );
  NAND2_X1 U6179 ( .A1(n6431), .A2(n7729), .ZN(n6421) );
  NAND2_X1 U6180 ( .A1(n5430), .A2(n5429), .ZN(n9609) );
  INV_X1 U6181 ( .A(n9609), .ZN(n4594) );
  INV_X1 U6182 ( .A(n5071), .ZN(n5477) );
  NOR3_X1 U6183 ( .A1(n7151), .A2(n9419), .A3(n4704), .ZN(n4701) );
  INV_X1 U6184 ( .A(n4702), .ZN(n9317) );
  NOR2_X1 U6185 ( .A1(n7151), .A2(n4704), .ZN(n4702) );
  NAND2_X1 U6186 ( .A1(n6797), .A2(n4693), .ZN(n4694) );
  INV_X1 U6187 ( .A(n6017), .ZN(n4564) );
  AND2_X1 U6188 ( .A1(n7642), .A2(SI_29_), .ZN(n4555) );
  INV_X1 U6189 ( .A(n4966), .ZN(n4965) );
  NAND2_X1 U6190 ( .A1(n4556), .A2(n7640), .ZN(n4966) );
  NAND2_X1 U6191 ( .A1(n7656), .A2(n10199), .ZN(n4556) );
  NAND2_X1 U6192 ( .A1(n5837), .A2(n5833), .ZN(n5836) );
  AND2_X1 U6193 ( .A1(n6948), .A2(n6947), .ZN(n4557) );
  NAND2_X1 U6194 ( .A1(n6242), .A2(n6234), .ZN(n9845) );
  INV_X1 U6195 ( .A(n9933), .ZN(n4592) );
  INV_X1 U6196 ( .A(n9926), .ZN(n4785) );
  AND2_X2 U6197 ( .A1(n6370), .A2(n6358), .ZN(n9979) );
  INV_X1 U6198 ( .A(n9979), .ZN(n4579) );
  AND2_X2 U6199 ( .A1(n6565), .A2(n9790), .ZN(n9767) );
  AND2_X1 U6200 ( .A1(n9565), .A2(n9618), .ZN(n9966) );
  INV_X1 U6201 ( .A(n6173), .ZN(n4874) );
  OR2_X1 U6202 ( .A1(n4579), .A2(n9966), .ZN(n4558) );
  INV_X1 U6203 ( .A(n6733), .ZN(n9001) );
  AND2_X1 U6204 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n4559) );
  INV_X1 U6205 ( .A(n4473), .ZN(n9785) );
  INV_X1 U6206 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n4770) );
  NAND2_X1 U6207 ( .A1(n4916), .A2(n5522), .ZN(n5536) );
  INV_X1 U6208 ( .A(n4667), .ZN(n5615) );
  NAND2_X1 U6209 ( .A1(n8283), .A2(n7814), .ZN(n8272) );
  OAI21_X2 U6210 ( .B1(n8303), .B2(n8263), .A(n7811), .ZN(n8285) );
  NOR2_X2 U6211 ( .A1(n7162), .A2(n7161), .ZN(n7164) );
  NAND2_X1 U6212 ( .A1(n9769), .A2(n6764), .ZN(n6793) );
  MUX2_X1 U6213 ( .A(n8837), .B(n8836), .S(n8921), .Z(n8842) );
  MUX2_X1 U6214 ( .A(n8866), .B(n8865), .S(n8901), .Z(n8884) );
  MUX2_X1 U6215 ( .A(n8804), .B(n8803), .S(n8901), .Z(n8811) );
  NAND2_X1 U6216 ( .A1(n4780), .A2(n4782), .ZN(n6146) );
  NAND3_X1 U6217 ( .A1(n4633), .A2(n8747), .A3(n6604), .ZN(n6605) );
  NAND2_X1 U6218 ( .A1(n4968), .A2(n9008), .ZN(P1_U3240) );
  NAND2_X2 U6219 ( .A1(n6150), .A2(n6151), .ZN(n6273) );
  NAND2_X1 U6220 ( .A1(n8998), .A2(n9785), .ZN(n4971) );
  NAND2_X2 U6221 ( .A1(n4519), .A2(n4564), .ZN(n6195) );
  NAND2_X1 U6222 ( .A1(n4828), .A2(n4500), .ZN(n4827) );
  NAND2_X2 U6223 ( .A1(n8636), .A2(n8635), .ZN(n7920) );
  NAND2_X1 U6224 ( .A1(n6207), .A2(n6255), .ZN(n6259) );
  NAND2_X1 U6225 ( .A1(n6777), .A2(n6776), .ZN(n6865) );
  OAI21_X1 U6226 ( .B1(n4868), .B2(n4867), .A(n6203), .ZN(n4866) );
  NAND3_X1 U6227 ( .A1(n7100), .A2(n7309), .A3(n7099), .ZN(n4846) );
  INV_X1 U6228 ( .A(n5038), .ZN(n5036) );
  NAND2_X1 U6229 ( .A1(n4675), .A2(n4674), .ZN(n4681) );
  INV_X1 U6230 ( .A(n5195), .ZN(n4875) );
  NOR2_X1 U6231 ( .A1(n8079), .A2(n5056), .ZN(n8074) );
  NAND2_X1 U6232 ( .A1(n4885), .A2(n4883), .ZN(n6934) );
  NAND2_X4 U6233 ( .A1(n6077), .A2(n7677), .ZN(n7681) );
  NAND2_X1 U6234 ( .A1(n9877), .A2(n9876), .ZN(n4567) );
  NAND2_X1 U6235 ( .A1(n6519), .A2(n5856), .ZN(n4568) );
  OAI21_X1 U6236 ( .B1(n4573), .B2(n4571), .A(n4569), .ZN(n6683) );
  INV_X2 U6237 ( .A(n8547), .ZN(n5084) );
  NAND2_X2 U6238 ( .A1(n4589), .A2(n5081), .ZN(n8547) );
  NAND2_X1 U6239 ( .A1(n8248), .A2(n4591), .ZN(n9567) );
  NAND2_X1 U6240 ( .A1(n4590), .A2(n4790), .ZN(n8405) );
  NAND3_X1 U6241 ( .A1(n9567), .A2(n4792), .A3(n8249), .ZN(n4590) );
  AND3_X2 U6242 ( .A1(n5069), .A2(n5068), .A3(n5184), .ZN(n5071) );
  INV_X1 U6243 ( .A(n4596), .ZN(n8410) );
  NAND2_X1 U6244 ( .A1(n4604), .A2(n4543), .ZN(n4603) );
  OAI21_X1 U6245 ( .B1(n7728), .B2(n7727), .A(n7726), .ZN(n4605) );
  NAND2_X2 U6246 ( .A1(n5083), .A2(n8547), .ZN(n5189) );
  OR2_X1 U6247 ( .A1(n7803), .A2(n4623), .ZN(n4622) );
  AOI21_X1 U6248 ( .B1(n4625), .B2(n8336), .A(n7834), .ZN(n4624) );
  NOR2_X2 U6249 ( .A1(n4630), .A2(n4629), .ZN(n6191) );
  NAND3_X1 U6250 ( .A1(n4824), .A2(n5815), .A3(n5001), .ZN(n4629) );
  NAND4_X1 U6251 ( .A1(n4632), .A2(n4631), .A3(n4522), .A4(n4480), .ZN(n4630)
         );
  AND2_X2 U6252 ( .A1(n5812), .A2(n5925), .ZN(n4632) );
  NOR2_X4 U6253 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5812) );
  NOR2_X4 U6254 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5925) );
  NAND2_X1 U6255 ( .A1(n6604), .A2(n6605), .ZN(n6810) );
  INV_X1 U6256 ( .A(n6575), .ZN(n4633) );
  NAND2_X1 U6257 ( .A1(n9326), .A2(n4638), .ZN(n4636) );
  INV_X1 U6258 ( .A(n8932), .ZN(n4645) );
  NAND2_X1 U6259 ( .A1(n4657), .A2(n4654), .ZN(P1_U3263) );
  NAND2_X1 U6260 ( .A1(n7634), .A2(n9786), .ZN(n4657) );
  NAND3_X1 U6261 ( .A1(n4709), .A2(n8234), .A3(n4658), .ZN(n4915) );
  MUX2_X1 U6262 ( .A(n5203), .B(n5204), .S(n5986), .Z(n5221) );
  MUX2_X1 U6263 ( .A(n5181), .B(n10179), .S(n5986), .Z(n5201) );
  MUX2_X1 U6264 ( .A(n5223), .B(n5994), .S(n4659), .Z(n5244) );
  MUX2_X1 U6265 ( .A(n5996), .B(n5248), .S(n4659), .Z(n5271) );
  MUX2_X1 U6266 ( .A(n5301), .B(n6015), .S(n4659), .Z(n5303) );
  MUX2_X1 U6267 ( .A(n5999), .B(n5998), .S(n4659), .Z(n5276) );
  MUX2_X1 U6268 ( .A(n6028), .B(n6027), .S(n4659), .Z(n5327) );
  MUX2_X1 U6269 ( .A(n5350), .B(n6031), .S(n4659), .Z(n5368) );
  NAND2_X1 U6270 ( .A1(n4899), .A2(n7459), .ZN(n4671) );
  NAND3_X1 U6271 ( .A1(n7459), .A2(n4673), .A3(n4476), .ZN(n4670) );
  NAND2_X1 U6272 ( .A1(n4672), .A2(n7335), .ZN(n4673) );
  NAND2_X1 U6273 ( .A1(n7276), .A2(n5518), .ZN(n4672) );
  NAND2_X1 U6274 ( .A1(n4678), .A2(n5654), .ZN(n4682) );
  INV_X1 U6275 ( .A(n4694), .ZN(n6999) );
  INV_X1 U6276 ( .A(n4700), .ZN(n9196) );
  INV_X1 U6277 ( .A(n4701), .ZN(n9316) );
  NOR2_X1 U6278 ( .A1(n9154), .A2(n9350), .ZN(n9112) );
  NOR2_X1 U6279 ( .A1(n9154), .A2(n4706), .ZN(n9136) );
  NOR2_X1 U6280 ( .A1(n9735), .A2(n4709), .ZN(n4755) );
  NAND2_X1 U6281 ( .A1(n5134), .A2(n5133), .ZN(n5137) );
  NAND2_X1 U6282 ( .A1(n6198), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4710) );
  NAND3_X1 U6283 ( .A1(n7873), .A2(n7869), .A3(n9895), .ZN(n4739) );
  MUX2_X1 U6284 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n5935), .S(n6251), .Z(n6052)
         );
  NAND2_X1 U6285 ( .A1(n9461), .A2(n6151), .ZN(n6274) );
  NAND3_X1 U6286 ( .A1(n6185), .A2(n6184), .A3(n4768), .ZN(n6235) );
  NAND2_X1 U6287 ( .A1(n9152), .A2(n4778), .ZN(n9129) );
  OAI211_X1 U6288 ( .C1(n9152), .C2(n4776), .A(n4772), .B(n4771), .ZN(n9134)
         );
  NAND2_X1 U6289 ( .A1(n9152), .A2(n4541), .ZN(n4771) );
  NAND2_X1 U6290 ( .A1(n8297), .A2(n8293), .ZN(n8267) );
  NAND2_X1 U6291 ( .A1(n8297), .A2(n4786), .ZN(n8240) );
  NOR2_X2 U6292 ( .A1(n7267), .A2(n7435), .ZN(n8235) );
  NOR2_X1 U6293 ( .A1(n8405), .A2(n4800), .ZN(n8256) );
  NAND2_X1 U6294 ( .A1(n4801), .A2(n4804), .ZN(n8265) );
  NAND2_X1 U6295 ( .A1(n8327), .A2(n4806), .ZN(n4801) );
  NAND2_X1 U6296 ( .A1(n7437), .A2(n4544), .ZN(n8248) );
  INV_X1 U6297 ( .A(n5501), .ZN(n4819) );
  NAND2_X1 U6298 ( .A1(n4820), .A2(n5046), .ZN(n5081) );
  OR2_X1 U6299 ( .A1(n5189), .A2(n5082), .ZN(n5089) );
  OAI21_X1 U6300 ( .B1(n6533), .B2(n6535), .A(n6353), .ZN(n5849) );
  OR2_X1 U6301 ( .A1(n5706), .A2(n6514), .ZN(n5088) );
  AND3_X2 U6302 ( .A1(n5925), .A2(n5812), .A3(n5815), .ZN(n4823) );
  NAND4_X1 U6303 ( .A1(n4829), .A2(n8016), .A3(n4827), .A4(n4825), .ZN(
        P1_U3218) );
  NAND3_X1 U6304 ( .A1(n4834), .A2(n4831), .A3(n4830), .ZN(n4829) );
  NAND2_X1 U6305 ( .A1(n7920), .A2(n4477), .ZN(n4840) );
  OAI21_X1 U6306 ( .B1(n7919), .B2(n4493), .A(n8687), .ZN(n4844) );
  OR2_X1 U6307 ( .A1(n4845), .A2(n4493), .ZN(n8685) );
  NAND2_X1 U6308 ( .A1(n4846), .A2(n4847), .ZN(n7349) );
  INV_X1 U6309 ( .A(n4850), .ZN(n6190) );
  INV_X1 U6310 ( .A(n4855), .ZN(n8636) );
  NAND3_X1 U6311 ( .A1(n7963), .A2(n8643), .A3(n7966), .ZN(n4864) );
  NAND3_X1 U6312 ( .A1(n4863), .A2(n4864), .A3(n7976), .ZN(n8614) );
  NAND2_X1 U6313 ( .A1(n8571), .A2(n4539), .ZN(n4863) );
  NAND2_X1 U6314 ( .A1(n7029), .A2(n7028), .ZN(n7033) );
  NAND2_X2 U6315 ( .A1(n6867), .A2(n6868), .ZN(n7029) );
  NAND3_X1 U6316 ( .A1(n4865), .A2(n6331), .A3(n6266), .ZN(n6332) );
  OR2_X1 U6317 ( .A1(n6264), .A2(n6265), .ZN(n4865) );
  NAND2_X1 U6318 ( .A1(n6264), .A2(n6265), .ZN(n6331) );
  INV_X2 U6319 ( .A(n4868), .ZN(n7998) );
  NAND2_X2 U6320 ( .A1(n6196), .A2(n6322), .ZN(n4868) );
  NAND2_X1 U6321 ( .A1(n7083), .A2(n4871), .ZN(n5491) );
  INV_X1 U6322 ( .A(n6140), .ZN(n5219) );
  NAND2_X1 U6323 ( .A1(n5889), .A2(n4879), .ZN(n4877) );
  NAND2_X1 U6324 ( .A1(n5360), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U6325 ( .A1(n4891), .A2(n7690), .ZN(n6349) );
  INV_X1 U6326 ( .A(n9895), .ZN(n4889) );
  NAND2_X1 U6327 ( .A1(n7277), .A2(n4896), .ZN(n4894) );
  INV_X1 U6328 ( .A(n5106), .ZN(n5107) );
  NAND2_X2 U6329 ( .A1(n4915), .A2(n4913), .ZN(n5164) );
  NAND3_X1 U6330 ( .A1(n4914), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U6331 ( .A1(n5499), .A2(n4917), .ZN(n4916) );
  NAND2_X1 U6332 ( .A1(n5200), .A2(n4923), .ZN(n4922) );
  NAND2_X1 U6333 ( .A1(n5300), .A2(n5299), .ZN(n5324) );
  NAND2_X1 U6334 ( .A1(n5300), .A2(n4932), .ZN(n4931) );
  NAND2_X1 U6335 ( .A1(n5641), .A2(n4942), .ZN(n4940) );
  NAND2_X1 U6336 ( .A1(n5641), .A2(n5640), .ZN(n4941) );
  NAND2_X1 U6337 ( .A1(n5562), .A2(n4489), .ZN(n4952) );
  OR2_X1 U6338 ( .A1(n5562), .A2(n5561), .ZN(n4957) );
  NAND3_X1 U6339 ( .A1(n4953), .A2(n4956), .A3(n5595), .ZN(n4951) );
  NAND3_X1 U6340 ( .A1(n8960), .A2(n8961), .A3(n9130), .ZN(n4962) );
  NAND2_X1 U6341 ( .A1(n7637), .A2(n7636), .ZN(n4967) );
  NAND3_X1 U6342 ( .A1(n4973), .A2(n4972), .A3(n4971), .ZN(n4970) );
  NAND2_X1 U6343 ( .A1(n6790), .A2(n6644), .ZN(n4976) );
  NAND2_X1 U6344 ( .A1(n6790), .A2(n4974), .ZN(n6736) );
  NAND2_X1 U6345 ( .A1(n6736), .A2(n4975), .ZN(n9817) );
  NAND2_X1 U6346 ( .A1(n4976), .A2(n6657), .ZN(n4975) );
  NAND2_X1 U6347 ( .A1(n4538), .A2(n4977), .ZN(n6764) );
  NAND2_X1 U6348 ( .A1(n9177), .A2(n4506), .ZN(n4980) );
  NAND2_X1 U6349 ( .A1(n7212), .A2(n4989), .ZN(n4987) );
  NAND3_X1 U6350 ( .A1(n5925), .A2(n5812), .A3(n5929), .ZN(n5922) );
  OAI21_X1 U6351 ( .B1(n6524), .B2(n5012), .A(n7706), .ZN(n5011) );
  NAND2_X1 U6352 ( .A1(n8285), .A2(n5017), .ZN(n5016) );
  NAND2_X1 U6353 ( .A1(n8285), .A2(n8284), .ZN(n8283) );
  NAND2_X1 U6354 ( .A1(n8416), .A2(n5022), .ZN(n5020) );
  NAND2_X1 U6355 ( .A1(n5020), .A2(n5021), .ZN(n8377) );
  NAND2_X1 U6356 ( .A1(n5025), .A2(n4482), .ZN(n7117) );
  NAND2_X1 U6357 ( .A1(n6830), .A2(n5027), .ZN(n5025) );
  NAND2_X1 U6358 ( .A1(n7648), .A2(n5031), .ZN(n7651) );
  XNOR2_X1 U6359 ( .A(n5735), .B(n6535), .ZN(n5129) );
  OR2_X1 U6360 ( .A1(n6495), .A2(n6535), .ZN(n7710) );
  NAND2_X1 U6361 ( .A1(n5423), .A2(n5062), .ZN(n5425) );
  NAND2_X1 U6362 ( .A1(n8968), .A2(n8967), .ZN(n6659) );
  OAI222_X1 U6363 ( .A1(n9509), .A2(n7633), .B1(n7632), .B2(n9771), .C1(n9166), 
        .C2(n9773), .ZN(n7634) );
  XNOR2_X1 U6364 ( .A(n7673), .B(SI_30_), .ZN(n8726) );
  XNOR2_X1 U6365 ( .A(n5639), .B(n5629), .ZN(n8028) );
  NAND4_X1 U6366 ( .A1(n6247), .A2(n6245), .A3(n6248), .A4(n6246), .ZN(n6570)
         );
  NAND2_X1 U6367 ( .A1(n5693), .A2(n5692), .ZN(n5695) );
  XNOR2_X1 U6368 ( .A(n5693), .B(n5692), .ZN(n7572) );
  XNOR2_X1 U6369 ( .A(n5674), .B(n5673), .ZN(n7563) );
  NAND2_X2 U6370 ( .A1(n7328), .A2(n5495), .ZN(n7277) );
  NAND2_X1 U6371 ( .A1(n6637), .A2(n4513), .ZN(n6639) );
  OR2_X1 U6372 ( .A1(n6273), .A2(n6229), .ZN(n6248) );
  XNOR2_X1 U6373 ( .A(n5615), .B(n5616), .ZN(n8079) );
  INV_X1 U6374 ( .A(n7954), .ZN(n7957) );
  OAI21_X1 U6375 ( .B1(n6492), .B2(n5850), .A(n7701), .ZN(n5866) );
  NAND2_X1 U6376 ( .A1(n5309), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5087) );
  XNOR2_X1 U6377 ( .A(n8272), .B(n8273), .ZN(n8278) );
  NAND4_X2 U6378 ( .A1(n5089), .A2(n5088), .A3(n5087), .A4(n5086), .ZN(n6157)
         );
  OR2_X1 U6379 ( .A1(n8298), .A2(n5706), .ZN(n5712) );
  INV_X1 U6380 ( .A(n5706), .ZN(n5791) );
  OR2_X1 U6381 ( .A1(n5706), .A2(n6534), .ZN(n5127) );
  NAND2_X1 U6382 ( .A1(n7502), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6200) );
  OAI211_X1 U6383 ( .C1(n6254), .C2(n6749), .A(n6253), .B(n6252), .ZN(n6279)
         );
  OR2_X1 U6384 ( .A1(n4479), .A2(n6250), .ZN(n6253) );
  INV_X1 U6385 ( .A(n5083), .ZN(n7643) );
  NAND2_X4 U6386 ( .A1(n5083), .A2(n5084), .ZN(n5706) );
  OAI21_X1 U6387 ( .B1(n5621), .B2(n5620), .A(n5619), .ZN(n5641) );
  AND2_X1 U6388 ( .A1(n8397), .A2(n7690), .ZN(n5056) );
  INV_X1 U6389 ( .A(n9593), .ZN(n8436) );
  OR2_X1 U6390 ( .A1(n9431), .A2(n9505), .ZN(n5057) );
  NAND2_X1 U6391 ( .A1(n7036), .A2(n7035), .ZN(n7100) );
  AND2_X1 U6392 ( .A1(n5348), .A2(n5329), .ZN(n5058) );
  INV_X1 U6393 ( .A(n8031), .ZN(n8364) );
  AND2_X1 U6394 ( .A1(n5653), .A2(n5652), .ZN(n8031) );
  AND2_X1 U6395 ( .A1(n5325), .A2(n5305), .ZN(n5061) );
  AND2_X1 U6396 ( .A1(n5424), .A2(n5405), .ZN(n5062) );
  NAND2_X1 U6397 ( .A1(n7654), .A2(n8326), .ZN(n8311) );
  NAND2_X1 U6398 ( .A1(n6579), .A2(n6578), .ZN(n9776) );
  AND2_X1 U6399 ( .A1(n6374), .A2(n8927), .ZN(n9504) );
  INV_X1 U6400 ( .A(n9504), .ZN(n9771) );
  INV_X1 U6401 ( .A(n9507), .ZN(n9773) );
  INV_X1 U6402 ( .A(n7834), .ZN(n7831) );
  NAND2_X1 U6403 ( .A1(n7866), .A2(n7831), .ZN(n7832) );
  NOR2_X1 U6404 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5067) );
  OR2_X1 U6405 ( .A1(n9426), .A2(n9328), .ZN(n7394) );
  INV_X1 U6406 ( .A(n9150), .ZN(n9124) );
  NAND2_X1 U6407 ( .A1(n9021), .A2(n9755), .ZN(n8968) );
  INV_X1 U6408 ( .A(n5616), .ZN(n5617) );
  INV_X1 U6409 ( .A(n5584), .ZN(n5583) );
  INV_X1 U6410 ( .A(n5570), .ZN(n5569) );
  INV_X1 U6411 ( .A(n8415), .ZN(n7653) );
  INV_X1 U6412 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5312) );
  INV_X1 U6413 ( .A(n7753), .ZN(n7161) );
  INV_X1 U6414 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5426) );
  INV_X1 U6415 ( .A(n7508), .ZN(n7477) );
  INV_X1 U6416 ( .A(n7072), .ZN(n7071) );
  AND2_X1 U6417 ( .A1(n6204), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6202) );
  INV_X1 U6418 ( .A(n6269), .ZN(n6266) );
  INV_X1 U6419 ( .A(n7544), .ZN(n7542) );
  INV_X1 U6420 ( .A(n7223), .ZN(n7221) );
  INV_X1 U6421 ( .A(n5890), .ZN(n5266) );
  OR2_X1 U6422 ( .A1(n5433), .A2(n5432), .ZN(n5464) );
  NOR2_X1 U6423 ( .A1(n4667), .A2(n5617), .ZN(n5618) );
  INV_X1 U6424 ( .A(n5647), .ZN(n5645) );
  NAND2_X1 U6425 ( .A1(n5569), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5584) );
  OR2_X1 U6426 ( .A1(n5607), .A2(n5606), .ZN(n5631) );
  OR2_X1 U6427 ( .A1(n5549), .A2(n5548), .ZN(n5570) );
  NAND2_X1 U6428 ( .A1(n5410), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5433) );
  AOI22_X1 U6429 ( .A1(n8304), .A2(n9864), .B1(n8275), .B2(n8274), .ZN(n8276)
         );
  NAND2_X1 U6430 ( .A1(n7477), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U6431 ( .A1(n7071), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7141) );
  INV_X1 U6432 ( .A(n7955), .ZN(n7956) );
  NAND2_X1 U6433 ( .A1(n7542), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7555) );
  OR2_X1 U6434 ( .A1(n7251), .A2(n7250), .ZN(n7409) );
  OR2_X1 U6435 ( .A1(n7520), .A2(n10225), .ZN(n7522) );
  OR2_X1 U6436 ( .A1(n7421), .A2(n7420), .ZN(n7486) );
  NAND2_X1 U6437 ( .A1(n7056), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7072) );
  INV_X1 U6438 ( .A(n9147), .ZN(n7620) );
  XNOR2_X1 U6439 ( .A(n9024), .B(n6819), .ZN(n6809) );
  NAND2_X1 U6440 ( .A1(n5327), .A2(n5326), .ZN(n5348) );
  INV_X1 U6441 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5929) );
  OR2_X1 U6442 ( .A1(n5631), .A2(n5630), .ZN(n5647) );
  OR2_X1 U6443 ( .A1(n5780), .A2(n5779), .ZN(n5781) );
  NAND2_X1 U6444 ( .A1(n5645), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U6445 ( .A1(n6161), .A2(n6160), .ZN(n6159) );
  OR2_X1 U6446 ( .A1(n5189), .A2(n6540), .ZN(n5126) );
  INV_X1 U6447 ( .A(n8471), .ZN(n8293) );
  INV_X1 U6448 ( .A(n8488), .ZN(n8260) );
  INV_X1 U6449 ( .A(n7858), .ZN(n7438) );
  NAND2_X1 U6450 ( .A1(n5285), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5313) );
  OR2_X1 U6451 ( .A1(n6157), .A2(n9894), .ZN(n6538) );
  INV_X1 U6452 ( .A(n9971), .ZN(n9962) );
  NAND2_X1 U6453 ( .A1(n6465), .A2(n6505), .ZN(n6506) );
  NAND2_X1 U6454 ( .A1(n7563), .A2(n4475), .ZN(n7565) );
  OR2_X1 U6455 ( .A1(n6270), .A2(n7456), .ZN(n8648) );
  NAND2_X1 U6456 ( .A1(n6271), .A2(n7456), .ZN(n8710) );
  NAND2_X1 U6457 ( .A1(n8614), .A2(n8615), .ZN(n8613) );
  OR2_X1 U6458 ( .A1(n8012), .A2(n7623), .ZN(n7609) );
  INV_X1 U6459 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7302) );
  AND2_X1 U6460 ( .A1(n8795), .A2(n8964), .ZN(n8927) );
  NAND2_X1 U6461 ( .A1(n8971), .A2(n8750), .ZN(n6634) );
  AND2_X1 U6462 ( .A1(n6566), .A2(n6733), .ZN(n9782) );
  INV_X1 U6463 ( .A(n9776), .ZN(n9509) );
  AND2_X1 U6464 ( .A1(n6470), .A2(n9793), .ZN(n6560) );
  OR2_X1 U6465 ( .A1(n8921), .A2(n9001), .ZN(n6787) );
  AND2_X1 U6466 ( .A1(n8088), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8051) );
  AND3_X1 U6467 ( .A1(n5553), .A2(n5552), .A3(n5551), .ZN(n8418) );
  INV_X1 U6468 ( .A(n9852), .ZN(n9477) );
  INV_X1 U6469 ( .A(n9854), .ZN(n9849) );
  INV_X1 U6470 ( .A(n9579), .ZN(n9864) );
  NOR2_X1 U6471 ( .A1(n5765), .A2(n9889), .ZN(n6369) );
  AND2_X1 U6472 ( .A1(n8453), .A2(n8452), .ZN(n8526) );
  AND2_X1 U6473 ( .A1(n6357), .A2(n6356), .ZN(n6370) );
  AND2_X1 U6474 ( .A1(n5768), .A2(n5754), .ZN(n9885) );
  AND2_X1 U6475 ( .A1(n5742), .A2(n5093), .ZN(n5768) );
  XNOR2_X1 U6476 ( .A(n5836), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7006) );
  AND2_X1 U6477 ( .A1(n7603), .A2(n7591), .ZN(n9156) );
  AND2_X1 U6478 ( .A1(n6476), .A2(n6475), .ZN(n8715) );
  AND2_X1 U6479 ( .A1(n7609), .A2(n7608), .ZN(n9150) );
  AND4_X1 U6480 ( .A1(n7484), .A2(n7483), .A3(n7482), .A4(n7481), .ZN(n9264)
         );
  AND2_X1 U6481 ( .A1(n5977), .A2(n7456), .ZN(n9740) );
  INV_X1 U6482 ( .A(n9740), .ZN(n9713) );
  INV_X1 U6483 ( .A(n9735), .ZN(n9749) );
  INV_X1 U6484 ( .A(n9252), .ZN(n9253) );
  AND2_X1 U6485 ( .A1(n7456), .A2(n8927), .ZN(n9507) );
  AND2_X1 U6486 ( .A1(n8828), .A2(n8829), .ZN(n8952) );
  AND2_X1 U6487 ( .A1(n9793), .A2(n8992), .ZN(n6222) );
  AND2_X1 U6488 ( .A1(n9455), .A2(n6559), .ZN(n6234) );
  AND2_X1 U6489 ( .A1(n9779), .A2(n6787), .ZN(n9434) );
  AND3_X1 U6490 ( .A1(n6560), .A2(n6233), .A3(n6232), .ZN(n6242) );
  AND2_X1 U6491 ( .A1(n7006), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6016) );
  INV_X1 U6492 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10090) );
  INV_X1 U6493 ( .A(n9488), .ZN(n9857) );
  AND2_X1 U6494 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  INV_X1 U6495 ( .A(n8106), .ZN(n8058) );
  INV_X1 U6496 ( .A(n8098), .ZN(n8063) );
  NAND2_X1 U6497 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  NAND2_X1 U6498 ( .A1(n5734), .A2(n5733), .ZN(n8304) );
  INV_X1 U6499 ( .A(n8038), .ZN(n8397) );
  INV_X1 U6500 ( .A(n9850), .ZN(n8227) );
  NAND2_X1 U6501 ( .A1(n5877), .A2(n9871), .ZN(n9591) );
  INV_X1 U6502 ( .A(n9591), .ZN(n9593) );
  INV_X1 U6503 ( .A(n9591), .ZN(n9884) );
  NAND2_X1 U6504 ( .A1(n9591), .A2(n6419), .ZN(n8458) );
  INV_X1 U6505 ( .A(n9995), .ZN(n9993) );
  NOR2_X1 U6506 ( .A1(n9886), .A2(n9885), .ZN(n9887) );
  INV_X1 U6507 ( .A(n9887), .ZN(n9890) );
  INV_X1 U6508 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10201) );
  INV_X1 U6509 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6417) );
  INV_X1 U6510 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6031) );
  INV_X1 U6511 ( .A(n7096), .ZN(n9829) );
  INV_X1 U6512 ( .A(n8692), .ZN(n8654) );
  INV_X1 U6513 ( .A(n8645), .ZN(n8719) );
  INV_X1 U6514 ( .A(n9166), .ZN(n9012) );
  INV_X1 U6515 ( .A(n8591), .ZN(n9277) );
  OR2_X1 U6516 ( .A1(P1_U3083), .A2(n5976), .ZN(n9735) );
  NAND2_X1 U6517 ( .A1(n9786), .A2(n6734), .ZN(n9335) );
  AND2_X1 U6519 ( .A1(n9793), .A2(n9792), .ZN(n9794) );
  INV_X1 U6520 ( .A(n9794), .ZN(n10024) );
  INV_X1 U6521 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10234) );
  INV_X1 U6522 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6028) );
  NOR2_X1 U6523 ( .A1(n10408), .A2(n10407), .ZN(n10406) );
  NOR2_X1 U6524 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  INV_X1 U6525 ( .A(n8123), .ZN(P2_U3966) );
  OR2_X1 U6526 ( .A1(n5811), .A2(n5810), .ZN(P2_U3242) );
  NOR2_X1 U6527 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5066) );
  INV_X2 U6528 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5378) );
  INV_X1 U6529 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5072) );
  NAND4_X1 U6530 ( .A1(n5101), .A2(n5751), .A3(n5739), .A4(n5072), .ZN(n5074)
         );
  NAND4_X1 U6531 ( .A1(n5747), .A2(n5104), .A3(n5771), .A4(n5100), .ZN(n5073)
         );
  INV_X1 U6532 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5077) );
  XNOR2_X2 U6533 ( .A(n5078), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U6534 ( .A1(n5079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5080) );
  INV_X1 U6535 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5082) );
  INV_X1 U6536 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6514) );
  NAND2_X2 U6537 ( .A1(n8547), .A2(n7643), .ZN(n5310) );
  INV_X1 U6538 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5085) );
  INV_X1 U6539 ( .A(n9861), .ZN(n5098) );
  INV_X1 U6540 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5090) );
  AND2_X1 U6541 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U6542 ( .A1(n5092), .A2(n5115), .ZN(n8549) );
  NAND2_X1 U6543 ( .A1(n5093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5094) );
  INV_X1 U6544 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5096) );
  MUX2_X1 U6545 ( .A(n5098), .B(n8549), .S(n6077), .Z(n9894) );
  INV_X1 U6546 ( .A(n9894), .ZN(n6516) );
  INV_X1 U6547 ( .A(n5101), .ZN(n5102) );
  OR2_X1 U6548 ( .A1(n5103), .A2(n8542), .ZN(n5105) );
  NAND2_X1 U6549 ( .A1(n5774), .A2(n7669), .ZN(n9895) );
  INV_X1 U6550 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6551 ( .A1(n5112), .A2(n5108), .ZN(n5109) );
  NAND2_X1 U6552 ( .A1(n5109), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5111) );
  INV_X1 U6553 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5110) );
  INV_X1 U6554 ( .A(n5774), .ZN(n7879) );
  NAND2_X1 U6555 ( .A1(n7879), .A2(n9573), .ZN(n7869) );
  NAND3_X1 U6556 ( .A1(n7869), .A2(n9895), .A3(n7669), .ZN(n5113) );
  NAND2_X1 U6557 ( .A1(n7871), .A2(n7840), .ZN(n5878) );
  AND2_X4 U6558 ( .A1(n5113), .A2(n5878), .ZN(n5735) );
  NAND2_X1 U6559 ( .A1(n5735), .A2(n9894), .ZN(n5114) );
  NAND2_X2 U6560 ( .A1(n6077), .A2(n4659), .ZN(n5279) );
  INV_X1 U6561 ( .A(SI_1_), .ZN(n5116) );
  MUX2_X1 U6562 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5164), .Z(n5133) );
  XNOR2_X1 U6563 ( .A(n5134), .B(n5133), .ZN(n6254) );
  OR2_X1 U6564 ( .A1(n5279), .A2(n6254), .ZN(n5123) );
  INV_X1 U6565 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5987) );
  OR2_X1 U6566 ( .A1(n7681), .A2(n5987), .ZN(n5122) );
  NAND2_X1 U6567 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n9861), .ZN(n5117) );
  MUX2_X1 U6568 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5117), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5120) );
  INV_X1 U6569 ( .A(n5118), .ZN(n5119) );
  NAND2_X1 U6570 ( .A1(n5120), .A2(n5119), .ZN(n6106) );
  OR2_X1 U6571 ( .A1(n6077), .A2(n6106), .ZN(n5121) );
  AND3_X2 U6572 ( .A1(n5123), .A2(n5122), .A3(n5121), .ZN(n6535) );
  NAND2_X1 U6573 ( .A1(n5309), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5128) );
  INV_X1 U6574 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6534) );
  INV_X1 U6575 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6540) );
  INV_X1 U6576 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5124) );
  OR2_X1 U6577 ( .A1(n5310), .A2(n5124), .ZN(n5125) );
  NAND4_X1 U6578 ( .A1(n5128), .A2(n5127), .A3(n5126), .A4(n5125), .ZN(n6495)
         );
  NAND2_X1 U6579 ( .A1(n6495), .A2(n7690), .ZN(n5131) );
  XNOR2_X1 U6580 ( .A(n5129), .B(n5131), .ZN(n6160) );
  INV_X1 U6581 ( .A(n5129), .ZN(n5130) );
  NAND2_X1 U6582 ( .A1(n5131), .A2(n5130), .ZN(n5132) );
  AND2_X1 U6583 ( .A1(n6159), .A2(n5132), .ZN(n8086) );
  NAND2_X1 U6584 ( .A1(n5135), .A2(SI_1_), .ZN(n5136) );
  NAND2_X1 U6585 ( .A1(n5137), .A2(n5136), .ZN(n5159) );
  INV_X1 U6586 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5990) );
  INV_X1 U6587 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5138) );
  MUX2_X1 U6588 ( .A(n5990), .B(n5138), .S(n5164), .Z(n5160) );
  XNOR2_X1 U6589 ( .A(n5160), .B(SI_2_), .ZN(n5158) );
  XNOR2_X1 U6590 ( .A(n5159), .B(n5158), .ZN(n6321) );
  OR2_X1 U6591 ( .A1(n5279), .A2(n6321), .ZN(n5143) );
  OR2_X1 U6592 ( .A1(n7681), .A2(n5990), .ZN(n5142) );
  OR2_X1 U6593 ( .A1(n5118), .A2(n8542), .ZN(n5140) );
  INV_X1 U6594 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5139) );
  XNOR2_X1 U6595 ( .A(n5140), .B(n5139), .ZN(n9492) );
  OR2_X1 U6596 ( .A1(n6077), .A2(n9492), .ZN(n5141) );
  XNOR2_X1 U6597 ( .A(n9908), .B(n5228), .ZN(n6171) );
  NAND2_X1 U6598 ( .A1(n5309), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5149) );
  INV_X1 U6599 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6105) );
  OR2_X1 U6600 ( .A1(n5189), .A2(n6105), .ZN(n5148) );
  INV_X1 U6601 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5144) );
  INV_X1 U6602 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5145) );
  OR2_X1 U6603 ( .A1(n5706), .A2(n5145), .ZN(n5146) );
  NAND2_X1 U6604 ( .A1(n6158), .A2(n7690), .ZN(n5150) );
  OR2_X1 U6605 ( .A1(n6171), .A2(n5150), .ZN(n5152) );
  NAND2_X1 U6606 ( .A1(n5150), .A2(n6171), .ZN(n5151) );
  NAND2_X1 U6607 ( .A1(n8086), .A2(n8085), .ZN(n6172) );
  NAND2_X1 U6608 ( .A1(n6172), .A2(n5152), .ZN(n5174) );
  NAND2_X1 U6609 ( .A1(n5309), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5157) );
  OR2_X1 U6610 ( .A1(n5706), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5156) );
  INV_X1 U6611 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6104) );
  OR2_X1 U6612 ( .A1(n5189), .A2(n6104), .ZN(n5155) );
  INV_X1 U6613 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5153) );
  OR2_X1 U6614 ( .A1(n5310), .A2(n5153), .ZN(n5154) );
  NAND4_X2 U6615 ( .A1(n5157), .A2(n5156), .A3(n5155), .A4(n5154), .ZN(n5855)
         );
  AND2_X1 U6616 ( .A1(n5855), .A2(n7690), .ZN(n5170) );
  NAND2_X1 U6617 ( .A1(n5159), .A2(n5158), .ZN(n5163) );
  INV_X1 U6618 ( .A(n5160), .ZN(n5161) );
  NAND2_X1 U6619 ( .A1(n5161), .A2(SI_2_), .ZN(n5162) );
  NAND2_X1 U6620 ( .A1(n5163), .A2(n5162), .ZN(n5176) );
  INV_X1 U6621 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5989) );
  INV_X1 U6622 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5165) );
  MUX2_X1 U6623 ( .A(n5989), .B(n5165), .S(n5164), .Z(n5177) );
  XNOR2_X1 U6624 ( .A(n5177), .B(SI_3_), .ZN(n5175) );
  XNOR2_X1 U6625 ( .A(n5176), .B(n5175), .ZN(n6458) );
  OR2_X1 U6626 ( .A1(n5279), .A2(n6458), .ZN(n5169) );
  OR2_X1 U6627 ( .A1(n7681), .A2(n5989), .ZN(n5168) );
  NAND2_X1 U6628 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4508), .ZN(n5166) );
  XNOR2_X1 U6629 ( .A(n5166), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8130) );
  INV_X1 U6630 ( .A(n8130), .ZN(n5988) );
  OR2_X1 U6631 ( .A1(n6077), .A2(n5988), .ZN(n5167) );
  AND3_X2 U6632 ( .A1(n5169), .A2(n5168), .A3(n5167), .ZN(n9914) );
  XNOR2_X1 U6633 ( .A(n5735), .B(n9914), .ZN(n5171) );
  NAND2_X1 U6634 ( .A1(n5170), .A2(n5171), .ZN(n5194) );
  INV_X1 U6635 ( .A(n5170), .ZN(n5172) );
  INV_X1 U6636 ( .A(n5171), .ZN(n8069) );
  NAND2_X1 U6637 ( .A1(n5172), .A2(n8069), .ZN(n5173) );
  AND2_X1 U6638 ( .A1(n5194), .A2(n5173), .ZN(n6173) );
  NAND2_X1 U6639 ( .A1(n5176), .A2(n5175), .ZN(n5180) );
  INV_X1 U6640 ( .A(n5177), .ZN(n5178) );
  NAND2_X1 U6641 ( .A1(n5178), .A2(SI_3_), .ZN(n5179) );
  INV_X1 U6642 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5181) );
  XNOR2_X1 U6643 ( .A(n5201), .B(SI_4_), .ZN(n5199) );
  XNOR2_X1 U6644 ( .A(n5200), .B(n5199), .ZN(n6452) );
  OR2_X1 U6645 ( .A1(n6452), .A2(n5279), .ZN(n5188) );
  INV_X2 U6646 ( .A(n7681), .ZN(n5543) );
  INV_X2 U6647 ( .A(n6077), .ZN(n6010) );
  NOR2_X1 U6648 ( .A1(n5184), .A2(n8542), .ZN(n5182) );
  MUX2_X1 U6649 ( .A(n8542), .B(n5182), .S(P2_IR_REG_4__SCAN_IN), .Z(n5186) );
  NAND2_X1 U6650 ( .A1(n5184), .A2(n5183), .ZN(n5224) );
  INV_X1 U6651 ( .A(n5224), .ZN(n5185) );
  NOR2_X1 U6652 ( .A1(n5186), .A2(n5185), .ZN(n8143) );
  AND2_X2 U6653 ( .A1(n5188), .A2(n5187), .ZN(n9919) );
  XNOR2_X1 U6654 ( .A(n9919), .B(n5735), .ZN(n5196) );
  INV_X2 U6655 ( .A(n5310), .ZN(n7664) );
  NAND2_X1 U6656 ( .A1(n7664), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5193) );
  INV_X1 U6657 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6079) );
  OR2_X1 U6658 ( .A1(n7668), .A2(n6079), .ZN(n5192) );
  INV_X1 U6659 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6109) );
  XNOR2_X1 U6660 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9872) );
  OR2_X1 U6661 ( .A1(n5706), .A2(n9872), .ZN(n5190) );
  NAND2_X1 U6662 ( .A1(n8122), .A2(n7690), .ZN(n5197) );
  XNOR2_X1 U6663 ( .A(n5196), .B(n5197), .ZN(n8068) );
  INV_X1 U6664 ( .A(n5196), .ZN(n5198) );
  INV_X1 U6665 ( .A(n5201), .ZN(n5202) );
  INV_X1 U6666 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5204) );
  INV_X1 U6667 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5203) );
  XNOR2_X1 U6668 ( .A(n5221), .B(SI_5_), .ZN(n5220) );
  OR2_X1 U6669 ( .A1(n6642), .A2(n5279), .ZN(n5207) );
  NAND2_X1 U6670 ( .A1(n5224), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5205) );
  XNOR2_X1 U6671 ( .A(n5205), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8155) );
  AOI22_X1 U6672 ( .A1(n5543), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6010), .B2(
        n8155), .ZN(n5206) );
  XNOR2_X1 U6673 ( .A(n5880), .B(n5735), .ZN(n5214) );
  NAND2_X1 U6674 ( .A1(n7664), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5213) );
  INV_X1 U6675 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5208) );
  OR2_X1 U6676 ( .A1(n7668), .A2(n5208), .ZN(n5212) );
  INV_X1 U6677 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6552) );
  NAND3_X1 U6678 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5230) );
  INV_X1 U6679 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U6680 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5209) );
  NAND2_X1 U6681 ( .A1(n6137), .A2(n5209), .ZN(n5210) );
  NAND2_X1 U6682 ( .A1(n5230), .A2(n5210), .ZN(n6553) );
  OR2_X1 U6683 ( .A1(n5706), .A2(n6553), .ZN(n5211) );
  AND2_X1 U6684 ( .A1(n9866), .A2(n7690), .ZN(n5215) );
  NAND2_X1 U6685 ( .A1(n5214), .A2(n5215), .ZN(n5236) );
  INV_X1 U6686 ( .A(n5214), .ZN(n8104) );
  INV_X1 U6687 ( .A(n5215), .ZN(n5216) );
  NAND2_X1 U6688 ( .A1(n8104), .A2(n5216), .ZN(n5217) );
  NAND2_X1 U6689 ( .A1(n5236), .A2(n5217), .ZN(n6139) );
  INV_X1 U6690 ( .A(n6139), .ZN(n5218) );
  INV_X1 U6691 ( .A(n5221), .ZN(n5222) );
  INV_X1 U6692 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5223) );
  XNOR2_X1 U6693 ( .A(n5244), .B(SI_6_), .ZN(n5242) );
  XNOR2_X1 U6694 ( .A(n5243), .B(n5242), .ZN(n6656) );
  OR2_X1 U6695 ( .A1(n6656), .A2(n5279), .ZN(n5227) );
  NAND2_X1 U6696 ( .A1(n5249), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5225) );
  XNOR2_X1 U6697 ( .A(n5225), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8167) );
  AOI22_X1 U6698 ( .A1(n5543), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6010), .B2(
        n8167), .ZN(n5226) );
  NAND2_X1 U6699 ( .A1(n5227), .A2(n5226), .ZN(n9926) );
  XNOR2_X1 U6700 ( .A(n9926), .B(n5702), .ZN(n5238) );
  NAND2_X1 U6701 ( .A1(n7664), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5235) );
  INV_X1 U6702 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6089) );
  OR2_X1 U6703 ( .A1(n7668), .A2(n6089), .ZN(n5234) );
  INV_X1 U6704 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6437) );
  OR2_X1 U6705 ( .A1(n5189), .A2(n6437), .ZN(n5233) );
  INV_X1 U6706 ( .A(n5230), .ZN(n5229) );
  NAND2_X1 U6707 ( .A1(n5229), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5256) );
  INV_X1 U6708 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10287) );
  NAND2_X1 U6709 ( .A1(n5230), .A2(n10287), .ZN(n5231) );
  NAND2_X1 U6710 ( .A1(n5256), .A2(n5231), .ZN(n8093) );
  OR2_X1 U6711 ( .A1(n5706), .A2(n8093), .ZN(n5232) );
  NAND4_X1 U6712 ( .A1(n5235), .A2(n5234), .A3(n5233), .A4(n5232), .ZN(n8121)
         );
  NAND2_X1 U6713 ( .A1(n8121), .A2(n7690), .ZN(n5239) );
  XNOR2_X1 U6714 ( .A(n5238), .B(n5239), .ZN(n8103) );
  AND2_X1 U6715 ( .A1(n8103), .A2(n5236), .ZN(n5237) );
  NAND2_X1 U6716 ( .A1(n8100), .A2(n5237), .ZN(n8099) );
  INV_X1 U6717 ( .A(n5238), .ZN(n5240) );
  NAND2_X1 U6718 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NAND2_X1 U6719 ( .A1(n8099), .A2(n5241), .ZN(n5891) );
  INV_X1 U6720 ( .A(n5891), .ZN(n5267) );
  NAND2_X1 U6721 ( .A1(n5243), .A2(n5242), .ZN(n5247) );
  INV_X1 U6722 ( .A(n5244), .ZN(n5245) );
  NAND2_X1 U6723 ( .A1(n5245), .A2(SI_6_), .ZN(n5246) );
  NAND2_X1 U6724 ( .A1(n5247), .A2(n5246), .ZN(n5270) );
  INV_X1 U6725 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5248) );
  XNOR2_X1 U6726 ( .A(n5271), .B(SI_7_), .ZN(n5269) );
  XNOR2_X1 U6727 ( .A(n5270), .B(n5269), .ZN(n6739) );
  OR2_X1 U6728 ( .A1(n6739), .A2(n5279), .ZN(n5252) );
  OR2_X1 U6729 ( .A1(n5281), .A2(n8542), .ZN(n5250) );
  XNOR2_X1 U6730 ( .A(n5250), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8179) );
  AOI22_X1 U6731 ( .A1(n5543), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6010), .B2(
        n8179), .ZN(n5251) );
  NAND2_X1 U6732 ( .A1(n5252), .A2(n5251), .ZN(n9933) );
  XNOR2_X1 U6733 ( .A(n9933), .B(n5702), .ZN(n6591) );
  NAND2_X1 U6734 ( .A1(n7664), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5261) );
  INV_X1 U6735 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5253) );
  OR2_X1 U6736 ( .A1(n7668), .A2(n5253), .ZN(n5260) );
  INV_X1 U6737 ( .A(n5256), .ZN(n5254) );
  NAND2_X1 U6738 ( .A1(n5254), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5287) );
  INV_X1 U6739 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6740 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  NAND2_X1 U6741 ( .A1(n5287), .A2(n5257), .ZN(n6426) );
  OR2_X1 U6742 ( .A1(n5706), .A2(n6426), .ZN(n5259) );
  INV_X1 U6743 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6425) );
  OR2_X1 U6744 ( .A1(n5189), .A2(n6425), .ZN(n5258) );
  NOR2_X1 U6745 ( .A1(n8095), .A2(n6170), .ZN(n5262) );
  NAND2_X1 U6746 ( .A1(n6591), .A2(n5262), .ZN(n5268) );
  INV_X1 U6747 ( .A(n6591), .ZN(n5264) );
  INV_X1 U6748 ( .A(n5262), .ZN(n5263) );
  NAND2_X1 U6749 ( .A1(n5264), .A2(n5263), .ZN(n5265) );
  NAND2_X1 U6750 ( .A1(n5268), .A2(n5265), .ZN(n5890) );
  NAND2_X1 U6751 ( .A1(n5270), .A2(n5269), .ZN(n5274) );
  INV_X1 U6752 ( .A(n5271), .ZN(n5272) );
  NAND2_X1 U6753 ( .A1(n5272), .A2(SI_7_), .ZN(n5273) );
  INV_X1 U6754 ( .A(SI_8_), .ZN(n5275) );
  INV_X1 U6755 ( .A(n5276), .ZN(n5277) );
  NAND2_X1 U6756 ( .A1(n5277), .A2(SI_8_), .ZN(n5278) );
  NAND2_X1 U6757 ( .A1(n5299), .A2(n5278), .ZN(n5297) );
  NAND2_X1 U6758 ( .A1(n6750), .A2(n7680), .ZN(n5284) );
  INV_X1 U6759 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6760 ( .A1(n5281), .A2(n5280), .ZN(n5306) );
  NAND2_X1 U6761 ( .A1(n5306), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5282) );
  XNOR2_X1 U6762 ( .A(n5282), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8192) );
  AOI22_X1 U6763 ( .A1(n5543), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6010), .B2(
        n8192), .ZN(n5283) );
  XNOR2_X1 U6764 ( .A(n6681), .B(n5702), .ZN(n5293) );
  NAND2_X1 U6765 ( .A1(n7664), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5292) );
  INV_X1 U6766 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6093) );
  OR2_X1 U6767 ( .A1(n7668), .A2(n6093), .ZN(n5291) );
  INV_X1 U6768 ( .A(n5287), .ZN(n5285) );
  INV_X1 U6769 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6770 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  NAND2_X1 U6771 ( .A1(n5313), .A2(n5288), .ZN(n6590) );
  OR2_X1 U6772 ( .A1(n5706), .A2(n6590), .ZN(n5290) );
  INV_X1 U6773 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6114) );
  OR2_X1 U6774 ( .A1(n5189), .A2(n6114), .ZN(n5289) );
  NOR2_X1 U6775 ( .A1(n6620), .A2(n6170), .ZN(n5294) );
  NAND2_X1 U6776 ( .A1(n5293), .A2(n5294), .ZN(n5319) );
  INV_X1 U6777 ( .A(n5293), .ZN(n6618) );
  INV_X1 U6778 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U6779 ( .A1(n6618), .A2(n5295), .ZN(n5296) );
  AND2_X1 U6780 ( .A1(n5319), .A2(n5296), .ZN(n6592) );
  INV_X1 U6781 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5301) );
  INV_X1 U6782 ( .A(SI_9_), .ZN(n5302) );
  INV_X1 U6783 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6784 ( .A1(n5304), .A2(SI_9_), .ZN(n5305) );
  XNOR2_X1 U6785 ( .A(n5324), .B(n5061), .ZN(n6980) );
  NAND2_X1 U6786 ( .A1(n6980), .A2(n7680), .ZN(n5308) );
  NAND2_X1 U6787 ( .A1(n5380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5330) );
  XNOR2_X1 U6788 ( .A(n5330), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6128) );
  AOI22_X1 U6789 ( .A1(n5543), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6010), .B2(
        n6128), .ZN(n5307) );
  NAND2_X1 U6790 ( .A1(n5308), .A2(n5307), .ZN(n6711) );
  XNOR2_X1 U6791 ( .A(n6711), .B(n5735), .ZN(n5323) );
  NAND2_X1 U6792 ( .A1(n5787), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5318) );
  INV_X1 U6793 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5311) );
  OR2_X1 U6794 ( .A1(n5310), .A2(n5311), .ZN(n5317) );
  NAND2_X1 U6795 ( .A1(n5313), .A2(n5312), .ZN(n5314) );
  NAND2_X1 U6796 ( .A1(n5334), .A2(n5314), .ZN(n6691) );
  OR2_X1 U6797 ( .A1(n5706), .A2(n6691), .ZN(n5316) );
  INV_X1 U6798 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6692) );
  OR2_X1 U6799 ( .A1(n5189), .A2(n6692), .ZN(n5315) );
  NOR2_X1 U6800 ( .A1(n6680), .A2(n6170), .ZN(n5321) );
  XNOR2_X1 U6801 ( .A(n5323), .B(n5321), .ZN(n6630) );
  AND2_X1 U6802 ( .A1(n6630), .A2(n5319), .ZN(n5320) );
  INV_X1 U6803 ( .A(n5321), .ZN(n5322) );
  INV_X1 U6804 ( .A(n5897), .ZN(n5345) );
  INV_X1 U6805 ( .A(SI_10_), .ZN(n5326) );
  INV_X1 U6806 ( .A(n5327), .ZN(n5328) );
  NAND2_X1 U6807 ( .A1(n5328), .A2(SI_10_), .ZN(n5329) );
  XNOR2_X1 U6808 ( .A(n5347), .B(n5058), .ZN(n7048) );
  NAND2_X1 U6809 ( .A1(n7048), .A2(n7680), .ZN(n5333) );
  NAND2_X1 U6810 ( .A1(n5330), .A2(n5378), .ZN(n5331) );
  NAND2_X1 U6811 ( .A1(n5331), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5351) );
  XNOR2_X1 U6812 ( .A(n5351), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6290) );
  AOI22_X1 U6813 ( .A1(n5543), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6290), .B2(
        n6010), .ZN(n5332) );
  XNOR2_X1 U6814 ( .A(n6825), .B(n5702), .ZN(n5340) );
  NAND2_X1 U6815 ( .A1(n7664), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5339) );
  INV_X1 U6816 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6123) );
  OR2_X1 U6817 ( .A1(n7668), .A2(n6123), .ZN(n5338) );
  NAND2_X1 U6818 ( .A1(n5334), .A2(n10102), .ZN(n5335) );
  NAND2_X1 U6819 ( .A1(n5388), .A2(n5335), .ZN(n6724) );
  OR2_X1 U6820 ( .A1(n5706), .A2(n6724), .ZN(n5337) );
  INV_X1 U6821 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6725) );
  OR2_X1 U6822 ( .A1(n5189), .A2(n6725), .ZN(n5336) );
  NOR2_X1 U6823 ( .A1(n6714), .A2(n6170), .ZN(n5341) );
  NAND2_X1 U6824 ( .A1(n5340), .A2(n5341), .ZN(n5346) );
  INV_X1 U6825 ( .A(n5340), .ZN(n6702) );
  INV_X1 U6826 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6827 ( .A1(n6702), .A2(n5342), .ZN(n5343) );
  NAND2_X1 U6828 ( .A1(n5346), .A2(n5343), .ZN(n5898) );
  INV_X1 U6829 ( .A(n5898), .ZN(n5344) );
  NAND2_X1 U6830 ( .A1(n6701), .A2(n5346), .ZN(n5360) );
  INV_X1 U6831 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6832 ( .A1(n7053), .A2(n7680), .ZN(n5355) );
  INV_X1 U6833 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6834 ( .A1(n5351), .A2(n5377), .ZN(n5352) );
  NAND2_X1 U6835 ( .A1(n5352), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5353) );
  XNOR2_X1 U6836 ( .A(n5353), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6306) );
  AOI22_X1 U6837 ( .A1(n6010), .A2(n6306), .B1(n5543), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5354) );
  XNOR2_X1 U6838 ( .A(n9961), .B(n5735), .ZN(n5361) );
  NAND2_X1 U6839 ( .A1(n7664), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5359) );
  INV_X1 U6840 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6288) );
  OR2_X1 U6841 ( .A1(n7668), .A2(n6288), .ZN(n5358) );
  INV_X1 U6842 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6706) );
  XNOR2_X1 U6843 ( .A(n5388), .B(n6706), .ZN(n6837) );
  OR2_X1 U6844 ( .A1(n5706), .A2(n6837), .ZN(n5357) );
  INV_X1 U6845 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6838) );
  OR2_X1 U6846 ( .A1(n5189), .A2(n6838), .ZN(n5356) );
  NOR2_X1 U6847 ( .A1(n6828), .A2(n6170), .ZN(n5362) );
  XNOR2_X1 U6848 ( .A(n5361), .B(n5362), .ZN(n6699) );
  INV_X1 U6849 ( .A(n5361), .ZN(n5363) );
  NAND2_X1 U6850 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  INV_X1 U6851 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6852 ( .A1(n5369), .A2(SI_11_), .ZN(n5370) );
  INV_X1 U6853 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5371) );
  MUX2_X1 U6854 ( .A(n6035), .B(n5371), .S(n7677), .Z(n5373) );
  INV_X1 U6855 ( .A(SI_12_), .ZN(n5372) );
  INV_X1 U6856 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6857 ( .A1(n5374), .A2(SI_12_), .ZN(n5375) );
  NAND2_X1 U6858 ( .A1(n5398), .A2(n5375), .ZN(n5399) );
  XNOR2_X1 U6859 ( .A(n5400), .B(n5399), .ZN(n7134) );
  NAND2_X1 U6860 ( .A1(n7134), .A2(n7680), .ZN(n5383) );
  INV_X1 U6861 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5376) );
  NAND3_X1 U6862 ( .A1(n5378), .A2(n5377), .A3(n5376), .ZN(n5379) );
  NAND2_X1 U6863 ( .A1(n5406), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5381) );
  XNOR2_X1 U6864 ( .A(n5381), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8207) );
  AOI22_X1 U6865 ( .A1(n5543), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6010), .B2(
        n8207), .ZN(n5382) );
  XNOR2_X1 U6866 ( .A(n7111), .B(n5735), .ZN(n5394) );
  NAND2_X1 U6867 ( .A1(n7665), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5393) );
  INV_X1 U6868 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5384) );
  OR2_X1 U6869 ( .A1(n5310), .A2(n5384), .ZN(n5392) );
  INV_X1 U6870 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6307) );
  OR2_X1 U6871 ( .A1(n7668), .A2(n6307), .ZN(n5391) );
  AND2_X1 U6872 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5385) );
  INV_X1 U6873 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5387) );
  OAI21_X1 U6874 ( .B1(n5388), .B2(n6706), .A(n5387), .ZN(n5389) );
  NAND2_X1 U6875 ( .A1(n5412), .A2(n5389), .ZN(n6952) );
  OR2_X1 U6876 ( .A1(n5706), .A2(n6952), .ZN(n5390) );
  OR2_X1 U6877 ( .A1(n7115), .A2(n6170), .ZN(n5395) );
  NAND2_X1 U6878 ( .A1(n5394), .A2(n5395), .ZN(n6844) );
  INV_X1 U6879 ( .A(n5394), .ZN(n5397) );
  INV_X1 U6880 ( .A(n5395), .ZN(n5396) );
  NAND2_X1 U6881 ( .A1(n5397), .A2(n5396), .ZN(n6843) );
  INV_X1 U6882 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5401) );
  MUX2_X1 U6883 ( .A(n6058), .B(n5401), .S(n7677), .Z(n5403) );
  INV_X1 U6884 ( .A(SI_13_), .ZN(n5402) );
  INV_X1 U6885 ( .A(n5403), .ZN(n5404) );
  NAND2_X1 U6886 ( .A1(n5404), .A2(SI_13_), .ZN(n5405) );
  XNOR2_X1 U6887 ( .A(n5423), .B(n5062), .ZN(n7213) );
  NAND2_X1 U6888 ( .A1(n7213), .A2(n7680), .ZN(n5408) );
  OAI21_X1 U6889 ( .B1(n5406), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5427) );
  XNOR2_X1 U6890 ( .A(n5427), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6407) );
  AOI22_X1 U6891 ( .A1(n6010), .A2(n6407), .B1(n5543), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5407) );
  XNOR2_X1 U6892 ( .A(n9615), .B(n5735), .ZN(n5418) );
  NAND2_X1 U6893 ( .A1(n7664), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5417) );
  INV_X1 U6894 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5409) );
  OR2_X1 U6895 ( .A1(n7668), .A2(n5409), .ZN(n5416) );
  INV_X1 U6896 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6897 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  NAND2_X1 U6898 ( .A1(n5433), .A2(n5413), .ZN(n7123) );
  OR2_X1 U6899 ( .A1(n5706), .A2(n7123), .ZN(n5415) );
  INV_X1 U6900 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7124) );
  OR2_X1 U6901 ( .A1(n5189), .A2(n7124), .ZN(n5414) );
  NOR2_X1 U6902 ( .A1(n7114), .A2(n6170), .ZN(n5419) );
  XNOR2_X1 U6903 ( .A(n5418), .B(n5419), .ZN(n6935) );
  NAND2_X1 U6904 ( .A1(n6934), .A2(n6935), .ZN(n5422) );
  INV_X1 U6905 ( .A(n5418), .ZN(n5420) );
  NAND2_X1 U6906 ( .A1(n5420), .A2(n5419), .ZN(n5421) );
  NAND2_X1 U6907 ( .A1(n5422), .A2(n5421), .ZN(n7085) );
  MUX2_X1 U6908 ( .A(n10243), .B(n6059), .S(n7677), .Z(n5449) );
  XNOR2_X1 U6909 ( .A(n5448), .B(n5446), .ZN(n7239) );
  NAND2_X1 U6910 ( .A1(n7239), .A2(n7680), .ZN(n5430) );
  NAND2_X1 U6911 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  NAND2_X1 U6912 ( .A1(n5428), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5457) );
  XNOR2_X1 U6913 ( .A(n5457), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6925) );
  AOI22_X1 U6914 ( .A1(n6925), .A2(n6010), .B1(n5543), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5429) );
  XNOR2_X1 U6915 ( .A(n9609), .B(n5735), .ZN(n5439) );
  NAND2_X1 U6916 ( .A1(n5787), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5438) );
  INV_X1 U6917 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5431) );
  OR2_X1 U6918 ( .A1(n5310), .A2(n5431), .ZN(n5437) );
  INV_X1 U6919 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6920 ( .A1(n5433), .A2(n5432), .ZN(n5434) );
  NAND2_X1 U6921 ( .A1(n5464), .A2(n5434), .ZN(n7173) );
  OR2_X1 U6922 ( .A1(n5706), .A2(n7173), .ZN(n5436) );
  INV_X1 U6923 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7174) );
  OR2_X1 U6924 ( .A1(n5189), .A2(n7174), .ZN(n5435) );
  OR2_X1 U6925 ( .A1(n7163), .A2(n6170), .ZN(n5440) );
  NAND2_X1 U6926 ( .A1(n5439), .A2(n5440), .ZN(n5445) );
  INV_X1 U6927 ( .A(n5439), .ZN(n5442) );
  INV_X1 U6928 ( .A(n5440), .ZN(n5441) );
  NAND2_X1 U6929 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  NAND2_X1 U6930 ( .A1(n5445), .A2(n5443), .ZN(n7086) );
  INV_X1 U6931 ( .A(n7086), .ZN(n5444) );
  INV_X1 U6932 ( .A(n5449), .ZN(n5450) );
  NAND2_X1 U6933 ( .A1(n5450), .A2(SI_14_), .ZN(n5451) );
  MUX2_X1 U6934 ( .A(n6181), .B(n6179), .S(n7677), .Z(n5453) );
  INV_X1 U6935 ( .A(SI_15_), .ZN(n5452) );
  NAND2_X1 U6936 ( .A1(n5453), .A2(n5452), .ZN(n5470) );
  INV_X1 U6937 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U6938 ( .A1(n5454), .A2(SI_15_), .ZN(n5455) );
  NAND2_X1 U6939 ( .A1(n5470), .A2(n5455), .ZN(n5471) );
  XNOR2_X1 U6940 ( .A(n5472), .B(n5471), .ZN(n7397) );
  NAND2_X1 U6941 ( .A1(n7397), .A2(n7680), .ZN(n5461) );
  NAND2_X1 U6942 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  NAND2_X1 U6943 ( .A1(n5458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5459) );
  XNOR2_X1 U6944 ( .A(n5459), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6967) );
  AOI22_X1 U6945 ( .A1(n6967), .A2(n6010), .B1(n5543), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5460) );
  XNOR2_X1 U6946 ( .A(n7435), .B(n5735), .ZN(n7289) );
  NAND2_X1 U6947 ( .A1(n7664), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5469) );
  INV_X1 U6948 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5462) );
  OR2_X1 U6949 ( .A1(n7668), .A2(n5462), .ZN(n5468) );
  INV_X1 U6950 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U6951 ( .A1(n5464), .A2(n10279), .ZN(n5465) );
  NAND2_X1 U6952 ( .A1(n5481), .A2(n5465), .ZN(n7296) );
  OR2_X1 U6953 ( .A1(n5706), .A2(n7296), .ZN(n5467) );
  INV_X1 U6954 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7270) );
  OR2_X1 U6955 ( .A1(n5189), .A2(n7270), .ZN(n5466) );
  OR2_X1 U6956 ( .A1(n7443), .A2(n6170), .ZN(n5488) );
  MUX2_X1 U6957 ( .A(n6399), .B(n6397), .S(n7677), .Z(n5474) );
  INV_X1 U6958 ( .A(SI_16_), .ZN(n5473) );
  NAND2_X1 U6959 ( .A1(n5474), .A2(n5473), .ZN(n5498) );
  INV_X1 U6960 ( .A(n5474), .ZN(n5475) );
  NAND2_X1 U6961 ( .A1(n5475), .A2(SI_16_), .ZN(n5476) );
  XNOR2_X1 U6962 ( .A(n5497), .B(n5496), .ZN(n7403) );
  NAND2_X1 U6963 ( .A1(n7403), .A2(n7680), .ZN(n5480) );
  NAND2_X1 U6964 ( .A1(n5477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5478) );
  XNOR2_X1 U6965 ( .A(n5478), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7190) );
  AOI22_X1 U6966 ( .A1(n5543), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6010), .B2(
        n7190), .ZN(n5479) );
  XNOR2_X1 U6967 ( .A(n9599), .B(n5735), .ZN(n5492) );
  INV_X1 U6968 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U6969 ( .A1(n5481), .A2(n6973), .ZN(n5482) );
  AND2_X1 U6970 ( .A1(n5509), .A2(n5482), .ZN(n7447) );
  NAND2_X1 U6971 ( .A1(n5791), .A2(n7447), .ZN(n5487) );
  INV_X1 U6972 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6962) );
  OR2_X1 U6973 ( .A1(n7668), .A2(n6962), .ZN(n5486) );
  INV_X1 U6974 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7449) );
  OR2_X1 U6975 ( .A1(n5189), .A2(n7449), .ZN(n5485) );
  INV_X1 U6976 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5483) );
  OR2_X1 U6977 ( .A1(n5310), .A2(n5483), .ZN(n5484) );
  NAND4_X1 U6978 ( .A1(n5487), .A2(n5486), .A3(n5485), .A4(n5484), .ZN(n8245)
         );
  NAND2_X1 U6979 ( .A1(n8245), .A2(n7690), .ZN(n5493) );
  XNOR2_X1 U6980 ( .A(n5492), .B(n5493), .ZN(n7325) );
  INV_X1 U6981 ( .A(n7289), .ZN(n7291) );
  INV_X1 U6982 ( .A(n5488), .ZN(n7293) );
  NAND2_X1 U6983 ( .A1(n7291), .A2(n7293), .ZN(n5489) );
  AND2_X1 U6984 ( .A1(n7325), .A2(n5489), .ZN(n5490) );
  NAND2_X1 U6985 ( .A1(n5491), .A2(n5490), .ZN(n7328) );
  INV_X1 U6986 ( .A(n5492), .ZN(n5494) );
  NAND2_X1 U6987 ( .A1(n5494), .A2(n5493), .ZN(n5495) );
  INV_X1 U6988 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5500) );
  MUX2_X1 U6989 ( .A(n6417), .B(n5500), .S(n7677), .Z(n5520) );
  NAND2_X1 U6990 ( .A1(n7497), .A2(n7680), .ZN(n5504) );
  NAND2_X1 U6991 ( .A1(n5501), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5502) );
  XNOR2_X1 U6992 ( .A(n5502), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7201) );
  AOI22_X1 U6993 ( .A1(n5543), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6010), .B2(
        n7201), .ZN(n5503) );
  XNOR2_X1 U6994 ( .A(n9568), .B(n5735), .ZN(n5514) );
  INV_X1 U6995 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5505) );
  OR2_X1 U6996 ( .A1(n5310), .A2(n5505), .ZN(n5507) );
  INV_X1 U6997 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7186) );
  OR2_X1 U6998 ( .A1(n7668), .A2(n7186), .ZN(n5506) );
  AND2_X1 U6999 ( .A1(n5507), .A2(n5506), .ZN(n5513) );
  INV_X1 U7000 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7278) );
  NAND2_X1 U7001 ( .A1(n5509), .A2(n7278), .ZN(n5510) );
  NAND2_X1 U7002 ( .A1(n5549), .A2(n5510), .ZN(n9585) );
  OR2_X1 U7003 ( .A1(n9585), .A2(n5706), .ZN(n5512) );
  NAND2_X1 U7004 ( .A1(n7665), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5511) );
  INV_X1 U7005 ( .A(n7649), .ZN(n8450) );
  NAND2_X1 U7006 ( .A1(n8450), .A2(n7690), .ZN(n5515) );
  XNOR2_X1 U7007 ( .A(n5514), .B(n5515), .ZN(n7276) );
  INV_X1 U7008 ( .A(n5514), .ZN(n5517) );
  INV_X1 U7009 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U7010 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  INV_X1 U7011 ( .A(n5520), .ZN(n5521) );
  NAND2_X1 U7012 ( .A1(n5521), .A2(SI_17_), .ZN(n5522) );
  MUX2_X1 U7013 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7677), .Z(n5537) );
  XNOR2_X1 U7014 ( .A(n5536), .B(n5534), .ZN(n7492) );
  NAND2_X1 U7015 ( .A1(n7492), .A2(n7680), .ZN(n5525) );
  OR2_X1 U7016 ( .A1(n5099), .A2(n8542), .ZN(n5523) );
  XNOR2_X1 U7017 ( .A(n5523), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8220) );
  AOI22_X1 U7018 ( .A1(n5543), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6010), .B2(
        n8220), .ZN(n5524) );
  XNOR2_X1 U7019 ( .A(n8523), .B(n5735), .ZN(n5531) );
  XNOR2_X1 U7020 ( .A(n5549), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U7021 ( .A1(n8445), .A2(n5791), .ZN(n5530) );
  INV_X1 U7022 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U7023 ( .A1(n7664), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7024 ( .A1(n7665), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5526) );
  OAI211_X1 U7025 ( .C1(n7668), .C2(n7202), .A(n5527), .B(n5526), .ZN(n5528)
         );
  INV_X1 U7026 ( .A(n5528), .ZN(n5529) );
  NOR2_X1 U7027 ( .A1(n9580), .A2(n6170), .ZN(n5532) );
  XNOR2_X1 U7028 ( .A(n5531), .B(n5532), .ZN(n7335) );
  INV_X1 U7029 ( .A(n5531), .ZN(n5533) );
  NAND2_X1 U7030 ( .A1(n5536), .A2(n5535), .ZN(n5539) );
  NAND2_X1 U7031 ( .A1(n5537), .A2(SI_18_), .ZN(n5538) );
  INV_X1 U7032 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6632) );
  MUX2_X1 U7033 ( .A(n6632), .B(n10234), .S(n7677), .Z(n5540) );
  INV_X1 U7034 ( .A(SI_19_), .ZN(n10158) );
  INV_X1 U7035 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7036 ( .A1(n5541), .A2(SI_19_), .ZN(n5542) );
  NAND2_X1 U7037 ( .A1(n5560), .A2(n5542), .ZN(n5561) );
  XNOR2_X1 U7038 ( .A(n5562), .B(n5561), .ZN(n7501) );
  NAND2_X1 U7039 ( .A1(n7501), .A2(n7680), .ZN(n5545) );
  AOI22_X1 U7040 ( .A1(n5543), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6010), .B2(
        n9573), .ZN(n5544) );
  XNOR2_X1 U7041 ( .A(n8519), .B(n5735), .ZN(n5554) );
  INV_X1 U7042 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5547) );
  INV_X1 U7043 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5546) );
  OAI21_X1 U7044 ( .B1(n5549), .B2(n5547), .A(n5546), .ZN(n5550) );
  NAND2_X1 U7045 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n5548) );
  NAND2_X1 U7046 ( .A1(n5550), .A2(n5570), .ZN(n8438) );
  OR2_X1 U7047 ( .A1(n8438), .A2(n5706), .ZN(n5553) );
  AOI22_X1 U7048 ( .A1(n7665), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n5787), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7049 ( .A1(n7664), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5551) );
  INV_X1 U7050 ( .A(n8418), .ZN(n8451) );
  NAND2_X1 U7051 ( .A1(n8451), .A2(n7690), .ZN(n5555) );
  NAND2_X1 U7052 ( .A1(n5554), .A2(n5555), .ZN(n5559) );
  INV_X1 U7053 ( .A(n5554), .ZN(n5557) );
  INV_X1 U7054 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U7055 ( .A1(n5557), .A2(n5556), .ZN(n5558) );
  INV_X1 U7056 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6942) );
  INV_X1 U7057 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6732) );
  MUX2_X1 U7058 ( .A(n6942), .B(n6732), .S(n7677), .Z(n5564) );
  INV_X1 U7059 ( .A(SI_20_), .ZN(n5563) );
  NAND2_X1 U7060 ( .A1(n5564), .A2(n5563), .ZN(n5580) );
  INV_X1 U7061 ( .A(n5564), .ZN(n5565) );
  NAND2_X1 U7062 ( .A1(n5565), .A2(SI_20_), .ZN(n5566) );
  XNOR2_X1 U7063 ( .A(n5579), .B(n5578), .ZN(n7517) );
  NAND2_X1 U7064 ( .A1(n7517), .A2(n7680), .ZN(n5568) );
  OR2_X1 U7065 ( .A1(n7681), .A2(n6942), .ZN(n5567) );
  XNOR2_X1 U7066 ( .A(n8513), .B(n5702), .ZN(n5576) );
  INV_X1 U7067 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U7068 ( .A1(n5570), .A2(n10290), .ZN(n5571) );
  NAND2_X1 U7069 ( .A1(n5584), .A2(n5571), .ZN(n8411) );
  OR2_X1 U7070 ( .A1(n8411), .A2(n5706), .ZN(n5574) );
  AOI22_X1 U7071 ( .A1(n5787), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n7664), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7072 ( .A1(n7665), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5572) );
  NOR2_X1 U7073 ( .A1(n8254), .A2(n6170), .ZN(n5575) );
  XNOR2_X1 U7074 ( .A(n5576), .B(n5575), .ZN(n7466) );
  NAND2_X1 U7075 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  INV_X1 U7076 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6852) );
  INV_X1 U7077 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6804) );
  MUX2_X1 U7078 ( .A(n6852), .B(n6804), .S(n7677), .Z(n5596) );
  XNOR2_X1 U7079 ( .A(n5596), .B(SI_21_), .ZN(n5595) );
  NAND2_X1 U7080 ( .A1(n7472), .A2(n7680), .ZN(n5582) );
  OR2_X1 U7081 ( .A1(n7681), .A2(n6852), .ZN(n5581) );
  XNOR2_X1 U7082 ( .A(n8508), .B(n5735), .ZN(n5591) );
  INV_X1 U7083 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U7084 ( .A1(n5584), .A2(n10273), .ZN(n5585) );
  NAND2_X1 U7085 ( .A1(n5607), .A2(n5585), .ZN(n8400) );
  OR2_X1 U7086 ( .A1(n8400), .A2(n5706), .ZN(n5590) );
  INV_X1 U7087 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10202) );
  NAND2_X1 U7088 ( .A1(n7665), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7089 ( .A1(n7664), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5586) );
  OAI211_X1 U7090 ( .C1(n7668), .C2(n10202), .A(n5587), .B(n5586), .ZN(n5588)
         );
  INV_X1 U7091 ( .A(n5588), .ZN(n5589) );
  NOR2_X1 U7092 ( .A1(n8419), .A2(n6170), .ZN(n5592) );
  XNOR2_X1 U7093 ( .A(n5591), .B(n5592), .ZN(n8036) );
  INV_X1 U7094 ( .A(n5591), .ZN(n5593) );
  AND2_X1 U7095 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  INV_X1 U7096 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7097 ( .A1(n5597), .A2(SI_21_), .ZN(n5598) );
  INV_X1 U7098 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7020) );
  MUX2_X1 U7099 ( .A(n10101), .B(n7020), .S(n7677), .Z(n5601) );
  INV_X1 U7100 ( .A(SI_22_), .ZN(n5600) );
  NAND2_X1 U7101 ( .A1(n5601), .A2(n5600), .ZN(n5619) );
  INV_X1 U7102 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7103 ( .A1(n5602), .A2(SI_22_), .ZN(n5603) );
  NAND2_X1 U7104 ( .A1(n5619), .A2(n5603), .ZN(n5620) );
  XNOR2_X1 U7105 ( .A(n5621), .B(n5620), .ZN(n7528) );
  NAND2_X1 U7106 ( .A1(n7528), .A2(n7680), .ZN(n5605) );
  OR2_X1 U7107 ( .A1(n7681), .A2(n10101), .ZN(n5604) );
  XNOR2_X1 U7108 ( .A(n8391), .B(n5702), .ZN(n5616) );
  INV_X1 U7109 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7110 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  NAND2_X1 U7111 ( .A1(n5631), .A2(n5608), .ZN(n8387) );
  OR2_X1 U7112 ( .A1(n8387), .A2(n5706), .ZN(n5614) );
  INV_X1 U7113 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7114 ( .A1(n7664), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7115 ( .A1(n5787), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5609) );
  OAI211_X1 U7116 ( .C1(n5611), .C2(n5189), .A(n5610), .B(n5609), .ZN(n5612)
         );
  INV_X1 U7117 ( .A(n5612), .ZN(n5613) );
  INV_X1 U7118 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7024) );
  INV_X1 U7119 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5622) );
  MUX2_X1 U7120 ( .A(n7024), .B(n5622), .S(n7677), .Z(n5624) );
  INV_X1 U7121 ( .A(SI_23_), .ZN(n5623) );
  NAND2_X1 U7122 ( .A1(n5624), .A2(n5623), .ZN(n5642) );
  INV_X1 U7123 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U7124 ( .A1(n5625), .A2(SI_23_), .ZN(n5626) );
  XNOR2_X1 U7125 ( .A(n5641), .B(n5640), .ZN(n7539) );
  NAND2_X1 U7126 ( .A1(n7539), .A2(n7680), .ZN(n5628) );
  OR2_X1 U7127 ( .A1(n7681), .A2(n7024), .ZN(n5627) );
  XNOR2_X1 U7128 ( .A(n8497), .B(n5702), .ZN(n5638) );
  INV_X1 U7129 ( .A(n5638), .ZN(n5629) );
  INV_X1 U7130 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7131 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  AND2_X1 U7132 ( .A1(n5647), .A2(n5632), .ZN(n8369) );
  NAND2_X1 U7133 ( .A1(n8369), .A2(n5791), .ZN(n5637) );
  INV_X1 U7134 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10260) );
  NAND2_X1 U7135 ( .A1(n7664), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7136 ( .A1(n7665), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5633) );
  OAI211_X1 U7137 ( .C1(n7668), .C2(n10260), .A(n5634), .B(n5633), .ZN(n5635)
         );
  INV_X1 U7138 ( .A(n5635), .ZN(n5636) );
  NOR2_X1 U7139 ( .A1(n8345), .A2(n6170), .ZN(n8027) );
  INV_X1 U7140 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7646) );
  MUX2_X1 U7141 ( .A(n10201), .B(n7646), .S(n7677), .Z(n5656) );
  XNOR2_X1 U7142 ( .A(n5656), .B(SI_24_), .ZN(n5655) );
  XNOR2_X1 U7143 ( .A(n5660), .B(n5655), .ZN(n7552) );
  NAND2_X1 U7144 ( .A1(n7552), .A2(n7680), .ZN(n5644) );
  OR2_X1 U7145 ( .A1(n7681), .A2(n10201), .ZN(n5643) );
  XNOR2_X1 U7146 ( .A(n8491), .B(n5702), .ZN(n5654) );
  INV_X1 U7147 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7148 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  NAND2_X1 U7149 ( .A1(n5682), .A2(n5648), .ZN(n8351) );
  OR2_X1 U7150 ( .A1(n8351), .A2(n5706), .ZN(n5653) );
  INV_X1 U7151 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U7152 ( .A1(n7665), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7153 ( .A1(n7664), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5649) );
  OAI211_X1 U7154 ( .C1(n7668), .C2(n10233), .A(n5650), .B(n5649), .ZN(n5651)
         );
  INV_X1 U7155 ( .A(n5651), .ZN(n5652) );
  NOR2_X1 U7156 ( .A1(n8031), .A2(n6170), .ZN(n8054) );
  INV_X1 U7157 ( .A(n5655), .ZN(n5659) );
  INV_X1 U7158 ( .A(n5656), .ZN(n5657) );
  NAND2_X1 U7159 ( .A1(n5657), .A2(SI_24_), .ZN(n5658) );
  INV_X1 U7160 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7287) );
  INV_X1 U7161 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10281) );
  MUX2_X1 U7162 ( .A(n7287), .B(n10281), .S(n7677), .Z(n5662) );
  INV_X1 U7163 ( .A(SI_25_), .ZN(n5661) );
  NAND2_X1 U7164 ( .A1(n5662), .A2(n5661), .ZN(n5672) );
  INV_X1 U7165 ( .A(n5662), .ZN(n5663) );
  NAND2_X1 U7166 ( .A1(n5663), .A2(SI_25_), .ZN(n5664) );
  NAND2_X1 U7167 ( .A1(n5672), .A2(n5664), .ZN(n5673) );
  NAND2_X1 U7168 ( .A1(n7563), .A2(n7680), .ZN(n5666) );
  OR2_X1 U7169 ( .A1(n7681), .A2(n7287), .ZN(n5665) );
  XNOR2_X1 U7170 ( .A(n8260), .B(n5702), .ZN(n8044) );
  XNOR2_X1 U7171 ( .A(n5682), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U7172 ( .A1(n8328), .A2(n5791), .ZN(n5671) );
  INV_X1 U7173 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U7174 ( .A1(n7665), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7175 ( .A1(n5787), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5667) );
  OAI211_X1 U7176 ( .C1(n5310), .C2(n10169), .A(n5668), .B(n5667), .ZN(n5669)
         );
  INV_X1 U7177 ( .A(n5669), .ZN(n5670) );
  NAND2_X1 U7178 ( .A1(n5671), .A2(n5670), .ZN(n8111) );
  NAND2_X1 U7179 ( .A1(n8111), .A2(n7690), .ZN(n8043) );
  INV_X1 U7180 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7343) );
  INV_X1 U7181 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5675) );
  MUX2_X1 U7182 ( .A(n7343), .B(n5675), .S(n7677), .Z(n5676) );
  INV_X1 U7183 ( .A(SI_26_), .ZN(n10213) );
  NAND2_X1 U7184 ( .A1(n5676), .A2(n10213), .ZN(n5694) );
  INV_X1 U7185 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U7186 ( .A1(n5677), .A2(SI_26_), .ZN(n5678) );
  NAND2_X1 U7187 ( .A1(n7572), .A2(n7680), .ZN(n5680) );
  OR2_X1 U7188 ( .A1(n7681), .A2(n7343), .ZN(n5679) );
  XNOR2_X1 U7189 ( .A(n8482), .B(n5702), .ZN(n8019) );
  INV_X1 U7190 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8047) );
  INV_X1 U7191 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5681) );
  OAI21_X1 U7192 ( .B1(n5682), .B2(n8047), .A(n5681), .ZN(n5683) );
  NAND2_X1 U7193 ( .A1(n5683), .A2(n5704), .ZN(n8322) );
  OR2_X1 U7194 ( .A1(n8322), .A2(n5706), .ZN(n5689) );
  INV_X1 U7195 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7196 ( .A1(n7664), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7197 ( .A1(n5787), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5684) );
  OAI211_X1 U7198 ( .C1(n5686), .C2(n5189), .A(n5685), .B(n5684), .ZN(n5687)
         );
  INV_X1 U7199 ( .A(n5687), .ZN(n5688) );
  NOR2_X1 U7200 ( .A1(n8018), .A2(n6170), .ZN(n5690) );
  NAND2_X1 U7201 ( .A1(n8019), .A2(n5690), .ZN(n5691) );
  OAI21_X1 U7202 ( .B1(n8019), .B2(n5690), .A(n5691), .ZN(n5805) );
  INV_X1 U7203 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7455) );
  INV_X1 U7204 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5696) );
  MUX2_X1 U7205 ( .A(n7455), .B(n5696), .S(n7677), .Z(n5697) );
  INV_X1 U7206 ( .A(SI_27_), .ZN(n10218) );
  NAND2_X1 U7207 ( .A1(n5697), .A2(n10218), .ZN(n5721) );
  INV_X1 U7208 ( .A(n5697), .ZN(n5698) );
  NAND2_X1 U7209 ( .A1(n5698), .A2(SI_27_), .ZN(n5699) );
  NAND2_X1 U7210 ( .A1(n7587), .A2(n7680), .ZN(n5701) );
  OR2_X1 U7211 ( .A1(n7681), .A2(n7455), .ZN(n5700) );
  XNOR2_X1 U7212 ( .A(n8476), .B(n5702), .ZN(n5713) );
  INV_X1 U7213 ( .A(n5704), .ZN(n5703) );
  NAND2_X1 U7214 ( .A1(n5703), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5727) );
  INV_X1 U7215 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U7216 ( .A1(n5704), .A2(n10305), .ZN(n5705) );
  NAND2_X1 U7217 ( .A1(n5727), .A2(n5705), .ZN(n8298) );
  INV_X1 U7218 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U7219 ( .A1(n7665), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U7220 ( .A1(n7664), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5707) );
  OAI211_X1 U7221 ( .C1(n7668), .C2(n5709), .A(n5708), .B(n5707), .ZN(n5710)
         );
  INV_X1 U7222 ( .A(n5710), .ZN(n5711) );
  NOR2_X1 U7223 ( .A1(n8262), .A2(n6170), .ZN(n5714) );
  NAND2_X1 U7224 ( .A1(n5713), .A2(n5714), .ZN(n5718) );
  INV_X1 U7225 ( .A(n5713), .ZN(n5716) );
  INV_X1 U7226 ( .A(n5714), .ZN(n5715) );
  NAND2_X1 U7227 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  INV_X1 U7228 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7645) );
  INV_X1 U7229 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5723) );
  MUX2_X1 U7230 ( .A(n7645), .B(n5723), .S(n7677), .Z(n7639) );
  XNOR2_X1 U7231 ( .A(n7639), .B(SI_28_), .ZN(n7636) );
  NAND2_X1 U7232 ( .A1(n7598), .A2(n7680), .ZN(n5725) );
  OR2_X1 U7233 ( .A1(n7681), .A2(n7645), .ZN(n5724) );
  INV_X1 U7234 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7235 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  NAND2_X1 U7236 ( .A1(n8290), .A2(n5791), .ZN(n5734) );
  INV_X1 U7237 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U7238 ( .A1(n7664), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U7239 ( .A1(n5787), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5729) );
  OAI211_X1 U7240 ( .C1(n5731), .C2(n5189), .A(n5730), .B(n5729), .ZN(n5732)
         );
  INV_X1 U7241 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U7242 ( .A1(n8304), .A2(n7690), .ZN(n5736) );
  XNOR2_X1 U7243 ( .A(n5736), .B(n5735), .ZN(n5777) );
  INV_X1 U7244 ( .A(n5777), .ZN(n5778) );
  NAND3_X1 U7245 ( .A1(n5747), .A2(n5771), .A3(n5751), .ZN(n5737) );
  NAND2_X1 U7246 ( .A1(n5740), .A2(n5739), .ZN(n5745) );
  NAND2_X1 U7247 ( .A1(n5745), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5741) );
  MUX2_X1 U7248 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5741), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5742) );
  NAND2_X1 U7249 ( .A1(n5743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5744) );
  MUX2_X1 U7250 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5744), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5746) );
  NAND2_X1 U7251 ( .A1(n5746), .A2(n5745), .ZN(n7285) );
  NAND2_X1 U7252 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  NAND2_X1 U7253 ( .A1(n5749), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7254 ( .A1(n5772), .A2(n5771), .ZN(n5750) );
  NAND2_X1 U7255 ( .A1(n5750), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5752) );
  XNOR2_X1 U7256 ( .A(n7092), .B(P2_B_REG_SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7257 ( .A1(n7285), .A2(n5753), .ZN(n5754) );
  INV_X1 U7258 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10293) );
  INV_X1 U7259 ( .A(n7285), .ZN(n5767) );
  NOR2_X1 U7260 ( .A1(n5767), .A2(n5768), .ZN(n9891) );
  NOR4_X1 U7261 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5758) );
  NOR4_X1 U7262 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5757) );
  NOR4_X1 U7263 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5756) );
  NOR4_X1 U7264 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5755) );
  NAND4_X1 U7265 ( .A1(n5758), .A2(n5757), .A3(n5756), .A4(n5755), .ZN(n5764)
         );
  NOR2_X1 U7266 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .ZN(
        n5762) );
  NOR4_X1 U7267 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5761) );
  NOR4_X1 U7268 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5760) );
  NOR4_X1 U7269 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5759) );
  NAND4_X1 U7270 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n5763)
         );
  OAI21_X1 U7271 ( .B1(n5764), .B2(n5763), .A(n9885), .ZN(n5876) );
  INV_X1 U7272 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9888) );
  AND2_X1 U7273 ( .A1(n9885), .A2(n9888), .ZN(n5765) );
  INV_X1 U7274 ( .A(n5768), .ZN(n7345) );
  AND2_X1 U7275 ( .A1(n7345), .A2(n7092), .ZN(n9889) );
  AND2_X1 U7276 ( .A1(n5876), .A2(n6369), .ZN(n5766) );
  NAND2_X1 U7277 ( .A1(n8386), .A2(n5766), .ZN(n5796) );
  AND2_X1 U7278 ( .A1(n5768), .A2(n5767), .ZN(n5770) );
  INV_X1 U7279 ( .A(n7092), .ZN(n5769) );
  XNOR2_X1 U7280 ( .A(n5772), .B(n5771), .ZN(n6009) );
  INV_X1 U7281 ( .A(n9892), .ZN(n5773) );
  NOR2_X1 U7282 ( .A1(n9895), .A2(n7840), .ZN(n9571) );
  NAND2_X1 U7283 ( .A1(n5793), .A2(n9571), .ZN(n5775) );
  AND2_X1 U7284 ( .A1(n5774), .A2(n9573), .ZN(n7714) );
  NAND2_X1 U7285 ( .A1(n7714), .A2(n7840), .ZN(n9618) );
  NOR3_X1 U7286 ( .A1(n8293), .A2(n5778), .A3(n8098), .ZN(n5776) );
  AOI21_X1 U7287 ( .B1(n8293), .B2(n5778), .A(n5776), .ZN(n5785) );
  NOR3_X1 U7288 ( .A1(n8293), .A2(n5777), .A3(n8098), .ZN(n5780) );
  NOR2_X1 U7289 ( .A1(n8471), .A2(n5778), .ZN(n5779) );
  NAND2_X1 U7290 ( .A1(n5786), .A2(n5781), .ZN(n5784) );
  NAND2_X1 U7291 ( .A1(n7879), .A2(n7871), .ZN(n6007) );
  AND2_X1 U7292 ( .A1(n9971), .A2(n6007), .ZN(n5782) );
  OAI21_X1 U7293 ( .B1(n8293), .B2(n8063), .A(n8082), .ZN(n5783) );
  OAI211_X1 U7294 ( .C1(n5786), .C2(n5785), .A(n5784), .B(n5783), .ZN(n5803)
         );
  INV_X1 U7295 ( .A(n8268), .ZN(n5792) );
  INV_X1 U7296 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8269) );
  NAND2_X1 U7297 ( .A1(n7664), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7298 ( .A1(n5787), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5788) );
  OAI211_X1 U7299 ( .C1(n8269), .C2(n5189), .A(n5789), .B(n5788), .ZN(n5790)
         );
  AOI21_X1 U7300 ( .B1(n5792), .B2(n5791), .A(n5790), .ZN(n7661) );
  INV_X1 U7301 ( .A(n7661), .ZN(n8287) );
  INV_X1 U7302 ( .A(n5794), .ZN(n6116) );
  INV_X1 U7303 ( .A(n8262), .ZN(n8286) );
  OR2_X1 U7304 ( .A1(n6007), .A2(n5794), .ZN(n9579) );
  AOI22_X1 U7305 ( .A1(n8287), .A2(n8084), .B1(n8286), .B2(n8106), .ZN(n5801)
         );
  INV_X1 U7306 ( .A(n6354), .ZN(n5795) );
  NAND2_X1 U7307 ( .A1(n5796), .A2(n5795), .ZN(n5799) );
  OR2_X1 U7308 ( .A1(n4890), .A2(n6007), .ZN(n5873) );
  NAND2_X1 U7309 ( .A1(n5873), .A2(n6009), .ZN(n5797) );
  NOR2_X1 U7310 ( .A1(n6074), .A2(n5797), .ZN(n5798) );
  NAND2_X1 U7311 ( .A1(n5799), .A2(n5798), .ZN(n8088) );
  AOI22_X1 U7312 ( .A1(n8290), .A2(n8051), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5800) );
  NAND2_X1 U7313 ( .A1(n5803), .A2(n5802), .ZN(P2_U3222) );
  AOI211_X1 U7314 ( .C1(n5805), .C2(n5804), .A(n8082), .B(n8017), .ZN(n5811)
         );
  NAND2_X1 U7315 ( .A1(n8482), .A2(n8098), .ZN(n5809) );
  INV_X1 U7316 ( .A(n8111), .ZN(n8346) );
  OAI22_X1 U7317 ( .A1(n8262), .A2(n9581), .B1(n8346), .B2(n9579), .ZN(n8317)
         );
  AOI22_X1 U7318 ( .A1(n8317), .A2(n8075), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n5806) );
  OAI21_X1 U7319 ( .B1(n8322), .B2(n8094), .A(n5806), .ZN(n5807) );
  INV_X1 U7320 ( .A(n5807), .ZN(n5808) );
  NAND2_X1 U7321 ( .A1(n6544), .A2(n5816), .ZN(n6188) );
  NAND2_X1 U7322 ( .A1(n6191), .A2(n6193), .ZN(n5826) );
  INV_X1 U7323 ( .A(n5826), .ZN(n5823) );
  INV_X1 U7324 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5820) );
  INV_X1 U7325 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7326 ( .A1(n5820), .A2(n5838), .ZN(n5832) );
  INV_X1 U7327 ( .A(n5832), .ZN(n5822) );
  NOR2_X1 U7328 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5821) );
  AND2_X1 U7329 ( .A1(n5822), .A2(n5821), .ZN(n5827) );
  NAND2_X1 U7330 ( .A1(n5823), .A2(n5827), .ZN(n5824) );
  NAND2_X1 U7331 ( .A1(n5824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5825) );
  XNOR2_X1 U7332 ( .A(n5825), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6019) );
  INV_X1 U7333 ( .A(n5827), .ZN(n5828) );
  NOR2_X1 U7334 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(n5828), .ZN(n5829) );
  NAND2_X1 U7335 ( .A1(n5842), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5831) );
  XNOR2_X1 U7336 ( .A(n5831), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7337 ( .A1(n5832), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5833) );
  INV_X1 U7338 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7339 ( .A1(n6204), .A2(n7006), .ZN(n5975) );
  NAND2_X2 U7340 ( .A1(n6074), .A2(n9892), .ZN(n8123) );
  NAND2_X1 U7341 ( .A1(n5837), .A2(n5838), .ZN(n5839) );
  NAND2_X1 U7342 ( .A1(n5839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7343 ( .A1(n8927), .A2(n7006), .ZN(n5841) );
  NAND2_X1 U7344 ( .A1(n5975), .A2(n5841), .ZN(n6038) );
  NOR2_X1 U7345 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5845) );
  INV_X1 U7346 ( .A(n5845), .ZN(n5847) );
  INV_X1 U7347 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5844) );
  INV_X1 U7348 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5843) );
  BUF_X4 U7349 ( .A(n6249), .Z(n7502) );
  OAI21_X1 U7350 ( .B1(n6038), .B2(n7502), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  INV_X1 U7351 ( .A(n6495), .ZN(n6353) );
  NAND2_X1 U7352 ( .A1(n6533), .A2(n6535), .ZN(n5848) );
  NAND2_X1 U7353 ( .A1(n5849), .A2(n5848), .ZN(n6491) );
  NOR2_X1 U7354 ( .A1(n6158), .A2(n9908), .ZN(n5850) );
  INV_X1 U7355 ( .A(n5850), .ZN(n7711) );
  NAND2_X1 U7356 ( .A1(n6158), .A2(n9908), .ZN(n7701) );
  NAND2_X1 U7357 ( .A1(n6491), .A2(n7839), .ZN(n5852) );
  INV_X1 U7358 ( .A(n9908), .ZN(n8087) );
  OR2_X1 U7359 ( .A1(n6158), .A2(n8087), .ZN(n5851) );
  NAND2_X1 U7360 ( .A1(n5852), .A2(n5851), .ZN(n6519) );
  NAND2_X1 U7361 ( .A1(n5855), .A2(n9914), .ZN(n7719) );
  INV_X1 U7362 ( .A(n7842), .ZN(n5856) );
  OR2_X1 U7363 ( .A1(n5855), .A2(n5853), .ZN(n5857) );
  NAND2_X1 U7364 ( .A1(n8122), .A2(n9919), .ZN(n7720) );
  NAND2_X1 U7365 ( .A1(n7705), .A2(n7720), .ZN(n9876) );
  INV_X1 U7366 ( .A(n9919), .ZN(n9869) );
  OR2_X1 U7367 ( .A1(n9869), .A2(n8122), .ZN(n5858) );
  AND2_X1 U7368 ( .A1(n8064), .A2(n5880), .ZN(n5860) );
  NAND2_X1 U7369 ( .A1(n7706), .A2(n7722), .ZN(n7844) );
  AND2_X1 U7370 ( .A1(n9926), .A2(n8121), .ZN(n5862) );
  OR2_X1 U7371 ( .A1(n9926), .A2(n8121), .ZN(n5861) );
  XNOR2_X1 U7372 ( .A(n9933), .B(n8095), .ZN(n7731) );
  INV_X1 U7373 ( .A(n8095), .ZN(n8120) );
  NOR2_X1 U7374 ( .A1(n9933), .A2(n8120), .ZN(n7733) );
  OR2_X1 U7375 ( .A1(n6681), .A2(n6620), .ZN(n7737) );
  NAND2_X1 U7376 ( .A1(n6681), .A2(n6620), .ZN(n7736) );
  OR2_X1 U7377 ( .A1(n5863), .A2(n7846), .ZN(n5864) );
  NAND2_X1 U7378 ( .A1(n6682), .A2(n5864), .ZN(n9940) );
  NAND2_X1 U7379 ( .A1(n5878), .A2(n5774), .ZN(n5865) );
  NAND3_X1 U7380 ( .A1(n5865), .A2(n7687), .A3(n6007), .ZN(n9565) );
  AND2_X1 U7381 ( .A1(n6495), .A2(n6535), .ZN(n7698) );
  OAI21_X2 U7382 ( .B1(n6538), .B2(n7698), .A(n7710), .ZN(n6492) );
  INV_X1 U7383 ( .A(n5866), .ZN(n6525) );
  XNOR2_X1 U7384 ( .A(n9926), .B(n8121), .ZN(n6433) );
  INV_X1 U7385 ( .A(n8121), .ZN(n7717) );
  NAND2_X1 U7386 ( .A1(n9926), .A2(n7717), .ZN(n7729) );
  NAND2_X1 U7387 ( .A1(n5867), .A2(n7846), .ZN(n5868) );
  NAND2_X1 U7388 ( .A1(n6687), .A2(n5868), .ZN(n5869) );
  INV_X1 U7389 ( .A(n7840), .ZN(n7870) );
  NAND2_X1 U7390 ( .A1(n7870), .A2(n7871), .ZN(n7689) );
  NAND2_X1 U7391 ( .A1(n5869), .A2(n9868), .ZN(n5872) );
  OAI22_X1 U7392 ( .A1(n8095), .A2(n9579), .B1(n6680), .B2(n9581), .ZN(n5870)
         );
  INV_X1 U7393 ( .A(n5870), .ZN(n5871) );
  OAI211_X1 U7394 ( .C1(n9940), .C2(n9565), .A(n5872), .B(n5871), .ZN(n9943)
         );
  INV_X1 U7395 ( .A(n5873), .ZN(n5874) );
  NOR2_X1 U7396 ( .A1(n9886), .A2(n5874), .ZN(n5875) );
  NAND2_X1 U7397 ( .A1(n5876), .A2(n5875), .ZN(n6355) );
  INV_X1 U7398 ( .A(n6355), .ZN(n8385) );
  NAND2_X1 U7399 ( .A1(n8385), .A2(n8386), .ZN(n5884) );
  OR2_X1 U7400 ( .A1(n5884), .A2(n6369), .ZN(n5877) );
  MUX2_X1 U7401 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9943), .S(n9591), .Z(n5888)
         );
  OR2_X1 U7402 ( .A1(n5878), .A2(n7687), .ZN(n6418) );
  INV_X1 U7403 ( .A(n6418), .ZN(n5879) );
  NAND2_X1 U7404 ( .A1(n9591), .A2(n5879), .ZN(n9584) );
  NOR2_X1 U7405 ( .A1(n9940), .A2(n9584), .ZN(n5887) );
  NAND2_X1 U7406 ( .A1(n9899), .A2(n9908), .ZN(n6520) );
  OR2_X1 U7407 ( .A1(n6520), .A2(n5853), .ZN(n9870) );
  INV_X1 U7408 ( .A(n6681), .ZN(n9941) );
  AND2_X1 U7409 ( .A1(n5881), .A2(n9941), .ZN(n6693) );
  NOR2_X1 U7410 ( .A1(n5881), .A2(n9941), .ZN(n5882) );
  OR2_X1 U7411 ( .A1(n6693), .A2(n5882), .ZN(n9942) );
  NOR2_X1 U7412 ( .A1(n6369), .A2(n9573), .ZN(n8384) );
  NAND2_X1 U7413 ( .A1(n8384), .A2(n9963), .ZN(n5883) );
  NOR2_X1 U7414 ( .A1(n9942), .A2(n9873), .ZN(n5886) );
  OAI22_X1 U7415 ( .A1(n9881), .A2(n9941), .B1(n9871), .B2(n6590), .ZN(n5885)
         );
  OR4_X1 U7416 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(P2_U3288)
         );
  INV_X1 U7417 ( .A(n5889), .ZN(n6593) );
  AOI211_X1 U7418 ( .C1(n5891), .C2(n5890), .A(n8082), .B(n6593), .ZN(n5895)
         );
  NOR2_X1 U7419 ( .A1(n8058), .A2(n7717), .ZN(n5894) );
  OAI22_X1 U7420 ( .A1(n8096), .A2(n6620), .B1(n4592), .B2(n8063), .ZN(n5893)
         );
  OAI22_X1 U7421 ( .A1(n8094), .A2(n6426), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5255), .ZN(n5892) );
  OR4_X1 U7422 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .ZN(P2_U3215)
         );
  INV_X1 U7423 ( .A(n6701), .ZN(n5896) );
  AOI211_X1 U7424 ( .C1(n5898), .C2(n5897), .A(n8082), .B(n5896), .ZN(n5902)
         );
  INV_X1 U7425 ( .A(n6825), .ZN(n9954) );
  NOR2_X1 U7426 ( .A1(n8063), .A2(n9954), .ZN(n5901) );
  OAI22_X1 U7427 ( .A1(n8094), .A2(n6724), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10102), .ZN(n5900) );
  OAI22_X1 U7428 ( .A1(n6828), .A2(n8096), .B1(n8058), .B2(n6680), .ZN(n5899)
         );
  OR4_X1 U7429 ( .A1(n5902), .A2(n5901), .A3(n5900), .A4(n5899), .ZN(P2_U3219)
         );
  OR2_X1 U7430 ( .A1(n5943), .A2(n9456), .ZN(n5903) );
  XNOR2_X1 U7431 ( .A(n5903), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U7432 ( .A1(n5904), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U7433 ( .A(n5905), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9049) );
  OR2_X1 U7434 ( .A1(n5906), .A2(n9456), .ZN(n5912) );
  NAND2_X1 U7435 ( .A1(n5912), .A2(n5907), .ZN(n5908) );
  NAND2_X1 U7436 ( .A1(n5908), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5909) );
  XNOR2_X1 U7437 ( .A(n5909), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9724) );
  INV_X1 U7438 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5910) );
  MUX2_X1 U7439 ( .A(n5910), .B(P1_REG2_REG_11__SCAN_IN), .S(n9724), .Z(n5911)
         );
  INV_X1 U7440 ( .A(n5911), .ZN(n9729) );
  XNOR2_X1 U7441 ( .A(n5912), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U7442 ( .A1(n5913), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5914) );
  XNOR2_X1 U7443 ( .A(n5914), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U7444 ( .A1(n9707), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5915) );
  OAI21_X1 U7445 ( .B1(n9707), .B2(P1_REG2_REG_9__SCAN_IN), .A(n5915), .ZN(
        n9702) );
  NAND2_X1 U7446 ( .A1(n4542), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5916) );
  XNOR2_X1 U7447 ( .A(n5916), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9682) );
  NOR2_X1 U7448 ( .A1(n9682), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5917) );
  AOI21_X1 U7449 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9682), .A(n5917), .ZN(
        n9694) );
  OR2_X1 U7450 ( .A1(n4551), .A2(n9456), .ZN(n5918) );
  XNOR2_X1 U7451 ( .A(n5918), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9027) );
  NOR2_X1 U7452 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9027), .ZN(n5919) );
  AOI21_X1 U7453 ( .B1(n9027), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5919), .ZN(
        n9035) );
  NAND2_X1 U7454 ( .A1(n5920), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5921) );
  XNOR2_X1 U7455 ( .A(n5921), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U7456 ( .A1(n5922), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5923) );
  XNOR2_X1 U7457 ( .A(n5923), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9663) );
  NOR2_X1 U7458 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9663), .ZN(n5924) );
  AOI21_X1 U7459 ( .B1(n9663), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5924), .ZN(
        n9666) );
  OR2_X1 U7460 ( .A1(n5925), .A2(n9456), .ZN(n5931) );
  OAI21_X1 U7461 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7462 ( .A1(n5931), .A2(n5926), .ZN(n5928) );
  INV_X1 U7463 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5927) );
  XNOR2_X1 U7464 ( .A(n5928), .B(n5927), .ZN(n9646) );
  NAND2_X1 U7465 ( .A1(n5931), .A2(n5929), .ZN(n5933) );
  NAND2_X1 U7466 ( .A1(n5933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U7467 ( .A(n5930), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6455) );
  INV_X1 U7468 ( .A(n5931), .ZN(n5932) );
  NAND2_X1 U7469 ( .A1(n5932), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5934) );
  AND2_X1 U7470 ( .A1(n5934), .A2(n5933), .ZN(n6391) );
  INV_X1 U7471 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6814) );
  MUX2_X1 U7472 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6814), .S(n6391), .Z(n6390)
         );
  INV_X1 U7473 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U7474 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6379) );
  INV_X1 U7475 ( .A(n6379), .ZN(n6051) );
  NAND2_X1 U7476 ( .A1(n6251), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7477 ( .A1(n6050), .A2(n5936), .ZN(n6389) );
  NAND2_X1 U7478 ( .A1(n6390), .A2(n6389), .ZN(n6388) );
  XNOR2_X1 U7479 ( .A(n6455), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6068) );
  NOR2_X1 U7480 ( .A1(n9646), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5937) );
  AOI21_X1 U7481 ( .B1(n9646), .B2(P1_REG2_REG_4__SCAN_IN), .A(n5937), .ZN(
        n9644) );
  NAND2_X1 U7482 ( .A1(n9645), .A2(n9644), .ZN(n9643) );
  OAI21_X1 U7483 ( .B1(n9646), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9643), .ZN(
        n9665) );
  NAND2_X1 U7484 ( .A1(n9666), .A2(n9665), .ZN(n9664) );
  OAI21_X1 U7485 ( .B1(n9663), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9664), .ZN(
        n9675) );
  NAND2_X1 U7486 ( .A1(n9679), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5938) );
  OAI21_X1 U7487 ( .B1(n9679), .B2(P1_REG2_REG_6__SCAN_IN), .A(n5938), .ZN(
        n9674) );
  NOR2_X1 U7488 ( .A1(n9675), .A2(n9674), .ZN(n9673) );
  AOI21_X1 U7489 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n9679), .A(n9673), .ZN(
        n9034) );
  NAND2_X1 U7490 ( .A1(n9035), .A2(n9034), .ZN(n9033) );
  OAI21_X1 U7491 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9027), .A(n9033), .ZN(
        n9693) );
  NAND2_X1 U7492 ( .A1(n9694), .A2(n9693), .ZN(n9692) );
  OAI21_X1 U7493 ( .B1(n9682), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9692), .ZN(
        n9703) );
  NAND2_X1 U7494 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n9720), .ZN(n5939) );
  OAI21_X1 U7495 ( .B1(n9720), .B2(P1_REG2_REG_10__SCAN_IN), .A(n5939), .ZN(
        n9715) );
  NAND2_X1 U7496 ( .A1(n9729), .A2(n9730), .ZN(n9728) );
  OAI21_X1 U7497 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9724), .A(n9728), .ZN(
        n9047) );
  NAND2_X1 U7498 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9049), .ZN(n5940) );
  OAI21_X1 U7499 ( .B1(n9049), .B2(P1_REG2_REG_12__SCAN_IN), .A(n5940), .ZN(
        n9046) );
  NOR2_X1 U7500 ( .A1(n9047), .A2(n9046), .ZN(n9045) );
  NAND2_X1 U7501 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9062), .ZN(n5941) );
  OAI21_X1 U7502 ( .B1(n9062), .B2(P1_REG2_REG_13__SCAN_IN), .A(n5941), .ZN(
        n9059) );
  NAND2_X1 U7503 ( .A1(n5943), .A2(n5942), .ZN(n6187) );
  NAND2_X1 U7504 ( .A1(n6187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5947) );
  XNOR2_X1 U7505 ( .A(n5947), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7240) );
  INV_X1 U7506 ( .A(n7240), .ZN(n6061) );
  NOR2_X1 U7507 ( .A1(n5944), .A2(n6061), .ZN(n5945) );
  NOR2_X1 U7508 ( .A1(n7245), .A2(n7010), .ZN(n7009) );
  NOR2_X1 U7509 ( .A1(n5945), .A2(n7009), .ZN(n9067) );
  NAND2_X1 U7510 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  NAND2_X1 U7511 ( .A1(n5948), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7512 ( .A(n5950), .B(n5949), .ZN(n9074) );
  XNOR2_X1 U7513 ( .A(n9067), .B(n9074), .ZN(n5955) );
  INV_X1 U7514 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5954) );
  NOR2_X1 U7515 ( .A1(n5954), .A2(n5955), .ZN(n9068) );
  NOR2_X1 U7516 ( .A1(n6038), .A2(P1_U3084), .ZN(n5972) );
  XNOR2_X1 U7517 ( .A(n5951), .B(P1_IR_REG_27__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U7518 ( .A1(n5972), .A2(n9113), .ZN(n9108) );
  INV_X1 U7519 ( .A(n9108), .ZN(n5977) );
  NAND2_X1 U7520 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5952) );
  NAND2_X1 U7521 ( .A1(n5951), .A2(n5952), .ZN(n5953) );
  XNOR2_X1 U7522 ( .A(n5953), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6374) );
  AOI211_X1 U7523 ( .C1(n5955), .C2(n5954), .A(n9068), .B(n9713), .ZN(n5982)
         );
  INV_X1 U7524 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7250) );
  NOR2_X1 U7525 ( .A1(n7250), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8712) );
  INV_X1 U7526 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5956) );
  XNOR2_X1 U7527 ( .A(n7240), .B(n5956), .ZN(n7014) );
  OR2_X1 U7528 ( .A1(n9062), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5971) );
  INV_X1 U7529 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5957) );
  MUX2_X1 U7530 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n5957), .S(n9062), .Z(n9055)
         );
  INV_X1 U7531 ( .A(n9720), .ZN(n6030) );
  INV_X1 U7532 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9531) );
  AOI22_X1 U7533 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n9720), .B1(n6030), .B2(
        n9531), .ZN(n9712) );
  OR2_X1 U7534 ( .A1(n9682), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7535 ( .A1(n9682), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7536 ( .A1(n5959), .A2(n5958), .ZN(n9684) );
  NOR2_X1 U7537 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9027), .ZN(n5967) );
  AOI21_X1 U7538 ( .B1(n9027), .B2(P1_REG1_REG_7__SCAN_IN), .A(n5967), .ZN(
        n9030) );
  NAND2_X1 U7539 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9663), .ZN(n5960) );
  OAI21_X1 U7540 ( .B1(n9663), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5960), .ZN(
        n9659) );
  INV_X1 U7541 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9839) );
  MUX2_X1 U7542 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9839), .S(n6391), .Z(n6385)
         );
  INV_X1 U7543 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9837) );
  MUX2_X1 U7544 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9837), .S(n6251), .Z(n6047)
         );
  AND2_X1 U7545 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6046) );
  NAND2_X1 U7546 ( .A1(n6047), .A2(n6046), .ZN(n6045) );
  NAND2_X1 U7547 ( .A1(n6251), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7548 ( .A1(n6045), .A2(n5961), .ZN(n6384) );
  NAND2_X1 U7549 ( .A1(n6385), .A2(n6384), .ZN(n6383) );
  NAND2_X1 U7550 ( .A1(n6391), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7551 ( .A1(n6383), .A2(n5962), .ZN(n6063) );
  INV_X1 U7552 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7553 ( .A(n6455), .B(n5963), .ZN(n6064) );
  NAND2_X1 U7554 ( .A1(n6063), .A2(n6064), .ZN(n6062) );
  NAND2_X1 U7555 ( .A1(n6455), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5964) );
  AND2_X1 U7556 ( .A1(n6062), .A2(n5964), .ZN(n9649) );
  NOR2_X1 U7557 ( .A1(n9646), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5965) );
  AOI21_X1 U7558 ( .B1(n9646), .B2(P1_REG1_REG_4__SCAN_IN), .A(n5965), .ZN(
        n9650) );
  NAND2_X1 U7559 ( .A1(n9649), .A2(n9650), .ZN(n9648) );
  OAI21_X1 U7560 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9646), .A(n9648), .ZN(
        n9660) );
  NOR2_X1 U7561 ( .A1(n9659), .A2(n9660), .ZN(n9658) );
  AOI21_X1 U7562 ( .B1(n9663), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9658), .ZN(
        n9672) );
  NOR2_X1 U7563 ( .A1(n9679), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5966) );
  AOI21_X1 U7564 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9679), .A(n5966), .ZN(
        n9671) );
  NAND2_X1 U7565 ( .A1(n9672), .A2(n9671), .ZN(n9670) );
  OAI21_X1 U7566 ( .B1(n9679), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9670), .ZN(
        n9029) );
  NAND2_X1 U7567 ( .A1(n9030), .A2(n9029), .ZN(n9028) );
  INV_X1 U7568 ( .A(n5967), .ZN(n5968) );
  NAND2_X1 U7569 ( .A1(n9028), .A2(n5968), .ZN(n9685) );
  NOR2_X1 U7570 ( .A1(n9684), .A2(n9685), .ZN(n9686) );
  AOI21_X1 U7571 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9682), .A(n9686), .ZN(
        n9700) );
  NOR2_X1 U7572 ( .A1(n9707), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5969) );
  AOI21_X1 U7573 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9707), .A(n5969), .ZN(
        n9699) );
  NAND2_X1 U7574 ( .A1(n9700), .A2(n9699), .ZN(n9698) );
  OAI21_X1 U7575 ( .B1(n9707), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9698), .ZN(
        n9711) );
  NAND2_X1 U7576 ( .A1(n9712), .A2(n9711), .ZN(n9710) );
  OAI21_X1 U7577 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9720), .A(n9710), .ZN(
        n9727) );
  INV_X1 U7578 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5970) );
  MUX2_X1 U7579 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n5970), .S(n9724), .Z(n9726)
         );
  NAND2_X1 U7580 ( .A1(n9727), .A2(n9726), .ZN(n9725) );
  OAI21_X1 U7581 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9724), .A(n9725), .ZN(
        n9041) );
  INV_X1 U7582 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7070) );
  MUX2_X1 U7583 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7070), .S(n9049), .Z(n9042)
         );
  NAND2_X1 U7584 ( .A1(n9041), .A2(n9042), .ZN(n9040) );
  OAI21_X1 U7585 ( .B1(n9049), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9040), .ZN(
        n9056) );
  NAND2_X1 U7586 ( .A1(n9055), .A2(n9056), .ZN(n9054) );
  NAND2_X1 U7587 ( .A1(n5971), .A2(n9054), .ZN(n7013) );
  NAND2_X1 U7588 ( .A1(n7014), .A2(n7013), .ZN(n7012) );
  OAI21_X1 U7589 ( .B1(n7240), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7012), .ZN(
        n9073) );
  XNOR2_X1 U7590 ( .A(n9074), .B(n9073), .ZN(n5974) );
  INV_X1 U7591 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5973) );
  NOR2_X1 U7592 ( .A1(n5973), .A2(n5974), .ZN(n9075) );
  OR2_X1 U7593 ( .A1(n6374), .A2(n9113), .ZN(n6037) );
  INV_X1 U7594 ( .A(n6037), .ZN(n6381) );
  INV_X1 U7595 ( .A(n9750), .ZN(n9657) );
  AOI211_X1 U7596 ( .C1(n5974), .C2(n5973), .A(n9075), .B(n9657), .ZN(n5981)
         );
  INV_X1 U7597 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n5979) );
  INV_X1 U7598 ( .A(n5975), .ZN(n5976) );
  INV_X1 U7599 ( .A(n9074), .ZN(n7398) );
  NAND2_X1 U7600 ( .A1(n9742), .A2(n7398), .ZN(n5978) );
  OAI21_X1 U7601 ( .B1(n5979), .B2(n9735), .A(n5978), .ZN(n5980) );
  OR4_X1 U7602 ( .A1(n5982), .A2(n8712), .A3(n5981), .A4(n5980), .ZN(P1_U3256)
         );
  NOR2_X2 U7603 ( .A1(n7677), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9465) );
  AOI22_X1 U7604 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n9465), .B1(n6391), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n5983) );
  OAI21_X1 U7605 ( .B1(n6321), .B2(n9463), .A(n5983), .ZN(P1_U3351) );
  AOI22_X1 U7606 ( .A1(n6455), .A2(P1_STATE_REG_SCAN_IN), .B1(n9465), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n5984) );
  OAI21_X1 U7607 ( .B1(n6458), .B2(n9463), .A(n5984), .ZN(P1_U3350) );
  AOI22_X1 U7608 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9646), .B1(n9465), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n5985) );
  OAI21_X1 U7609 ( .B1(n6452), .B2(n9463), .A(n5985), .ZN(P1_U3349) );
  AND2_X1 U7610 ( .A1(n7677), .A2(P2_U3152), .ZN(n8544) );
  INV_X2 U7611 ( .A(n8544), .ZN(n8546) );
  AND2_X1 U7612 ( .A1(n5986), .A2(P2_U3152), .ZN(n7022) );
  INV_X2 U7613 ( .A(n7022), .ZN(n8548) );
  OAI222_X1 U7614 ( .A1(n8546), .A2(n5987), .B1(n8548), .B2(n6254), .C1(
        P2_U3152), .C2(n6106), .ZN(P2_U3357) );
  OAI222_X1 U7615 ( .A1(n8546), .A2(n5989), .B1(n8548), .B2(n6458), .C1(
        P2_U3152), .C2(n5988), .ZN(P2_U3355) );
  INV_X1 U7616 ( .A(n8143), .ZN(n6108) );
  OAI222_X1 U7617 ( .A1(n8546), .A2(n10179), .B1(n8548), .B2(n6452), .C1(
        P2_U3152), .C2(n6108), .ZN(P2_U3354) );
  OAI222_X1 U7618 ( .A1(n8546), .A2(n5990), .B1(n8548), .B2(n6321), .C1(
        P2_U3152), .C2(n9492), .ZN(P2_U3356) );
  INV_X1 U7619 ( .A(n9465), .ZN(n7885) );
  INV_X1 U7620 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6250) );
  INV_X1 U7621 ( .A(n6251), .ZN(n6055) );
  OAI222_X1 U7622 ( .A1(n7885), .A2(n6250), .B1(n9463), .B2(n6254), .C1(n6055), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  AOI22_X1 U7623 ( .A1(n8155), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8544), .ZN(n5991) );
  OAI21_X1 U7624 ( .B1(n6642), .B2(n8548), .A(n5991), .ZN(P2_U3353) );
  AOI22_X1 U7625 ( .A1(n9663), .A2(P1_STATE_REG_SCAN_IN), .B1(n9465), .B2(
        P2_DATAO_REG_5__SCAN_IN), .ZN(n5992) );
  OAI21_X1 U7626 ( .B1(n6642), .B2(n9463), .A(n5992), .ZN(P1_U3348) );
  AOI22_X1 U7627 ( .A1(n9679), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9465), .ZN(n5993) );
  OAI21_X1 U7628 ( .B1(n6656), .B2(n9463), .A(n5993), .ZN(P1_U3347) );
  INV_X1 U7629 ( .A(n8167), .ZN(n6111) );
  OAI222_X1 U7630 ( .A1(n8546), .A2(n5994), .B1(n8548), .B2(n6656), .C1(
        P2_U3152), .C2(n6111), .ZN(P2_U3352) );
  AOI22_X1 U7631 ( .A1(n8179), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8544), .ZN(n5995) );
  OAI21_X1 U7632 ( .B1(n6739), .B2(n8548), .A(n5995), .ZN(P2_U3351) );
  INV_X1 U7633 ( .A(n9027), .ZN(n5997) );
  OAI222_X1 U7634 ( .A1(n5997), .A2(P1_U3084), .B1(n9463), .B2(n6739), .C1(
        n5996), .C2(n7885), .ZN(P1_U3346) );
  INV_X1 U7635 ( .A(n6750), .ZN(n6000) );
  INV_X1 U7636 ( .A(n8192), .ZN(n6113) );
  OAI222_X1 U7637 ( .A1(n8546), .A2(n5998), .B1(n8548), .B2(n6000), .C1(
        P2_U3152), .C2(n6113), .ZN(P2_U3350) );
  INV_X1 U7638 ( .A(n9682), .ZN(n6753) );
  OAI222_X1 U7639 ( .A1(n6753), .A2(P1_U3084), .B1(n9463), .B2(n6000), .C1(
        n5999), .C2(n7885), .ZN(P1_U3345) );
  INV_X1 U7640 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6005) );
  INV_X1 U7641 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7642 ( .A1(n7664), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7643 ( .A1(n7665), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6001) );
  OAI211_X1 U7644 ( .C1(n7668), .C2(n6003), .A(n6002), .B(n6001), .ZN(n8237)
         );
  NAND2_X1 U7645 ( .A1(n8237), .A2(P2_U3966), .ZN(n6004) );
  OAI21_X1 U7646 ( .B1(n6005), .B2(P2_U3966), .A(n6004), .ZN(P2_U3583) );
  INV_X1 U7647 ( .A(n6980), .ZN(n6014) );
  AOI22_X1 U7648 ( .A1(n9707), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9465), .ZN(n6006) );
  OAI21_X1 U7649 ( .B1(n6014), .B2(n9463), .A(n6006), .ZN(P1_U3344) );
  INV_X1 U7650 ( .A(n6007), .ZN(n6076) );
  NAND2_X1 U7651 ( .A1(n6008), .A2(n6076), .ZN(n6013) );
  OR2_X1 U7652 ( .A1(n6009), .A2(P2_U3152), .ZN(n7882) );
  NAND2_X1 U7653 ( .A1(n9886), .A2(n7882), .ZN(n6011) );
  NAND2_X1 U7654 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  AND2_X1 U7655 ( .A1(n6013), .A2(n6012), .ZN(n9488) );
  NOR2_X1 U7656 ( .A1(n9857), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7657 ( .A(n6128), .ZN(n6121) );
  OAI222_X1 U7658 ( .A1(n8546), .A2(n6015), .B1(n8548), .B2(n6014), .C1(n6121), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7659 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10291) );
  INV_X1 U7660 ( .A(P1_B_REG_SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7661 ( .A1(n4564), .A2(n6018), .ZN(n6022) );
  INV_X1 U7662 ( .A(n6019), .ZN(n7283) );
  NAND3_X1 U7663 ( .A1(n6017), .A2(P1_B_REG_SCAN_IN), .A3(n7283), .ZN(n6021)
         );
  NAND3_X1 U7664 ( .A1(n6022), .A2(n6021), .A3(n6020), .ZN(n9792) );
  OR2_X1 U7665 ( .A1(n9792), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6024) );
  INV_X1 U7666 ( .A(n6020), .ZN(n6208) );
  NAND2_X1 U7667 ( .A1(n6208), .A2(n7283), .ZN(n6023) );
  NAND2_X1 U7668 ( .A1(n6024), .A2(n6023), .ZN(n6233) );
  INV_X1 U7669 ( .A(n6233), .ZN(n6561) );
  NAND2_X1 U7670 ( .A1(n6561), .A2(n9793), .ZN(n6025) );
  OAI21_X1 U7671 ( .B1(n9793), .B2(n10291), .A(n6025), .ZN(P1_U3441) );
  INV_X1 U7672 ( .A(n7053), .ZN(n6032) );
  AOI22_X1 U7673 ( .A1(n9724), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9465), .ZN(n6026) );
  OAI21_X1 U7674 ( .B1(n6032), .B2(n9463), .A(n6026), .ZN(P1_U3342) );
  INV_X1 U7675 ( .A(n7048), .ZN(n6029) );
  INV_X1 U7676 ( .A(n6290), .ZN(n6136) );
  OAI222_X1 U7677 ( .A1(n8546), .A2(n6027), .B1(n8548), .B2(n6029), .C1(n6136), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  OAI222_X1 U7678 ( .A1(P1_U3084), .A2(n6030), .B1(n9463), .B2(n6029), .C1(
        n6028), .C2(n7885), .ZN(P1_U3343) );
  INV_X1 U7679 ( .A(n6306), .ZN(n6300) );
  OAI222_X1 U7680 ( .A1(P2_U3152), .A2(n6300), .B1(n8548), .B2(n6032), .C1(
        n6031), .C2(n8546), .ZN(P2_U3347) );
  INV_X1 U7681 ( .A(n7134), .ZN(n6034) );
  AOI22_X1 U7682 ( .A1(n9049), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9465), .ZN(n6033) );
  OAI21_X1 U7683 ( .B1(n6034), .B2(n9463), .A(n6033), .ZN(P1_U3341) );
  INV_X1 U7684 ( .A(n8207), .ZN(n6308) );
  OAI222_X1 U7685 ( .A1(n8546), .A2(n6035), .B1(n8548), .B2(n6034), .C1(
        P2_U3152), .C2(n6308), .ZN(P2_U3346) );
  INV_X1 U7686 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6044) );
  INV_X1 U7687 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6183) );
  AND2_X1 U7688 ( .A1(n9113), .A2(n6183), .ZN(n6036) );
  OR2_X1 U7689 ( .A1(n6036), .A2(n6374), .ZN(n6377) );
  INV_X1 U7690 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6376) );
  XNOR2_X1 U7691 ( .A(n6377), .B(n6376), .ZN(n6040) );
  OAI211_X1 U7692 ( .C1(n6037), .C2(P1_REG1_REG_0__SCAN_IN), .A(n6754), .B(
        P1_STATE_REG_SCAN_IN), .ZN(n6039) );
  NOR3_X1 U7693 ( .A1(n6040), .A2(n6039), .A3(n6038), .ZN(n6042) );
  INV_X1 U7694 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10135) );
  AND3_X1 U7695 ( .A1(n9750), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10135), .ZN(
        n6041) );
  AOI211_X1 U7696 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6042), .B(
        n6041), .ZN(n6043) );
  OAI21_X1 U7697 ( .B1(n9735), .B2(n6044), .A(n6043), .ZN(P1_U3241) );
  INV_X1 U7698 ( .A(n9742), .ZN(n9082) );
  INV_X1 U7699 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6585) );
  OAI211_X1 U7700 ( .C1(n6047), .C2(n6046), .A(n9750), .B(n6045), .ZN(n6048)
         );
  OAI21_X1 U7701 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6585), .A(n6048), .ZN(n6049) );
  AOI21_X1 U7702 ( .B1(n9749), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n6049), .ZN(
        n6054) );
  OAI211_X1 U7703 ( .C1(n6052), .C2(n6051), .A(n9740), .B(n6050), .ZN(n6053)
         );
  OAI211_X1 U7704 ( .C1(n9082), .C2(n6055), .A(n6054), .B(n6053), .ZN(P1_U3242) );
  INV_X1 U7705 ( .A(n7213), .ZN(n6057) );
  AOI22_X1 U7706 ( .A1(n9062), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9465), .ZN(n6056) );
  OAI21_X1 U7707 ( .B1(n6057), .B2(n9463), .A(n6056), .ZN(P1_U3340) );
  INV_X1 U7708 ( .A(n6407), .ZN(n6317) );
  OAI222_X1 U7709 ( .A1(n8546), .A2(n6058), .B1(n8548), .B2(n6057), .C1(n6317), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7710 ( .A(n7239), .ZN(n6060) );
  INV_X1 U7711 ( .A(n6925), .ZN(n6411) );
  OAI222_X1 U7712 ( .A1(n8546), .A2(n10243), .B1(n8548), .B2(n6060), .C1(n6411), .C2(P2_U3152), .ZN(P2_U3344) );
  OAI222_X1 U7713 ( .A1(P1_U3084), .A2(n6061), .B1(n9463), .B2(n6060), .C1(
        n6059), .C2(n7885), .ZN(P1_U3339) );
  INV_X1 U7714 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10263) );
  OAI211_X1 U7715 ( .C1(n6064), .C2(n6063), .A(n9750), .B(n6062), .ZN(n6066)
         );
  INV_X1 U7716 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10240) );
  NOR2_X1 U7717 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10240), .ZN(n6510) );
  INV_X1 U7718 ( .A(n6510), .ZN(n6065) );
  OAI211_X1 U7719 ( .C1(n10263), .C2(n9735), .A(n6066), .B(n6065), .ZN(n6071)
         );
  AOI211_X1 U7720 ( .C1(n6069), .C2(n6068), .A(n6067), .B(n9713), .ZN(n6070)
         );
  AOI211_X1 U7721 ( .C1(n9742), .C2(n6455), .A(n6071), .B(n6070), .ZN(n6072)
         );
  INV_X1 U7722 ( .A(n6072), .ZN(P1_U3244) );
  INV_X1 U7723 ( .A(n7882), .ZN(n6073) );
  AOI21_X1 U7724 ( .B1(n6074), .B2(P2_STATE_REG_SCAN_IN), .A(n6073), .ZN(n6075) );
  OAI21_X1 U7725 ( .B1(n9886), .B2(n6076), .A(n6075), .ZN(n6078) );
  NAND2_X1 U7726 ( .A1(n6078), .A2(n6077), .ZN(n6095) );
  NAND2_X1 U7727 ( .A1(n6095), .A2(n8123), .ZN(n6115) );
  NAND2_X1 U7728 ( .A1(n6115), .A2(n5794), .ZN(n9852) );
  NAND2_X1 U7729 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6623) );
  INV_X1 U7730 ( .A(n6623), .ZN(n6100) );
  XNOR2_X1 U7731 ( .A(n8143), .B(n6079), .ZN(n8146) );
  NAND2_X1 U7732 ( .A1(n8130), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6085) );
  INV_X1 U7733 ( .A(n9492), .ZN(n6082) );
  INV_X1 U7734 ( .A(n6106), .ZN(n9476) );
  NAND2_X1 U7735 ( .A1(n9861), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9474) );
  INV_X1 U7736 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6080) );
  MUX2_X1 U7737 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6080), .S(n6106), .Z(n9473)
         );
  NOR2_X1 U7738 ( .A1(n9474), .A2(n9473), .ZN(n9472) );
  AOI21_X1 U7739 ( .B1(n9476), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9472), .ZN(
        n9485) );
  INV_X1 U7740 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6081) );
  MUX2_X1 U7741 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6081), .S(n9492), .Z(n9486)
         );
  NOR2_X1 U7742 ( .A1(n9485), .A2(n9486), .ZN(n9484) );
  AOI21_X1 U7743 ( .B1(n6082), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9484), .ZN(
        n8133) );
  OR2_X1 U7744 ( .A1(n8130), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7745 ( .A1(n6083), .A2(n6085), .ZN(n8132) );
  NOR2_X1 U7746 ( .A1(n8133), .A2(n8132), .ZN(n8131) );
  INV_X1 U7747 ( .A(n8131), .ZN(n6084) );
  NAND2_X1 U7748 ( .A1(n6085), .A2(n6084), .ZN(n8145) );
  NAND2_X1 U7749 ( .A1(n8146), .A2(n8145), .ZN(n8144) );
  NAND2_X1 U7750 ( .A1(n8143), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7751 ( .A1(n8144), .A2(n6086), .ZN(n8157) );
  OR2_X1 U7752 ( .A1(n8155), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7753 ( .A1(n8155), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6088) );
  AND2_X1 U7754 ( .A1(n6087), .A2(n6088), .ZN(n8158) );
  NAND2_X1 U7755 ( .A1(n8157), .A2(n8158), .ZN(n8156) );
  NAND2_X1 U7756 ( .A1(n8156), .A2(n6088), .ZN(n8169) );
  XNOR2_X1 U7757 ( .A(n8167), .B(n6089), .ZN(n8170) );
  NAND2_X1 U7758 ( .A1(n8169), .A2(n8170), .ZN(n8168) );
  NAND2_X1 U7759 ( .A1(n8167), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7760 ( .A1(n8168), .A2(n6090), .ZN(n8181) );
  OR2_X1 U7761 ( .A1(n8179), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7762 ( .A1(n8179), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6092) );
  AND2_X1 U7763 ( .A1(n6091), .A2(n6092), .ZN(n8182) );
  NAND2_X1 U7764 ( .A1(n8181), .A2(n8182), .ZN(n8180) );
  NAND2_X1 U7765 ( .A1(n8180), .A2(n6092), .ZN(n8195) );
  XNOR2_X1 U7766 ( .A(n8192), .B(n6093), .ZN(n8196) );
  AND2_X1 U7767 ( .A1(n8195), .A2(n8196), .ZN(n8193) );
  AOI21_X1 U7768 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n8192), .A(n8193), .ZN(
        n6098) );
  INV_X1 U7769 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6094) );
  MUX2_X1 U7770 ( .A(n6094), .B(P2_REG1_REG_9__SCAN_IN), .S(n6128), .Z(n6097)
         );
  NOR2_X1 U7771 ( .A1(n6098), .A2(n6097), .ZN(n6122) );
  INV_X1 U7772 ( .A(n6095), .ZN(n6096) );
  NAND2_X1 U7773 ( .A1(n6096), .A2(n7878), .ZN(n9854) );
  AOI211_X1 U7774 ( .C1(n6098), .C2(n6097), .A(n6122), .B(n9854), .ZN(n6099)
         );
  AOI211_X1 U7775 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9857), .A(n6100), .B(
        n6099), .ZN(n6120) );
  MUX2_X1 U7776 ( .A(n6692), .B(P2_REG2_REG_9__SCAN_IN), .S(n6128), .Z(n6101)
         );
  INV_X1 U7777 ( .A(n6101), .ZN(n6118) );
  NAND2_X1 U7778 ( .A1(n8179), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6112) );
  MUX2_X1 U7779 ( .A(n6425), .B(P2_REG2_REG_7__SCAN_IN), .S(n8179), .Z(n6102)
         );
  INV_X1 U7780 ( .A(n6102), .ZN(n8176) );
  NAND2_X1 U7781 ( .A1(n8155), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6110) );
  MUX2_X1 U7782 ( .A(n6552), .B(P2_REG2_REG_5__SCAN_IN), .S(n8155), .Z(n6103)
         );
  INV_X1 U7783 ( .A(n6103), .ZN(n8152) );
  NAND2_X1 U7784 ( .A1(n8130), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6107) );
  MUX2_X1 U7785 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6104), .S(n8130), .Z(n8126)
         );
  MUX2_X1 U7786 ( .A(n6105), .B(P2_REG2_REG_2__SCAN_IN), .S(n9492), .Z(n9495)
         );
  MUX2_X1 U7787 ( .A(n6540), .B(P2_REG2_REG_1__SCAN_IN), .S(n6106), .Z(n9479)
         );
  NAND3_X1 U7788 ( .A1(n9861), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n9479), .ZN(
        n9478) );
  OAI21_X1 U7789 ( .B1(n6106), .B2(n6540), .A(n9478), .ZN(n9496) );
  NAND2_X1 U7790 ( .A1(n9495), .A2(n9496), .ZN(n9494) );
  OAI21_X1 U7791 ( .B1(n9492), .B2(n6105), .A(n9494), .ZN(n8127) );
  NAND2_X1 U7792 ( .A1(n8126), .A2(n8127), .ZN(n8125) );
  NAND2_X1 U7793 ( .A1(n6107), .A2(n8125), .ZN(n8141) );
  MUX2_X1 U7794 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6109), .S(n8143), .Z(n8140)
         );
  NAND2_X1 U7795 ( .A1(n8141), .A2(n8140), .ZN(n8139) );
  OAI21_X1 U7796 ( .B1(n6109), .B2(n6108), .A(n8139), .ZN(n8153) );
  NAND2_X1 U7797 ( .A1(n8152), .A2(n8153), .ZN(n8151) );
  NAND2_X1 U7798 ( .A1(n6110), .A2(n8151), .ZN(n8165) );
  MUX2_X1 U7799 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6437), .S(n8167), .Z(n8164)
         );
  NAND2_X1 U7800 ( .A1(n8165), .A2(n8164), .ZN(n8163) );
  OAI21_X1 U7801 ( .B1(n6437), .B2(n6111), .A(n8163), .ZN(n8177) );
  NAND2_X1 U7802 ( .A1(n8176), .A2(n8177), .ZN(n8175) );
  NAND2_X1 U7803 ( .A1(n6112), .A2(n8175), .ZN(n8189) );
  MUX2_X1 U7804 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6114), .S(n8192), .Z(n8188)
         );
  NAND2_X1 U7805 ( .A1(n8189), .A2(n8188), .ZN(n8187) );
  OAI21_X1 U7806 ( .B1(n6114), .B2(n6113), .A(n8187), .ZN(n6117) );
  INV_X1 U7807 ( .A(n7878), .ZN(n8236) );
  AND2_X1 U7808 ( .A1(n6115), .A2(n8236), .ZN(n9851) );
  NAND2_X1 U7809 ( .A1(n6118), .A2(n6117), .ZN(n6129) );
  OAI211_X1 U7810 ( .C1(n6118), .C2(n6117), .A(n9850), .B(n6129), .ZN(n6119)
         );
  OAI211_X1 U7811 ( .C1(n9852), .C2(n6121), .A(n6120), .B(n6119), .ZN(P2_U3254) );
  NOR2_X1 U7812 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10102), .ZN(n6127) );
  AOI21_X1 U7813 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n6128), .A(n6122), .ZN(
        n6125) );
  MUX2_X1 U7814 ( .A(n6123), .B(P2_REG1_REG_10__SCAN_IN), .S(n6290), .Z(n6124)
         );
  NOR2_X1 U7815 ( .A1(n6125), .A2(n6124), .ZN(n6289) );
  AOI211_X1 U7816 ( .C1(n6125), .C2(n6124), .A(n6289), .B(n9854), .ZN(n6126)
         );
  AOI211_X1 U7817 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9857), .A(n6127), .B(
        n6126), .ZN(n6135) );
  NAND2_X1 U7818 ( .A1(n6128), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7819 ( .A1(n6130), .A2(n6129), .ZN(n6133) );
  MUX2_X1 U7820 ( .A(n6725), .B(P2_REG2_REG_10__SCAN_IN), .S(n6290), .Z(n6131)
         );
  INV_X1 U7821 ( .A(n6131), .ZN(n6132) );
  NAND2_X1 U7822 ( .A1(n6132), .A2(n6133), .ZN(n6283) );
  OAI211_X1 U7823 ( .C1(n6133), .C2(n6132), .A(n9850), .B(n6283), .ZN(n6134)
         );
  OAI211_X1 U7824 ( .C1(n9852), .C2(n6136), .A(n6135), .B(n6134), .ZN(P2_U3255) );
  INV_X1 U7825 ( .A(n8075), .ZN(n8048) );
  AOI22_X1 U7826 ( .A1(n9864), .A2(n8122), .B1(n8121), .B2(n9865), .ZN(n6364)
         );
  OAI22_X1 U7827 ( .A1(n8048), .A2(n6364), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6137), .ZN(n6138) );
  AOI21_X1 U7828 ( .B1(n6555), .B2(n8098), .A(n6138), .ZN(n6143) );
  AOI21_X1 U7829 ( .B1(n6140), .B2(n6139), .A(n8082), .ZN(n6141) );
  NAND2_X1 U7830 ( .A1(n6141), .A2(n8100), .ZN(n6142) );
  OAI211_X1 U7831 ( .C1(n8094), .C2(n6553), .A(n6143), .B(n6142), .ZN(P2_U3229) );
  CLKBUF_X2 U7832 ( .A(P1_U4006), .Z(n9025) );
  INV_X1 U7833 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6156) );
  INV_X1 U7834 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7835 ( .A1(n6146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6147) );
  MUX2_X1 U7836 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6147), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n6149) );
  INV_X1 U7837 ( .A(n6148), .ZN(n9457) );
  INV_X1 U7838 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6154) );
  AND2_X2 U7839 ( .A1(n6150), .A2(n9466), .ZN(n6444) );
  NAND2_X1 U7840 ( .A1(n8721), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6153) );
  INV_X1 U7841 ( .A(n6274), .ZN(n7069) );
  INV_X1 U7842 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9116) );
  OR2_X1 U7843 ( .A1(n7549), .A2(n9116), .ZN(n6152) );
  OAI211_X1 U7844 ( .C1(n6273), .C2(n6154), .A(n6153), .B(n6152), .ZN(n8917)
         );
  NAND2_X1 U7845 ( .A1(n8917), .A2(n9025), .ZN(n6155) );
  OAI21_X1 U7846 ( .B1(n9025), .B2(n6156), .A(n6155), .ZN(P1_U3586) );
  INV_X1 U7847 ( .A(n6157), .ZN(n6348) );
  INV_X1 U7848 ( .A(n6535), .ZN(n9902) );
  AOI22_X1 U7849 ( .A1(n8084), .A2(n6158), .B1(n9902), .B2(n8098), .ZN(n6166)
         );
  INV_X1 U7850 ( .A(n8082), .ZN(n8101) );
  OAI21_X1 U7851 ( .B1(n6161), .B2(n6160), .A(n6159), .ZN(n6164) );
  INV_X1 U7852 ( .A(n8088), .ZN(n6162) );
  NAND2_X1 U7853 ( .A1(P2_U3152), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9470) );
  OAI21_X1 U7854 ( .B1(n6162), .B2(n6534), .A(n9470), .ZN(n6163) );
  AOI21_X1 U7855 ( .B1(n8101), .B2(n6164), .A(n6163), .ZN(n6165) );
  OAI211_X1 U7856 ( .C1(n8058), .C2(n6348), .A(n6166), .B(n6165), .ZN(P2_U3224) );
  INV_X1 U7857 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U7858 ( .A1(n8098), .A2(n5853), .ZN(n6167) );
  OAI21_X1 U7859 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n8128), .A(n6167), .ZN(n6169) );
  INV_X1 U7860 ( .A(n8122), .ZN(n6526) );
  OAI22_X1 U7861 ( .A1(n8096), .A2(n6526), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8094), .ZN(n6168) );
  AOI211_X1 U7862 ( .C1(n8106), .C2(n6158), .A(n6169), .B(n6168), .ZN(n6178)
         );
  NOR2_X1 U7863 ( .A1(n8082), .A2(n6170), .ZN(n8078) );
  INV_X1 U7864 ( .A(n8078), .ZN(n8105) );
  INV_X1 U7865 ( .A(n6158), .ZN(n6527) );
  NOR3_X1 U7866 ( .A1(n8105), .A2(n6171), .A3(n6527), .ZN(n6176) );
  AOI21_X1 U7867 ( .B1(n6172), .B2(n4874), .A(n8082), .ZN(n6175) );
  OAI21_X1 U7868 ( .B1(n6176), .B2(n6175), .A(n6174), .ZN(n6177) );
  NAND2_X1 U7869 ( .A1(n6178), .A2(n6177), .ZN(P2_U3220) );
  INV_X1 U7870 ( .A(n7397), .ZN(n6180) );
  OAI222_X1 U7871 ( .A1(n7885), .A2(n6179), .B1(n9463), .B2(n6180), .C1(n9074), 
        .C2(P1_U3084), .ZN(P1_U3338) );
  INV_X1 U7872 ( .A(n6967), .ZN(n6959) );
  OAI222_X1 U7873 ( .A1(n8546), .A2(n6181), .B1(n8548), .B2(n6180), .C1(
        P2_U3152), .C2(n6959), .ZN(P2_U3343) );
  INV_X1 U7874 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7875 ( .A1(n6444), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7876 ( .A1(n6188), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7877 ( .A1(n6192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6194) );
  INV_X2 U7878 ( .A(n6261), .ZN(n6322) );
  INV_X1 U7879 ( .A(n6572), .ZN(n6197) );
  NAND2_X4 U7880 ( .A1(n6195), .A2(n6197), .ZN(n8003) );
  INV_X1 U7881 ( .A(n8003), .ZN(n6318) );
  INV_X1 U7882 ( .A(n6198), .ZN(n6199) );
  XNOR2_X1 U7883 ( .A(n6199), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9469) );
  INV_X1 U7884 ( .A(n9469), .ZN(n6201) );
  OAI21_X2 U7885 ( .B1(n7502), .B2(n6201), .A(n6200), .ZN(n6583) );
  NAND2_X1 U7886 ( .A1(n6235), .A2(n6318), .ZN(n6206) );
  AOI22_X1 U7887 ( .A1(n6583), .A2(n6322), .B1(n6204), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7888 ( .A1(n6206), .A2(n6205), .ZN(n6255) );
  OAI21_X1 U7889 ( .B1(n6207), .B2(n6255), .A(n6259), .ZN(n6373) );
  OR2_X1 U7890 ( .A1(n9792), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7891 ( .A1(n6017), .A2(n6208), .ZN(n6209) );
  NOR2_X1 U7892 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .ZN(
        n6214) );
  NOR4_X1 U7893 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6213) );
  NOR4_X1 U7894 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6212) );
  NOR4_X1 U7895 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6211) );
  NAND4_X1 U7896 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n6220)
         );
  NOR4_X1 U7897 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6218) );
  NOR4_X1 U7898 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6217) );
  NOR4_X1 U7899 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6216) );
  NOR4_X1 U7900 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6215) );
  NAND4_X1 U7901 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n6219)
         );
  NOR2_X1 U7902 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  NAND2_X1 U7903 ( .A1(n6234), .A2(n6561), .ZN(n6473) );
  INV_X1 U7904 ( .A(n9793), .ZN(n9454) );
  OR2_X1 U7905 ( .A1(n6473), .A2(n9454), .ZN(n6223) );
  OR2_X1 U7906 ( .A1(n9524), .A2(n8927), .ZN(n6469) );
  NOR2_X2 U7907 ( .A1(n6223), .A2(n6469), .ZN(n8645) );
  NAND2_X1 U7908 ( .A1(n6566), .A2(n9001), .ZN(n9784) );
  AOI22_X1 U7909 ( .A1(n6373), .A2(n8645), .B1(n6583), .B2(n8692), .ZN(n6231)
         );
  INV_X1 U7910 ( .A(n6473), .ZN(n6228) );
  NAND2_X1 U7911 ( .A1(n6224), .A2(n8927), .ZN(n6470) );
  NOR2_X1 U7912 ( .A1(n9003), .A2(n6572), .ZN(n6225) );
  NAND2_X1 U7913 ( .A1(n4473), .A2(n6225), .ZN(n6574) );
  NAND2_X1 U7914 ( .A1(n6574), .A2(n9784), .ZN(n6226) );
  AND2_X1 U7915 ( .A1(n6226), .A2(n9793), .ZN(n6227) );
  NAND2_X1 U7916 ( .A1(n6473), .A2(n6227), .ZN(n6475) );
  OAI211_X1 U7917 ( .C1(n6228), .C2(n9524), .A(n6560), .B(n6475), .ZN(n6343)
         );
  INV_X1 U7918 ( .A(n6574), .ZN(n6236) );
  NAND2_X1 U7919 ( .A1(n6236), .A2(n9793), .ZN(n9007) );
  OR2_X1 U7920 ( .A1(n6473), .A2(n9007), .ZN(n6270) );
  INV_X2 U7921 ( .A(n8648), .ZN(n8713) );
  OR2_X1 U7922 ( .A1(n6338), .A2(n6585), .ZN(n6247) );
  OR2_X1 U7923 ( .A1(n6274), .A2(n5935), .ZN(n6245) );
  INV_X1 U7924 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7925 ( .A1(n6444), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6246) );
  AOI22_X1 U7926 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n6343), .B1(n8713), .B2(
        n6570), .ZN(n6230) );
  NAND2_X1 U7927 ( .A1(n6231), .A2(n6230), .ZN(P1_U3230) );
  OR2_X1 U7928 ( .A1(n6787), .A2(n8964), .ZN(n6232) );
  INV_X2 U7929 ( .A(n9845), .ZN(n9848) );
  INV_X1 U7930 ( .A(n6583), .ZN(n6584) );
  INV_X1 U7931 ( .A(n6566), .ZN(n6238) );
  NAND2_X1 U7932 ( .A1(n4867), .A2(n6583), .ZN(n6575) );
  NAND2_X1 U7933 ( .A1(n9026), .A2(n6584), .ZN(n8746) );
  NAND2_X1 U7934 ( .A1(n6575), .A2(n8746), .ZN(n8935) );
  NOR2_X1 U7935 ( .A1(n6236), .A2(n6566), .ZN(n6237) );
  AOI22_X1 U7936 ( .A1(n8935), .A2(n6237), .B1(n9504), .B2(n6570), .ZN(n6563)
         );
  OAI21_X1 U7937 ( .B1(n6584), .B2(n6238), .A(n6563), .ZN(n6243) );
  NAND2_X1 U7938 ( .A1(n6243), .A2(n9848), .ZN(n6239) );
  OAI21_X1 U7939 ( .B1(n9848), .B2(n10135), .A(n6239), .ZN(P1_U3523) );
  INV_X1 U7940 ( .A(n6559), .ZN(n6240) );
  NOR2_X1 U7941 ( .A1(n9455), .A2(n6240), .ZN(n6241) );
  NAND2_X1 U7942 ( .A1(n6243), .A2(n4474), .ZN(n6244) );
  OAI21_X1 U7943 ( .B1(n4474), .B2(n6182), .A(n6244), .ZN(P1_U3454) );
  NAND2_X1 U7944 ( .A1(n7502), .A2(n6251), .ZN(n6252) );
  INV_X1 U7945 ( .A(n6279), .ZN(n9797) );
  OAI22_X1 U7946 ( .A1(n6262), .A2(n4868), .B1(n9797), .B2(n8003), .ZN(n6269)
         );
  INV_X1 U7947 ( .A(n6255), .ZN(n6258) );
  NAND2_X1 U7948 ( .A1(n4473), .A2(n8795), .ZN(n6257) );
  NAND2_X4 U7949 ( .A1(n6257), .A2(n6572), .ZN(n8001) );
  NAND2_X1 U7950 ( .A1(n6258), .A2(n8001), .ZN(n6260) );
  NAND2_X1 U7951 ( .A1(n6260), .A2(n6259), .ZN(n6264) );
  OAI22_X1 U7952 ( .A1(n6262), .A2(n8003), .B1(n9797), .B2(n7985), .ZN(n6263)
         );
  XNOR2_X1 U7953 ( .A(n6263), .B(n7996), .ZN(n6265) );
  INV_X1 U7954 ( .A(n6332), .ZN(n6267) );
  AOI21_X1 U7955 ( .B1(n6269), .B2(n6268), .A(n6267), .ZN(n6282) );
  INV_X1 U7956 ( .A(n6270), .ZN(n6271) );
  INV_X1 U7957 ( .A(n8710), .ZN(n7390) );
  INV_X1 U7958 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7959 ( .A1(n6444), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6277) );
  OR2_X1 U7960 ( .A1(n6274), .A2(n6814), .ZN(n6276) );
  INV_X1 U7961 ( .A(n6338), .ZN(n6646) );
  NAND2_X1 U7962 ( .A1(n6646), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6275) );
  NAND4_X2 U7963 ( .A1(n6278), .A2(n6277), .A3(n6276), .A4(n6275), .ZN(n9024)
         );
  AOI22_X1 U7964 ( .A1(n7390), .A2(n9026), .B1(n8713), .B2(n9024), .ZN(n6281)
         );
  AOI22_X1 U7965 ( .A1(n6599), .A2(n8692), .B1(n6343), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6280) );
  OAI211_X1 U7966 ( .C1(n6282), .C2(n8719), .A(n6281), .B(n6280), .ZN(P1_U3220) );
  NAND2_X1 U7967 ( .A1(n6290), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7968 ( .A1(n6284), .A2(n6283), .ZN(n6286) );
  MUX2_X1 U7969 ( .A(n6838), .B(P2_REG2_REG_11__SCAN_IN), .S(n6306), .Z(n6285)
         );
  NOR2_X1 U7970 ( .A1(n6286), .A2(n6285), .ZN(n6299) );
  AOI21_X1 U7971 ( .B1(n6286), .B2(n6285), .A(n6299), .ZN(n6298) );
  AND2_X1 U7972 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6287) );
  AOI21_X1 U7973 ( .B1(n9857), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6287), .ZN(
        n6295) );
  MUX2_X1 U7974 ( .A(n6288), .B(P2_REG1_REG_11__SCAN_IN), .S(n6306), .Z(n6292)
         );
  AOI21_X1 U7975 ( .B1(n6290), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6289), .ZN(
        n6291) );
  NOR2_X1 U7976 ( .A1(n6291), .A2(n6292), .ZN(n6305) );
  AOI21_X1 U7977 ( .B1(n6292), .B2(n6291), .A(n6305), .ZN(n6293) );
  NAND2_X1 U7978 ( .A1(n9849), .A2(n6293), .ZN(n6294) );
  OAI211_X1 U7979 ( .C1(n9852), .C2(n6300), .A(n6295), .B(n6294), .ZN(n6296)
         );
  INV_X1 U7980 ( .A(n6296), .ZN(n6297) );
  OAI21_X1 U7981 ( .B1(n6298), .B2(n8227), .A(n6297), .ZN(P2_U3256) );
  NAND2_X1 U7982 ( .A1(n8207), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6301) );
  INV_X1 U7983 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8201) );
  AOI21_X1 U7984 ( .B1(n6300), .B2(n6838), .A(n6299), .ZN(n8204) );
  OAI211_X1 U7985 ( .C1(n8207), .C2(P2_REG2_REG_12__SCAN_IN), .A(n8204), .B(
        n6301), .ZN(n8202) );
  NAND2_X1 U7986 ( .A1(n6301), .A2(n8202), .ZN(n6303) );
  AOI22_X1 U7987 ( .A1(n6407), .A2(n7124), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6317), .ZN(n6302) );
  NOR2_X1 U7988 ( .A1(n6303), .A2(n6302), .ZN(n6402) );
  AOI21_X1 U7989 ( .B1(n6303), .B2(n6302), .A(n6402), .ZN(n6304) );
  OR2_X1 U7990 ( .A1(n6304), .A2(n8227), .ZN(n6316) );
  AOI22_X1 U7991 ( .A1(n6407), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5409), .B2(
        n6317), .ZN(n6311) );
  AOI21_X1 U7992 ( .B1(n6306), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6305), .ZN(
        n8210) );
  MUX2_X1 U7993 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6307), .S(n8207), .Z(n8209)
         );
  NAND2_X1 U7994 ( .A1(n8210), .A2(n8209), .ZN(n8208) );
  NAND2_X1 U7995 ( .A1(n6308), .A2(n6307), .ZN(n6309) );
  NAND2_X1 U7996 ( .A1(n8208), .A2(n6309), .ZN(n6310) );
  NAND2_X1 U7997 ( .A1(n6311), .A2(n6310), .ZN(n6406) );
  OAI21_X1 U7998 ( .B1(n6311), .B2(n6310), .A(n6406), .ZN(n6314) );
  INV_X1 U7999 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U8000 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6936) );
  OAI21_X1 U8001 ( .B1(n9488), .B2(n6312), .A(n6936), .ZN(n6313) );
  AOI21_X1 U8002 ( .B1(n9849), .B2(n6314), .A(n6313), .ZN(n6315) );
  OAI211_X1 U8003 ( .C1(n9852), .C2(n6317), .A(n6316), .B(n6315), .ZN(P2_U3258) );
  INV_X1 U8004 ( .A(n6331), .ZN(n6330) );
  NAND2_X1 U8005 ( .A1(n9024), .A2(n7893), .ZN(n6324) );
  INV_X2 U8006 ( .A(n4479), .ZN(n7473) );
  NAND2_X1 U8007 ( .A1(n7473), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U8008 ( .A1(n7502), .A2(n6391), .ZN(n6319) );
  OAI211_X2 U8009 ( .C1(n6321), .C2(n6749), .A(n6320), .B(n6319), .ZN(n6819)
         );
  NAND2_X1 U8010 ( .A1(n6819), .A2(n8005), .ZN(n6323) );
  NAND2_X1 U8011 ( .A1(n6324), .A2(n6323), .ZN(n6325) );
  XNOR2_X1 U8012 ( .A(n6325), .B(n7996), .ZN(n6328) );
  AND2_X1 U8013 ( .A1(n6819), .A2(n7893), .ZN(n6326) );
  AOI21_X1 U8014 ( .B1(n9024), .B2(n7998), .A(n6326), .ZN(n6327) );
  OR2_X1 U8015 ( .A1(n6328), .A2(n6327), .ZN(n6329) );
  NAND2_X1 U8016 ( .A1(n6328), .A2(n6327), .ZN(n6503) );
  AND2_X1 U8017 ( .A1(n6329), .A2(n6503), .ZN(n6333) );
  NOR2_X1 U8018 ( .A1(n6330), .A2(n6333), .ZN(n6336) );
  NAND2_X1 U8019 ( .A1(n6332), .A2(n6331), .ZN(n6334) );
  NAND2_X1 U8020 ( .A1(n6334), .A2(n6333), .ZN(n6454) );
  INV_X1 U8021 ( .A(n6454), .ZN(n6335) );
  AOI21_X1 U8022 ( .B1(n6336), .B2(n6332), .A(n6335), .ZN(n6346) );
  NAND2_X1 U8023 ( .A1(n6444), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6342) );
  INV_X1 U8024 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6337) );
  OR2_X1 U8025 ( .A1(n6273), .A2(n6337), .ZN(n6341) );
  INV_X1 U8026 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6902) );
  OR2_X1 U8027 ( .A1(n6274), .A2(n6902), .ZN(n6340) );
  OR2_X1 U8028 ( .A1(n6338), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6339) );
  INV_X1 U8029 ( .A(n9774), .ZN(n9023) );
  AOI22_X1 U8030 ( .A1(n7390), .A2(n6570), .B1(n8713), .B2(n9023), .ZN(n6345)
         );
  AOI22_X1 U8031 ( .A1(n6819), .A2(n8692), .B1(n6343), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6344) );
  OAI211_X1 U8032 ( .C1(n6346), .C2(n8719), .A(n6345), .B(n6344), .ZN(P1_U3235) );
  NOR2_X1 U8033 ( .A1(n6514), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9856) );
  NOR2_X1 U8034 ( .A1(n8063), .A2(n9894), .ZN(n6347) );
  AOI211_X1 U8035 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n8088), .A(n9856), .B(
        n6347), .ZN(n6352) );
  OAI22_X1 U8036 ( .A1(n8105), .A2(n6348), .B1(n9894), .B2(n8082), .ZN(n6350)
         );
  NAND2_X1 U8037 ( .A1(n6350), .A2(n6349), .ZN(n6351) );
  OAI211_X1 U8038 ( .C1(n6353), .C2(n8096), .A(n6352), .B(n6351), .ZN(P2_U3234) );
  NOR2_X1 U8039 ( .A1(n6355), .A2(n6354), .ZN(n6357) );
  INV_X1 U8040 ( .A(n8386), .ZN(n6356) );
  INV_X1 U8041 ( .A(n6369), .ZN(n6358) );
  INV_X1 U8042 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6368) );
  XOR2_X1 U8043 ( .A(n6359), .B(n7844), .Z(n6558) );
  INV_X1 U8044 ( .A(n6360), .ZN(n6362) );
  INV_X1 U8045 ( .A(n6438), .ZN(n6361) );
  AOI211_X1 U8046 ( .C1(n6555), .C2(n6362), .A(n9973), .B(n6361), .ZN(n6550)
         );
  XOR2_X1 U8047 ( .A(n7844), .B(n6363), .Z(n6365) );
  INV_X1 U8048 ( .A(n9868), .ZN(n9576) );
  OAI21_X1 U8049 ( .B1(n6365), .B2(n9576), .A(n6364), .ZN(n6549) );
  AOI211_X1 U8050 ( .C1(n9962), .C2(n6555), .A(n6550), .B(n6549), .ZN(n6366)
         );
  OAI21_X1 U8051 ( .B1(n9966), .B2(n6558), .A(n6366), .ZN(n6371) );
  NAND2_X1 U8052 ( .A1(n6371), .A2(n9979), .ZN(n6367) );
  OAI21_X1 U8053 ( .B1(n9979), .B2(n6368), .A(n6367), .ZN(P2_U3466) );
  NAND2_X1 U8054 ( .A1(n6371), .A2(n9995), .ZN(n6372) );
  OAI21_X1 U8055 ( .B1(n9995), .B2(n5208), .A(n6372), .ZN(P2_U3525) );
  INV_X1 U8056 ( .A(n6373), .ZN(n6382) );
  INV_X1 U8057 ( .A(n9113), .ZN(n6375) );
  OR2_X1 U8058 ( .A1(n6375), .A2(n6374), .ZN(n9006) );
  NAND2_X1 U8059 ( .A1(n6377), .A2(n6376), .ZN(n6378) );
  OAI211_X1 U8060 ( .C1(n6379), .C2(n9006), .A(n9025), .B(n6378), .ZN(n6380)
         );
  AOI21_X1 U8061 ( .B1(n6382), .B2(n6381), .A(n6380), .ZN(n9651) );
  OAI211_X1 U8062 ( .C1(n6385), .C2(n6384), .A(n9750), .B(n6383), .ZN(n6387)
         );
  NAND2_X1 U8063 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6386) );
  OAI211_X1 U8064 ( .C1(n10090), .C2(n9735), .A(n6387), .B(n6386), .ZN(n6395)
         );
  OAI211_X1 U8065 ( .C1(n6390), .C2(n6389), .A(n9740), .B(n6388), .ZN(n6393)
         );
  NAND2_X1 U8066 ( .A1(n9742), .A2(n6391), .ZN(n6392) );
  NAND2_X1 U8067 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  OR3_X1 U8068 ( .A1(n9651), .A2(n6395), .A3(n6394), .ZN(P1_U3243) );
  NAND2_X1 U8069 ( .A1(n4548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6396) );
  XNOR2_X1 U8070 ( .A(n6396), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9091) );
  INV_X1 U8071 ( .A(n9091), .ZN(n9081) );
  INV_X1 U8072 ( .A(n7403), .ZN(n6398) );
  OAI222_X1 U8073 ( .A1(P1_U3084), .A2(n9081), .B1(n9463), .B2(n6398), .C1(
        n6397), .C2(n7885), .ZN(P1_U3337) );
  INV_X1 U8074 ( .A(n7190), .ZN(n6976) );
  OAI222_X1 U8075 ( .A1(n8546), .A2(n6399), .B1(n8548), .B2(n6398), .C1(n6976), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8076 ( .A(n7497), .ZN(n6416) );
  XNOR2_X1 U8077 ( .A(n6400), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9105) );
  AOI22_X1 U8078 ( .A1(n9105), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9465), .ZN(n6401) );
  OAI21_X1 U8079 ( .B1(n6416), .B2(n9463), .A(n6401), .ZN(P1_U3336) );
  NOR2_X1 U8080 ( .A1(n6407), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6403) );
  NOR2_X1 U8081 ( .A1(n6403), .A2(n6402), .ZN(n6405) );
  AOI22_X1 U8082 ( .A1(n6925), .A2(n7174), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n6411), .ZN(n6404) );
  NOR2_X1 U8083 ( .A1(n6405), .A2(n6404), .ZN(n6921) );
  AOI21_X1 U8084 ( .B1(n6405), .B2(n6404), .A(n6921), .ZN(n6415) );
  INV_X1 U8085 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9614) );
  AOI22_X1 U8086 ( .A1(n6925), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9614), .B2(
        n6411), .ZN(n6409) );
  OAI21_X1 U8087 ( .B1(n6407), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6406), .ZN(
        n6408) );
  NAND2_X1 U8088 ( .A1(n6409), .A2(n6408), .ZN(n6924) );
  OAI21_X1 U8089 ( .B1(n6409), .B2(n6408), .A(n6924), .ZN(n6413) );
  NAND2_X1 U8090 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7087) );
  NAND2_X1 U8091 ( .A1(n9857), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6410) );
  OAI211_X1 U8092 ( .C1(n9852), .C2(n6411), .A(n7087), .B(n6410), .ZN(n6412)
         );
  AOI21_X1 U8093 ( .B1(n6413), .B2(n9849), .A(n6412), .ZN(n6414) );
  OAI21_X1 U8094 ( .B1(n6415), .B2(n8227), .A(n6414), .ZN(P2_U3259) );
  INV_X1 U8095 ( .A(n7201), .ZN(n7198) );
  OAI222_X1 U8096 ( .A1(n8546), .A2(n6417), .B1(n8548), .B2(n6416), .C1(n7198), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U8097 ( .A1(n9565), .A2(n6418), .ZN(n6419) );
  INV_X1 U8098 ( .A(n7731), .ZN(n7848) );
  XNOR2_X1 U8099 ( .A(n6420), .B(n7848), .ZN(n9937) );
  XNOR2_X1 U8100 ( .A(n6421), .B(n7848), .ZN(n6424) );
  NAND2_X1 U8101 ( .A1(n8121), .A2(n9864), .ZN(n6422) );
  OAI21_X1 U8102 ( .B1(n6620), .B2(n9581), .A(n6422), .ZN(n6423) );
  AOI21_X1 U8103 ( .B1(n6424), .B2(n9868), .A(n6423), .ZN(n9936) );
  MUX2_X1 U8104 ( .A(n6425), .B(n9936), .S(n9591), .Z(n6429) );
  XOR2_X1 U8105 ( .A(n9933), .B(n6440), .Z(n9934) );
  OAI22_X1 U8106 ( .A1(n9881), .A2(n4592), .B1(n9871), .B2(n6426), .ZN(n6427)
         );
  AOI21_X1 U8107 ( .B1(n8456), .B2(n9934), .A(n6427), .ZN(n6428) );
  OAI211_X1 U8108 ( .C1(n8458), .C2(n9937), .A(n6429), .B(n6428), .ZN(P2_U3289) );
  INV_X1 U8109 ( .A(n6433), .ZN(n7845) );
  XNOR2_X1 U8110 ( .A(n6430), .B(n7845), .ZN(n9928) );
  OAI21_X1 U8111 ( .B1(n6433), .B2(n6432), .A(n6431), .ZN(n6436) );
  NAND2_X1 U8112 ( .A1(n9866), .A2(n9864), .ZN(n6434) );
  OAI21_X1 U8113 ( .B1(n8095), .B2(n9581), .A(n6434), .ZN(n6435) );
  AOI21_X1 U8114 ( .B1(n6436), .B2(n9868), .A(n6435), .ZN(n9931) );
  MUX2_X1 U8115 ( .A(n6437), .B(n9931), .S(n9591), .Z(n6443) );
  NAND2_X1 U8116 ( .A1(n6438), .A2(n9926), .ZN(n6439) );
  AND2_X1 U8117 ( .A1(n6440), .A2(n6439), .ZN(n9927) );
  OAI22_X1 U8118 ( .A1(n9881), .A2(n4785), .B1(n9871), .B2(n8093), .ZN(n6441)
         );
  AOI21_X1 U8119 ( .B1(n8456), .B2(n9927), .A(n6441), .ZN(n6442) );
  OAI211_X1 U8120 ( .C1(n9928), .C2(n8458), .A(n6443), .B(n6442), .ZN(P2_U3290) );
  NAND2_X1 U8121 ( .A1(n6444), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6449) );
  INV_X1 U8122 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6445) );
  OR2_X1 U8123 ( .A1(n6274), .A2(n6445), .ZN(n6448) );
  XNOR2_X1 U8124 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9791) );
  OR2_X1 U8125 ( .A1(n6338), .A2(n9791), .ZN(n6446) );
  NAND2_X1 U8126 ( .A1(n7473), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U8127 ( .A1(n7502), .A2(n9646), .ZN(n6450) );
  OAI211_X1 U8128 ( .C1(n6452), .C2(n6749), .A(n6451), .B(n6450), .ZN(n6673)
         );
  INV_X1 U8129 ( .A(n6673), .ZN(n9808) );
  OAI22_X1 U8130 ( .A1(n6633), .A2(n8003), .B1(n9808), .B2(n7985), .ZN(n6453)
         );
  XNOR2_X1 U8131 ( .A(n6453), .B(n7996), .ZN(n6775) );
  OAI22_X1 U8132 ( .A1(n6633), .A2(n4868), .B1(n9808), .B2(n8003), .ZN(n6773)
         );
  XNOR2_X1 U8133 ( .A(n6775), .B(n6773), .ZN(n6468) );
  NAND2_X1 U8134 ( .A1(n6454), .A2(n6503), .ZN(n6465) );
  NAND2_X1 U8135 ( .A1(n7473), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U8136 ( .A1(n7502), .A2(n6455), .ZN(n6456) );
  OAI22_X1 U8137 ( .A1(n9774), .A2(n8003), .B1(n6903), .B2(n7985), .ZN(n6459)
         );
  XNOR2_X1 U8138 ( .A(n6459), .B(n7996), .ZN(n6461) );
  OAI22_X1 U8139 ( .A1(n9774), .A2(n4868), .B1(n6903), .B2(n8003), .ZN(n6462)
         );
  INV_X1 U8140 ( .A(n6462), .ZN(n6460) );
  NAND2_X1 U8141 ( .A1(n6461), .A2(n6460), .ZN(n6466) );
  INV_X1 U8142 ( .A(n6461), .ZN(n6463) );
  NAND2_X1 U8143 ( .A1(n6463), .A2(n6462), .ZN(n6464) );
  AND2_X1 U8144 ( .A1(n6466), .A2(n6464), .ZN(n6505) );
  NAND2_X1 U8145 ( .A1(n6506), .A2(n6466), .ZN(n6467) );
  NAND2_X1 U8146 ( .A1(n6467), .A2(n6468), .ZN(n6777) );
  OAI21_X1 U8147 ( .B1(n6468), .B2(n6467), .A(n6777), .ZN(n6489) );
  INV_X1 U8148 ( .A(n6469), .ZN(n6472) );
  NAND3_X1 U8149 ( .A1(n6470), .A2(n7006), .A3(n6195), .ZN(n6471) );
  AOI21_X1 U8150 ( .B1(n6473), .B2(n6472), .A(n6471), .ZN(n6474) );
  OR2_X1 U8151 ( .A1(n6474), .A2(P1_U3084), .ZN(n6476) );
  AOI22_X1 U8152 ( .A1(n7390), .A2(n9023), .B1(n8692), .B2(n6673), .ZN(n6487)
         );
  NAND2_X1 U8153 ( .A1(n7624), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6485) );
  INV_X1 U8154 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6477) );
  OR2_X1 U8155 ( .A1(n7628), .A2(n6477), .ZN(n6484) );
  NAND3_X1 U8156 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6648) );
  INV_X1 U8157 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8158 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6478) );
  NAND2_X1 U8159 ( .A1(n6479), .A2(n6478), .ZN(n6480) );
  NAND2_X1 U8160 ( .A1(n6648), .A2(n6480), .ZN(n9754) );
  OR2_X1 U8161 ( .A1(n7623), .A2(n9754), .ZN(n6483) );
  INV_X1 U8162 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6481) );
  OR2_X1 U8163 ( .A1(n6274), .A2(n6481), .ZN(n6482) );
  AND2_X1 U8164 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9652) );
  AOI21_X1 U8165 ( .B1(n8713), .B2(n9021), .A(n9652), .ZN(n6486) );
  OAI211_X1 U8166 ( .C1(n8715), .C2(n9791), .A(n6487), .B(n6486), .ZN(n6488)
         );
  AOI21_X1 U8167 ( .B1(n6489), .B2(n8645), .A(n6488), .ZN(n6490) );
  INV_X1 U8168 ( .A(n6490), .ZN(P1_U3228) );
  INV_X1 U8169 ( .A(n7839), .ZN(n6493) );
  XNOR2_X1 U8170 ( .A(n6491), .B(n6493), .ZN(n9907) );
  OAI21_X1 U8171 ( .B1(n9899), .B2(n9908), .A(n6520), .ZN(n9909) );
  XNOR2_X1 U8172 ( .A(n6492), .B(n6493), .ZN(n6494) );
  NAND2_X1 U8173 ( .A1(n6494), .A2(n9868), .ZN(n6497) );
  AOI22_X1 U8174 ( .A1(n9864), .A2(n8124), .B1(n5855), .B2(n9865), .ZN(n6496)
         );
  NAND2_X1 U8175 ( .A1(n6497), .A2(n6496), .ZN(n9912) );
  NAND2_X1 U8176 ( .A1(n8436), .A2(n9912), .ZN(n6500) );
  OAI22_X1 U8177 ( .A1(n9871), .A2(n5145), .B1(n6105), .B2(n9591), .ZN(n6498)
         );
  INV_X1 U8178 ( .A(n6498), .ZN(n6499) );
  OAI211_X1 U8179 ( .C1(n9873), .C2(n9909), .A(n6500), .B(n6499), .ZN(n6501)
         );
  AOI21_X1 U8180 ( .B1(n8440), .B2(n8087), .A(n6501), .ZN(n6502) );
  OAI21_X1 U8181 ( .B1(n9907), .B2(n8458), .A(n6502), .ZN(P2_U3294) );
  INV_X1 U8182 ( .A(n6503), .ZN(n6504) );
  NOR2_X1 U8183 ( .A1(n6505), .A2(n6504), .ZN(n6508) );
  INV_X1 U8184 ( .A(n6506), .ZN(n6507) );
  AOI21_X1 U8185 ( .B1(n6508), .B2(n6454), .A(n6507), .ZN(n6513) );
  AOI22_X1 U8186 ( .A1(n6612), .A2(n8717), .B1(n8713), .B2(n9022), .ZN(n6512)
         );
  NOR2_X1 U8187 ( .A1(n8715), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6509) );
  AOI211_X1 U8188 ( .C1(n7390), .C2(n9024), .A(n6510), .B(n6509), .ZN(n6511)
         );
  OAI211_X1 U8189 ( .C1(n6513), .C2(n8719), .A(n6512), .B(n6511), .ZN(P1_U3216) );
  NAND2_X1 U8190 ( .A1(n6157), .A2(n9894), .ZN(n7699) );
  NAND2_X1 U8191 ( .A1(n6538), .A2(n7699), .ZN(n7838) );
  INV_X1 U8192 ( .A(n7838), .ZN(n9896) );
  AOI22_X1 U8193 ( .A1(n7838), .A2(n9868), .B1(n9865), .B2(n8124), .ZN(n9893)
         );
  OAI22_X1 U8194 ( .A1(n9593), .A2(n9893), .B1(n6514), .B2(n9871), .ZN(n6515)
         );
  AOI21_X1 U8195 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9593), .A(n6515), .ZN(
        n6518) );
  OAI21_X1 U8196 ( .B1(n8440), .B2(n8456), .A(n6516), .ZN(n6517) );
  OAI211_X1 U8197 ( .C1(n9896), .C2(n8458), .A(n6518), .B(n6517), .ZN(P2_U3296) );
  XNOR2_X1 U8198 ( .A(n6519), .B(n7842), .ZN(n9913) );
  NAND2_X1 U8199 ( .A1(n6520), .A2(n5853), .ZN(n6521) );
  NAND2_X1 U8200 ( .A1(n9870), .A2(n6521), .ZN(n9915) );
  OAI22_X1 U8201 ( .A1(n9873), .A2(n9915), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9871), .ZN(n6523) );
  NOR2_X1 U8202 ( .A1(n8436), .A2(n6104), .ZN(n6522) );
  AOI211_X1 U8203 ( .C1(n8440), .C2(n5853), .A(n6523), .B(n6522), .ZN(n6532)
         );
  OAI21_X1 U8204 ( .B1(n6525), .B2(n7842), .A(n6524), .ZN(n6529) );
  OAI22_X1 U8205 ( .A1(n6527), .A2(n9579), .B1(n6526), .B2(n9581), .ZN(n6528)
         );
  AOI21_X1 U8206 ( .B1(n6529), .B2(n9868), .A(n6528), .ZN(n6530) );
  OAI21_X1 U8207 ( .B1(n9913), .B2(n9565), .A(n6530), .ZN(n9916) );
  NAND2_X1 U8208 ( .A1(n9916), .A2(n8436), .ZN(n6531) );
  OAI211_X1 U8209 ( .C1(n9913), .C2(n9584), .A(n6532), .B(n6531), .ZN(P2_U3293) );
  XOR2_X1 U8210 ( .A(n9902), .B(n8124), .Z(n7841) );
  XOR2_X1 U8211 ( .A(n6533), .B(n7841), .Z(n9905) );
  NOR2_X1 U8212 ( .A1(n9871), .A2(n6534), .ZN(n6537) );
  NOR2_X1 U8213 ( .A1(n6535), .A2(n9894), .ZN(n9900) );
  NOR3_X1 U8214 ( .A1(n9873), .A2(n9899), .A3(n9900), .ZN(n6536) );
  AOI211_X1 U8215 ( .C1(n8440), .C2(n9902), .A(n6537), .B(n6536), .ZN(n6542)
         );
  XNOR2_X1 U8216 ( .A(n7841), .B(n6538), .ZN(n6539) );
  AOI222_X1 U8217 ( .A1(n9868), .A2(n6539), .B1(n6158), .B2(n9865), .C1(n6157), 
        .C2(n9864), .ZN(n9904) );
  MUX2_X1 U8218 ( .A(n6540), .B(n9904), .S(n9591), .Z(n6541) );
  OAI211_X1 U8219 ( .C1(n8458), .C2(n9905), .A(n6542), .B(n6541), .ZN(P2_U3295) );
  INV_X1 U8220 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6543) );
  INV_X1 U8221 ( .A(n7492), .ZN(n6548) );
  INV_X1 U8222 ( .A(n8220), .ZN(n7205) );
  OAI222_X1 U8223 ( .A1(n8546), .A2(n6543), .B1(n8548), .B2(n6548), .C1(
        P2_U3152), .C2(n7205), .ZN(P2_U3340) );
  NAND2_X1 U8224 ( .A1(n6400), .A2(n6544), .ZN(n6545) );
  NAND2_X1 U8225 ( .A1(n6545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6546) );
  XNOR2_X1 U8226 ( .A(n6546), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9741) );
  INV_X1 U8227 ( .A(n9741), .ZN(n9103) );
  INV_X1 U8228 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6547) );
  OAI222_X1 U8229 ( .A1(n9103), .A2(P1_U3084), .B1(n9463), .B2(n6548), .C1(
        n6547), .C2(n7885), .ZN(P1_U3335) );
  AOI21_X1 U8230 ( .B1(n6550), .B2(n7687), .A(n6549), .ZN(n6551) );
  MUX2_X1 U8231 ( .A(n6552), .B(n6551), .S(n9591), .Z(n6557) );
  INV_X1 U8232 ( .A(n9871), .ZN(n9586) );
  INV_X1 U8233 ( .A(n6553), .ZN(n6554) );
  AOI22_X1 U8234 ( .A1(n8440), .A2(n6555), .B1(n9586), .B2(n6554), .ZN(n6556)
         );
  OAI211_X1 U8235 ( .C1(n6558), .C2(n8458), .A(n6557), .B(n6556), .ZN(P2_U3291) );
  INV_X1 U8236 ( .A(n9455), .ZN(n6562) );
  NAND4_X1 U8237 ( .A1(n6562), .A2(n6561), .A3(n6560), .A4(n6559), .ZN(n6565)
         );
  OAI21_X1 U8238 ( .B1(n4770), .B2(n9790), .A(n6563), .ZN(n6564) );
  NAND2_X1 U8239 ( .A1(n6564), .A2(n9786), .ZN(n6569) );
  NOR2_X1 U8240 ( .A1(n6565), .A2(n9785), .ZN(n9521) );
  INV_X1 U8241 ( .A(n9521), .ZN(n7157) );
  INV_X1 U8242 ( .A(n9784), .ZN(n6567) );
  OAI21_X1 U8243 ( .B1(n9333), .B2(n9516), .A(n6583), .ZN(n6568) );
  OAI211_X1 U8244 ( .C1(n6183), .C2(n9786), .A(n6569), .B(n6568), .ZN(P1_U3291) );
  NAND2_X1 U8245 ( .A1(n6570), .A2(n9797), .ZN(n8747) );
  AND2_X1 U8246 ( .A1(n9026), .A2(n6583), .ZN(n6571) );
  NAND2_X1 U8247 ( .A1(n6576), .A2(n6571), .ZN(n6601) );
  OAI21_X1 U8248 ( .B1(n6576), .B2(n6571), .A(n6601), .ZN(n9795) );
  NOR2_X1 U8249 ( .A1(n4473), .A2(n6572), .ZN(n6573) );
  NAND2_X1 U8250 ( .A1(n9786), .A2(n6573), .ZN(n7005) );
  NAND2_X1 U8251 ( .A1(n8001), .A2(n6574), .ZN(n9761) );
  OR2_X1 U8252 ( .A1(n9761), .A2(n9785), .ZN(n9779) );
  INV_X1 U8253 ( .A(n6576), .ZN(n6577) );
  OAI21_X1 U8254 ( .B1(n6577), .B2(n4633), .A(n6605), .ZN(n6581) );
  NAND2_X1 U8255 ( .A1(n9785), .A2(n8795), .ZN(n6579) );
  NAND2_X1 U8256 ( .A1(n8964), .A2(n9001), .ZN(n6578) );
  INV_X1 U8257 ( .A(n9024), .ZN(n6606) );
  OAI22_X1 U8258 ( .A1(n4867), .A2(n9773), .B1(n6606), .B2(n9771), .ZN(n6580)
         );
  AOI21_X1 U8259 ( .B1(n6581), .B2(n9776), .A(n6580), .ZN(n6582) );
  OAI21_X1 U8260 ( .B1(n9779), .B2(n9795), .A(n6582), .ZN(n9798) );
  OR2_X1 U8261 ( .A1(n6599), .A2(n6583), .ZN(n6816) );
  OAI211_X1 U8262 ( .C1(n9797), .C2(n6584), .A(n9782), .B(n6816), .ZN(n9796)
         );
  OAI22_X1 U8263 ( .A1(n9796), .A2(n9785), .B1(n6585), .B2(n9790), .ZN(n6586)
         );
  OAI21_X1 U8264 ( .B1(n9798), .B2(n6586), .A(n9786), .ZN(n6588) );
  AOI22_X1 U8265 ( .A1(n9516), .A2(n6599), .B1(n9767), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6587) );
  OAI211_X1 U8266 ( .C1(n9795), .C2(n7005), .A(n6588), .B(n6587), .ZN(P1_U3290) );
  INV_X1 U8267 ( .A(n6680), .ZN(n8118) );
  AOI22_X1 U8268 ( .A1(n8106), .A2(n8120), .B1(n8084), .B2(n8118), .ZN(n6589)
         );
  NAND2_X1 U8269 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8190) );
  OAI211_X1 U8270 ( .C1(n6590), .C2(n8094), .A(n6589), .B(n8190), .ZN(n6597)
         );
  NAND3_X1 U8271 ( .A1(n8078), .A2(n6591), .A3(n8120), .ZN(n6595) );
  OAI21_X1 U8272 ( .B1(n6593), .B2(n6592), .A(n8101), .ZN(n6594) );
  AOI21_X1 U8273 ( .B1(n6595), .B2(n6594), .A(n4554), .ZN(n6596) );
  AOI211_X1 U8274 ( .C1(n6681), .C2(n8098), .A(n6597), .B(n6596), .ZN(n6598)
         );
  INV_X1 U8275 ( .A(n6598), .ZN(P2_U3223) );
  NAND2_X1 U8276 ( .A1(n6570), .A2(n6599), .ZN(n6600) );
  NAND2_X1 U8277 ( .A1(n6601), .A2(n6600), .ZN(n6807) );
  INV_X1 U8278 ( .A(n6807), .ZN(n6602) );
  INV_X1 U8279 ( .A(n6809), .ZN(n8940) );
  NAND2_X1 U8280 ( .A1(n6602), .A2(n8940), .ZN(n6805) );
  INV_X1 U8281 ( .A(n6819), .ZN(n9802) );
  NAND2_X1 U8282 ( .A1(n6606), .A2(n9802), .ZN(n6603) );
  NAND2_X1 U8283 ( .A1(n6805), .A2(n6603), .ZN(n6635) );
  NAND2_X1 U8284 ( .A1(n9774), .A2(n6612), .ZN(n8971) );
  NAND2_X1 U8285 ( .A1(n9023), .A2(n6903), .ZN(n8750) );
  NAND2_X1 U8286 ( .A1(n6635), .A2(n6634), .ZN(n9765) );
  OAI21_X1 U8287 ( .B1(n6635), .B2(n6634), .A(n9765), .ZN(n6907) );
  INV_X1 U8288 ( .A(n6907), .ZN(n6614) );
  INV_X1 U8289 ( .A(n9779), .ZN(n9512) );
  OAI22_X1 U8290 ( .A1(n6606), .A2(n9773), .B1(n6633), .B2(n9771), .ZN(n6610)
         );
  NAND2_X1 U8291 ( .A1(n6810), .A2(n6809), .ZN(n6808) );
  NAND2_X1 U8292 ( .A1(n6606), .A2(n6819), .ZN(n6607) );
  INV_X1 U8293 ( .A(n8979), .ZN(n8749) );
  NAND2_X1 U8294 ( .A1(n8749), .A2(n6634), .ZN(n6608) );
  INV_X1 U8295 ( .A(n6634), .ZN(n8937) );
  AOI21_X1 U8296 ( .B1(n6608), .B2(n6658), .A(n9509), .ZN(n6609) );
  AOI211_X1 U8297 ( .C1(n9512), .C2(n6907), .A(n6610), .B(n6609), .ZN(n6910)
         );
  NOR2_X1 U8298 ( .A1(n6816), .A2(n6819), .ZN(n6611) );
  INV_X1 U8299 ( .A(n6611), .ZN(n6817) );
  AOI21_X1 U8300 ( .B1(n6612), .B2(n6817), .A(n9783), .ZN(n6906) );
  AOI22_X1 U8301 ( .A1(n6906), .A2(n9782), .B1(n9524), .B2(n6612), .ZN(n6613)
         );
  OAI211_X1 U8302 ( .C1(n6614), .C2(n6787), .A(n6910), .B(n6613), .ZN(n6616)
         );
  NAND2_X1 U8303 ( .A1(n6616), .A2(n4474), .ZN(n6615) );
  OAI21_X1 U8304 ( .B1(n4474), .B2(n6337), .A(n6615), .ZN(P1_U3463) );
  NAND2_X1 U8305 ( .A1(n6616), .A2(n9848), .ZN(n6617) );
  OAI21_X1 U8306 ( .B1(n9848), .B2(n5963), .A(n6617), .ZN(P1_U3526) );
  NOR3_X1 U8307 ( .A1(n8105), .A2(n6618), .A3(n6620), .ZN(n6619) );
  AOI21_X1 U8308 ( .B1(n4554), .B2(n8101), .A(n6619), .ZN(n6631) );
  INV_X1 U8309 ( .A(n6620), .ZN(n8119) );
  NAND2_X1 U8310 ( .A1(n8106), .A2(n8119), .ZN(n6625) );
  INV_X1 U8311 ( .A(n6714), .ZN(n8117) );
  NAND2_X1 U8312 ( .A1(n8084), .A2(n8117), .ZN(n6624) );
  INV_X1 U8313 ( .A(n6691), .ZN(n6621) );
  NAND2_X1 U8314 ( .A1(n8051), .A2(n6621), .ZN(n6622) );
  NAND4_X1 U8315 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6628)
         );
  NOR2_X1 U8316 ( .A1(n6626), .A2(n8082), .ZN(n6627) );
  AOI211_X1 U8317 ( .C1(n6711), .C2(n8098), .A(n6628), .B(n6627), .ZN(n6629)
         );
  OAI21_X1 U8318 ( .B1(n6631), .B2(n6630), .A(n6629), .ZN(P2_U3233) );
  INV_X1 U8319 ( .A(n7501), .ZN(n7884) );
  OAI222_X1 U8320 ( .A1(n8546), .A2(n6632), .B1(n8548), .B2(n7884), .C1(n7687), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U8321 ( .A1(n6633), .A2(n9808), .ZN(n6637) );
  AND2_X1 U8322 ( .A1(n6639), .A2(n6634), .ZN(n6636) );
  NAND2_X1 U8323 ( .A1(n6636), .A2(n6635), .ZN(n6789) );
  NAND2_X1 U8324 ( .A1(n9774), .A2(n6903), .ZN(n9764) );
  NAND2_X1 U8325 ( .A1(n9764), .A2(n6637), .ZN(n6638) );
  NAND2_X1 U8326 ( .A1(n6639), .A2(n6638), .ZN(n6788) );
  NAND2_X1 U8327 ( .A1(n7473), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U8328 ( .A1(n7502), .A2(n9663), .ZN(n6640) );
  INV_X1 U8329 ( .A(n6798), .ZN(n9755) );
  NAND2_X1 U8330 ( .A1(n9772), .A2(n6798), .ZN(n8967) );
  AND2_X1 U8331 ( .A1(n6788), .A2(n6659), .ZN(n6643) );
  NAND2_X1 U8332 ( .A1(n6789), .A2(n6643), .ZN(n6790) );
  NAND2_X1 U8333 ( .A1(n9021), .A2(n6798), .ZN(n6644) );
  NAND2_X1 U8334 ( .A1(n7624), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6653) );
  INV_X1 U8335 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6645) );
  OR2_X1 U8336 ( .A1(n7628), .A2(n6645), .ZN(n6652) );
  INV_X1 U8337 ( .A(n6648), .ZN(n6647) );
  NAND2_X1 U8338 ( .A1(n6647), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6663) );
  INV_X1 U8339 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U8340 ( .A1(n6648), .A2(n6883), .ZN(n6649) );
  NAND2_X1 U8341 ( .A1(n6663), .A2(n6649), .ZN(n6886) );
  OR2_X1 U8342 ( .A1(n7623), .A2(n6886), .ZN(n6651) );
  INV_X1 U8343 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6672) );
  OR2_X1 U8344 ( .A1(n6274), .A2(n6672), .ZN(n6650) );
  NAND2_X1 U8345 ( .A1(n7473), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U8346 ( .A1(n7502), .A2(n9679), .ZN(n6654) );
  NAND2_X1 U8347 ( .A1(n6895), .A2(n6882), .ZN(n8973) );
  INV_X1 U8348 ( .A(n6895), .ZN(n9020) );
  NAND2_X1 U8349 ( .A1(n9020), .A2(n9813), .ZN(n8799) );
  AND2_X1 U8350 ( .A1(n8973), .A2(n8799), .ZN(n6657) );
  INV_X1 U8351 ( .A(n6657), .ZN(n8941) );
  INV_X1 U8352 ( .A(n9817), .ZN(n6679) );
  INV_X1 U8353 ( .A(n6659), .ZN(n8936) );
  NAND2_X1 U8354 ( .A1(n6793), .A2(n8936), .ZN(n6792) );
  NAND2_X1 U8355 ( .A1(n6792), .A2(n8967), .ZN(n8798) );
  XNOR2_X1 U8356 ( .A(n8798), .B(n8941), .ZN(n6671) );
  NAND2_X1 U8357 ( .A1(n7624), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6668) );
  INV_X1 U8358 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6660) );
  OR2_X1 U8359 ( .A1(n7628), .A2(n6660), .ZN(n6667) );
  INV_X1 U8360 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6914) );
  OR2_X1 U8361 ( .A1(n7549), .A2(n6914), .ZN(n6666) );
  INV_X1 U8362 ( .A(n6663), .ZN(n6661) );
  NAND2_X1 U8363 ( .A1(n6661), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6743) );
  INV_X1 U8364 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U8365 ( .A1(n6663), .A2(n6662), .ZN(n6664) );
  NAND2_X1 U8366 ( .A1(n6743), .A2(n6664), .ZN(n6913) );
  OR2_X1 U8367 ( .A1(n7623), .A2(n6913), .ZN(n6665) );
  OAI22_X1 U8368 ( .A1(n7040), .A2(n9771), .B1(n9772), .B2(n9773), .ZN(n6669)
         );
  AOI21_X1 U8369 ( .B1(n9817), .B2(n9512), .A(n6669), .ZN(n6670) );
  OAI21_X1 U8370 ( .B1(n9509), .B2(n6671), .A(n6670), .ZN(n9815) );
  NAND2_X1 U8371 ( .A1(n9815), .A2(n9786), .ZN(n6678) );
  OAI22_X1 U8372 ( .A1(n9786), .A2(n6672), .B1(n6886), .B2(n9790), .ZN(n6676)
         );
  OR2_X1 U8373 ( .A1(n6797), .A2(n9813), .ZN(n6674) );
  NAND2_X1 U8374 ( .A1(n6892), .A2(n6674), .ZN(n9814) );
  NOR2_X1 U8375 ( .A1(n9814), .A2(n9139), .ZN(n6675) );
  AOI211_X1 U8376 ( .C1(n9516), .C2(n6882), .A(n6676), .B(n6675), .ZN(n6677)
         );
  OAI211_X1 U8377 ( .C1(n6679), .C2(n7005), .A(n6678), .B(n6677), .ZN(P1_U3285) );
  OR2_X1 U8378 ( .A1(n6711), .A2(n6680), .ZN(n7742) );
  AND2_X1 U8379 ( .A1(n6711), .A2(n6680), .ZN(n7740) );
  INV_X1 U8380 ( .A(n7740), .ZN(n7744) );
  INV_X1 U8381 ( .A(n6683), .ZN(n6685) );
  INV_X1 U8382 ( .A(n6713), .ZN(n6686) );
  AOI21_X1 U8383 ( .B1(n7849), .B2(n6683), .A(n6686), .ZN(n9947) );
  AOI22_X1 U8384 ( .A1(n9864), .A2(n8119), .B1(n8117), .B2(n9865), .ZN(n6690)
         );
  XNOR2_X1 U8385 ( .A(n6718), .B(n7849), .ZN(n6688) );
  NAND2_X1 U8386 ( .A1(n6688), .A2(n9868), .ZN(n6689) );
  OAI211_X1 U8387 ( .C1(n9947), .C2(n9565), .A(n6690), .B(n6689), .ZN(n9950)
         );
  NAND2_X1 U8388 ( .A1(n9950), .A2(n8436), .ZN(n6698) );
  OAI22_X1 U8389 ( .A1(n9591), .A2(n6692), .B1(n6691), .B2(n9871), .ZN(n6696)
         );
  INV_X1 U8390 ( .A(n6711), .ZN(n9948) );
  OR2_X1 U8391 ( .A1(n6693), .A2(n9948), .ZN(n6694) );
  NAND2_X1 U8392 ( .A1(n6726), .A2(n6694), .ZN(n9949) );
  NOR2_X1 U8393 ( .A1(n9949), .A2(n9873), .ZN(n6695) );
  AOI211_X1 U8394 ( .C1(n8440), .C2(n6711), .A(n6696), .B(n6695), .ZN(n6697)
         );
  OAI211_X1 U8395 ( .C1(n9947), .C2(n9584), .A(n6698), .B(n6697), .ZN(P2_U3287) );
  INV_X1 U8396 ( .A(n6699), .ZN(n6700) );
  AOI21_X1 U8397 ( .B1(n6701), .B2(n6700), .A(n8082), .ZN(n6705) );
  NOR3_X1 U8398 ( .A1(n8105), .A2(n6702), .A3(n6714), .ZN(n6704) );
  OAI21_X1 U8399 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6710) );
  OAI22_X1 U8400 ( .A1(n8094), .A2(n6837), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6706), .ZN(n6708) );
  OAI22_X1 U8401 ( .A1(n7115), .A2(n8096), .B1(n8058), .B2(n6714), .ZN(n6707)
         );
  AOI211_X1 U8402 ( .C1(n9961), .C2(n8098), .A(n6708), .B(n6707), .ZN(n6709)
         );
  NAND2_X1 U8403 ( .A1(n6710), .A2(n6709), .ZN(P2_U3238) );
  OR2_X1 U8404 ( .A1(n6711), .A2(n8118), .ZN(n6712) );
  NAND2_X1 U8405 ( .A1(n6825), .A2(n6714), .ZN(n7746) );
  NAND2_X1 U8406 ( .A1(n6716), .A2(n7851), .ZN(n6717) );
  NAND2_X1 U8407 ( .A1(n6827), .A2(n6717), .ZN(n9953) );
  INV_X1 U8408 ( .A(n6718), .ZN(n6719) );
  NAND2_X1 U8409 ( .A1(n6719), .A2(n7744), .ZN(n6720) );
  NAND2_X1 U8410 ( .A1(n6720), .A2(n7742), .ZN(n6721) );
  NAND2_X1 U8411 ( .A1(n6721), .A2(n7851), .ZN(n6830) );
  OAI211_X1 U8412 ( .C1(n6721), .C2(n7851), .A(n6830), .B(n9868), .ZN(n6723)
         );
  INV_X1 U8413 ( .A(n6828), .ZN(n8116) );
  AOI22_X1 U8414 ( .A1(n9865), .A2(n8116), .B1(n8118), .B2(n9864), .ZN(n6722)
         );
  OAI211_X1 U8415 ( .C1(n9953), .C2(n9565), .A(n6723), .B(n6722), .ZN(n9956)
         );
  NAND2_X1 U8416 ( .A1(n9956), .A2(n8436), .ZN(n6731) );
  OAI22_X1 U8417 ( .A1(n9591), .A2(n6725), .B1(n6724), .B2(n9871), .ZN(n6729)
         );
  NAND2_X1 U8418 ( .A1(n6726), .A2(n6825), .ZN(n6727) );
  NAND2_X1 U8419 ( .A1(n6835), .A2(n6727), .ZN(n9955) );
  NOR2_X1 U8420 ( .A1(n9955), .A2(n9873), .ZN(n6728) );
  AOI211_X1 U8421 ( .C1(n8440), .C2(n6825), .A(n6729), .B(n6728), .ZN(n6730)
         );
  OAI211_X1 U8422 ( .C1(n9953), .C2(n9584), .A(n6731), .B(n6730), .ZN(P2_U3286) );
  INV_X1 U8423 ( .A(n7517), .ZN(n6941) );
  OAI222_X1 U8424 ( .A1(P1_U3084), .A2(n6733), .B1(n9463), .B2(n6941), .C1(
        n6732), .C2(n7885), .ZN(P1_U3333) );
  INV_X1 U8425 ( .A(n9761), .ZN(n6734) );
  NAND2_X1 U8426 ( .A1(n6895), .A2(n9813), .ZN(n6735) );
  NAND2_X1 U8427 ( .A1(n6736), .A2(n6735), .ZN(n6890) );
  NAND2_X1 U8428 ( .A1(n7473), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n6738) );
  NAND2_X1 U8429 ( .A1(n7502), .A2(n9027), .ZN(n6737) );
  NAND2_X1 U8430 ( .A1(n7040), .A2(n6896), .ZN(n8801) );
  INV_X1 U8431 ( .A(n7040), .ZN(n9019) );
  INV_X1 U8432 ( .A(n6896), .ZN(n6912) );
  NAND2_X1 U8433 ( .A1(n9019), .A2(n6912), .ZN(n8800) );
  NAND2_X1 U8434 ( .A1(n6890), .A2(n8939), .ZN(n6889) );
  NAND2_X1 U8435 ( .A1(n7040), .A2(n6912), .ZN(n6740) );
  NAND2_X1 U8436 ( .A1(n7624), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6748) );
  INV_X1 U8437 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6741) );
  OR2_X1 U8438 ( .A1(n7628), .A2(n6741), .ZN(n6747) );
  INV_X1 U8439 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6768) );
  OR2_X1 U8440 ( .A1(n7549), .A2(n6768), .ZN(n6746) );
  INV_X1 U8441 ( .A(n6743), .ZN(n6742) );
  INV_X1 U8442 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7039) );
  NAND2_X1 U8443 ( .A1(n6743), .A2(n7039), .ZN(n6744) );
  NAND2_X1 U8444 ( .A1(n6757), .A2(n6744), .ZN(n7043) );
  OR2_X1 U8445 ( .A1(n7623), .A2(n7043), .ZN(n6745) );
  NAND2_X1 U8446 ( .A1(n6750), .A2(n4475), .ZN(n6752) );
  NAND2_X1 U8447 ( .A1(n7473), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n6751) );
  OAI211_X1 U8448 ( .C1(n6754), .C2(n6753), .A(n6752), .B(n6751), .ZN(n6984)
         );
  NAND2_X1 U8449 ( .A1(n7104), .A2(n6984), .ZN(n8981) );
  INV_X1 U8450 ( .A(n6984), .ZN(n9820) );
  NAND2_X1 U8451 ( .A1(n9018), .A2(n9820), .ZN(n8810) );
  NAND2_X1 U8452 ( .A1(n8981), .A2(n8810), .ZN(n8943) );
  OAI21_X1 U8453 ( .B1(n6755), .B2(n8943), .A(n6986), .ZN(n9819) );
  NAND2_X1 U8454 ( .A1(n6757), .A2(n6756), .ZN(n6758) );
  NAND2_X1 U8455 ( .A1(n6987), .A2(n6758), .ZN(n7107) );
  OR2_X1 U8456 ( .A1(n7623), .A2(n7107), .ZN(n6763) );
  NAND2_X1 U8457 ( .A1(n8721), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6762) );
  INV_X1 U8458 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6998) );
  OR2_X1 U8459 ( .A1(n7549), .A2(n6998), .ZN(n6761) );
  INV_X1 U8460 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6759) );
  OR2_X1 U8461 ( .A1(n6273), .A2(n6759), .ZN(n6760) );
  NAND4_X1 U8462 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n9506)
         );
  INV_X1 U8463 ( .A(n9506), .ZN(n7303) );
  AND3_X1 U8464 ( .A1(n8973), .A2(n8967), .A3(n6764), .ZN(n8972) );
  NAND2_X1 U8465 ( .A1(n8799), .A2(n8968), .ZN(n6765) );
  NAND2_X1 U8466 ( .A1(n8973), .A2(n6765), .ZN(n8753) );
  XNOR2_X1 U8467 ( .A(n8804), .B(n8943), .ZN(n6767) );
  OAI222_X1 U8468 ( .A1(n9771), .A2(n7303), .B1(n9773), .B2(n7040), .C1(n6767), 
        .C2(n9509), .ZN(n9822) );
  OAI21_X1 U8469 ( .B1(n9820), .B2(n4492), .A(n4694), .ZN(n9821) );
  OAI22_X1 U8470 ( .A1(n9786), .A2(n6768), .B1(n7043), .B2(n9790), .ZN(n6769)
         );
  AOI21_X1 U8471 ( .B1(n9516), .B2(n6984), .A(n6769), .ZN(n6770) );
  OAI21_X1 U8472 ( .B1(n9821), .B2(n9139), .A(n6770), .ZN(n6771) );
  AOI21_X1 U8473 ( .B1(n9822), .B2(n9786), .A(n6771), .ZN(n6772) );
  OAI21_X1 U8474 ( .B1(n9335), .B2(n9819), .A(n6772), .ZN(P1_U3283) );
  OAI22_X1 U8475 ( .A1(n9772), .A2(n4868), .B1(n9755), .B2(n8003), .ZN(n6860)
         );
  INV_X1 U8476 ( .A(n6860), .ZN(n6781) );
  INV_X1 U8477 ( .A(n6773), .ZN(n6774) );
  NAND2_X1 U8478 ( .A1(n6775), .A2(n6774), .ZN(n6776) );
  INV_X1 U8479 ( .A(n6865), .ZN(n6779) );
  OAI22_X1 U8480 ( .A1(n9772), .A2(n8003), .B1(n9755), .B2(n7985), .ZN(n6778)
         );
  XNOR2_X1 U8481 ( .A(n6778), .B(n8001), .ZN(n6861) );
  NOR2_X1 U8482 ( .A1(n6779), .A2(n6861), .ZN(n6876) );
  AOI21_X1 U8483 ( .B1(n6779), .B2(n6861), .A(n6876), .ZN(n6780) );
  NAND2_X1 U8484 ( .A1(n6780), .A2(n6781), .ZN(n6879) );
  OAI21_X1 U8485 ( .B1(n6781), .B2(n6780), .A(n6879), .ZN(n6785) );
  AOI22_X1 U8486 ( .A1(n7390), .A2(n9022), .B1(n8717), .B2(n6798), .ZN(n6783)
         );
  AND2_X1 U8487 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9662) );
  AOI21_X1 U8488 ( .B1(n8713), .B2(n9020), .A(n9662), .ZN(n6782) );
  OAI211_X1 U8489 ( .C1(n8715), .C2(n9754), .A(n6783), .B(n6782), .ZN(n6784)
         );
  AOI21_X1 U8490 ( .B1(n6785), .B2(n8645), .A(n6784), .ZN(n6786) );
  INV_X1 U8491 ( .A(n6786), .ZN(P1_U3225) );
  AND2_X1 U8492 ( .A1(n6789), .A2(n6788), .ZN(n6791) );
  OAI21_X1 U8493 ( .B1(n6791), .B2(n6659), .A(n6790), .ZN(n9760) );
  OAI21_X1 U8494 ( .B1(n8936), .B2(n6793), .A(n6792), .ZN(n6794) );
  AOI222_X1 U8495 ( .A1(n9776), .A2(n6794), .B1(n9020), .B2(n9504), .C1(n9022), 
        .C2(n9507), .ZN(n9759) );
  NAND2_X1 U8496 ( .A1(n9781), .A2(n6798), .ZN(n6795) );
  NAND2_X1 U8497 ( .A1(n6795), .A2(n9782), .ZN(n6796) );
  NOR2_X1 U8498 ( .A1(n6797), .A2(n6796), .ZN(n9757) );
  AOI21_X1 U8499 ( .B1(n9524), .B2(n6798), .A(n9757), .ZN(n6799) );
  OAI211_X1 U8500 ( .C1(n9434), .C2(n9760), .A(n9759), .B(n6799), .ZN(n6801)
         );
  NAND2_X1 U8501 ( .A1(n6801), .A2(n9848), .ZN(n6800) );
  OAI21_X1 U8502 ( .B1(n9848), .B2(n6477), .A(n6800), .ZN(P1_U3528) );
  INV_X1 U8503 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U8504 ( .A1(n6801), .A2(n4474), .ZN(n6802) );
  OAI21_X1 U8505 ( .B1(n4474), .B2(n6803), .A(n6802), .ZN(P1_U3469) );
  INV_X1 U8506 ( .A(n7472), .ZN(n6851) );
  OAI222_X1 U8507 ( .A1(P1_U3084), .A2(n8992), .B1(n9463), .B2(n6851), .C1(
        n6804), .C2(n7885), .ZN(P1_U3332) );
  INV_X1 U8508 ( .A(n6805), .ZN(n6806) );
  AOI21_X1 U8509 ( .B1(n6809), .B2(n6807), .A(n6806), .ZN(n9801) );
  OAI21_X1 U8510 ( .B1(n6810), .B2(n6809), .A(n6808), .ZN(n6812) );
  OAI22_X1 U8511 ( .A1(n9774), .A2(n9771), .B1(n6262), .B2(n9773), .ZN(n6811)
         );
  AOI21_X1 U8512 ( .B1(n6812), .B2(n9776), .A(n6811), .ZN(n6813) );
  OAI21_X1 U8513 ( .B1(n9801), .B2(n9779), .A(n6813), .ZN(n9804) );
  INV_X1 U8514 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6815) );
  OAI22_X1 U8515 ( .A1(n9790), .A2(n6815), .B1(n6814), .B2(n9786), .ZN(n6823)
         );
  INV_X1 U8516 ( .A(n6816), .ZN(n6818) );
  OAI21_X1 U8517 ( .B1(n9802), .B2(n6818), .A(n6817), .ZN(n9803) );
  INV_X1 U8518 ( .A(n9803), .ZN(n6820) );
  AOI22_X1 U8519 ( .A1(n6820), .A2(n9333), .B1(n9516), .B2(n6819), .ZN(n6821)
         );
  OAI21_X1 U8520 ( .B1(n9801), .B2(n7005), .A(n6821), .ZN(n6822) );
  AOI211_X1 U8521 ( .C1(n9786), .C2(n9804), .A(n6823), .B(n6822), .ZN(n6824)
         );
  INV_X1 U8522 ( .A(n6824), .ZN(P1_U3289) );
  NAND2_X1 U8523 ( .A1(n6825), .A2(n8117), .ZN(n6826) );
  NAND2_X1 U8524 ( .A1(n6827), .A2(n6826), .ZN(n6829) );
  NAND2_X1 U8525 ( .A1(n9961), .A2(n6828), .ZN(n7751) );
  OAI21_X1 U8526 ( .B1(n6829), .B2(n5030), .A(n6948), .ZN(n9967) );
  OAI211_X1 U8527 ( .C1(n6832), .C2(n6831), .A(n6943), .B(n9868), .ZN(n6834)
         );
  INV_X1 U8528 ( .A(n7115), .ZN(n8115) );
  AOI22_X1 U8529 ( .A1(n9865), .A2(n8115), .B1(n8117), .B2(n9864), .ZN(n6833)
         );
  NAND2_X1 U8530 ( .A1(n6834), .A2(n6833), .ZN(n9969) );
  NAND2_X1 U8531 ( .A1(n9969), .A2(n8436), .ZN(n6842) );
  AOI21_X1 U8532 ( .B1(n9961), .B2(n6835), .A(n6951), .ZN(n9964) );
  INV_X1 U8533 ( .A(n9961), .ZN(n6836) );
  NOR2_X1 U8534 ( .A1(n6836), .A2(n9881), .ZN(n6840) );
  OAI22_X1 U8535 ( .A1(n9591), .A2(n6838), .B1(n6837), .B2(n9871), .ZN(n6839)
         );
  AOI211_X1 U8536 ( .C1(n9964), .C2(n8456), .A(n6840), .B(n6839), .ZN(n6841)
         );
  OAI211_X1 U8537 ( .C1(n8458), .C2(n9967), .A(n6842), .B(n6841), .ZN(P2_U3285) );
  NAND2_X1 U8538 ( .A1(n6844), .A2(n6843), .ZN(n6846) );
  XOR2_X1 U8539 ( .A(n6846), .B(n6845), .Z(n6850) );
  INV_X1 U8540 ( .A(n7114), .ZN(n8114) );
  AOI22_X1 U8541 ( .A1(n8106), .A2(n8116), .B1(n8084), .B2(n8114), .ZN(n6847)
         );
  NAND2_X1 U8542 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8205) );
  OAI211_X1 U8543 ( .C1(n6952), .C2(n8094), .A(n6847), .B(n8205), .ZN(n6848)
         );
  AOI21_X1 U8544 ( .B1(n7111), .B2(n8098), .A(n6848), .ZN(n6849) );
  OAI21_X1 U8545 ( .B1(n6850), .B2(n8082), .A(n6849), .ZN(P2_U3226) );
  OAI222_X1 U8546 ( .A1(n8546), .A2(n6852), .B1(P2_U3152), .B2(n7669), .C1(
        n8548), .C2(n6851), .ZN(P2_U3337) );
  OAI22_X1 U8547 ( .A1(n7040), .A2(n8003), .B1(n6912), .B2(n7985), .ZN(n6853)
         );
  XNOR2_X1 U8548 ( .A(n6853), .B(n7996), .ZN(n7027) );
  OAI22_X1 U8549 ( .A1(n7040), .A2(n4868), .B1(n6912), .B2(n8003), .ZN(n7025)
         );
  XNOR2_X1 U8550 ( .A(n7027), .B(n7025), .ZN(n6868) );
  NOR2_X1 U8551 ( .A1(n6861), .A2(n6860), .ZN(n6864) );
  OAI22_X1 U8552 ( .A1(n6895), .A2(n8003), .B1(n9813), .B2(n7985), .ZN(n6854)
         );
  XNOR2_X1 U8553 ( .A(n6854), .B(n7996), .ZN(n6856) );
  OAI22_X1 U8554 ( .A1(n6895), .A2(n4868), .B1(n9813), .B2(n8003), .ZN(n6857)
         );
  INV_X1 U8555 ( .A(n6857), .ZN(n6855) );
  NAND2_X1 U8556 ( .A1(n6856), .A2(n6855), .ZN(n6866) );
  INV_X1 U8557 ( .A(n6856), .ZN(n6858) );
  NAND2_X1 U8558 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  NAND2_X1 U8559 ( .A1(n6866), .A2(n6859), .ZN(n6878) );
  AND2_X1 U8560 ( .A1(n6861), .A2(n6860), .ZN(n6862) );
  NOR2_X1 U8561 ( .A1(n6878), .A2(n6862), .ZN(n6863) );
  OAI21_X2 U8562 ( .B1(n6865), .B2(n6864), .A(n6863), .ZN(n6880) );
  NAND2_X1 U8563 ( .A1(n6880), .A2(n6866), .ZN(n6867) );
  OAI21_X1 U8564 ( .B1(n6868), .B2(n6867), .A(n7029), .ZN(n6874) );
  NAND2_X1 U8565 ( .A1(n8713), .A2(n9018), .ZN(n6870) );
  AND2_X1 U8566 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9031) );
  INV_X1 U8567 ( .A(n9031), .ZN(n6869) );
  OAI211_X1 U8568 ( .C1(n8710), .C2(n6895), .A(n6870), .B(n6869), .ZN(n6873)
         );
  NAND2_X1 U8569 ( .A1(n8717), .A2(n6896), .ZN(n6871) );
  OAI21_X1 U8570 ( .B1(n8715), .B2(n6913), .A(n6871), .ZN(n6872) );
  AOI211_X1 U8571 ( .C1(n6874), .C2(n8645), .A(n6873), .B(n6872), .ZN(n6875)
         );
  INV_X1 U8572 ( .A(n6875), .ZN(P1_U3211) );
  INV_X1 U8573 ( .A(n6876), .ZN(n6877) );
  NAND3_X1 U8574 ( .A1(n6879), .A2(n6878), .A3(n6877), .ZN(n6881) );
  AOI21_X1 U8575 ( .B1(n6881), .B2(n6880), .A(n8719), .ZN(n6888) );
  AOI22_X1 U8576 ( .A1(n7390), .A2(n9021), .B1(n8717), .B2(n6882), .ZN(n6885)
         );
  NOR2_X1 U8577 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6883), .ZN(n9677) );
  AOI21_X1 U8578 ( .B1(n8713), .B2(n9019), .A(n9677), .ZN(n6884) );
  OAI211_X1 U8579 ( .C1(n8715), .C2(n6886), .A(n6885), .B(n6884), .ZN(n6887)
         );
  OR2_X1 U8580 ( .A1(n6888), .A2(n6887), .ZN(P1_U3237) );
  INV_X1 U8581 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6899) );
  OAI21_X1 U8582 ( .B1(n6890), .B2(n8939), .A(n6889), .ZN(n6891) );
  INV_X1 U8583 ( .A(n6891), .ZN(n6920) );
  AOI211_X1 U8584 ( .C1(n6896), .C2(n6892), .A(n9830), .B(n4492), .ZN(n6917)
         );
  XOR2_X1 U8585 ( .A(n8939), .B(n6893), .Z(n6894) );
  OAI222_X1 U8586 ( .A1(n9773), .A2(n6895), .B1(n9771), .B2(n7104), .C1(n9509), 
        .C2(n6894), .ZN(n6911) );
  AOI211_X1 U8587 ( .C1(n9524), .C2(n6896), .A(n6917), .B(n6911), .ZN(n6897)
         );
  OAI21_X1 U8588 ( .B1(n9434), .B2(n6920), .A(n6897), .ZN(n6900) );
  NAND2_X1 U8589 ( .A1(n6900), .A2(n4474), .ZN(n6898) );
  OAI21_X1 U8590 ( .B1(n4474), .B2(n6899), .A(n6898), .ZN(P1_U3475) );
  NAND2_X1 U8591 ( .A1(n6900), .A2(n9848), .ZN(n6901) );
  OAI21_X1 U8592 ( .B1(n9848), .B2(n6660), .A(n6901), .ZN(P1_U3530) );
  OAI22_X1 U8593 ( .A1(n9786), .A2(n6902), .B1(n9790), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n6905) );
  NOR2_X1 U8594 ( .A1(n9321), .A2(n6903), .ZN(n6904) );
  AOI211_X1 U8595 ( .C1(n6906), .C2(n9333), .A(n6905), .B(n6904), .ZN(n6909)
         );
  INV_X1 U8596 ( .A(n7005), .ZN(n9768) );
  NAND2_X1 U8597 ( .A1(n6907), .A2(n9768), .ZN(n6908) );
  OAI211_X1 U8598 ( .C1(n6910), .C2(n9767), .A(n6909), .B(n6908), .ZN(P1_U3288) );
  NAND2_X1 U8599 ( .A1(n6911), .A2(n9786), .ZN(n6919) );
  NOR2_X1 U8600 ( .A1(n9321), .A2(n6912), .ZN(n6916) );
  OAI22_X1 U8601 ( .A1(n9786), .A2(n6914), .B1(n6913), .B2(n9790), .ZN(n6915)
         );
  AOI211_X1 U8602 ( .C1(n6917), .C2(n9521), .A(n6916), .B(n6915), .ZN(n6918)
         );
  OAI211_X1 U8603 ( .C1(n6920), .C2(n9335), .A(n6919), .B(n6918), .ZN(P1_U3284) );
  NOR2_X1 U8604 ( .A1(n6925), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6922) );
  NOR2_X1 U8605 ( .A1(n6922), .A2(n6921), .ZN(n6966) );
  XNOR2_X1 U8606 ( .A(n6966), .B(n6967), .ZN(n6923) );
  NOR2_X1 U8607 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n6923), .ZN(n6968) );
  AOI21_X1 U8608 ( .B1(n6923), .B2(P2_REG2_REG_15__SCAN_IN), .A(n6968), .ZN(
        n6933) );
  OAI21_X1 U8609 ( .B1(n6925), .B2(P2_REG1_REG_14__SCAN_IN), .A(n6924), .ZN(
        n6958) );
  XNOR2_X1 U8610 ( .A(n6958), .B(n6959), .ZN(n6926) );
  NOR2_X1 U8611 ( .A1(n5462), .A2(n6926), .ZN(n6960) );
  AOI211_X1 U8612 ( .C1(n6926), .C2(n5462), .A(n6960), .B(n9854), .ZN(n6931)
         );
  NOR2_X1 U8613 ( .A1(n9852), .A2(n6959), .ZN(n6930) );
  NAND2_X1 U8614 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n7294) );
  INV_X1 U8615 ( .A(n7294), .ZN(n6929) );
  INV_X1 U8616 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6927) );
  NOR2_X1 U8617 ( .A1(n9488), .A2(n6927), .ZN(n6928) );
  NOR4_X1 U8618 ( .A1(n6931), .A2(n6930), .A3(n6929), .A4(n6928), .ZN(n6932)
         );
  OAI21_X1 U8619 ( .B1(n6933), .B2(n8227), .A(n6932), .ZN(P2_U3260) );
  XNOR2_X1 U8620 ( .A(n6934), .B(n6935), .ZN(n6940) );
  INV_X1 U8621 ( .A(n7163), .ZN(n8113) );
  AOI22_X1 U8622 ( .A1(n8106), .A2(n8115), .B1(n8084), .B2(n8113), .ZN(n6937)
         );
  OAI211_X1 U8623 ( .C1(n8094), .C2(n7123), .A(n6937), .B(n6936), .ZN(n6938)
         );
  AOI21_X1 U8624 ( .B1(n9615), .B2(n8098), .A(n6938), .ZN(n6939) );
  OAI21_X1 U8625 ( .B1(n6940), .B2(n8082), .A(n6939), .ZN(P2_U3236) );
  OAI222_X1 U8626 ( .A1(n8546), .A2(n6942), .B1(P2_U3152), .B2(n7840), .C1(
        n8548), .C2(n6941), .ZN(P2_U3338) );
  NAND2_X1 U8627 ( .A1(n7111), .A2(n7115), .ZN(n7757) );
  INV_X1 U8628 ( .A(n6949), .ZN(n7853) );
  NAND3_X1 U8629 ( .A1(n6943), .A2(n7756), .A3(n7853), .ZN(n6944) );
  NAND3_X1 U8630 ( .A1(n7117), .A2(n9868), .A3(n6944), .ZN(n6946) );
  AOI22_X1 U8631 ( .A1(n9864), .A2(n8116), .B1(n8114), .B2(n9865), .ZN(n6945)
         );
  NAND2_X1 U8632 ( .A1(n6946), .A2(n6945), .ZN(n9975) );
  INV_X1 U8633 ( .A(n9975), .ZN(n6957) );
  NAND2_X1 U8634 ( .A1(n9961), .A2(n8116), .ZN(n6947) );
  OAI21_X1 U8635 ( .B1(n4557), .B2(n7853), .A(n7113), .ZN(n9977) );
  INV_X1 U8636 ( .A(n8458), .ZN(n9878) );
  INV_X1 U8637 ( .A(n7111), .ZN(n9972) );
  INV_X1 U8638 ( .A(n7121), .ZN(n6950) );
  OAI21_X1 U8639 ( .B1(n9972), .B2(n6951), .A(n6950), .ZN(n9974) );
  OAI22_X1 U8640 ( .A1(n9591), .A2(n8201), .B1(n6952), .B2(n9871), .ZN(n6953)
         );
  AOI21_X1 U8641 ( .B1(n7111), .B2(n8440), .A(n6953), .ZN(n6954) );
  OAI21_X1 U8642 ( .B1(n9974), .B2(n9873), .A(n6954), .ZN(n6955) );
  AOI21_X1 U8643 ( .B1(n9977), .B2(n9878), .A(n6955), .ZN(n6956) );
  OAI21_X1 U8644 ( .B1(n6957), .B2(n9884), .A(n6956), .ZN(P2_U3284) );
  NOR2_X1 U8645 ( .A1(n6959), .A2(n6958), .ZN(n6961) );
  NOR2_X1 U8646 ( .A1(n6961), .A2(n6960), .ZN(n6965) );
  NOR2_X1 U8647 ( .A1(n6976), .A2(n6962), .ZN(n6963) );
  AOI21_X1 U8648 ( .B1(n6962), .B2(n6976), .A(n6963), .ZN(n6964) );
  NAND2_X1 U8649 ( .A1(n6964), .A2(n6965), .ZN(n7189) );
  OAI21_X1 U8650 ( .B1(n6965), .B2(n6964), .A(n7189), .ZN(n6978) );
  NOR2_X1 U8651 ( .A1(n6967), .A2(n6966), .ZN(n6969) );
  NOR2_X1 U8652 ( .A1(n6969), .A2(n6968), .ZN(n6972) );
  NAND2_X1 U8653 ( .A1(n7190), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7181) );
  INV_X1 U8654 ( .A(n7181), .ZN(n6970) );
  AOI21_X1 U8655 ( .B1(n7449), .B2(n6976), .A(n6970), .ZN(n6971) );
  NAND2_X1 U8656 ( .A1(n6971), .A2(n6972), .ZN(n7180) );
  OAI211_X1 U8657 ( .C1(n6972), .C2(n6971), .A(n9850), .B(n7180), .ZN(n6975)
         );
  NOR2_X1 U8658 ( .A1(n6973), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7332) );
  AOI21_X1 U8659 ( .B1(n9857), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7332), .ZN(
        n6974) );
  OAI211_X1 U8660 ( .C1(n9852), .C2(n6976), .A(n6975), .B(n6974), .ZN(n6977)
         );
  AOI21_X1 U8661 ( .B1(n9849), .B2(n6978), .A(n6977), .ZN(n6979) );
  INV_X1 U8662 ( .A(n6979), .ZN(P2_U3261) );
  NAND2_X1 U8663 ( .A1(n6980), .A2(n4475), .ZN(n6982) );
  AOI22_X1 U8664 ( .A1(n8730), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9707), .B2(
        n7502), .ZN(n6981) );
  NAND2_X1 U8665 ( .A1(n6982), .A2(n6981), .ZN(n7096) );
  NOR2_X1 U8666 ( .A1(n9829), .A2(n9506), .ZN(n8812) );
  NAND2_X1 U8667 ( .A1(n9829), .A2(n9506), .ZN(n9500) );
  INV_X1 U8668 ( .A(n9500), .ZN(n6983) );
  NOR2_X1 U8669 ( .A1(n8812), .A2(n6983), .ZN(n8945) );
  NAND2_X1 U8670 ( .A1(n9018), .A2(n6984), .ZN(n6985) );
  XOR2_X1 U8671 ( .A(n8945), .B(n7047), .Z(n9827) );
  XNOR2_X1 U8672 ( .A(n7079), .B(n8945), .ZN(n6996) );
  NAND2_X1 U8673 ( .A1(n6987), .A2(n7302), .ZN(n6988) );
  NAND2_X1 U8674 ( .A1(n7058), .A2(n6988), .ZN(n9513) );
  OR2_X1 U8675 ( .A1(n7623), .A2(n9513), .ZN(n6994) );
  NAND2_X1 U8676 ( .A1(n8721), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6993) );
  INV_X1 U8677 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6989) );
  OR2_X1 U8678 ( .A1(n6273), .A2(n6989), .ZN(n6992) );
  INV_X1 U8679 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6990) );
  OR2_X1 U8680 ( .A1(n7549), .A2(n6990), .ZN(n6991) );
  NAND4_X1 U8681 ( .A1(n6994), .A2(n6993), .A3(n6992), .A4(n6991), .ZN(n9017)
         );
  OAI22_X1 U8682 ( .A1(n8675), .A2(n9771), .B1(n7104), .B2(n9773), .ZN(n6995)
         );
  AOI21_X1 U8683 ( .B1(n6996), .B2(n9776), .A(n6995), .ZN(n6997) );
  OAI21_X1 U8684 ( .B1(n9827), .B2(n9779), .A(n6997), .ZN(n9832) );
  NAND2_X1 U8685 ( .A1(n9832), .A2(n9786), .ZN(n7004) );
  OAI22_X1 U8687 ( .A1(n9786), .A2(n6998), .B1(n7107), .B2(n9790), .ZN(n7002)
         );
  NOR2_X1 U8688 ( .A1(n6999), .A2(n9829), .ZN(n7000) );
  OR2_X1 U8689 ( .A1(n9519), .A2(n7000), .ZN(n9831) );
  NOR2_X1 U8690 ( .A1(n9831), .A2(n9139), .ZN(n7001) );
  AOI211_X1 U8691 ( .C1(n9516), .C2(n7096), .A(n7002), .B(n7001), .ZN(n7003)
         );
  OAI211_X1 U8692 ( .C1(n9827), .C2(n7005), .A(n7004), .B(n7003), .ZN(P1_U3282) );
  INV_X1 U8693 ( .A(n7539), .ZN(n7008) );
  NOR2_X1 U8694 ( .A1(n7006), .A2(P1_U3084), .ZN(n9004) );
  AOI21_X1 U8695 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9465), .A(n9004), .ZN(
        n7007) );
  OAI21_X1 U8696 ( .B1(n7008), .B2(n9463), .A(n7007), .ZN(P1_U3330) );
  INV_X1 U8697 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7019) );
  AOI211_X1 U8698 ( .C1(n7010), .C2(n7245), .A(n7009), .B(n9713), .ZN(n7011)
         );
  AOI21_X1 U8699 ( .B1(n9742), .B2(n7240), .A(n7011), .ZN(n7018) );
  OAI21_X1 U8700 ( .B1(n7014), .B2(n7013), .A(n7012), .ZN(n7016) );
  NAND2_X1 U8701 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8563) );
  INV_X1 U8702 ( .A(n8563), .ZN(n7015) );
  AOI21_X1 U8703 ( .B1(n9750), .B2(n7016), .A(n7015), .ZN(n7017) );
  OAI211_X1 U8704 ( .C1(n9735), .C2(n7019), .A(n7018), .B(n7017), .ZN(P1_U3255) );
  INV_X1 U8705 ( .A(n7528), .ZN(n7021) );
  OAI222_X1 U8706 ( .A1(n8546), .A2(n10101), .B1(n8548), .B2(n7021), .C1(n5774), .C2(P2_U3152), .ZN(P2_U3336) );
  OAI222_X1 U8707 ( .A1(n9003), .A2(P1_U3084), .B1(n9463), .B2(n7021), .C1(
        n7020), .C2(n7885), .ZN(P1_U3331) );
  NAND2_X1 U8708 ( .A1(n7539), .A2(n7022), .ZN(n7023) );
  OAI211_X1 U8709 ( .C1(n7024), .C2(n8546), .A(n7023), .B(n7882), .ZN(P2_U3335) );
  INV_X1 U8710 ( .A(n7025), .ZN(n7026) );
  NAND2_X1 U8711 ( .A1(n7027), .A2(n7026), .ZN(n7028) );
  OAI22_X1 U8712 ( .A1(n7104), .A2(n4868), .B1(n9820), .B2(n8003), .ZN(n7030)
         );
  INV_X1 U8713 ( .A(n7030), .ZN(n7032) );
  OAI22_X1 U8714 ( .A1(n7104), .A2(n8003), .B1(n9820), .B2(n7985), .ZN(n7031)
         );
  XNOR2_X1 U8715 ( .A(n7031), .B(n7996), .ZN(n7035) );
  NAND2_X1 U8716 ( .A1(n7033), .A2(n7032), .ZN(n7099) );
  INV_X1 U8717 ( .A(n7099), .ZN(n7034) );
  NOR2_X1 U8718 ( .A1(n7100), .A2(n7034), .ZN(n7038) );
  AOI21_X1 U8719 ( .B1(n7036), .B2(n7099), .A(n7035), .ZN(n7037) );
  OAI21_X1 U8720 ( .B1(n7038), .B2(n7037), .A(n8645), .ZN(n7046) );
  NOR2_X1 U8721 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7039), .ZN(n9683) );
  AOI21_X1 U8722 ( .B1(n8713), .B2(n9506), .A(n9683), .ZN(n7042) );
  OR2_X1 U8723 ( .A1(n8710), .A2(n7040), .ZN(n7041) );
  OAI211_X1 U8724 ( .C1(n8715), .C2(n7043), .A(n7042), .B(n7041), .ZN(n7044)
         );
  INV_X1 U8725 ( .A(n7044), .ZN(n7045) );
  OAI211_X1 U8726 ( .C1(n9820), .C2(n8654), .A(n7046), .B(n7045), .ZN(P1_U3219) );
  NAND2_X1 U8727 ( .A1(n7048), .A2(n4475), .ZN(n7050) );
  AOI22_X1 U8728 ( .A1(n8730), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9720), .B2(
        n7502), .ZN(n7049) );
  NAND2_X1 U8729 ( .A1(n9526), .A2(n9017), .ZN(n8738) );
  INV_X1 U8730 ( .A(n9526), .ZN(n9517) );
  NAND2_X1 U8731 ( .A1(n9517), .A2(n8675), .ZN(n8815) );
  NAND2_X1 U8732 ( .A1(n8738), .A2(n8815), .ZN(n9503) );
  NAND2_X1 U8733 ( .A1(n9499), .A2(n9503), .ZN(n7052) );
  NAND2_X1 U8734 ( .A1(n9526), .A2(n8675), .ZN(n7051) );
  NAND2_X1 U8735 ( .A1(n7052), .A2(n7051), .ZN(n7130) );
  NAND2_X1 U8736 ( .A1(n7053), .A2(n4475), .ZN(n7055) );
  AOI22_X1 U8737 ( .A1(n8730), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9724), .B2(
        n7502), .ZN(n7054) );
  INV_X1 U8738 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7057) );
  NAND2_X1 U8739 ( .A1(n7058), .A2(n7057), .ZN(n7059) );
  NAND2_X1 U8740 ( .A1(n7072), .A2(n7059), .ZN(n8678) );
  OR2_X1 U8741 ( .A1(n7623), .A2(n8678), .ZN(n7064) );
  NAND2_X1 U8742 ( .A1(n8721), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7063) );
  INV_X1 U8743 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7060) );
  OR2_X1 U8744 ( .A1(n6273), .A2(n7060), .ZN(n7062) );
  OR2_X1 U8745 ( .A1(n7549), .A2(n5910), .ZN(n7061) );
  NAND4_X1 U8746 ( .A1(n7064), .A2(n7063), .A3(n7062), .A4(n7061), .ZN(n9505)
         );
  INV_X1 U8747 ( .A(n9505), .ZN(n8599) );
  XNOR2_X1 U8748 ( .A(n9431), .B(n8599), .ZN(n8948) );
  INV_X1 U8749 ( .A(n8948), .ZN(n8821) );
  XNOR2_X1 U8750 ( .A(n7130), .B(n8821), .ZN(n9433) );
  NAND2_X1 U8751 ( .A1(n9519), .A2(n9526), .ZN(n9518) );
  INV_X1 U8752 ( .A(n7151), .ZN(n7065) );
  AOI211_X1 U8753 ( .C1(n9431), .C2(n9518), .A(n9830), .B(n7065), .ZN(n9430)
         );
  INV_X1 U8754 ( .A(n9431), .ZN(n7066) );
  NOR2_X1 U8755 ( .A1(n7066), .A2(n9321), .ZN(n7068) );
  OAI22_X1 U8756 ( .A1(n9786), .A2(n5910), .B1(n8678), .B2(n9790), .ZN(n7067)
         );
  AOI211_X1 U8757 ( .C1(n9430), .C2(n9521), .A(n7068), .B(n7067), .ZN(n7082)
         );
  NAND2_X1 U8758 ( .A1(n7069), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7078) );
  OR2_X1 U8759 ( .A1(n7628), .A2(n7070), .ZN(n7077) );
  INV_X1 U8760 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U8761 ( .A1(n7072), .A2(n8598), .ZN(n7073) );
  NAND2_X1 U8762 ( .A1(n7141), .A2(n7073), .ZN(n8602) );
  OR2_X1 U8763 ( .A1(n7623), .A2(n8602), .ZN(n7076) );
  INV_X1 U8764 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7074) );
  OR2_X1 U8765 ( .A1(n6273), .A2(n7074), .ZN(n7075) );
  AND2_X1 U8766 ( .A1(n8738), .A2(n9500), .ZN(n8818) );
  XNOR2_X1 U8767 ( .A(n7137), .B(n8948), .ZN(n7080) );
  OAI222_X1 U8768 ( .A1(n9771), .A2(n7357), .B1(n9773), .B2(n8675), .C1(n9509), 
        .C2(n7080), .ZN(n9429) );
  NAND2_X1 U8769 ( .A1(n9429), .A2(n9786), .ZN(n7081) );
  OAI211_X1 U8770 ( .C1(n9433), .C2(n9335), .A(n7082), .B(n7081), .ZN(P1_U3280) );
  INV_X1 U8771 ( .A(n7083), .ZN(n7084) );
  AOI21_X1 U8772 ( .B1(n7086), .B2(n7085), .A(n7084), .ZN(n7091) );
  INV_X1 U8773 ( .A(n7443), .ZN(n8112) );
  AOI22_X1 U8774 ( .A1(n8106), .A2(n8114), .B1(n8084), .B2(n8112), .ZN(n7088)
         );
  OAI211_X1 U8775 ( .C1(n8094), .C2(n7173), .A(n7088), .B(n7087), .ZN(n7089)
         );
  AOI21_X1 U8776 ( .B1(n9609), .B2(n8098), .A(n7089), .ZN(n7090) );
  OAI21_X1 U8777 ( .B1(n7091), .B2(n8082), .A(n7090), .ZN(P2_U3217) );
  INV_X1 U8778 ( .A(n7552), .ZN(n7647) );
  OAI222_X1 U8779 ( .A1(P2_U3152), .A2(n7092), .B1(n8548), .B2(n7647), .C1(
        n10201), .C2(n8546), .ZN(P2_U3334) );
  NAND2_X1 U8780 ( .A1(n9506), .A2(n7893), .ZN(n7094) );
  NAND2_X1 U8781 ( .A1(n7096), .A2(n8005), .ZN(n7093) );
  NAND2_X1 U8782 ( .A1(n7094), .A2(n7093), .ZN(n7095) );
  XNOR2_X1 U8783 ( .A(n7095), .B(n7996), .ZN(n7308) );
  NAND2_X1 U8784 ( .A1(n9506), .A2(n7998), .ZN(n7098) );
  NAND2_X1 U8785 ( .A1(n7096), .A2(n7893), .ZN(n7097) );
  NAND2_X1 U8786 ( .A1(n7098), .A2(n7097), .ZN(n7306) );
  XNOR2_X1 U8787 ( .A(n7308), .B(n7306), .ZN(n7102) );
  OAI21_X1 U8788 ( .B1(n7102), .B2(n7101), .A(n7310), .ZN(n7103) );
  NAND2_X1 U8789 ( .A1(n7103), .A2(n8645), .ZN(n7110) );
  AND2_X1 U8790 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9705) );
  AOI21_X1 U8791 ( .B1(n8713), .B2(n9017), .A(n9705), .ZN(n7106) );
  OR2_X1 U8792 ( .A1(n8710), .A2(n7104), .ZN(n7105) );
  OAI211_X1 U8793 ( .C1(n8715), .C2(n7107), .A(n7106), .B(n7105), .ZN(n7108)
         );
  INV_X1 U8794 ( .A(n7108), .ZN(n7109) );
  OAI211_X1 U8795 ( .C1(n9829), .C2(n8654), .A(n7110), .B(n7109), .ZN(P1_U3229) );
  OR2_X1 U8796 ( .A1(n7111), .A2(n8115), .ZN(n7112) );
  OR2_X1 U8797 ( .A1(n9615), .A2(n7114), .ZN(n7758) );
  NAND2_X1 U8798 ( .A1(n9615), .A2(n7114), .ZN(n7753) );
  NAND2_X1 U8799 ( .A1(n7758), .A2(n7753), .ZN(n7854) );
  OAI21_X1 U8800 ( .B1(n4553), .B2(n7854), .A(n7168), .ZN(n9619) );
  OAI22_X1 U8801 ( .A1(n7115), .A2(n9579), .B1(n7163), .B2(n9581), .ZN(n7116)
         );
  INV_X1 U8802 ( .A(n7116), .ZN(n7120) );
  NAND2_X1 U8803 ( .A1(n7117), .A2(n7755), .ZN(n7160) );
  XNOR2_X1 U8804 ( .A(n7160), .B(n7854), .ZN(n7118) );
  NAND2_X1 U8805 ( .A1(n7118), .A2(n9868), .ZN(n7119) );
  OAI211_X1 U8806 ( .C1(n9619), .C2(n9565), .A(n7120), .B(n7119), .ZN(n9621)
         );
  NAND2_X1 U8807 ( .A1(n9621), .A2(n8436), .ZN(n7129) );
  INV_X1 U8808 ( .A(n9615), .ZN(n7125) );
  OR2_X1 U8809 ( .A1(n7121), .A2(n7125), .ZN(n7122) );
  AND2_X1 U8810 ( .A1(n7171), .A2(n7122), .ZN(n9616) );
  OAI22_X1 U8811 ( .A1(n9591), .A2(n7124), .B1(n7123), .B2(n9871), .ZN(n7127)
         );
  NOR2_X1 U8812 ( .A1(n7125), .A2(n9881), .ZN(n7126) );
  AOI211_X1 U8813 ( .C1(n9616), .C2(n8456), .A(n7127), .B(n7126), .ZN(n7128)
         );
  OAI211_X1 U8814 ( .C1(n9619), .C2(n9584), .A(n7129), .B(n7128), .ZN(P2_U3283) );
  INV_X1 U8815 ( .A(n7130), .ZN(n7131) );
  NAND2_X1 U8816 ( .A1(n7131), .A2(n5057), .ZN(n7133) );
  NAND2_X1 U8817 ( .A1(n9431), .A2(n9505), .ZN(n7132) );
  NAND2_X1 U8818 ( .A1(n7134), .A2(n4475), .ZN(n7136) );
  AOI22_X1 U8819 ( .A1(n8730), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9049), .B2(
        n7502), .ZN(n7135) );
  OR2_X1 U8820 ( .A1(n9634), .A2(n7357), .ZN(n8824) );
  NAND2_X1 U8821 ( .A1(n9634), .A2(n7357), .ZN(n8816) );
  NAND2_X1 U8822 ( .A1(n8824), .A2(n8816), .ZN(n8947) );
  INV_X1 U8823 ( .A(n8947), .ZN(n7138) );
  XNOR2_X1 U8824 ( .A(n7212), .B(n7138), .ZN(n9638) );
  OR2_X1 U8825 ( .A1(n9431), .A2(n8599), .ZN(n7217) );
  NAND2_X1 U8826 ( .A1(n7218), .A2(n7217), .ZN(n7139) );
  XNOR2_X1 U8827 ( .A(n7139), .B(n7138), .ZN(n7149) );
  INV_X1 U8828 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7140) );
  NAND2_X1 U8829 ( .A1(n7141), .A2(n7140), .ZN(n7142) );
  NAND2_X1 U8830 ( .A1(n7223), .A2(n7142), .ZN(n7387) );
  OR2_X1 U8831 ( .A1(n7623), .A2(n7387), .ZN(n7147) );
  NAND2_X1 U8832 ( .A1(n8721), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7146) );
  INV_X1 U8833 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7234) );
  OR2_X1 U8834 ( .A1(n7549), .A2(n7234), .ZN(n7145) );
  INV_X1 U8835 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7143) );
  OR2_X1 U8836 ( .A1(n6273), .A2(n7143), .ZN(n7144) );
  NAND4_X1 U8837 ( .A1(n7147), .A2(n7146), .A3(n7145), .A4(n7144), .ZN(n9015)
         );
  AOI22_X1 U8838 ( .A1(n9504), .A2(n9015), .B1(n9505), .B2(n9507), .ZN(n7148)
         );
  OAI21_X1 U8839 ( .B1(n7149), .B2(n9509), .A(n7148), .ZN(n7150) );
  AOI21_X1 U8840 ( .B1(n9638), .B2(n9512), .A(n7150), .ZN(n9640) );
  NAND2_X1 U8841 ( .A1(n7151), .A2(n9634), .ZN(n7152) );
  NAND2_X1 U8842 ( .A1(n7152), .A2(n9782), .ZN(n7153) );
  OR2_X1 U8843 ( .A1(n7232), .A2(n7153), .ZN(n9635) );
  INV_X1 U8844 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7154) );
  OAI22_X1 U8845 ( .A1(n9786), .A2(n7154), .B1(n8602), .B2(n9790), .ZN(n7155)
         );
  AOI21_X1 U8846 ( .B1(n9634), .B2(n9516), .A(n7155), .ZN(n7156) );
  OAI21_X1 U8847 ( .B1(n9635), .B2(n7157), .A(n7156), .ZN(n7158) );
  AOI21_X1 U8848 ( .B1(n9638), .B2(n9768), .A(n7158), .ZN(n7159) );
  OAI21_X1 U8849 ( .B1(n9640), .B2(n9767), .A(n7159), .ZN(P1_U3279) );
  NOR2_X1 U8850 ( .A1(n7160), .A2(n7854), .ZN(n7162) );
  NAND2_X1 U8851 ( .A1(n9609), .A2(n7163), .ZN(n7761) );
  NAND2_X1 U8852 ( .A1(n7760), .A2(n7761), .ZN(n7169) );
  INV_X1 U8853 ( .A(n7169), .ZN(n7857) );
  NAND2_X1 U8854 ( .A1(n7164), .A2(n7857), .ZN(n7263) );
  OAI211_X1 U8855 ( .C1(n7164), .C2(n7857), .A(n9868), .B(n7263), .ZN(n7166)
         );
  AOI22_X1 U8856 ( .A1(n9864), .A2(n8114), .B1(n8112), .B2(n9865), .ZN(n7165)
         );
  NAND2_X1 U8857 ( .A1(n7166), .A2(n7165), .ZN(n9611) );
  INV_X1 U8858 ( .A(n9611), .ZN(n7179) );
  NAND2_X1 U8859 ( .A1(n9615), .A2(n8114), .ZN(n7167) );
  OAI21_X1 U8860 ( .B1(n7170), .B2(n7169), .A(n7262), .ZN(n9613) );
  NAND2_X1 U8861 ( .A1(n7171), .A2(n9609), .ZN(n7172) );
  NAND2_X1 U8862 ( .A1(n7267), .A2(n7172), .ZN(n9610) );
  OAI22_X1 U8863 ( .A1(n9591), .A2(n7174), .B1(n7173), .B2(n9871), .ZN(n7175)
         );
  AOI21_X1 U8864 ( .B1(n9609), .B2(n8440), .A(n7175), .ZN(n7176) );
  OAI21_X1 U8865 ( .B1(n9610), .B2(n9873), .A(n7176), .ZN(n7177) );
  AOI21_X1 U8866 ( .B1(n9613), .B2(n9878), .A(n7177), .ZN(n7178) );
  OAI21_X1 U8867 ( .B1(n7179), .B2(n9593), .A(n7178), .ZN(P2_U3282) );
  NAND2_X1 U8868 ( .A1(n7181), .A2(n7180), .ZN(n7185) );
  OR2_X1 U8869 ( .A1(n7201), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7183) );
  NAND2_X1 U8870 ( .A1(n7201), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7182) );
  AND2_X1 U8871 ( .A1(n7183), .A2(n7182), .ZN(n7184) );
  NAND2_X1 U8872 ( .A1(n7184), .A2(n7185), .ZN(n7197) );
  OAI211_X1 U8873 ( .C1(n7185), .C2(n7184), .A(n9850), .B(n7197), .ZN(n7196)
         );
  NOR2_X1 U8874 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7278), .ZN(n7194) );
  OR2_X1 U8875 ( .A1(n7201), .A2(n7186), .ZN(n7188) );
  NAND2_X1 U8876 ( .A1(n7201), .A2(n7186), .ZN(n7187) );
  AND2_X1 U8877 ( .A1(n7188), .A2(n7187), .ZN(n7192) );
  OAI21_X1 U8878 ( .B1(n7190), .B2(P2_REG1_REG_16__SCAN_IN), .A(n7189), .ZN(
        n7191) );
  NOR2_X1 U8879 ( .A1(n7192), .A2(n7191), .ZN(n7200) );
  AOI211_X1 U8880 ( .C1(n7192), .C2(n7191), .A(n7200), .B(n9854), .ZN(n7193)
         );
  AOI211_X1 U8881 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9857), .A(n7194), .B(
        n7193), .ZN(n7195) );
  OAI211_X1 U8882 ( .C1(n9852), .C2(n7198), .A(n7196), .B(n7195), .ZN(P2_U3262) );
  INV_X1 U8883 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9590) );
  OAI21_X1 U8884 ( .B1(n9590), .B2(n7198), .A(n7197), .ZN(n8219) );
  XOR2_X1 U8885 ( .A(n7205), .B(n8219), .Z(n7199) );
  NOR2_X1 U8886 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n7199), .ZN(n8222) );
  AOI21_X1 U8887 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n7199), .A(n8222), .ZN(
        n7210) );
  AOI21_X1 U8888 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n7201), .A(n7200), .ZN(
        n7204) );
  AOI22_X1 U8889 ( .A1(n8220), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n7202), .B2(
        n7205), .ZN(n7203) );
  NAND2_X1 U8890 ( .A1(n7204), .A2(n7203), .ZN(n8216) );
  OAI21_X1 U8891 ( .B1(n7204), .B2(n7203), .A(n8216), .ZN(n7208) );
  NOR2_X1 U8892 ( .A1(n9852), .A2(n7205), .ZN(n7207) );
  INV_X1 U8893 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10404) );
  NAND2_X1 U8894 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7337) );
  OAI21_X1 U8895 ( .B1(n9488), .B2(n10404), .A(n7337), .ZN(n7206) );
  AOI211_X1 U8896 ( .C1(n7208), .C2(n9849), .A(n7207), .B(n7206), .ZN(n7209)
         );
  OAI21_X1 U8897 ( .B1(n7210), .B2(n8227), .A(n7209), .ZN(P2_U3263) );
  AND2_X1 U8898 ( .A1(n9634), .A2(n9016), .ZN(n7211) );
  NAND2_X1 U8899 ( .A1(n7213), .A2(n4475), .ZN(n7215) );
  AOI22_X1 U8900 ( .A1(n8730), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9062), .B2(
        n7502), .ZN(n7214) );
  XNOR2_X1 U8901 ( .A(n8762), .B(n9015), .ZN(n8950) );
  INV_X1 U8902 ( .A(n8950), .ZN(n7216) );
  XNOR2_X1 U8903 ( .A(n4552), .B(n7216), .ZN(n9631) );
  AND2_X1 U8904 ( .A1(n8824), .A2(n7217), .ZN(n8760) );
  NAND2_X1 U8905 ( .A1(n7219), .A2(n8816), .ZN(n7248) );
  XNOR2_X1 U8906 ( .A(n7248), .B(n8950), .ZN(n7220) );
  NAND2_X1 U8907 ( .A1(n7220), .A2(n9776), .ZN(n7230) );
  INV_X1 U8908 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7222) );
  NAND2_X1 U8909 ( .A1(n7223), .A2(n7222), .ZN(n7224) );
  NAND2_X1 U8910 ( .A1(n7251), .A2(n7224), .ZN(n8566) );
  OR2_X1 U8911 ( .A1(n7623), .A2(n8566), .ZN(n7228) );
  NAND2_X1 U8912 ( .A1(n8721), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7227) );
  INV_X1 U8913 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7245) );
  OR2_X1 U8914 ( .A1(n7549), .A2(n7245), .ZN(n7226) );
  INV_X1 U8915 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10121) );
  OR2_X1 U8916 ( .A1(n6273), .A2(n10121), .ZN(n7225) );
  NAND4_X1 U8917 ( .A1(n7228), .A2(n7227), .A3(n7226), .A4(n7225), .ZN(n9328)
         );
  AOI22_X1 U8918 ( .A1(n9016), .A2(n9507), .B1(n9504), .B2(n9328), .ZN(n7229)
         );
  NAND2_X1 U8919 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  AOI21_X1 U8920 ( .B1(n9631), .B2(n9512), .A(n7231), .ZN(n9633) );
  NOR2_X1 U8921 ( .A1(n7232), .A2(n9628), .ZN(n7233) );
  OR2_X1 U8922 ( .A1(n7243), .A2(n7233), .ZN(n9629) );
  OAI22_X1 U8923 ( .A1(n9786), .A2(n7234), .B1(n7387), .B2(n9790), .ZN(n7235)
         );
  AOI21_X1 U8924 ( .B1(n8762), .B2(n9516), .A(n7235), .ZN(n7236) );
  OAI21_X1 U8925 ( .B1(n9629), .B2(n9139), .A(n7236), .ZN(n7237) );
  AOI21_X1 U8926 ( .B1(n9631), .B2(n9768), .A(n7237), .ZN(n7238) );
  OAI21_X1 U8927 ( .B1(n9633), .B2(n9767), .A(n7238), .ZN(P1_U3278) );
  NAND2_X1 U8928 ( .A1(n7239), .A2(n4475), .ZN(n7242) );
  AOI22_X1 U8929 ( .A1(n8730), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7240), .B2(
        n7502), .ZN(n7241) );
  OR2_X1 U8930 ( .A1(n9426), .A2(n8709), .ZN(n8828) );
  NAND2_X1 U8931 ( .A1(n9426), .A2(n8709), .ZN(n8829) );
  INV_X1 U8932 ( .A(n9015), .ZN(n8761) );
  XOR2_X1 U8933 ( .A(n8952), .B(n7395), .Z(n9428) );
  INV_X1 U8934 ( .A(n7243), .ZN(n7244) );
  INV_X1 U8935 ( .A(n9426), .ZN(n7396) );
  AOI211_X1 U8936 ( .C1(n9426), .C2(n7244), .A(n9830), .B(n4702), .ZN(n9425)
         );
  NOR2_X1 U8937 ( .A1(n7396), .A2(n9321), .ZN(n7247) );
  OAI22_X1 U8938 ( .A1(n9786), .A2(n7245), .B1(n8566), .B2(n9790), .ZN(n7246)
         );
  AOI211_X1 U8939 ( .C1(n9425), .C2(n9521), .A(n7247), .B(n7246), .ZN(n7260)
         );
  AND2_X1 U8940 ( .A1(n8762), .A2(n8761), .ZN(n8743) );
  NAND2_X1 U8941 ( .A1(n7249), .A2(n8952), .ZN(n7429) );
  OAI211_X1 U8942 ( .C1(n7249), .C2(n8952), .A(n7429), .B(n9776), .ZN(n7258)
         );
  NAND2_X1 U8943 ( .A1(n7251), .A2(n7250), .ZN(n7252) );
  NAND2_X1 U8944 ( .A1(n7409), .A2(n7252), .ZN(n9318) );
  OR2_X1 U8945 ( .A1(n7623), .A2(n9318), .ZN(n7256) );
  NAND2_X1 U8946 ( .A1(n8721), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7255) );
  INV_X1 U8947 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10149) );
  OR2_X1 U8948 ( .A1(n6273), .A2(n10149), .ZN(n7254) );
  OR2_X1 U8949 ( .A1(n7549), .A2(n5954), .ZN(n7253) );
  NAND4_X1 U8950 ( .A1(n7256), .A2(n7255), .A3(n7254), .A4(n7253), .ZN(n9014)
         );
  AOI22_X1 U8951 ( .A1(n9507), .A2(n9015), .B1(n9014), .B2(n9504), .ZN(n7257)
         );
  NAND2_X1 U8952 ( .A1(n7258), .A2(n7257), .ZN(n9424) );
  NAND2_X1 U8953 ( .A1(n9424), .A2(n9786), .ZN(n7259) );
  OAI211_X1 U8954 ( .C1(n9428), .C2(n9335), .A(n7260), .B(n7259), .ZN(P1_U3277) );
  OR2_X1 U8955 ( .A1(n9609), .A2(n8113), .ZN(n7261) );
  NAND2_X1 U8956 ( .A1(n7262), .A2(n7261), .ZN(n7434) );
  NAND2_X1 U8957 ( .A1(n7435), .A2(n7443), .ZN(n7765) );
  XNOR2_X1 U8958 ( .A(n7434), .B(n7433), .ZN(n9608) );
  INV_X1 U8959 ( .A(n9608), .ZN(n7275) );
  NAND2_X1 U8960 ( .A1(n7263), .A2(n7760), .ZN(n7264) );
  NAND2_X1 U8961 ( .A1(n7264), .A2(n7856), .ZN(n7441) );
  OAI211_X1 U8962 ( .C1(n7264), .C2(n7856), .A(n7441), .B(n9868), .ZN(n7266)
         );
  AOI22_X1 U8963 ( .A1(n8113), .A2(n9864), .B1(n9865), .B2(n8245), .ZN(n7265)
         );
  NAND2_X1 U8964 ( .A1(n7266), .A2(n7265), .ZN(n9606) );
  INV_X1 U8965 ( .A(n7435), .ZN(n9604) );
  INV_X1 U8966 ( .A(n7267), .ZN(n7269) );
  INV_X1 U8967 ( .A(n8235), .ZN(n7268) );
  OAI21_X1 U8968 ( .B1(n9604), .B2(n7269), .A(n7268), .ZN(n9605) );
  OAI22_X1 U8969 ( .A1(n9591), .A2(n7270), .B1(n7296), .B2(n9871), .ZN(n7271)
         );
  AOI21_X1 U8970 ( .B1(n7435), .B2(n8440), .A(n7271), .ZN(n7272) );
  OAI21_X1 U8971 ( .B1(n9605), .B2(n9873), .A(n7272), .ZN(n7273) );
  AOI21_X1 U8972 ( .B1(n9606), .B2(n8436), .A(n7273), .ZN(n7274) );
  OAI21_X1 U8973 ( .B1(n7275), .B2(n8458), .A(n7274), .ZN(P2_U3281) );
  XNOR2_X1 U8974 ( .A(n7277), .B(n7276), .ZN(n7282) );
  OAI22_X1 U8975 ( .A1(n8094), .A2(n9585), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7278), .ZN(n7280) );
  INV_X1 U8976 ( .A(n8245), .ZN(n9578) );
  OAI22_X1 U8977 ( .A1(n9578), .A2(n8058), .B1(n8096), .B2(n9580), .ZN(n7279)
         );
  AOI211_X1 U8978 ( .C1(n9568), .C2(n8098), .A(n7280), .B(n7279), .ZN(n7281)
         );
  OAI21_X1 U8979 ( .B1(n7282), .B2(n8082), .A(n7281), .ZN(P2_U3230) );
  INV_X1 U8980 ( .A(n7563), .ZN(n7286) );
  OAI222_X1 U8981 ( .A1(P1_U3084), .A2(n7283), .B1(n9463), .B2(n7286), .C1(
        n10281), .C2(n7885), .ZN(P1_U3328) );
  OAI222_X1 U8982 ( .A1(n8546), .A2(n7287), .B1(n8548), .B2(n7286), .C1(
        P2_U3152), .C2(n7285), .ZN(P2_U3333) );
  INV_X1 U8983 ( .A(n7288), .ZN(n7290) );
  NAND2_X1 U8984 ( .A1(n7290), .A2(n7289), .ZN(n7324) );
  NAND2_X1 U8985 ( .A1(n7288), .A2(n7291), .ZN(n7292) );
  NAND2_X1 U8986 ( .A1(n7324), .A2(n7292), .ZN(n7298) );
  NOR2_X1 U8987 ( .A1(n7298), .A2(n7293), .ZN(n7327) );
  INV_X1 U8988 ( .A(n7327), .ZN(n7301) );
  AOI22_X1 U8989 ( .A1(n8084), .A2(n8245), .B1(n8106), .B2(n8113), .ZN(n7295)
         );
  OAI211_X1 U8990 ( .C1(n7296), .C2(n8094), .A(n7295), .B(n7294), .ZN(n7297)
         );
  AOI21_X1 U8991 ( .B1(n7435), .B2(n8098), .A(n7297), .ZN(n7300) );
  NAND3_X1 U8992 ( .A1(n7298), .A2(n8078), .A3(n8112), .ZN(n7299) );
  OAI211_X1 U8993 ( .C1(n7301), .C2(n8082), .A(n7300), .B(n7299), .ZN(P2_U3243) );
  NOR2_X1 U8994 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7302), .ZN(n9718) );
  AOI21_X1 U8995 ( .B1(n8713), .B2(n9505), .A(n9718), .ZN(n7305) );
  OR2_X1 U8996 ( .A1(n8710), .A2(n7303), .ZN(n7304) );
  OAI211_X1 U8997 ( .C1(n8715), .C2(n9513), .A(n7305), .B(n7304), .ZN(n7321)
         );
  INV_X1 U8998 ( .A(n7306), .ZN(n7307) );
  NAND2_X1 U8999 ( .A1(n7308), .A2(n7307), .ZN(n7309) );
  OAI22_X1 U9000 ( .A1(n9526), .A2(n7985), .B1(n8675), .B2(n8003), .ZN(n7311)
         );
  XNOR2_X1 U9001 ( .A(n7311), .B(n8001), .ZN(n7314) );
  OR2_X1 U9002 ( .A1(n9526), .A2(n8003), .ZN(n7313) );
  NAND2_X1 U9003 ( .A1(n9017), .A2(n7998), .ZN(n7312) );
  NAND2_X1 U9004 ( .A1(n7313), .A2(n7312), .ZN(n7315) );
  NAND2_X1 U9005 ( .A1(n7314), .A2(n7315), .ZN(n7346) );
  INV_X1 U9006 ( .A(n7314), .ZN(n7317) );
  INV_X1 U9007 ( .A(n7315), .ZN(n7316) );
  NAND2_X1 U9008 ( .A1(n7317), .A2(n7316), .ZN(n7348) );
  NAND2_X1 U9009 ( .A1(n7346), .A2(n7348), .ZN(n7318) );
  XNOR2_X1 U9010 ( .A(n7347), .B(n7318), .ZN(n7319) );
  NOR2_X1 U9011 ( .A1(n7319), .A2(n8719), .ZN(n7320) );
  AOI211_X1 U9012 ( .C1(n9517), .C2(n8717), .A(n7321), .B(n7320), .ZN(n7322)
         );
  INV_X1 U9013 ( .A(n7322), .ZN(P1_U3215) );
  INV_X1 U9014 ( .A(n7572), .ZN(n7344) );
  AOI22_X1 U9015 ( .A1(n6020), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9465), .ZN(n7323) );
  OAI21_X1 U9016 ( .B1(n7344), .B2(n9463), .A(n7323), .ZN(P1_U3327) );
  INV_X1 U9017 ( .A(n7324), .ZN(n7326) );
  NOR3_X1 U9018 ( .A1(n7327), .A2(n7326), .A3(n7325), .ZN(n7330) );
  INV_X1 U9019 ( .A(n7328), .ZN(n7329) );
  OAI21_X1 U9020 ( .B1(n7330), .B2(n7329), .A(n8101), .ZN(n7334) );
  OAI22_X1 U9021 ( .A1(n7443), .A2(n8058), .B1(n8096), .B2(n7649), .ZN(n7331)
         );
  AOI211_X1 U9022 ( .C1(n8051), .C2(n7447), .A(n7332), .B(n7331), .ZN(n7333)
         );
  OAI211_X1 U9023 ( .C1(n9599), .C2(n8063), .A(n7334), .B(n7333), .ZN(P2_U3228) );
  XNOR2_X1 U9024 ( .A(n7336), .B(n7335), .ZN(n7342) );
  INV_X1 U9025 ( .A(n8445), .ZN(n7339) );
  AOI22_X1 U9026 ( .A1(n8106), .A2(n8450), .B1(n8084), .B2(n8451), .ZN(n7338)
         );
  OAI211_X1 U9027 ( .C1(n8094), .C2(n7339), .A(n7338), .B(n7337), .ZN(n7340)
         );
  AOI21_X1 U9028 ( .B1(n8523), .B2(n8098), .A(n7340), .ZN(n7341) );
  OAI21_X1 U9029 ( .B1(n7342), .B2(n8082), .A(n7341), .ZN(P2_U3240) );
  OAI222_X1 U9030 ( .A1(P2_U3152), .A2(n7345), .B1(n8548), .B2(n7344), .C1(
        n7343), .C2(n8546), .ZN(P2_U3332) );
  NAND2_X1 U9031 ( .A1(n7349), .A2(n7348), .ZN(n8603) );
  NAND2_X1 U9032 ( .A1(n9431), .A2(n8005), .ZN(n7351) );
  NAND2_X1 U9033 ( .A1(n9505), .A2(n7893), .ZN(n7350) );
  NAND2_X1 U9034 ( .A1(n7351), .A2(n7350), .ZN(n7352) );
  XNOR2_X1 U9035 ( .A(n7352), .B(n7996), .ZN(n7365) );
  AND2_X1 U9036 ( .A1(n9505), .A2(n7998), .ZN(n7353) );
  AOI21_X1 U9037 ( .B1(n9431), .B2(n8011), .A(n7353), .ZN(n7366) );
  XNOR2_X1 U9038 ( .A(n7365), .B(n7366), .ZN(n8681) );
  NAND2_X1 U9039 ( .A1(n9634), .A2(n8005), .ZN(n7355) );
  NAND2_X1 U9040 ( .A1(n9016), .A2(n7893), .ZN(n7354) );
  NAND2_X1 U9041 ( .A1(n7355), .A2(n7354), .ZN(n7356) );
  XNOR2_X1 U9042 ( .A(n7356), .B(n7996), .ZN(n8606) );
  NOR2_X1 U9043 ( .A1(n7357), .A2(n4868), .ZN(n7358) );
  AOI21_X1 U9044 ( .B1(n9634), .B2(n8011), .A(n7358), .ZN(n7369) );
  AND2_X1 U9045 ( .A1(n8606), .A2(n7369), .ZN(n7373) );
  OR2_X1 U9046 ( .A1(n8681), .A2(n7373), .ZN(n7359) );
  OR2_X2 U9047 ( .A1(n8603), .A2(n7359), .ZN(n7381) );
  NAND2_X1 U9048 ( .A1(n8762), .A2(n8005), .ZN(n7361) );
  NAND2_X1 U9049 ( .A1(n9015), .A2(n7893), .ZN(n7360) );
  NAND2_X1 U9050 ( .A1(n7361), .A2(n7360), .ZN(n7362) );
  XNOR2_X1 U9051 ( .A(n7362), .B(n8001), .ZN(n7376) );
  NAND2_X1 U9052 ( .A1(n8762), .A2(n7893), .ZN(n7364) );
  NAND2_X1 U9053 ( .A1(n9015), .A2(n7998), .ZN(n7363) );
  NAND2_X1 U9054 ( .A1(n7364), .A2(n7363), .ZN(n7377) );
  AND2_X1 U9055 ( .A1(n7376), .A2(n7377), .ZN(n7383) );
  INV_X1 U9056 ( .A(n7383), .ZN(n7374) );
  INV_X1 U9057 ( .A(n7365), .ZN(n7368) );
  INV_X1 U9058 ( .A(n7366), .ZN(n7367) );
  NAND2_X1 U9059 ( .A1(n7368), .A2(n7367), .ZN(n8604) );
  INV_X1 U9060 ( .A(n8606), .ZN(n7370) );
  INV_X1 U9061 ( .A(n7369), .ZN(n8605) );
  NAND2_X1 U9062 ( .A1(n7370), .A2(n8605), .ZN(n7371) );
  AND2_X1 U9063 ( .A1(n8604), .A2(n7371), .ZN(n7372) );
  OR2_X1 U9064 ( .A1(n7373), .A2(n7372), .ZN(n7380) );
  AND2_X1 U9065 ( .A1(n7374), .A2(n7380), .ZN(n7375) );
  NAND2_X2 U9066 ( .A1(n7381), .A2(n7375), .ZN(n7887) );
  INV_X1 U9067 ( .A(n7376), .ZN(n7379) );
  INV_X1 U9068 ( .A(n7377), .ZN(n7378) );
  NAND2_X1 U9069 ( .A1(n7379), .A2(n7378), .ZN(n7886) );
  INV_X1 U9070 ( .A(n7886), .ZN(n7385) );
  NAND2_X1 U9071 ( .A1(n7381), .A2(n7380), .ZN(n7382) );
  OAI21_X1 U9072 ( .B1(n7385), .B2(n7383), .A(n7382), .ZN(n7384) );
  OAI21_X1 U9073 ( .B1(n7887), .B2(n7385), .A(n7384), .ZN(n7386) );
  NAND2_X1 U9074 ( .A1(n7386), .A2(n8645), .ZN(n7392) );
  NOR2_X1 U9075 ( .A1(n8715), .A2(n7387), .ZN(n7389) );
  NAND2_X1 U9076 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9064) );
  OAI21_X1 U9077 ( .B1(n8648), .B2(n8709), .A(n9064), .ZN(n7388) );
  AOI211_X1 U9078 ( .C1(n7390), .C2(n9016), .A(n7389), .B(n7388), .ZN(n7391)
         );
  OAI211_X1 U9079 ( .C1(n9628), .C2(n8654), .A(n7392), .B(n7391), .ZN(P1_U3232) );
  INV_X1 U9080 ( .A(n7587), .ZN(n7454) );
  AOI22_X1 U9081 ( .A1(n9113), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n9465), .ZN(n7393) );
  OAI21_X1 U9082 ( .B1(n7454), .B2(n9463), .A(n7393), .ZN(P1_U3326) );
  NAND2_X1 U9083 ( .A1(n7397), .A2(n4475), .ZN(n7400) );
  AOI22_X1 U9084 ( .A1(n8730), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7398), .B2(
        n7502), .ZN(n7399) );
  NAND2_X1 U9085 ( .A1(n9315), .A2(n7401), .ZN(n7402) );
  INV_X1 U9086 ( .A(n9419), .ZN(n9322) );
  NAND2_X1 U9087 ( .A1(n7402), .A2(n5060), .ZN(n7496) );
  NAND2_X1 U9088 ( .A1(n7403), .A2(n4475), .ZN(n7405) );
  AOI22_X1 U9089 ( .A1(n8730), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9091), .B2(
        n7502), .ZN(n7404) );
  NAND2_X1 U9090 ( .A1(n8721), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7414) );
  INV_X1 U9091 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7406) );
  OR2_X1 U9092 ( .A1(n6273), .A2(n7406), .ZN(n7413) );
  INV_X1 U9093 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7408) );
  NAND2_X1 U9094 ( .A1(n7409), .A2(n7408), .ZN(n7410) );
  NAND2_X1 U9095 ( .A1(n7421), .A2(n7410), .ZN(n8628) );
  OR2_X1 U9096 ( .A1(n7623), .A2(n8628), .ZN(n7412) );
  INV_X1 U9097 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7417) );
  OR2_X1 U9098 ( .A1(n6274), .A2(n7417), .ZN(n7411) );
  NAND2_X1 U9099 ( .A1(n9416), .A2(n9311), .ZN(n8844) );
  NAND2_X1 U9100 ( .A1(n8845), .A2(n8844), .ZN(n8956) );
  XNOR2_X1 U9101 ( .A(n7496), .B(n8956), .ZN(n9418) );
  INV_X1 U9102 ( .A(n9301), .ZN(n7415) );
  AOI211_X1 U9103 ( .C1(n9416), .C2(n9316), .A(n9830), .B(n7415), .ZN(n9415)
         );
  INV_X1 U9104 ( .A(n9416), .ZN(n7416) );
  NOR2_X1 U9105 ( .A1(n7416), .A2(n9321), .ZN(n7419) );
  OAI22_X1 U9106 ( .A1(n9786), .A2(n7417), .B1(n8628), .B2(n9790), .ZN(n7418)
         );
  AOI211_X1 U9107 ( .C1(n9415), .C2(n9521), .A(n7419), .B(n7418), .ZN(n7432)
         );
  INV_X1 U9108 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7420) );
  NAND2_X1 U9109 ( .A1(n7421), .A2(n7420), .ZN(n7422) );
  NAND2_X1 U9110 ( .A1(n7486), .A2(n7422), .ZN(n9303) );
  OR2_X1 U9111 ( .A1(n7623), .A2(n9303), .ZN(n7427) );
  NAND2_X1 U9112 ( .A1(n8721), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7426) );
  INV_X1 U9113 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7423) );
  OR2_X1 U9114 ( .A1(n6273), .A2(n7423), .ZN(n7425) );
  INV_X1 U9115 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9304) );
  OR2_X1 U9116 ( .A1(n6274), .A2(n9304), .ZN(n7424) );
  NAND4_X1 U9117 ( .A1(n7427), .A2(n7426), .A3(n7425), .A4(n7424), .ZN(n9283)
         );
  OR2_X1 U9118 ( .A1(n9419), .A2(n8630), .ZN(n8839) );
  NAND2_X1 U9119 ( .A1(n9419), .A2(n8630), .ZN(n8838) );
  NAND2_X1 U9120 ( .A1(n8839), .A2(n8838), .ZN(n9323) );
  INV_X1 U9121 ( .A(n8828), .ZN(n9324) );
  NOR2_X1 U9122 ( .A1(n9323), .A2(n9324), .ZN(n7428) );
  NAND2_X1 U9123 ( .A1(n7429), .A2(n7428), .ZN(n9326) );
  XNOR2_X1 U9124 ( .A(n7614), .B(n8956), .ZN(n7430) );
  OAI222_X1 U9125 ( .A1(n9771), .A2(n8689), .B1(n9773), .B2(n8630), .C1(n7430), 
        .C2(n9509), .ZN(n9414) );
  NAND2_X1 U9126 ( .A1(n9414), .A2(n9786), .ZN(n7431) );
  OAI211_X1 U9127 ( .C1(n9418), .C2(n9335), .A(n7432), .B(n7431), .ZN(P1_U3275) );
  NAND2_X1 U9128 ( .A1(n7434), .A2(n7433), .ZN(n7437) );
  OR2_X1 U9129 ( .A1(n7435), .A2(n8112), .ZN(n7436) );
  NAND2_X1 U9130 ( .A1(n9599), .A2(n8245), .ZN(n7772) );
  NAND2_X1 U9131 ( .A1(n8246), .A2(n9578), .ZN(n7771) );
  NAND2_X1 U9132 ( .A1(n7439), .A2(n7858), .ZN(n7440) );
  NAND2_X1 U9133 ( .A1(n8248), .A2(n7440), .ZN(n9598) );
  AND2_X2 U9134 ( .A1(n7441), .A2(n7766), .ZN(n7442) );
  OAI21_X1 U9135 ( .B1(n7858), .B2(n7442), .A(n7648), .ZN(n7445) );
  OAI22_X1 U9136 ( .A1(n7649), .A2(n9581), .B1(n7443), .B2(n9579), .ZN(n7444)
         );
  AOI21_X1 U9137 ( .B1(n7445), .B2(n9868), .A(n7444), .ZN(n7446) );
  OAI21_X1 U9138 ( .B1(n9565), .B2(n9598), .A(n7446), .ZN(n9601) );
  NAND2_X1 U9139 ( .A1(n9601), .A2(n8436), .ZN(n7453) );
  INV_X1 U9140 ( .A(n7447), .ZN(n7448) );
  OAI22_X1 U9141 ( .A1(n9591), .A2(n7449), .B1(n7448), .B2(n9871), .ZN(n7451)
         );
  XNOR2_X1 U9142 ( .A(n8235), .B(n9599), .ZN(n9600) );
  NOR2_X1 U9143 ( .A1(n9600), .A2(n9873), .ZN(n7450) );
  AOI211_X1 U9144 ( .C1(n8440), .C2(n8246), .A(n7451), .B(n7450), .ZN(n7452)
         );
  OAI211_X1 U9145 ( .C1(n9598), .C2(n9584), .A(n7453), .B(n7452), .ZN(P2_U3280) );
  OAI222_X1 U9146 ( .A1(n8546), .A2(n7455), .B1(n8548), .B2(n7454), .C1(n7878), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9147 ( .A(n7598), .ZN(n7644) );
  AOI22_X1 U9148 ( .A1(n7456), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9465), .ZN(n7457) );
  OAI21_X1 U9149 ( .B1(n7644), .B2(n9463), .A(n7457), .ZN(P1_U3325) );
  INV_X1 U9150 ( .A(n8519), .ZN(n8252) );
  OAI21_X1 U9151 ( .B1(n7460), .B2(n7459), .A(n7458), .ZN(n7461) );
  NAND2_X1 U9152 ( .A1(n7461), .A2(n8101), .ZN(n7465) );
  OAI22_X1 U9153 ( .A1(n8254), .A2(n9581), .B1(n9580), .B2(n9579), .ZN(n8432)
         );
  NAND2_X1 U9154 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8232) );
  INV_X1 U9155 ( .A(n8232), .ZN(n7463) );
  NOR2_X1 U9156 ( .A1(n8094), .A2(n8438), .ZN(n7462) );
  AOI211_X1 U9157 ( .C1(n8075), .C2(n8432), .A(n7463), .B(n7462), .ZN(n7464)
         );
  OAI211_X1 U9158 ( .C1(n8252), .C2(n8063), .A(n7465), .B(n7464), .ZN(P2_U3221) );
  XNOR2_X1 U9159 ( .A(n4566), .B(n7466), .ZN(n7471) );
  OAI22_X1 U9160 ( .A1(n8094), .A2(n8411), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10290), .ZN(n7469) );
  OAI22_X1 U9161 ( .A1(n8418), .A2(n8058), .B1(n8096), .B2(n8419), .ZN(n7468)
         );
  AOI211_X1 U9162 ( .C1(n8513), .C2(n8098), .A(n7469), .B(n7468), .ZN(n7470)
         );
  OAI21_X1 U9163 ( .B1(n7471), .B2(n8082), .A(n7470), .ZN(P2_U3235) );
  NAND2_X1 U9164 ( .A1(n7472), .A2(n4475), .ZN(n7475) );
  NAND2_X1 U9165 ( .A1(n8730), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7474) );
  INV_X1 U9166 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10225) );
  INV_X1 U9167 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U9168 ( .A1(n7522), .A2(n8590), .ZN(n7478) );
  AND2_X1 U9169 ( .A1(n7532), .A2(n7478), .ZN(n9244) );
  NAND2_X1 U9170 ( .A1(n9244), .A2(n6646), .ZN(n7484) );
  NAND2_X1 U9171 ( .A1(n8721), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7483) );
  INV_X1 U9172 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n7479) );
  OR2_X1 U9173 ( .A1(n6273), .A2(n7479), .ZN(n7482) );
  INV_X1 U9174 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n7480) );
  OR2_X1 U9175 ( .A1(n7549), .A2(n7480), .ZN(n7481) );
  NAND2_X1 U9176 ( .A1(n7624), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7491) );
  INV_X1 U9177 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10262) );
  OR2_X1 U9178 ( .A1(n7628), .A2(n10262), .ZN(n7490) );
  INV_X1 U9179 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7485) );
  NAND2_X1 U9180 ( .A1(n7486), .A2(n7485), .ZN(n7487) );
  NAND2_X1 U9181 ( .A1(n7508), .A2(n7487), .ZN(n9293) );
  OR2_X1 U9182 ( .A1(n7623), .A2(n9293), .ZN(n7489) );
  INV_X1 U9183 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9294) );
  OR2_X1 U9184 ( .A1(n7549), .A2(n9294), .ZN(n7488) );
  NAND2_X1 U9185 ( .A1(n7492), .A2(n4475), .ZN(n7494) );
  AOI22_X1 U9186 ( .A1(n8730), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9741), .B2(
        n7502), .ZN(n7493) );
  INV_X1 U9187 ( .A(n9404), .ZN(n9292) );
  NAND2_X1 U9188 ( .A1(n7497), .A2(n4475), .ZN(n7499) );
  AOI22_X1 U9189 ( .A1(n8730), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9105), .B2(
        n7502), .ZN(n7498) );
  NAND2_X1 U9190 ( .A1(n9411), .A2(n9283), .ZN(n7500) );
  INV_X1 U9191 ( .A(n9411), .ZN(n9302) );
  AOI22_X1 U9192 ( .A1(n9299), .A2(n7500), .B1(n8689), .B2(n9302), .ZN(n9287)
         );
  NAND2_X1 U9193 ( .A1(n9404), .A2(n9312), .ZN(n8849) );
  NAND2_X1 U9194 ( .A1(n8860), .A2(n8849), .ZN(n9286) );
  NAND2_X1 U9195 ( .A1(n9287), .A2(n9286), .ZN(n9402) );
  OAI21_X1 U9196 ( .B1(n9312), .B2(n9292), .A(n9402), .ZN(n9267) );
  NAND2_X1 U9197 ( .A1(n7501), .A2(n4475), .ZN(n7504) );
  AOI22_X1 U9198 ( .A1(n8730), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9785), .B2(
        n7502), .ZN(n7503) );
  NAND2_X1 U9199 ( .A1(n7624), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7513) );
  INV_X1 U9200 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n7505) );
  OR2_X1 U9201 ( .A1(n7628), .A2(n7505), .ZN(n7512) );
  INV_X1 U9202 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7506) );
  OR2_X1 U9203 ( .A1(n6274), .A2(n7506), .ZN(n7511) );
  INV_X1 U9204 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U9205 ( .A1(n7508), .A2(n7507), .ZN(n7509) );
  NAND2_X1 U9206 ( .A1(n7520), .A2(n7509), .ZN(n8582) );
  OR2_X1 U9207 ( .A1(n7623), .A2(n8582), .ZN(n7510) );
  NAND2_X1 U9208 ( .A1(n9272), .A2(n9263), .ZN(n7514) );
  NAND2_X1 U9209 ( .A1(n9267), .A2(n7514), .ZN(n7516) );
  NAND2_X1 U9210 ( .A1(n9398), .A2(n9284), .ZN(n7515) );
  NAND2_X1 U9211 ( .A1(n7516), .A2(n7515), .ZN(n9252) );
  NAND2_X1 U9212 ( .A1(n7517), .A2(n4475), .ZN(n7519) );
  NAND2_X1 U9213 ( .A1(n8730), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U9214 ( .A1(n7624), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7526) );
  INV_X1 U9215 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10265) );
  OR2_X1 U9216 ( .A1(n7628), .A2(n10265), .ZN(n7525) );
  NAND2_X1 U9217 ( .A1(n7520), .A2(n10225), .ZN(n7521) );
  NAND2_X1 U9218 ( .A1(n7522), .A2(n7521), .ZN(n9256) );
  OR2_X1 U9219 ( .A1(n7623), .A2(n9256), .ZN(n7524) );
  INV_X1 U9220 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9257) );
  OR2_X1 U9221 ( .A1(n7549), .A2(n9257), .ZN(n7523) );
  NAND2_X1 U9222 ( .A1(n9387), .A2(n9264), .ZN(n8736) );
  NAND2_X1 U9223 ( .A1(n7528), .A2(n4475), .ZN(n7530) );
  NAND2_X1 U9224 ( .A1(n8730), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7529) );
  INV_X1 U9225 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10219) );
  INV_X1 U9226 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U9227 ( .A1(n7532), .A2(n8669), .ZN(n7533) );
  NAND2_X1 U9228 ( .A1(n7544), .A2(n7533), .ZN(n9224) );
  OR2_X1 U9229 ( .A1(n9224), .A2(n7623), .ZN(n7537) );
  NAND2_X1 U9230 ( .A1(n8721), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7535) );
  NAND2_X1 U9231 ( .A1(n7069), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7534) );
  AND2_X1 U9232 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  OAI211_X1 U9233 ( .C1(n6273), .C2(n10219), .A(n7537), .B(n7536), .ZN(n9240)
         );
  NOR2_X1 U9234 ( .A1(n9380), .A2(n9240), .ZN(n7538) );
  INV_X1 U9235 ( .A(n9240), .ZN(n8592) );
  NAND2_X1 U9236 ( .A1(n7539), .A2(n4475), .ZN(n7541) );
  NAND2_X1 U9237 ( .A1(n8730), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7540) );
  INV_X1 U9238 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n7548) );
  INV_X1 U9239 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7543) );
  NAND2_X1 U9240 ( .A1(n7544), .A2(n7543), .ZN(n7545) );
  NAND2_X1 U9241 ( .A1(n7555), .A2(n7545), .ZN(n9206) );
  OR2_X1 U9242 ( .A1(n9206), .A2(n7623), .ZN(n7547) );
  AOI22_X1 U9243 ( .A1(n7624), .A2(P1_REG0_REG_23__SCAN_IN), .B1(n8721), .B2(
        P1_REG1_REG_23__SCAN_IN), .ZN(n7546) );
  OAI211_X1 U9244 ( .C1(n7549), .C2(n7548), .A(n7547), .B(n7546), .ZN(n9230)
         );
  INV_X1 U9245 ( .A(n9375), .ZN(n9209) );
  INV_X1 U9246 ( .A(n9230), .ZN(n9194) );
  NAND2_X1 U9247 ( .A1(n7552), .A2(n4475), .ZN(n7554) );
  NAND2_X1 U9248 ( .A1(n8730), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7553) );
  INV_X1 U9249 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U9250 ( .A1(n7555), .A2(n8647), .ZN(n7556) );
  AND2_X1 U9251 ( .A1(n7579), .A2(n7556), .ZN(n9197) );
  NAND2_X1 U9252 ( .A1(n9197), .A2(n6646), .ZN(n7562) );
  INV_X1 U9253 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U9254 ( .A1(n8721), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9255 ( .A1(n7069), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7557) );
  OAI211_X1 U9256 ( .C1(n6273), .C2(n7559), .A(n7558), .B(n7557), .ZN(n7560)
         );
  INV_X1 U9257 ( .A(n7560), .ZN(n7561) );
  NAND2_X1 U9258 ( .A1(n8730), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7564) );
  XNOR2_X1 U9259 ( .A(n7579), .B(P1_REG3_REG_25__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U9260 ( .A1(n9179), .A2(n6646), .ZN(n7571) );
  INV_X1 U9261 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U9262 ( .A1(n8721), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7567) );
  NAND2_X1 U9263 ( .A1(n7069), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7566) );
  OAI211_X1 U9264 ( .C1(n7568), .C2(n6273), .A(n7567), .B(n7566), .ZN(n7569)
         );
  INV_X1 U9265 ( .A(n7569), .ZN(n7570) );
  NAND2_X1 U9266 ( .A1(n9365), .A2(n9195), .ZN(n8877) );
  INV_X1 U9267 ( .A(n9195), .ZN(n9013) );
  NAND2_X1 U9268 ( .A1(n7572), .A2(n4475), .ZN(n7574) );
  NAND2_X1 U9269 ( .A1(n8730), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7573) );
  INV_X1 U9270 ( .A(n7579), .ZN(n7576) );
  AND2_X1 U9271 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n7575) );
  NAND2_X1 U9272 ( .A1(n7576), .A2(n7575), .ZN(n7590) );
  INV_X1 U9273 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7578) );
  INV_X1 U9274 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7577) );
  OAI21_X1 U9275 ( .B1(n7579), .B2(n7578), .A(n7577), .ZN(n7580) );
  NAND2_X1 U9276 ( .A1(n7590), .A2(n7580), .ZN(n9170) );
  OR2_X1 U9277 ( .A1(n9170), .A2(n7623), .ZN(n7585) );
  INV_X1 U9278 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U9279 ( .A1(n7069), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7582) );
  NAND2_X1 U9280 ( .A1(n8721), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7581) );
  OAI211_X1 U9281 ( .C1(n6273), .C2(n10288), .A(n7582), .B(n7581), .ZN(n7583)
         );
  INV_X1 U9282 ( .A(n7583), .ZN(n7584) );
  NAND2_X1 U9283 ( .A1(n9174), .A2(n9149), .ZN(n7586) );
  NAND2_X1 U9284 ( .A1(n8730), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7588) );
  INV_X1 U9285 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10138) );
  NAND2_X1 U9286 ( .A1(n7590), .A2(n10138), .ZN(n7591) );
  NAND2_X1 U9287 ( .A1(n9156), .A2(n6646), .ZN(n7597) );
  INV_X1 U9288 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n7594) );
  NAND2_X1 U9289 ( .A1(n8721), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9290 ( .A1(n7069), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7592) );
  OAI211_X1 U9291 ( .C1(n6273), .C2(n7594), .A(n7593), .B(n7592), .ZN(n7595)
         );
  INV_X1 U9292 ( .A(n7595), .ZN(n7596) );
  NAND2_X1 U9293 ( .A1(n9356), .A2(n9166), .ZN(n8881) );
  INV_X1 U9294 ( .A(n9356), .ZN(n9146) );
  NAND2_X1 U9295 ( .A1(n7598), .A2(n4475), .ZN(n7600) );
  NAND2_X1 U9296 ( .A1(n8730), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7599) );
  INV_X1 U9297 ( .A(n7603), .ZN(n7601) );
  NAND2_X1 U9298 ( .A1(n7601), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9135) );
  INV_X1 U9299 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9300 ( .A1(n7603), .A2(n7602), .ZN(n7604) );
  NAND2_X1 U9301 ( .A1(n9135), .A2(n7604), .ZN(n8012) );
  INV_X1 U9302 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10137) );
  NAND2_X1 U9303 ( .A1(n7069), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U9304 ( .A1(n8721), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7605) );
  OAI211_X1 U9305 ( .C1(n6273), .C2(n10137), .A(n7606), .B(n7605), .ZN(n7607)
         );
  INV_X1 U9306 ( .A(n7607), .ZN(n7608) );
  NAND2_X1 U9307 ( .A1(n9350), .A2(n9150), .ZN(n9128) );
  NAND2_X1 U9308 ( .A1(n8896), .A2(n9128), .ZN(n7621) );
  OR2_X1 U9309 ( .A1(n7610), .A2(n7621), .ZN(n7611) );
  INV_X1 U9310 ( .A(n7621), .ZN(n8961) );
  NAND2_X1 U9311 ( .A1(n7611), .A2(n9126), .ZN(n9354) );
  NAND2_X1 U9312 ( .A1(n9300), .A2(n9292), .ZN(n9289) );
  INV_X1 U9313 ( .A(n9387), .ZN(n8597) );
  INV_X1 U9314 ( .A(n9365), .ZN(n9181) );
  NAND2_X1 U9315 ( .A1(n9178), .A2(n9174), .ZN(n9167) );
  AOI21_X1 U9316 ( .B1(n9350), .B2(n9154), .A(n9112), .ZN(n9351) );
  INV_X1 U9317 ( .A(n9350), .ZN(n9123) );
  INV_X1 U9318 ( .A(n8012), .ZN(n7612) );
  INV_X1 U9319 ( .A(n9790), .ZN(n9514) );
  AOI22_X1 U9320 ( .A1(n7612), .A2(n9514), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9767), .ZN(n7613) );
  OAI21_X1 U9321 ( .B1(n9123), .B2(n9321), .A(n7613), .ZN(n7635) );
  NAND2_X1 U9322 ( .A1(n9411), .A2(n8689), .ZN(n8848) );
  OR2_X1 U9323 ( .A1(n9411), .A2(n8689), .ZN(n8843) );
  INV_X1 U9324 ( .A(n8860), .ZN(n7615) );
  OR2_X1 U9325 ( .A1(n9398), .A2(n9263), .ZN(n8861) );
  NAND2_X1 U9326 ( .A1(n9398), .A2(n9263), .ZN(n8863) );
  INV_X1 U9327 ( .A(n9246), .ZN(n7617) );
  NOR2_X1 U9328 ( .A1(n7617), .A2(n8934), .ZN(n7618) );
  NAND2_X1 U9329 ( .A1(n9238), .A2(n8736), .ZN(n9229) );
  NAND2_X1 U9330 ( .A1(n9380), .A2(n8592), .ZN(n8931) );
  NAND2_X1 U9331 ( .A1(n9375), .A2(n9194), .ZN(n8888) );
  NAND2_X1 U9332 ( .A1(n9190), .A2(n8888), .ZN(n9213) );
  INV_X1 U9333 ( .A(n9213), .ZN(n7619) );
  INV_X1 U9334 ( .A(n9216), .ZN(n8618) );
  OR2_X1 U9335 ( .A1(n9372), .A2(n8618), .ZN(n8871) );
  NAND2_X1 U9336 ( .A1(n9183), .A2(n8877), .ZN(n9162) );
  AND2_X1 U9337 ( .A1(n8894), .A2(n9161), .ZN(n8779) );
  NAND2_X1 U9338 ( .A1(n9362), .A2(n9149), .ZN(n8880) );
  OAI21_X1 U9339 ( .B1(n4515), .B2(n8961), .A(n9129), .ZN(n7622) );
  INV_X1 U9340 ( .A(n7622), .ZN(n7633) );
  OR2_X1 U9341 ( .A1(n9135), .A2(n7623), .ZN(n7631) );
  INV_X1 U9342 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7627) );
  NAND2_X1 U9343 ( .A1(n7624), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U9344 ( .A1(n7069), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7625) );
  OAI211_X1 U9345 ( .C1(n7628), .C2(n7627), .A(n7626), .B(n7625), .ZN(n7629)
         );
  INV_X1 U9346 ( .A(n7629), .ZN(n7630) );
  NAND2_X1 U9347 ( .A1(n7631), .A2(n7630), .ZN(n9011) );
  INV_X1 U9348 ( .A(n9011), .ZN(n7632) );
  INV_X1 U9349 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10212) );
  INV_X1 U9350 ( .A(SI_28_), .ZN(n7638) );
  NAND2_X1 U9351 ( .A1(n7639), .A2(n7638), .ZN(n7640) );
  INV_X1 U9352 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10184) );
  INV_X1 U9353 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7641) );
  MUX2_X1 U9354 ( .A(n10184), .B(n7641), .S(n7677), .Z(n7656) );
  INV_X1 U9355 ( .A(SI_29_), .ZN(n10199) );
  INV_X1 U9356 ( .A(n7656), .ZN(n7642) );
  MUX2_X1 U9357 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7677), .Z(n7674) );
  INV_X1 U9358 ( .A(n8726), .ZN(n9464) );
  OAI222_X1 U9359 ( .A1(n8546), .A2(n10212), .B1(n8548), .B2(n9464), .C1(n7643), .C2(P2_U3152), .ZN(P2_U3328) );
  OAI222_X1 U9360 ( .A1(n8546), .A2(n7645), .B1(P2_U3152), .B2(n5794), .C1(
        n8548), .C2(n7644), .ZN(P2_U3330) );
  OAI222_X1 U9361 ( .A1(n6017), .A2(P1_U3084), .B1(n9463), .B2(n7647), .C1(
        n7646), .C2(n7885), .ZN(P1_U3329) );
  NAND2_X1 U9362 ( .A1(n9568), .A2(n7649), .ZN(n7693) );
  INV_X1 U9363 ( .A(n9574), .ZN(n7650) );
  NAND2_X1 U9364 ( .A1(n7651), .A2(n7695), .ZN(n8448) );
  NAND2_X1 U9365 ( .A1(n8523), .A2(n9580), .ZN(n7777) );
  NAND2_X1 U9366 ( .A1(n8448), .A2(n8449), .ZN(n8426) );
  OR2_X1 U9367 ( .A1(n8519), .A2(n8418), .ZN(n7786) );
  NAND2_X1 U9368 ( .A1(n8519), .A2(n8418), .ZN(n7782) );
  NAND2_X1 U9369 ( .A1(n7786), .A2(n7782), .ZN(n8427) );
  INV_X1 U9370 ( .A(n7784), .ZN(n8428) );
  NOR2_X1 U9371 ( .A1(n8427), .A2(n8428), .ZN(n7652) );
  NAND2_X1 U9372 ( .A1(n8513), .A2(n8254), .ZN(n7789) );
  NAND2_X1 U9373 ( .A1(n7780), .A2(n7789), .ZN(n8415) );
  OR2_X1 U9374 ( .A1(n8508), .A2(n8419), .ZN(n7791) );
  NAND2_X1 U9375 ( .A1(n8508), .A2(n8419), .ZN(n7790) );
  NAND2_X1 U9376 ( .A1(n7791), .A2(n7790), .ZN(n8404) );
  NAND2_X1 U9377 ( .A1(n8504), .A2(n8038), .ZN(n7781) );
  NAND2_X1 U9378 ( .A1(n7793), .A2(n7781), .ZN(n8376) );
  OR2_X2 U9379 ( .A1(n8377), .A2(n8376), .ZN(n8379) );
  OR2_X1 U9380 ( .A1(n8497), .A2(n8345), .ZN(n7799) );
  NAND2_X1 U9381 ( .A1(n8497), .A2(n8345), .ZN(n7795) );
  NAND2_X1 U9382 ( .A1(n7799), .A2(n7795), .ZN(n8362) );
  NAND2_X1 U9383 ( .A1(n8491), .A2(n8031), .ZN(n7804) );
  NAND2_X1 U9384 ( .A1(n8335), .A2(n7804), .ZN(n8356) );
  NAND2_X1 U9385 ( .A1(n8482), .A2(n8018), .ZN(n7812) );
  NOR2_X1 U9386 ( .A1(n8488), .A2(n8346), .ZN(n8313) );
  NOR2_X1 U9387 ( .A1(n8312), .A2(n8313), .ZN(n7655) );
  NAND2_X1 U9388 ( .A1(n8311), .A2(n7655), .ZN(n8315) );
  NAND2_X1 U9389 ( .A1(n8315), .A2(n7812), .ZN(n8303) );
  NAND2_X1 U9390 ( .A1(n8476), .A2(n8262), .ZN(n7808) );
  INV_X1 U9391 ( .A(n8304), .ZN(n8022) );
  OR2_X1 U9392 ( .A1(n8471), .A2(n8022), .ZN(n7814) );
  XNOR2_X1 U9393 ( .A(n7656), .B(SI_29_), .ZN(n7657) );
  NAND2_X1 U9394 ( .A1(n8729), .A2(n7680), .ZN(n7660) );
  OR2_X1 U9395 ( .A1(n7681), .A2(n10184), .ZN(n7659) );
  NAND2_X1 U9396 ( .A1(n8466), .A2(n7661), .ZN(n7822) );
  INV_X1 U9397 ( .A(n7670), .ZN(n7672) );
  NAND2_X1 U9398 ( .A1(n8726), .A2(n7680), .ZN(n7663) );
  OR2_X1 U9399 ( .A1(n7681), .A2(n10212), .ZN(n7662) );
  INV_X1 U9400 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U9401 ( .A1(n7664), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U9402 ( .A1(n7665), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7666) );
  OAI211_X1 U9403 ( .C1(n7668), .C2(n10245), .A(n7667), .B(n7666), .ZN(n8274)
         );
  AND2_X1 U9404 ( .A1(n8241), .A2(n8274), .ZN(n7828) );
  OAI22_X1 U9405 ( .A1(n7670), .A2(n7828), .B1(n7669), .B2(n8237), .ZN(n7671)
         );
  OAI21_X1 U9406 ( .B1(n7672), .B2(n8462), .A(n7671), .ZN(n7686) );
  NAND2_X1 U9407 ( .A1(n7675), .A2(n7674), .ZN(n7676) );
  MUX2_X1 U9408 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7677), .Z(n7678) );
  XNOR2_X1 U9409 ( .A(n7678), .B(SI_31_), .ZN(n7679) );
  NAND2_X1 U9410 ( .A1(n8789), .A2(n7680), .ZN(n7683) );
  OR2_X1 U9411 ( .A1(n7681), .A2(n6156), .ZN(n7682) );
  INV_X1 U9412 ( .A(n8237), .ZN(n7685) );
  INV_X1 U9413 ( .A(n8274), .ZN(n7684) );
  NAND2_X1 U9414 ( .A1(n8462), .A2(n7684), .ZN(n7826) );
  AOI21_X1 U9415 ( .B1(n7686), .B2(n7691), .A(n7692), .ZN(n7688) );
  XNOR2_X1 U9416 ( .A(n7688), .B(n7687), .ZN(n7876) );
  INV_X1 U9417 ( .A(n7691), .ZN(n7867) );
  INV_X1 U9418 ( .A(n7692), .ZN(n7830) );
  NAND3_X1 U9419 ( .A1(n7867), .A2(n7834), .A3(n7830), .ZN(n7833) );
  INV_X1 U9420 ( .A(n8362), .ZN(n8366) );
  AND2_X1 U9421 ( .A1(n7777), .A2(n7693), .ZN(n7694) );
  MUX2_X1 U9422 ( .A(n7695), .B(n7694), .S(n7834), .Z(n7776) );
  NAND2_X1 U9423 ( .A1(n7705), .A2(n7696), .ZN(n7697) );
  NAND2_X1 U9424 ( .A1(n7697), .A2(n7831), .ZN(n7704) );
  INV_X1 U9425 ( .A(n7698), .ZN(n7700) );
  NAND2_X1 U9426 ( .A1(n7700), .A2(n7699), .ZN(n7712) );
  NAND2_X1 U9427 ( .A1(n7701), .A2(n7871), .ZN(n7713) );
  OAI21_X1 U9428 ( .B1(n7712), .B2(n7713), .A(n7831), .ZN(n7702) );
  NAND2_X1 U9429 ( .A1(n7702), .A2(n7842), .ZN(n7703) );
  NAND3_X1 U9430 ( .A1(n6524), .A2(n7704), .A3(n7703), .ZN(n7709) );
  INV_X1 U9431 ( .A(n7724), .ZN(n7708) );
  AOI21_X1 U9432 ( .B1(n7729), .B2(n7706), .A(n7834), .ZN(n7707) );
  AOI21_X1 U9433 ( .B1(n7709), .B2(n7708), .A(n7707), .ZN(n7728) );
  NAND3_X1 U9434 ( .A1(n7712), .A2(n7711), .A3(n7710), .ZN(n7716) );
  INV_X1 U9435 ( .A(n7713), .ZN(n7715) );
  NAND3_X1 U9436 ( .A1(n7716), .A2(n7715), .A3(n7714), .ZN(n7718) );
  OR2_X1 U9437 ( .A1(n9926), .A2(n7717), .ZN(n7721) );
  NAND2_X1 U9438 ( .A1(n7718), .A2(n7721), .ZN(n7727) );
  AND2_X1 U9439 ( .A1(n7720), .A2(n7719), .ZN(n7723) );
  OAI211_X1 U9440 ( .C1(n7724), .C2(n7723), .A(n7722), .B(n7721), .ZN(n7725)
         );
  NAND2_X1 U9441 ( .A1(n7725), .A2(n7834), .ZN(n7726) );
  NOR2_X1 U9442 ( .A1(n7729), .A2(n7831), .ZN(n7730) );
  NOR2_X1 U9443 ( .A1(n7731), .A2(n7730), .ZN(n7735) );
  MUX2_X1 U9444 ( .A(n8120), .B(n9933), .S(n7834), .Z(n7732) );
  NOR2_X1 U9445 ( .A1(n7733), .A2(n7732), .ZN(n7734) );
  INV_X1 U9446 ( .A(n7737), .ZN(n7738) );
  MUX2_X1 U9447 ( .A(n5034), .B(n7738), .S(n7831), .Z(n7739) );
  NAND3_X1 U9448 ( .A1(n7745), .A2(n7742), .A3(n7747), .ZN(n7741) );
  NAND3_X1 U9449 ( .A1(n7741), .A2(n7746), .A3(n7751), .ZN(n7750) );
  INV_X1 U9450 ( .A(n7742), .ZN(n7743) );
  INV_X1 U9451 ( .A(n7746), .ZN(n7748) );
  INV_X1 U9452 ( .A(n7755), .ZN(n7752) );
  NOR2_X1 U9453 ( .A1(n7854), .A2(n7752), .ZN(n7754) );
  NOR2_X1 U9454 ( .A1(n7854), .A2(n4735), .ZN(n7759) );
  MUX2_X1 U9455 ( .A(n7761), .B(n7760), .S(n7831), .Z(n7762) );
  NAND2_X1 U9456 ( .A1(n7856), .A2(n7762), .ZN(n7763) );
  AOI21_X1 U9457 ( .B1(n7764), .B2(n7857), .A(n7763), .ZN(n7770) );
  INV_X1 U9458 ( .A(n7765), .ZN(n7768) );
  INV_X1 U9459 ( .A(n7766), .ZN(n7767) );
  MUX2_X1 U9460 ( .A(n7768), .B(n7767), .S(n7834), .Z(n7769) );
  OAI21_X1 U9461 ( .B1(n7770), .B2(n7769), .A(n7858), .ZN(n7774) );
  MUX2_X1 U9462 ( .A(n7772), .B(n7771), .S(n7831), .Z(n7773) );
  NAND3_X1 U9463 ( .A1(n7774), .A2(n7650), .A3(n7773), .ZN(n7775) );
  NAND3_X1 U9464 ( .A1(n7776), .A2(n7784), .A3(n7775), .ZN(n7785) );
  NAND3_X1 U9465 ( .A1(n7785), .A2(n7782), .A3(n7777), .ZN(n7779) );
  INV_X1 U9466 ( .A(n7789), .ZN(n7778) );
  NAND2_X1 U9467 ( .A1(n7791), .A2(n7780), .ZN(n7788) );
  INV_X1 U9468 ( .A(n7782), .ZN(n7783) );
  INV_X1 U9469 ( .A(n7786), .ZN(n7787) );
  NAND2_X1 U9470 ( .A1(n7790), .A2(n7789), .ZN(n7792) );
  INV_X1 U9471 ( .A(n7793), .ZN(n7794) );
  OR2_X1 U9472 ( .A1(n7795), .A2(n7834), .ZN(n7796) );
  OAI211_X1 U9473 ( .C1(n7798), .C2(n7797), .A(n7796), .B(n7804), .ZN(n7801)
         );
  AOI21_X1 U9474 ( .B1(n8335), .B2(n7799), .A(n7831), .ZN(n7800) );
  AOI21_X1 U9475 ( .B1(n7801), .B2(n8335), .A(n7800), .ZN(n7803) );
  INV_X1 U9476 ( .A(n8312), .ZN(n8261) );
  NAND2_X1 U9477 ( .A1(n8488), .A2(n8346), .ZN(n7802) );
  INV_X1 U9478 ( .A(n8313), .ZN(n7805) );
  AOI21_X1 U9479 ( .B1(n7806), .B2(n7805), .A(n7831), .ZN(n7807) );
  NAND2_X1 U9480 ( .A1(n8471), .A2(n8022), .ZN(n7809) );
  NAND2_X1 U9481 ( .A1(n7809), .A2(n7808), .ZN(n7810) );
  INV_X1 U9482 ( .A(n7812), .ZN(n7813) );
  NOR2_X1 U9483 ( .A1(n8263), .A2(n7813), .ZN(n7815) );
  AOI21_X1 U9484 ( .B1(n7816), .B2(n7815), .A(n5019), .ZN(n7817) );
  NAND2_X1 U9485 ( .A1(n7818), .A2(n7817), .ZN(n7821) );
  MUX2_X1 U9486 ( .A(n8304), .B(n8471), .S(n7834), .Z(n7819) );
  OAI21_X1 U9487 ( .B1(n8293), .B2(n8022), .A(n7819), .ZN(n7820) );
  NAND2_X1 U9488 ( .A1(n7823), .A2(n7822), .ZN(n8273) );
  INV_X1 U9489 ( .A(n7822), .ZN(n7825) );
  INV_X1 U9490 ( .A(n7823), .ZN(n7824) );
  MUX2_X1 U9491 ( .A(n7825), .B(n7824), .S(n7831), .Z(n7827) );
  INV_X1 U9492 ( .A(n7828), .ZN(n7829) );
  NAND2_X1 U9493 ( .A1(n7830), .A2(n7829), .ZN(n7866) );
  AOI21_X1 U9494 ( .B1(n7837), .B2(n7836), .A(n7870), .ZN(n7873) );
  INV_X1 U9495 ( .A(n8284), .ZN(n8281) );
  INV_X1 U9496 ( .A(n8273), .ZN(n8264) );
  INV_X1 U9497 ( .A(n8376), .ZN(n8257) );
  INV_X1 U9498 ( .A(n8404), .ZN(n7862) );
  INV_X1 U9499 ( .A(n8449), .ZN(n7860) );
  NOR4_X1 U9500 ( .A1(n7841), .A2(n7840), .A3(n7839), .A4(n7838), .ZN(n7843)
         );
  INV_X1 U9501 ( .A(n9876), .ZN(n9862) );
  NAND3_X1 U9502 ( .A1(n7843), .A2(n7842), .A3(n9862), .ZN(n7847) );
  NOR4_X1 U9503 ( .A1(n7847), .A2(n7846), .A3(n7845), .A4(n7844), .ZN(n7850)
         );
  NAND4_X1 U9504 ( .A1(n7851), .A2(n7850), .A3(n7849), .A4(n7848), .ZN(n7852)
         );
  NOR4_X1 U9505 ( .A1(n7854), .A2(n7853), .A3(n5030), .A4(n7852), .ZN(n7855)
         );
  NAND4_X1 U9506 ( .A1(n7858), .A2(n7857), .A3(n7856), .A4(n7855), .ZN(n7859)
         );
  NOR4_X1 U9507 ( .A1(n8427), .A2(n7860), .A3(n9574), .A4(n7859), .ZN(n7861)
         );
  NAND4_X1 U9508 ( .A1(n8257), .A2(n7862), .A3(n7653), .A4(n7861), .ZN(n7863)
         );
  NOR4_X1 U9509 ( .A1(n8312), .A2(n8362), .A3(n8356), .A4(n7863), .ZN(n7864)
         );
  NAND4_X1 U9510 ( .A1(n8264), .A2(n8302), .A3(n7864), .A4(n8326), .ZN(n7865)
         );
  XNOR2_X1 U9511 ( .A(n7868), .B(n9573), .ZN(n7872) );
  OAI22_X1 U9512 ( .A1(n7872), .A2(n7871), .B1(n7870), .B2(n7869), .ZN(n7874)
         );
  NOR4_X1 U9513 ( .A1(n9886), .A2(n7878), .A3(n7877), .A4(n9579), .ZN(n7881)
         );
  OAI21_X1 U9514 ( .B1(n7882), .B2(n7879), .A(P2_B_REG_SCAN_IN), .ZN(n7880) );
  OAI22_X1 U9515 ( .A1(n7883), .A2(n7882), .B1(n7881), .B2(n7880), .ZN(
        P2_U3244) );
  OAI222_X1 U9516 ( .A1(n7885), .A2(n10234), .B1(n9463), .B2(n7884), .C1(
        P1_U3084), .C2(n4473), .ZN(P1_U3334) );
  NAND2_X1 U9517 ( .A1(n9426), .A2(n8005), .ZN(n7889) );
  NAND2_X1 U9518 ( .A1(n9328), .A2(n7893), .ZN(n7888) );
  NAND2_X1 U9519 ( .A1(n7889), .A2(n7888), .ZN(n7890) );
  XNOR2_X1 U9520 ( .A(n7890), .B(n7996), .ZN(n7905) );
  NAND2_X1 U9521 ( .A1(n9426), .A2(n7893), .ZN(n7892) );
  NAND2_X1 U9522 ( .A1(n9328), .A2(n7998), .ZN(n7891) );
  NAND2_X1 U9523 ( .A1(n7892), .A2(n7891), .ZN(n8562) );
  NAND2_X1 U9524 ( .A1(n9416), .A2(n8005), .ZN(n7895) );
  NAND2_X1 U9525 ( .A1(n9329), .A2(n7893), .ZN(n7894) );
  NAND2_X1 U9526 ( .A1(n7895), .A2(n7894), .ZN(n7896) );
  XNOR2_X1 U9527 ( .A(n7896), .B(n8001), .ZN(n8625) );
  NAND2_X1 U9528 ( .A1(n9416), .A2(n8011), .ZN(n7898) );
  NAND2_X1 U9529 ( .A1(n9329), .A2(n7998), .ZN(n7897) );
  NAND2_X1 U9530 ( .A1(n7898), .A2(n7897), .ZN(n8624) );
  NAND2_X1 U9531 ( .A1(n9419), .A2(n8011), .ZN(n7900) );
  NAND2_X1 U9532 ( .A1(n9014), .A2(n7998), .ZN(n7899) );
  NAND2_X1 U9533 ( .A1(n7900), .A2(n7899), .ZN(n8707) );
  NAND2_X1 U9534 ( .A1(n9419), .A2(n8005), .ZN(n7902) );
  NAND2_X1 U9535 ( .A1(n9014), .A2(n8011), .ZN(n7901) );
  NAND2_X1 U9536 ( .A1(n7902), .A2(n7901), .ZN(n7903) );
  XNOR2_X1 U9537 ( .A(n7903), .B(n8001), .ZN(n7907) );
  AOI22_X1 U9538 ( .A1(n8625), .A2(n8624), .B1(n8707), .B2(n7907), .ZN(n7904)
         );
  INV_X1 U9539 ( .A(n8625), .ZN(n7910) );
  OAI21_X1 U9540 ( .B1(n7907), .B2(n8707), .A(n8624), .ZN(n7909) );
  NOR2_X1 U9541 ( .A1(n8624), .A2(n8707), .ZN(n7908) );
  INV_X1 U9542 ( .A(n7907), .ZN(n8622) );
  AOI22_X1 U9543 ( .A1(n7910), .A2(n7909), .B1(n7908), .B2(n8622), .ZN(n7911)
         );
  NAND2_X1 U9544 ( .A1(n9411), .A2(n8005), .ZN(n7913) );
  NAND2_X1 U9545 ( .A1(n9283), .A2(n8011), .ZN(n7912) );
  NAND2_X1 U9546 ( .A1(n7913), .A2(n7912), .ZN(n7914) );
  XNOR2_X1 U9547 ( .A(n7914), .B(n8001), .ZN(n7916) );
  AND2_X1 U9548 ( .A1(n9283), .A2(n7998), .ZN(n7915) );
  AOI21_X1 U9549 ( .B1(n9411), .B2(n8011), .A(n7915), .ZN(n7917) );
  XNOR2_X1 U9550 ( .A(n7916), .B(n7917), .ZN(n8635) );
  INV_X1 U9551 ( .A(n7916), .ZN(n7918) );
  NAND2_X1 U9552 ( .A1(n7918), .A2(n7917), .ZN(n7919) );
  NAND2_X1 U9553 ( .A1(n9404), .A2(n8005), .ZN(n7922) );
  INV_X1 U9554 ( .A(n9312), .ZN(n9276) );
  NAND2_X1 U9555 ( .A1(n9276), .A2(n8011), .ZN(n7921) );
  NAND2_X1 U9556 ( .A1(n7922), .A2(n7921), .ZN(n7923) );
  NAND2_X1 U9557 ( .A1(n9404), .A2(n8011), .ZN(n7925) );
  NAND2_X1 U9558 ( .A1(n9276), .A2(n7998), .ZN(n7924) );
  NAND2_X1 U9559 ( .A1(n7925), .A2(n7924), .ZN(n8687) );
  OAI22_X1 U9560 ( .A1(n9272), .A2(n7985), .B1(n9263), .B2(n8003), .ZN(n7926)
         );
  XNOR2_X1 U9561 ( .A(n7926), .B(n7996), .ZN(n7931) );
  OR2_X1 U9562 ( .A1(n9272), .A2(n8003), .ZN(n7928) );
  NAND2_X1 U9563 ( .A1(n9284), .A2(n7998), .ZN(n7927) );
  NAND2_X1 U9564 ( .A1(n7928), .A2(n7927), .ZN(n7929) );
  XNOR2_X1 U9565 ( .A(n7931), .B(n7929), .ZN(n8580) );
  INV_X1 U9566 ( .A(n7929), .ZN(n7930) );
  NAND2_X1 U9567 ( .A1(n7931), .A2(n7930), .ZN(n7932) );
  NAND2_X1 U9568 ( .A1(n8578), .A2(n7932), .ZN(n8659) );
  OAI22_X1 U9569 ( .A1(n9255), .A2(n7985), .B1(n8591), .B2(n8003), .ZN(n7933)
         );
  XNOR2_X1 U9570 ( .A(n7933), .B(n8001), .ZN(n7936) );
  OR2_X1 U9571 ( .A1(n9255), .A2(n8003), .ZN(n7935) );
  NAND2_X1 U9572 ( .A1(n9277), .A2(n7998), .ZN(n7934) );
  NAND2_X1 U9573 ( .A1(n7935), .A2(n7934), .ZN(n7937) );
  NAND2_X1 U9574 ( .A1(n7936), .A2(n7937), .ZN(n8656) );
  NAND2_X1 U9575 ( .A1(n8659), .A2(n8656), .ZN(n7940) );
  INV_X1 U9576 ( .A(n7936), .ZN(n7939) );
  INV_X1 U9577 ( .A(n7937), .ZN(n7938) );
  NAND2_X1 U9578 ( .A1(n7939), .A2(n7938), .ZN(n8657) );
  NAND2_X1 U9579 ( .A1(n7940), .A2(n8657), .ZN(n8587) );
  NAND2_X1 U9580 ( .A1(n9387), .A2(n8005), .ZN(n7942) );
  NAND2_X1 U9581 ( .A1(n9231), .A2(n8011), .ZN(n7941) );
  NAND2_X1 U9582 ( .A1(n7942), .A2(n7941), .ZN(n7943) );
  XNOR2_X1 U9583 ( .A(n7943), .B(n8001), .ZN(n7945) );
  NOR2_X1 U9584 ( .A1(n9264), .A2(n4868), .ZN(n7944) );
  AOI21_X1 U9585 ( .B1(n9387), .B2(n8011), .A(n7944), .ZN(n7946) );
  XNOR2_X1 U9586 ( .A(n7945), .B(n7946), .ZN(n8588) );
  NAND2_X1 U9587 ( .A1(n8587), .A2(n8588), .ZN(n7949) );
  INV_X1 U9588 ( .A(n7945), .ZN(n7947) );
  NAND2_X1 U9589 ( .A1(n7947), .A2(n7946), .ZN(n7948) );
  NAND2_X1 U9590 ( .A1(n7949), .A2(n7948), .ZN(n7954) );
  AND2_X1 U9591 ( .A1(n9240), .A2(n7998), .ZN(n7950) );
  AOI21_X1 U9592 ( .B1(n9380), .B2(n8011), .A(n7950), .ZN(n7955) );
  NAND2_X1 U9593 ( .A1(n7954), .A2(n7955), .ZN(n8665) );
  NAND2_X1 U9594 ( .A1(n9380), .A2(n8005), .ZN(n7952) );
  NAND2_X1 U9595 ( .A1(n9240), .A2(n8011), .ZN(n7951) );
  NAND2_X1 U9596 ( .A1(n7952), .A2(n7951), .ZN(n7953) );
  XNOR2_X1 U9597 ( .A(n7953), .B(n8001), .ZN(n8668) );
  NAND2_X1 U9598 ( .A1(n8665), .A2(n8668), .ZN(n7963) );
  NAND2_X1 U9599 ( .A1(n7963), .A2(n8666), .ZN(n7961) );
  NAND2_X1 U9600 ( .A1(n9375), .A2(n8005), .ZN(n7959) );
  NAND2_X1 U9601 ( .A1(n9230), .A2(n8011), .ZN(n7958) );
  NAND2_X1 U9602 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  XNOR2_X1 U9603 ( .A(n7960), .B(n8001), .ZN(n7964) );
  NAND2_X1 U9604 ( .A1(n7961), .A2(n7964), .ZN(n8571) );
  AND2_X1 U9605 ( .A1(n7998), .A2(n9230), .ZN(n7962) );
  AOI21_X1 U9606 ( .B1(n9375), .B2(n8011), .A(n7962), .ZN(n8570) );
  INV_X1 U9607 ( .A(n7964), .ZN(n7965) );
  AND2_X1 U9608 ( .A1(n8666), .A2(n7965), .ZN(n7966) );
  NAND2_X1 U9609 ( .A1(n9372), .A2(n8005), .ZN(n7968) );
  NAND2_X1 U9610 ( .A1(n9216), .A2(n8011), .ZN(n7967) );
  NAND2_X1 U9611 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  XNOR2_X1 U9612 ( .A(n7969), .B(n7996), .ZN(n7971) );
  AND2_X1 U9613 ( .A1(n9216), .A2(n7998), .ZN(n7970) );
  AOI21_X1 U9614 ( .B1(n9372), .B2(n8011), .A(n7970), .ZN(n7972) );
  NAND2_X1 U9615 ( .A1(n7971), .A2(n7972), .ZN(n7976) );
  INV_X1 U9616 ( .A(n7971), .ZN(n7974) );
  INV_X1 U9617 ( .A(n7972), .ZN(n7973) );
  NAND2_X1 U9618 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  AND2_X1 U9619 ( .A1(n7976), .A2(n7975), .ZN(n8643) );
  NAND2_X1 U9620 ( .A1(n9365), .A2(n8005), .ZN(n7978) );
  NAND2_X1 U9621 ( .A1(n9013), .A2(n8011), .ZN(n7977) );
  NAND2_X1 U9622 ( .A1(n7978), .A2(n7977), .ZN(n7979) );
  XNOR2_X1 U9623 ( .A(n7979), .B(n8001), .ZN(n7981) );
  NOR2_X1 U9624 ( .A1(n9195), .A2(n4868), .ZN(n7980) );
  AOI21_X1 U9625 ( .B1(n9365), .B2(n8011), .A(n7980), .ZN(n7982) );
  XNOR2_X1 U9626 ( .A(n7981), .B(n7982), .ZN(n8615) );
  INV_X1 U9627 ( .A(n7981), .ZN(n7983) );
  NAND2_X1 U9628 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  NAND2_X1 U9629 ( .A1(n8613), .A2(n7984), .ZN(n8698) );
  OAI22_X1 U9630 ( .A1(n9174), .A2(n7985), .B1(n9149), .B2(n8003), .ZN(n7986)
         );
  XNOR2_X1 U9631 ( .A(n7986), .B(n8001), .ZN(n7989) );
  OR2_X1 U9632 ( .A1(n9174), .A2(n8003), .ZN(n7988) );
  NAND2_X1 U9633 ( .A1(n9184), .A2(n7998), .ZN(n7987) );
  NAND2_X1 U9634 ( .A1(n7988), .A2(n7987), .ZN(n7990) );
  NAND2_X1 U9635 ( .A1(n7989), .A2(n7990), .ZN(n8695) );
  NAND2_X1 U9636 ( .A1(n8698), .A2(n8695), .ZN(n7993) );
  INV_X1 U9637 ( .A(n7989), .ZN(n7992) );
  INV_X1 U9638 ( .A(n7990), .ZN(n7991) );
  NAND2_X1 U9639 ( .A1(n7992), .A2(n7991), .ZN(n8696) );
  NAND2_X1 U9640 ( .A1(n7993), .A2(n8696), .ZN(n8554) );
  NAND2_X1 U9641 ( .A1(n9356), .A2(n8005), .ZN(n7995) );
  NAND2_X1 U9642 ( .A1(n9012), .A2(n8011), .ZN(n7994) );
  NAND2_X1 U9643 ( .A1(n7995), .A2(n7994), .ZN(n7997) );
  XNOR2_X1 U9644 ( .A(n7997), .B(n7996), .ZN(n8552) );
  NAND2_X1 U9645 ( .A1(n9350), .A2(n8011), .ZN(n8000) );
  NAND2_X1 U9646 ( .A1(n9124), .A2(n7998), .ZN(n7999) );
  NAND2_X1 U9647 ( .A1(n8000), .A2(n7999), .ZN(n8002) );
  XNOR2_X1 U9648 ( .A(n8002), .B(n8001), .ZN(n8007) );
  NOR2_X1 U9649 ( .A1(n9150), .A2(n8003), .ZN(n8004) );
  AOI21_X1 U9650 ( .B1(n9350), .B2(n8005), .A(n8004), .ZN(n8006) );
  XNOR2_X1 U9651 ( .A(n8007), .B(n8006), .ZN(n8009) );
  INV_X1 U9652 ( .A(n8009), .ZN(n8008) );
  NOR2_X1 U9653 ( .A1(n9166), .A2(n4868), .ZN(n8010) );
  AOI21_X1 U9654 ( .B1(n9356), .B2(n8011), .A(n8010), .ZN(n8551) );
  NOR2_X1 U9655 ( .A1(n8012), .A2(n8715), .ZN(n8015) );
  AOI22_X1 U9656 ( .A1(n9011), .A2(n8713), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8013) );
  OAI21_X1 U9657 ( .B1(n9166), .B2(n8710), .A(n8013), .ZN(n8014) );
  AOI211_X1 U9658 ( .C1(n9350), .C2(n8717), .A(n8015), .B(n8014), .ZN(n8016)
         );
  INV_X1 U9659 ( .A(n8476), .ZN(n8301) );
  NAND3_X1 U9660 ( .A1(n8019), .A2(n8078), .A3(n8305), .ZN(n8020) );
  OAI22_X1 U9661 ( .A1(n8094), .A2(n8298), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10305), .ZN(n8024) );
  NOR2_X1 U9662 ( .A1(n8022), .A2(n8096), .ZN(n8023) );
  AOI211_X1 U9663 ( .C1(n8106), .C2(n8305), .A(n8024), .B(n8023), .ZN(n8025)
         );
  OAI211_X1 U9664 ( .C1(n8301), .C2(n8063), .A(n8026), .B(n8025), .ZN(P2_U3216) );
  INV_X1 U9665 ( .A(n8345), .ZN(n8258) );
  NAND2_X1 U9666 ( .A1(n8078), .A2(n8258), .ZN(n8030) );
  OR2_X1 U9667 ( .A1(n8082), .A2(n8027), .ZN(n8029) );
  MUX2_X1 U9668 ( .A(n8030), .B(n8029), .S(n8028), .Z(n8035) );
  AOI22_X1 U9669 ( .A1(n8051), .A2(n8369), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8034) );
  AOI22_X1 U9670 ( .A1(n8084), .A2(n8364), .B1(n8106), .B2(n8397), .ZN(n8033)
         );
  NAND2_X1 U9671 ( .A1(n8497), .A2(n8098), .ZN(n8032) );
  NAND4_X1 U9672 ( .A1(n8035), .A2(n8034), .A3(n8033), .A4(n8032), .ZN(
        P2_U3218) );
  XNOR2_X1 U9673 ( .A(n8037), .B(n8036), .ZN(n8042) );
  OAI22_X1 U9674 ( .A1(n8094), .A2(n8400), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10273), .ZN(n8040) );
  OAI22_X1 U9675 ( .A1(n8254), .A2(n8058), .B1(n8096), .B2(n8038), .ZN(n8039)
         );
  AOI211_X1 U9676 ( .C1(n8508), .C2(n8098), .A(n8040), .B(n8039), .ZN(n8041)
         );
  OAI21_X1 U9677 ( .B1(n8042), .B2(n8082), .A(n8041), .ZN(P2_U3225) );
  XNOR2_X1 U9678 ( .A(n8044), .B(n8043), .ZN(n8045) );
  XNOR2_X1 U9679 ( .A(n8046), .B(n8045), .ZN(n8053) );
  AOI22_X1 U9680 ( .A1(n8305), .A2(n9865), .B1(n9864), .B2(n8364), .ZN(n8338)
         );
  OAI22_X1 U9681 ( .A1(n8338), .A2(n8048), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8047), .ZN(n8050) );
  NOR2_X1 U9682 ( .A1(n8260), .A2(n8063), .ZN(n8049) );
  AOI211_X1 U9683 ( .C1(n8051), .C2(n8328), .A(n8050), .B(n8049), .ZN(n8052)
         );
  OAI21_X1 U9684 ( .B1(n8053), .B2(n8082), .A(n8052), .ZN(P2_U3227) );
  INV_X1 U9685 ( .A(n8491), .ZN(n8354) );
  NAND2_X1 U9686 ( .A1(n8078), .A2(n8364), .ZN(n8057) );
  OR2_X1 U9687 ( .A1(n8082), .A2(n8054), .ZN(n8056) );
  MUX2_X1 U9688 ( .A(n8057), .B(n8056), .S(n8055), .Z(n8062) );
  NOR2_X1 U9689 ( .A1(n8094), .A2(n8351), .ZN(n8060) );
  OAI22_X1 U9690 ( .A1(n8345), .A2(n8058), .B1(n8096), .B2(n8346), .ZN(n8059)
         );
  AOI211_X1 U9691 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3152), .A(n8060), 
        .B(n8059), .ZN(n8061) );
  OAI211_X1 U9692 ( .C1(n8354), .C2(n8063), .A(n8062), .B(n8061), .ZN(P2_U3231) );
  AND2_X1 U9693 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8142) );
  OAI22_X1 U9694 ( .A1(n8096), .A2(n8064), .B1(n8094), .B2(n9872), .ZN(n8065)
         );
  AOI211_X1 U9695 ( .C1(n9869), .C2(n8098), .A(n8142), .B(n8065), .ZN(n8073)
         );
  OAI21_X1 U9696 ( .B1(n6174), .B2(n8068), .A(n8066), .ZN(n8067) );
  NAND2_X1 U9697 ( .A1(n8067), .A2(n8101), .ZN(n8072) );
  NOR3_X1 U9698 ( .A1(n8105), .A2(n8069), .A3(n8068), .ZN(n8070) );
  OAI21_X1 U9699 ( .B1(n8070), .B2(n8106), .A(n5855), .ZN(n8071) );
  NAND3_X1 U9700 ( .A1(n8073), .A2(n8072), .A3(n8071), .ZN(P2_U3232) );
  INV_X1 U9701 ( .A(n8074), .ZN(n8083) );
  OAI22_X1 U9702 ( .A1(n8345), .A2(n9581), .B1(n8419), .B2(n9579), .ZN(n8378)
         );
  AOI22_X1 U9703 ( .A1(n8075), .A2(n8378), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8076) );
  OAI21_X1 U9704 ( .B1(n8387), .B2(n8094), .A(n8076), .ZN(n8077) );
  AOI21_X1 U9705 ( .B1(n8504), .B2(n8098), .A(n8077), .ZN(n8081) );
  NAND3_X1 U9706 ( .A1(n8079), .A2(n8078), .A3(n8397), .ZN(n8080) );
  OAI211_X1 U9707 ( .C1(n8083), .C2(n8082), .A(n8081), .B(n8080), .ZN(P2_U3237) );
  AOI22_X1 U9708 ( .A1(n8106), .A2(n8124), .B1(n8084), .B2(n5855), .ZN(n8092)
         );
  OAI211_X1 U9709 ( .C1(n8086), .C2(n8085), .A(n8101), .B(n6172), .ZN(n8091)
         );
  NAND2_X1 U9710 ( .A1(n8098), .A2(n8087), .ZN(n8090) );
  OAI21_X1 U9711 ( .B1(n8088), .B2(P2_U3152), .A(P2_REG3_REG_2__SCAN_IN), .ZN(
        n8089) );
  NAND4_X1 U9712 ( .A1(n8092), .A2(n8091), .A3(n8090), .A4(n8089), .ZN(
        P2_U3239) );
  AND2_X1 U9713 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8166) );
  OAI22_X1 U9714 ( .A1(n8096), .A2(n8095), .B1(n8094), .B2(n8093), .ZN(n8097)
         );
  AOI211_X1 U9715 ( .C1(n9926), .C2(n8098), .A(n8166), .B(n8097), .ZN(n8110)
         );
  OAI21_X1 U9716 ( .B1(n8103), .B2(n8100), .A(n8099), .ZN(n8102) );
  NAND2_X1 U9717 ( .A1(n8102), .A2(n8101), .ZN(n8109) );
  NOR3_X1 U9718 ( .A1(n8105), .A2(n8104), .A3(n8103), .ZN(n8107) );
  OAI21_X1 U9719 ( .B1(n8107), .B2(n8106), .A(n9866), .ZN(n8108) );
  NAND3_X1 U9720 ( .A1(n8110), .A2(n8109), .A3(n8108), .ZN(P2_U3241) );
  MUX2_X1 U9721 ( .A(n8274), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8123), .Z(
        P2_U3582) );
  MUX2_X1 U9722 ( .A(n8287), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8123), .Z(
        P2_U3581) );
  MUX2_X1 U9723 ( .A(n8304), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8123), .Z(
        P2_U3580) );
  MUX2_X1 U9724 ( .A(n8286), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8123), .Z(
        P2_U3579) );
  MUX2_X1 U9725 ( .A(n8305), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8123), .Z(
        P2_U3578) );
  MUX2_X1 U9726 ( .A(n8111), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8123), .Z(
        P2_U3577) );
  MUX2_X1 U9727 ( .A(n8364), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8123), .Z(
        P2_U3576) );
  MUX2_X1 U9728 ( .A(n8258), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8123), .Z(
        P2_U3575) );
  MUX2_X1 U9729 ( .A(n8397), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8123), .Z(
        P2_U3574) );
  INV_X1 U9730 ( .A(n8419), .ZN(n8255) );
  MUX2_X1 U9731 ( .A(n8255), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8123), .Z(
        P2_U3573) );
  INV_X1 U9732 ( .A(n8254), .ZN(n8396) );
  MUX2_X1 U9733 ( .A(n8396), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8123), .Z(
        P2_U3572) );
  MUX2_X1 U9734 ( .A(n8451), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8123), .Z(
        P2_U3571) );
  INV_X1 U9735 ( .A(n9580), .ZN(n8250) );
  MUX2_X1 U9736 ( .A(n8250), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8123), .Z(
        P2_U3570) );
  MUX2_X1 U9737 ( .A(n8450), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8123), .Z(
        P2_U3569) );
  MUX2_X1 U9738 ( .A(n8245), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8123), .Z(
        P2_U3568) );
  MUX2_X1 U9739 ( .A(n8112), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8123), .Z(
        P2_U3567) );
  MUX2_X1 U9740 ( .A(n8113), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8123), .Z(
        P2_U3566) );
  MUX2_X1 U9741 ( .A(n8114), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8123), .Z(
        P2_U3565) );
  MUX2_X1 U9742 ( .A(n8115), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8123), .Z(
        P2_U3564) );
  MUX2_X1 U9743 ( .A(n8116), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8123), .Z(
        P2_U3563) );
  MUX2_X1 U9744 ( .A(n8117), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8123), .Z(
        P2_U3562) );
  MUX2_X1 U9745 ( .A(n8118), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8123), .Z(
        P2_U3561) );
  MUX2_X1 U9746 ( .A(n8119), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8123), .Z(
        P2_U3560) );
  MUX2_X1 U9747 ( .A(n8120), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8123), .Z(
        P2_U3559) );
  MUX2_X1 U9748 ( .A(n8121), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8123), .Z(
        P2_U3558) );
  MUX2_X1 U9749 ( .A(n9866), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8123), .Z(
        P2_U3557) );
  MUX2_X1 U9750 ( .A(n8122), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8123), .Z(
        P2_U3556) );
  MUX2_X1 U9751 ( .A(n5855), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8123), .Z(
        P2_U3555) );
  MUX2_X1 U9752 ( .A(n6158), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8123), .Z(
        P2_U3554) );
  MUX2_X1 U9753 ( .A(n8124), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8123), .Z(
        P2_U3553) );
  MUX2_X1 U9754 ( .A(n6157), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8123), .Z(
        P2_U3552) );
  OAI211_X1 U9755 ( .C1(n8127), .C2(n8126), .A(n9850), .B(n8125), .ZN(n8138)
         );
  NOR2_X1 U9756 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8128), .ZN(n8129) );
  AOI21_X1 U9757 ( .B1(n9857), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8129), .ZN(
        n8137) );
  NAND2_X1 U9758 ( .A1(n9477), .A2(n8130), .ZN(n8136) );
  AOI21_X1 U9759 ( .B1(n8133), .B2(n8132), .A(n8131), .ZN(n8134) );
  NAND2_X1 U9760 ( .A1(n9849), .A2(n8134), .ZN(n8135) );
  NAND4_X1 U9761 ( .A1(n8138), .A2(n8137), .A3(n8136), .A4(n8135), .ZN(
        P2_U3248) );
  OAI211_X1 U9762 ( .C1(n8141), .C2(n8140), .A(n9850), .B(n8139), .ZN(n8150)
         );
  AOI21_X1 U9763 ( .B1(n9857), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8142), .ZN(
        n8149) );
  NAND2_X1 U9764 ( .A1(n9477), .A2(n8143), .ZN(n8148) );
  OAI211_X1 U9765 ( .C1(n8146), .C2(n8145), .A(n9849), .B(n8144), .ZN(n8147)
         );
  NAND4_X1 U9766 ( .A1(n8150), .A2(n8149), .A3(n8148), .A4(n8147), .ZN(
        P2_U3249) );
  OAI211_X1 U9767 ( .C1(n8153), .C2(n8152), .A(n9850), .B(n8151), .ZN(n8162)
         );
  NOR2_X1 U9768 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6137), .ZN(n8154) );
  AOI21_X1 U9769 ( .B1(n9857), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8154), .ZN(
        n8161) );
  NAND2_X1 U9770 ( .A1(n9477), .A2(n8155), .ZN(n8160) );
  OAI211_X1 U9771 ( .C1(n8158), .C2(n8157), .A(n9849), .B(n8156), .ZN(n8159)
         );
  NAND4_X1 U9772 ( .A1(n8162), .A2(n8161), .A3(n8160), .A4(n8159), .ZN(
        P2_U3250) );
  OAI211_X1 U9773 ( .C1(n8165), .C2(n8164), .A(n9850), .B(n8163), .ZN(n8174)
         );
  AOI21_X1 U9774 ( .B1(n9857), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8166), .ZN(
        n8173) );
  NAND2_X1 U9775 ( .A1(n9477), .A2(n8167), .ZN(n8172) );
  OAI211_X1 U9776 ( .C1(n8170), .C2(n8169), .A(n9849), .B(n8168), .ZN(n8171)
         );
  NAND4_X1 U9777 ( .A1(n8174), .A2(n8173), .A3(n8172), .A4(n8171), .ZN(
        P2_U3251) );
  OAI211_X1 U9778 ( .C1(n8177), .C2(n8176), .A(n9850), .B(n8175), .ZN(n8186)
         );
  NOR2_X1 U9779 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5255), .ZN(n8178) );
  AOI21_X1 U9780 ( .B1(n9857), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8178), .ZN(
        n8185) );
  NAND2_X1 U9781 ( .A1(n9477), .A2(n8179), .ZN(n8184) );
  OAI211_X1 U9782 ( .C1(n8182), .C2(n8181), .A(n9849), .B(n8180), .ZN(n8183)
         );
  NAND4_X1 U9783 ( .A1(n8186), .A2(n8185), .A3(n8184), .A4(n8183), .ZN(
        P2_U3252) );
  OAI211_X1 U9784 ( .C1(n8189), .C2(n8188), .A(n9850), .B(n8187), .ZN(n8200)
         );
  INV_X1 U9785 ( .A(n8190), .ZN(n8191) );
  AOI21_X1 U9786 ( .B1(n9857), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8191), .ZN(
        n8199) );
  NAND2_X1 U9787 ( .A1(n9477), .A2(n8192), .ZN(n8198) );
  INV_X1 U9788 ( .A(n8193), .ZN(n8194) );
  OAI211_X1 U9789 ( .C1(n8196), .C2(n8195), .A(n9849), .B(n8194), .ZN(n8197)
         );
  NAND4_X1 U9790 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n8197), .ZN(
        P2_U3253) );
  MUX2_X1 U9791 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8201), .S(n8207), .Z(n8203)
         );
  OAI211_X1 U9792 ( .C1(n8204), .C2(n8203), .A(n9850), .B(n8202), .ZN(n8215)
         );
  INV_X1 U9793 ( .A(n8205), .ZN(n8206) );
  AOI21_X1 U9794 ( .B1(n9857), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8206), .ZN(
        n8214) );
  NAND2_X1 U9795 ( .A1(n9477), .A2(n8207), .ZN(n8213) );
  OAI21_X1 U9796 ( .B1(n8210), .B2(n8209), .A(n8208), .ZN(n8211) );
  NAND2_X1 U9797 ( .A1(n9849), .A2(n8211), .ZN(n8212) );
  NAND4_X1 U9798 ( .A1(n8215), .A2(n8214), .A3(n8213), .A4(n8212), .ZN(
        P2_U3257) );
  OAI21_X1 U9799 ( .B1(n8220), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8216), .ZN(
        n8218) );
  INV_X1 U9800 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8217) );
  XNOR2_X1 U9801 ( .A(n8218), .B(n8217), .ZN(n8226) );
  INV_X1 U9802 ( .A(n8226), .ZN(n8225) );
  NOR2_X1 U9803 ( .A1(n8220), .A2(n8219), .ZN(n8221) );
  NOR2_X1 U9804 ( .A1(n8222), .A2(n8221), .ZN(n8223) );
  XNOR2_X1 U9805 ( .A(n8223), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U9806 ( .A1(n8228), .A2(n9850), .ZN(n8224) );
  OAI211_X1 U9807 ( .C1(n9854), .C2(n8225), .A(n8224), .B(n9852), .ZN(n8230)
         );
  OAI22_X1 U9808 ( .A1(n8228), .A2(n8227), .B1(n8226), .B2(n9854), .ZN(n8229)
         );
  MUX2_X1 U9809 ( .A(n8230), .B(n8229), .S(n7687), .Z(n8231) );
  INV_X1 U9810 ( .A(n8231), .ZN(n8233) );
  OAI211_X1 U9811 ( .C1(n9488), .C2(n8234), .A(n8233), .B(n8232), .ZN(P2_U3264) );
  INV_X1 U9812 ( .A(n8523), .ZN(n8447) );
  AOI21_X1 U9813 ( .B1(n8236), .B2(P2_B_REG_SCAN_IN), .A(n9581), .ZN(n8275) );
  NAND2_X1 U9814 ( .A1(n8275), .A2(n8237), .ZN(n8464) );
  NOR2_X1 U9815 ( .A1(n9593), .A2(n8464), .ZN(n8243) );
  AOI21_X1 U9816 ( .B1(n9884), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8243), .ZN(
        n8239) );
  NAND2_X1 U9817 ( .A1(n8459), .A2(n8440), .ZN(n8238) );
  OAI211_X1 U9818 ( .C1(n8461), .C2(n9873), .A(n8239), .B(n8238), .ZN(P2_U3265) );
  OAI21_X1 U9819 ( .B1(n8241), .B2(n8266), .A(n8240), .ZN(n8465) );
  NOR2_X1 U9820 ( .A1(n8241), .A2(n9881), .ZN(n8242) );
  AOI211_X1 U9821 ( .C1(n9593), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8243), .B(
        n8242), .ZN(n8244) );
  OAI21_X1 U9822 ( .B1(n8465), .B2(n9873), .A(n8244), .ZN(P2_U3266) );
  INV_X1 U9823 ( .A(n8508), .ZN(n8403) );
  NAND2_X1 U9824 ( .A1(n8246), .A2(n8245), .ZN(n8247) );
  OR2_X1 U9825 ( .A1(n9568), .A2(n8450), .ZN(n8249) );
  NAND2_X1 U9826 ( .A1(n8523), .A2(n8250), .ZN(n8251) );
  NAND2_X1 U9827 ( .A1(n8252), .A2(n8418), .ZN(n8253) );
  INV_X1 U9828 ( .A(n8513), .ZN(n8414) );
  AOI21_X1 U9829 ( .B1(n8419), .B2(n8403), .A(n8256), .ZN(n8375) );
  OAI22_X1 U9830 ( .A1(n8375), .A2(n8257), .B1(n8397), .B2(n8504), .ZN(n8367)
         );
  NAND2_X1 U9831 ( .A1(n8354), .A2(n8031), .ZN(n8259) );
  XNOR2_X1 U9832 ( .A(n8265), .B(n8264), .ZN(n8470) );
  NOR2_X1 U9833 ( .A1(n4788), .A2(n9881), .ZN(n8271) );
  OAI22_X1 U9834 ( .A1(n8269), .A2(n8436), .B1(n8268), .B2(n9871), .ZN(n8270)
         );
  AOI211_X1 U9835 ( .C1(n8467), .C2(n8456), .A(n8271), .B(n8270), .ZN(n8280)
         );
  OR2_X1 U9836 ( .A1(n8469), .A2(n9593), .ZN(n8279) );
  OAI211_X1 U9837 ( .C1(n8470), .C2(n8458), .A(n8280), .B(n8279), .ZN(P2_U3267) );
  XNOR2_X1 U9838 ( .A(n8282), .B(n8281), .ZN(n8475) );
  OAI211_X1 U9839 ( .C1(n8285), .C2(n8284), .A(n8283), .B(n9868), .ZN(n8289)
         );
  AOI22_X1 U9840 ( .A1(n8287), .A2(n9865), .B1(n8286), .B2(n9864), .ZN(n8288)
         );
  INV_X1 U9841 ( .A(n8474), .ZN(n8295) );
  XNOR2_X1 U9842 ( .A(n8297), .B(n8471), .ZN(n8472) );
  NAND2_X1 U9843 ( .A1(n8472), .A2(n8456), .ZN(n8292) );
  AOI22_X1 U9844 ( .A1(n8290), .A2(n9586), .B1(n9593), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8291) );
  OAI211_X1 U9845 ( .C1(n8293), .C2(n9881), .A(n8292), .B(n8291), .ZN(n8294)
         );
  AOI21_X1 U9846 ( .B1(n8295), .B2(n8436), .A(n8294), .ZN(n8296) );
  OAI21_X1 U9847 ( .B1(n8475), .B2(n8458), .A(n8296), .ZN(P2_U3268) );
  AOI21_X1 U9848 ( .B1(n8476), .B2(n8319), .A(n8297), .ZN(n8477) );
  INV_X1 U9849 ( .A(n8298), .ZN(n8299) );
  AOI22_X1 U9850 ( .A1(n9593), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8299), .B2(
        n9586), .ZN(n8300) );
  OAI21_X1 U9851 ( .B1(n8301), .B2(n9881), .A(n8300), .ZN(n8308) );
  XNOR2_X1 U9852 ( .A(n8303), .B(n8302), .ZN(n8306) );
  AOI222_X1 U9853 ( .A1(n9868), .A2(n8306), .B1(n8305), .B2(n9864), .C1(n8304), 
        .C2(n9865), .ZN(n8479) );
  NOR2_X1 U9854 ( .A1(n8479), .A2(n9593), .ZN(n8307) );
  AOI211_X1 U9855 ( .C1(n8477), .C2(n8456), .A(n8308), .B(n8307), .ZN(n8309)
         );
  OAI21_X1 U9856 ( .B1(n8480), .B2(n8458), .A(n8309), .ZN(P2_U3269) );
  XNOR2_X1 U9857 ( .A(n8310), .B(n8312), .ZN(n8485) );
  AOI22_X1 U9858 ( .A1(n8482), .A2(n8440), .B1(n9593), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8325) );
  INV_X1 U9859 ( .A(n8311), .ZN(n8314) );
  OAI21_X1 U9860 ( .B1(n8314), .B2(n8313), .A(n8312), .ZN(n8316) );
  NAND2_X1 U9861 ( .A1(n8316), .A2(n8315), .ZN(n8318) );
  AOI21_X1 U9862 ( .B1(n8318), .B2(n9868), .A(n8317), .ZN(n8484) );
  AOI21_X1 U9863 ( .B1(n8331), .B2(n8482), .A(n9973), .ZN(n8320) );
  AND2_X1 U9864 ( .A1(n8320), .A2(n8319), .ZN(n8481) );
  NAND2_X1 U9865 ( .A1(n8481), .A2(n7687), .ZN(n8321) );
  OAI211_X1 U9866 ( .C1(n9871), .C2(n8322), .A(n8484), .B(n8321), .ZN(n8323)
         );
  NAND2_X1 U9867 ( .A1(n8323), .A2(n8436), .ZN(n8324) );
  OAI211_X1 U9868 ( .C1(n8485), .C2(n8458), .A(n8325), .B(n8324), .ZN(P2_U3270) );
  XNOR2_X1 U9869 ( .A(n8327), .B(n8326), .ZN(n8490) );
  INV_X1 U9870 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8330) );
  INV_X1 U9871 ( .A(n8328), .ZN(n8329) );
  OAI22_X1 U9872 ( .A1(n9591), .A2(n8330), .B1(n8329), .B2(n9871), .ZN(n8342)
         );
  INV_X1 U9873 ( .A(n8349), .ZN(n8333) );
  INV_X1 U9874 ( .A(n8331), .ZN(n8332) );
  AOI211_X1 U9875 ( .C1(n8488), .C2(n8333), .A(n9973), .B(n8332), .ZN(n8487)
         );
  NAND3_X1 U9876 ( .A1(n8334), .A2(n8336), .A3(n8335), .ZN(n8337) );
  NAND3_X1 U9877 ( .A1(n8311), .A2(n9868), .A3(n8337), .ZN(n8339) );
  NAND2_X1 U9878 ( .A1(n8339), .A2(n8338), .ZN(n8486) );
  AOI21_X1 U9879 ( .B1(n8487), .B2(n7687), .A(n8486), .ZN(n8340) );
  NOR2_X1 U9880 ( .A1(n8340), .A2(n9593), .ZN(n8341) );
  AOI211_X1 U9881 ( .C1(n8440), .C2(n8488), .A(n8342), .B(n8341), .ZN(n8343)
         );
  OAI21_X1 U9882 ( .B1(n8490), .B2(n8458), .A(n8343), .ZN(P2_U3271) );
  AOI21_X1 U9883 ( .B1(n8344), .B2(n8356), .A(n9576), .ZN(n8348) );
  OAI22_X1 U9884 ( .A1(n8346), .A2(n9581), .B1(n8345), .B2(n9579), .ZN(n8347)
         );
  AOI21_X1 U9885 ( .B1(n8348), .B2(n8334), .A(n8347), .ZN(n8494) );
  AOI21_X1 U9886 ( .B1(n8491), .B2(n8350), .A(n8349), .ZN(n8492) );
  INV_X1 U9887 ( .A(n8351), .ZN(n8352) );
  AOI22_X1 U9888 ( .A1(n9593), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8352), .B2(
        n9586), .ZN(n8353) );
  OAI21_X1 U9889 ( .B1(n8354), .B2(n9881), .A(n8353), .ZN(n8360) );
  OAI21_X1 U9890 ( .B1(n8357), .B2(n8356), .A(n8355), .ZN(n8358) );
  INV_X1 U9891 ( .A(n8358), .ZN(n8495) );
  NOR2_X1 U9892 ( .A1(n8495), .A2(n8458), .ZN(n8359) );
  AOI211_X1 U9893 ( .C1(n8492), .C2(n8456), .A(n8360), .B(n8359), .ZN(n8361)
         );
  OAI21_X1 U9894 ( .B1(n9593), .B2(n8494), .A(n8361), .ZN(P2_U3272) );
  XNOR2_X1 U9895 ( .A(n8363), .B(n8362), .ZN(n8365) );
  AOI222_X1 U9896 ( .A1(n9868), .A2(n8365), .B1(n8397), .B2(n9864), .C1(n8364), 
        .C2(n9865), .ZN(n8500) );
  INV_X1 U9897 ( .A(n8502), .ZN(n8368) );
  NAND2_X1 U9898 ( .A1(n8367), .A2(n8366), .ZN(n8496) );
  NAND3_X1 U9899 ( .A1(n8368), .A2(n9878), .A3(n8496), .ZN(n8374) );
  XOR2_X1 U9900 ( .A(n8381), .B(n8497), .Z(n8498) );
  INV_X1 U9901 ( .A(n8497), .ZN(n8371) );
  AOI22_X1 U9902 ( .A1(n9593), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8369), .B2(
        n9586), .ZN(n8370) );
  OAI21_X1 U9903 ( .B1(n8371), .B2(n9881), .A(n8370), .ZN(n8372) );
  AOI21_X1 U9904 ( .B1(n8498), .B2(n8456), .A(n8372), .ZN(n8373) );
  OAI211_X1 U9905 ( .C1(n9593), .C2(n8500), .A(n8374), .B(n8373), .ZN(P2_U3273) );
  XNOR2_X1 U9906 ( .A(n8375), .B(n8376), .ZN(n8507) );
  AOI21_X1 U9907 ( .B1(n8377), .B2(n8376), .A(n9576), .ZN(n8380) );
  AOI21_X1 U9908 ( .B1(n8380), .B2(n8379), .A(n8378), .ZN(n8506) );
  INV_X1 U9909 ( .A(n8506), .ZN(n8393) );
  INV_X1 U9910 ( .A(n8399), .ZN(n8383) );
  INV_X1 U9911 ( .A(n8381), .ZN(n8382) );
  AOI211_X1 U9912 ( .C1(n8504), .C2(n8383), .A(n9973), .B(n8382), .ZN(n8503)
         );
  NAND4_X1 U9913 ( .A1(n8503), .A2(n8386), .A3(n8385), .A4(n8384), .ZN(n8390)
         );
  INV_X1 U9914 ( .A(n8387), .ZN(n8388) );
  AOI22_X1 U9915 ( .A1(n9593), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8388), .B2(
        n9586), .ZN(n8389) );
  OAI211_X1 U9916 ( .C1(n8391), .C2(n9881), .A(n8390), .B(n8389), .ZN(n8392)
         );
  AOI21_X1 U9917 ( .B1(n8393), .B2(n8436), .A(n8392), .ZN(n8394) );
  OAI21_X1 U9918 ( .B1(n8507), .B2(n8458), .A(n8394), .ZN(P2_U3274) );
  XNOR2_X1 U9919 ( .A(n8395), .B(n8404), .ZN(n8398) );
  AOI222_X1 U9920 ( .A1(n9868), .A2(n8398), .B1(n8397), .B2(n9865), .C1(n8396), 
        .C2(n9864), .ZN(n8511) );
  AOI21_X1 U9921 ( .B1(n8508), .B2(n8410), .A(n8399), .ZN(n8509) );
  INV_X1 U9922 ( .A(n8400), .ZN(n8401) );
  AOI22_X1 U9923 ( .A1(n9593), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8401), .B2(
        n9586), .ZN(n8402) );
  OAI21_X1 U9924 ( .B1(n8403), .B2(n9881), .A(n8402), .ZN(n8407) );
  XNOR2_X1 U9925 ( .A(n8405), .B(n8404), .ZN(n8512) );
  NOR2_X1 U9926 ( .A1(n8512), .A2(n8458), .ZN(n8406) );
  AOI211_X1 U9927 ( .C1(n8509), .C2(n8456), .A(n8407), .B(n8406), .ZN(n8408)
         );
  OAI21_X1 U9928 ( .B1(n9884), .B2(n8511), .A(n8408), .ZN(P2_U3275) );
  XNOR2_X1 U9929 ( .A(n8409), .B(n7653), .ZN(n8517) );
  AOI21_X1 U9930 ( .B1(n8513), .B2(n8434), .A(n4596), .ZN(n8514) );
  INV_X1 U9931 ( .A(n8411), .ZN(n8412) );
  AOI22_X1 U9932 ( .A1(n9593), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8412), .B2(
        n9586), .ZN(n8413) );
  OAI21_X1 U9933 ( .B1(n8414), .B2(n9881), .A(n8413), .ZN(n8423) );
  AOI21_X1 U9934 ( .B1(n8416), .B2(n8415), .A(n9576), .ZN(n8421) );
  OAI22_X1 U9935 ( .A1(n8419), .A2(n9581), .B1(n8418), .B2(n9579), .ZN(n8420)
         );
  AOI21_X1 U9936 ( .B1(n8421), .B2(n8417), .A(n8420), .ZN(n8516) );
  NOR2_X1 U9937 ( .A1(n8516), .A2(n9593), .ZN(n8422) );
  AOI211_X1 U9938 ( .C1(n8514), .C2(n8456), .A(n8423), .B(n8422), .ZN(n8424)
         );
  OAI21_X1 U9939 ( .B1(n8458), .B2(n8517), .A(n8424), .ZN(P2_U3276) );
  XNOR2_X1 U9940 ( .A(n8425), .B(n8427), .ZN(n8522) );
  INV_X1 U9941 ( .A(n8426), .ZN(n8429) );
  OAI21_X1 U9942 ( .B1(n8429), .B2(n8428), .A(n8427), .ZN(n8431) );
  AOI21_X1 U9943 ( .B1(n8431), .B2(n8430), .A(n9576), .ZN(n8433) );
  NOR2_X1 U9944 ( .A1(n8433), .A2(n8432), .ZN(n8521) );
  AOI211_X1 U9945 ( .C1(n8519), .C2(n8444), .A(n9973), .B(n4789), .ZN(n8518)
         );
  NAND2_X1 U9946 ( .A1(n8518), .A2(n7687), .ZN(n8435) );
  OAI211_X1 U9947 ( .C1(n8522), .C2(n9565), .A(n8521), .B(n8435), .ZN(n8437)
         );
  NAND2_X1 U9948 ( .A1(n8437), .A2(n8436), .ZN(n8442) );
  INV_X1 U9949 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10230) );
  OAI22_X1 U9950 ( .A1(n9591), .A2(n10230), .B1(n8438), .B2(n9871), .ZN(n8439)
         );
  AOI21_X1 U9951 ( .B1(n8519), .B2(n8440), .A(n8439), .ZN(n8441) );
  OAI211_X1 U9952 ( .C1(n8522), .C2(n9584), .A(n8442), .B(n8441), .ZN(P2_U3277) );
  XNOR2_X1 U9953 ( .A(n8443), .B(n8449), .ZN(n8527) );
  AOI21_X1 U9954 ( .B1(n8523), .B2(n4491), .A(n4600), .ZN(n8524) );
  AOI22_X1 U9955 ( .A1(n9593), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8445), .B2(
        n9586), .ZN(n8446) );
  OAI21_X1 U9956 ( .B1(n8447), .B2(n9881), .A(n8446), .ZN(n8455) );
  OAI211_X1 U9957 ( .C1(n8449), .C2(n8448), .A(n8426), .B(n9868), .ZN(n8453)
         );
  AOI22_X1 U9958 ( .A1(n8451), .A2(n9865), .B1(n9864), .B2(n8450), .ZN(n8452)
         );
  NOR2_X1 U9959 ( .A1(n8526), .A2(n9593), .ZN(n8454) );
  AOI211_X1 U9960 ( .C1(n8524), .C2(n8456), .A(n8455), .B(n8454), .ZN(n8457)
         );
  OAI21_X1 U9961 ( .B1(n8527), .B2(n8458), .A(n8457), .ZN(P2_U3278) );
  NAND2_X1 U9962 ( .A1(n8459), .A2(n9962), .ZN(n8460) );
  OAI211_X1 U9963 ( .C1(n8461), .C2(n9973), .A(n8464), .B(n8460), .ZN(n8528)
         );
  MUX2_X1 U9964 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8528), .S(n9995), .Z(
        P2_U3551) );
  NAND2_X1 U9965 ( .A1(n8462), .A2(n9962), .ZN(n8463) );
  OAI211_X1 U9966 ( .C1(n8465), .C2(n9973), .A(n8464), .B(n8463), .ZN(n8529)
         );
  MUX2_X1 U9967 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8529), .S(n9995), .Z(
        P2_U3550) );
  OAI211_X1 U9968 ( .C1(n8470), .C2(n9966), .A(n8469), .B(n8468), .ZN(n8530)
         );
  MUX2_X1 U9969 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8530), .S(n9995), .Z(
        P2_U3549) );
  AOI22_X1 U9970 ( .A1(n8472), .A2(n9963), .B1(n9962), .B2(n8471), .ZN(n8473)
         );
  OAI211_X1 U9971 ( .C1(n8475), .C2(n9966), .A(n8474), .B(n8473), .ZN(n8531)
         );
  MUX2_X1 U9972 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8531), .S(n9995), .Z(
        P2_U3548) );
  AOI22_X1 U9973 ( .A1(n8477), .A2(n9963), .B1(n9962), .B2(n8476), .ZN(n8478)
         );
  MUX2_X1 U9974 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8532), .S(n9995), .Z(
        P2_U3547) );
  AOI21_X1 U9975 ( .B1(n9962), .B2(n8482), .A(n8481), .ZN(n8483) );
  OAI211_X1 U9976 ( .C1(n8485), .C2(n9966), .A(n8484), .B(n8483), .ZN(n8533)
         );
  MUX2_X1 U9977 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8533), .S(n9995), .Z(
        P2_U3546) );
  AOI211_X1 U9978 ( .C1(n9962), .C2(n8488), .A(n8487), .B(n8486), .ZN(n8489)
         );
  OAI21_X1 U9979 ( .B1(n8490), .B2(n9966), .A(n8489), .ZN(n8534) );
  MUX2_X1 U9980 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8534), .S(n9995), .Z(
        P2_U3545) );
  AOI22_X1 U9981 ( .A1(n8492), .A2(n9963), .B1(n9962), .B2(n8491), .ZN(n8493)
         );
  OAI211_X1 U9982 ( .C1(n8495), .C2(n9966), .A(n8494), .B(n8493), .ZN(n8535)
         );
  MUX2_X1 U9983 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8535), .S(n9995), .Z(
        P2_U3544) );
  INV_X1 U9984 ( .A(n9966), .ZN(n9978) );
  NAND2_X1 U9985 ( .A1(n8496), .A2(n9978), .ZN(n8501) );
  AOI22_X1 U9986 ( .A1(n8498), .A2(n9963), .B1(n9962), .B2(n8497), .ZN(n8499)
         );
  OAI211_X1 U9987 ( .C1(n8502), .C2(n8501), .A(n8500), .B(n8499), .ZN(n8536)
         );
  MUX2_X1 U9988 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8536), .S(n9995), .Z(
        P2_U3543) );
  AOI21_X1 U9989 ( .B1(n9962), .B2(n8504), .A(n8503), .ZN(n8505) );
  OAI211_X1 U9990 ( .C1(n8507), .C2(n9966), .A(n8506), .B(n8505), .ZN(n8537)
         );
  MUX2_X1 U9991 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8537), .S(n9995), .Z(
        P2_U3542) );
  AOI22_X1 U9992 ( .A1(n8509), .A2(n9963), .B1(n9962), .B2(n8508), .ZN(n8510)
         );
  OAI211_X1 U9993 ( .C1(n9966), .C2(n8512), .A(n8511), .B(n8510), .ZN(n8538)
         );
  MUX2_X1 U9994 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8538), .S(n9995), .Z(
        P2_U3541) );
  AOI22_X1 U9995 ( .A1(n8514), .A2(n9963), .B1(n9962), .B2(n8513), .ZN(n8515)
         );
  OAI211_X1 U9996 ( .C1(n8517), .C2(n9966), .A(n8516), .B(n8515), .ZN(n8539)
         );
  MUX2_X1 U9997 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8539), .S(n9995), .Z(
        P2_U3540) );
  AOI21_X1 U9998 ( .B1(n9962), .B2(n8519), .A(n8518), .ZN(n8520) );
  OAI211_X1 U9999 ( .C1(n9966), .C2(n8522), .A(n8521), .B(n8520), .ZN(n8540)
         );
  MUX2_X1 U10000 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8540), .S(n9995), .Z(
        P2_U3539) );
  AOI22_X1 U10001 ( .A1(n8524), .A2(n9963), .B1(n9962), .B2(n8523), .ZN(n8525)
         );
  OAI211_X1 U10002 ( .C1(n9966), .C2(n8527), .A(n8526), .B(n8525), .ZN(n8541)
         );
  MUX2_X1 U10003 ( .A(n8541), .B(P2_REG1_REG_18__SCAN_IN), .S(n9993), .Z(
        P2_U3538) );
  MUX2_X1 U10004 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8528), .S(n9979), .Z(
        P2_U3519) );
  MUX2_X1 U10005 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8529), .S(n9979), .Z(
        P2_U3518) );
  MUX2_X1 U10006 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8530), .S(n9979), .Z(
        P2_U3517) );
  MUX2_X1 U10007 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8531), .S(n9979), .Z(
        P2_U3516) );
  MUX2_X1 U10008 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8533), .S(n9979), .Z(
        P2_U3514) );
  MUX2_X1 U10009 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8534), .S(n9979), .Z(
        P2_U3513) );
  MUX2_X1 U10010 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8535), .S(n9979), .Z(
        P2_U3512) );
  MUX2_X1 U10011 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8536), .S(n9979), .Z(
        P2_U3511) );
  MUX2_X1 U10012 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8537), .S(n9979), .Z(
        P2_U3510) );
  MUX2_X1 U10013 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8538), .S(n9979), .Z(
        P2_U3509) );
  MUX2_X1 U10014 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8539), .S(n9979), .Z(
        P2_U3508) );
  MUX2_X1 U10015 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8540), .S(n9979), .Z(
        P2_U3507) );
  MUX2_X1 U10016 ( .A(n8541), .B(P2_REG0_REG_18__SCAN_IN), .S(n4579), .Z(
        P2_U3505) );
  INV_X1 U10017 ( .A(n8789), .ZN(n9460) );
  NOR4_X1 U10018 ( .A1(n5081), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8542), .A4(
        P2_U3152), .ZN(n8543) );
  AOI21_X1 U10019 ( .B1(n8544), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8543), .ZN(
        n8545) );
  OAI21_X1 U10020 ( .B1(n9460), .B2(n8548), .A(n8545), .ZN(P2_U3327) );
  INV_X1 U10021 ( .A(n8729), .ZN(n9468) );
  OAI222_X1 U10022 ( .A1(n8548), .A2(n9468), .B1(P2_U3152), .B2(n8547), .C1(
        n10184), .C2(n8546), .ZN(P2_U3329) );
  INV_X1 U10023 ( .A(n8549), .ZN(n8550) );
  MUX2_X1 U10024 ( .A(n8550), .B(n9861), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10025 ( .A(n8552), .B(n8551), .ZN(n8553) );
  XNOR2_X1 U10026 ( .A(n8554), .B(n8553), .ZN(n8559) );
  INV_X1 U10027 ( .A(n8715), .ZN(n8651) );
  OAI22_X1 U10028 ( .A1(n9149), .A2(n8710), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10138), .ZN(n8556) );
  NOR2_X1 U10029 ( .A1(n9150), .A2(n8648), .ZN(n8555) );
  AOI211_X1 U10030 ( .C1(n9156), .C2(n8651), .A(n8556), .B(n8555), .ZN(n8558)
         );
  NAND2_X1 U10031 ( .A1(n9356), .A2(n8717), .ZN(n8557) );
  OAI211_X1 U10032 ( .C1(n8559), .C2(n8719), .A(n8558), .B(n8557), .ZN(
        P1_U3212) );
  NAND2_X1 U10033 ( .A1(n4547), .A2(n8560), .ZN(n8561) );
  XOR2_X1 U10034 ( .A(n8562), .B(n8561), .Z(n8569) );
  OAI21_X1 U10035 ( .B1(n8710), .B2(n8761), .A(n8563), .ZN(n8564) );
  AOI21_X1 U10036 ( .B1(n8713), .B2(n9014), .A(n8564), .ZN(n8565) );
  OAI21_X1 U10037 ( .B1(n8715), .B2(n8566), .A(n8565), .ZN(n8567) );
  AOI21_X1 U10038 ( .B1(n9426), .B2(n8717), .A(n8567), .ZN(n8568) );
  OAI21_X1 U10039 ( .B1(n8569), .B2(n8719), .A(n8568), .ZN(P1_U3213) );
  AOI21_X1 U10040 ( .B1(n8571), .B2(n8642), .A(n8570), .ZN(n8572) );
  AOI21_X1 U10041 ( .B1(n4496), .B2(n8642), .A(n8572), .ZN(n8577) );
  NOR2_X1 U10042 ( .A1(n8715), .A2(n9206), .ZN(n8575) );
  AOI22_X1 U10043 ( .A1(n9216), .A2(n8713), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8573) );
  OAI21_X1 U10044 ( .B1(n8592), .B2(n8710), .A(n8573), .ZN(n8574) );
  AOI211_X1 U10045 ( .C1(n9375), .C2(n8717), .A(n8575), .B(n8574), .ZN(n8576)
         );
  OAI21_X1 U10046 ( .B1(n8577), .B2(n8719), .A(n8576), .ZN(P1_U3214) );
  OAI21_X1 U10047 ( .B1(n8580), .B2(n8579), .A(n8578), .ZN(n8581) );
  NAND2_X1 U10048 ( .A1(n8581), .A2(n8645), .ZN(n8586) );
  INV_X1 U10049 ( .A(n8582), .ZN(n9270) );
  AOI22_X1 U10050 ( .A1(n8713), .A2(n9277), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3084), .ZN(n8583) );
  OAI21_X1 U10051 ( .B1(n9312), .B2(n8710), .A(n8583), .ZN(n8584) );
  AOI21_X1 U10052 ( .B1(n9270), .B2(n8651), .A(n8584), .ZN(n8585) );
  OAI211_X1 U10053 ( .C1(n9272), .C2(n8654), .A(n8586), .B(n8585), .ZN(
        P1_U3217) );
  XNOR2_X1 U10054 ( .A(n8587), .B(n8588), .ZN(n8589) );
  NAND2_X1 U10055 ( .A1(n8589), .A2(n8645), .ZN(n8596) );
  OAI22_X1 U10056 ( .A1(n8710), .A2(n8591), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8590), .ZN(n8594) );
  NOR2_X1 U10057 ( .A1(n8648), .A2(n8592), .ZN(n8593) );
  AOI211_X1 U10058 ( .C1(n9244), .C2(n8651), .A(n8594), .B(n8593), .ZN(n8595)
         );
  OAI211_X1 U10059 ( .C1(n8597), .C2(n8654), .A(n8596), .B(n8595), .ZN(
        P1_U3221) );
  NOR2_X1 U10060 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8598), .ZN(n9044) );
  AOI21_X1 U10061 ( .B1(n8713), .B2(n9015), .A(n9044), .ZN(n8601) );
  OR2_X1 U10062 ( .A1(n8710), .A2(n8599), .ZN(n8600) );
  OAI211_X1 U10063 ( .C1(n8715), .C2(n8602), .A(n8601), .B(n8600), .ZN(n8611)
         );
  OR2_X1 U10064 ( .A1(n8603), .A2(n8681), .ZN(n8679) );
  NAND2_X1 U10065 ( .A1(n8679), .A2(n8604), .ZN(n8608) );
  XNOR2_X1 U10066 ( .A(n8606), .B(n8605), .ZN(n8607) );
  XNOR2_X1 U10067 ( .A(n8608), .B(n8607), .ZN(n8609) );
  NOR2_X1 U10068 ( .A1(n8609), .A2(n8719), .ZN(n8610) );
  AOI211_X1 U10069 ( .C1(n9634), .C2(n8692), .A(n8611), .B(n8610), .ZN(n8612)
         );
  INV_X1 U10070 ( .A(n8612), .ZN(P1_U3222) );
  OAI21_X1 U10071 ( .B1(n8615), .B2(n8614), .A(n8613), .ZN(n8616) );
  NAND2_X1 U10072 ( .A1(n8616), .A2(n8645), .ZN(n8621) );
  AOI22_X1 U10073 ( .A1(n9184), .A2(n8713), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8617) );
  OAI21_X1 U10074 ( .B1(n8618), .B2(n8710), .A(n8617), .ZN(n8619) );
  AOI21_X1 U10075 ( .B1(n9179), .B2(n8651), .A(n8619), .ZN(n8620) );
  OAI211_X1 U10076 ( .C1(n9181), .C2(n8654), .A(n8621), .B(n8620), .ZN(
        P1_U3223) );
  NAND3_X1 U10077 ( .A1(n8623), .A2(n8622), .A3(n4547), .ZN(n8704) );
  AOI21_X1 U10078 ( .B1(n8623), .B2(n4547), .A(n8622), .ZN(n8705) );
  AOI21_X1 U10079 ( .B1(n8707), .B2(n8704), .A(n8705), .ZN(n8627) );
  XNOR2_X1 U10080 ( .A(n8625), .B(n8624), .ZN(n8626) );
  XNOR2_X1 U10081 ( .A(n8627), .B(n8626), .ZN(n8634) );
  NOR2_X1 U10082 ( .A1(n8715), .A2(n8628), .ZN(n8632) );
  AOI22_X1 U10083 ( .A1(n8713), .A2(n9283), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8629) );
  OAI21_X1 U10084 ( .B1(n8630), .B2(n8710), .A(n8629), .ZN(n8631) );
  AOI211_X1 U10085 ( .C1(n9416), .C2(n8692), .A(n8632), .B(n8631), .ZN(n8633)
         );
  OAI21_X1 U10086 ( .B1(n8634), .B2(n8719), .A(n8633), .ZN(P1_U3224) );
  XOR2_X1 U10087 ( .A(n8636), .B(n8635), .Z(n8641) );
  NOR2_X1 U10088 ( .A1(n8715), .A2(n9303), .ZN(n8639) );
  AOI22_X1 U10089 ( .A1(n8713), .A2(n9276), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n8637) );
  OAI21_X1 U10090 ( .B1(n9311), .B2(n8710), .A(n8637), .ZN(n8638) );
  AOI211_X1 U10091 ( .C1(n9411), .C2(n8692), .A(n8639), .B(n8638), .ZN(n8640)
         );
  OAI21_X1 U10092 ( .B1(n8641), .B2(n8719), .A(n8640), .ZN(P1_U3226) );
  INV_X1 U10093 ( .A(n9372), .ZN(n8655) );
  INV_X1 U10094 ( .A(n8642), .ZN(n8644) );
  NOR3_X1 U10095 ( .A1(n4496), .A2(n8644), .A3(n8643), .ZN(n8646) );
  OAI21_X1 U10096 ( .B1(n8646), .B2(n4530), .A(n8645), .ZN(n8653) );
  OAI22_X1 U10097 ( .A1(n9194), .A2(n8710), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8647), .ZN(n8650) );
  NOR2_X1 U10098 ( .A1(n9195), .A2(n8648), .ZN(n8649) );
  AOI211_X1 U10099 ( .C1(n9197), .C2(n8651), .A(n8650), .B(n8649), .ZN(n8652)
         );
  OAI211_X1 U10100 ( .C1(n8655), .C2(n8654), .A(n8653), .B(n8652), .ZN(
        P1_U3227) );
  NAND2_X1 U10101 ( .A1(n8657), .A2(n8656), .ZN(n8658) );
  XNOR2_X1 U10102 ( .A(n8659), .B(n8658), .ZN(n8664) );
  NOR2_X1 U10103 ( .A1(n8715), .A2(n9256), .ZN(n8662) );
  AOI22_X1 U10104 ( .A1(n8713), .A2(n9231), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8660) );
  OAI21_X1 U10105 ( .B1(n9263), .B2(n8710), .A(n8660), .ZN(n8661) );
  AOI211_X1 U10106 ( .C1(n9394), .C2(n8717), .A(n8662), .B(n8661), .ZN(n8663)
         );
  OAI21_X1 U10107 ( .B1(n8664), .B2(n8719), .A(n8663), .ZN(P1_U3231) );
  NAND2_X1 U10108 ( .A1(n8666), .A2(n8665), .ZN(n8667) );
  XOR2_X1 U10109 ( .A(n8668), .B(n8667), .Z(n8674) );
  OAI22_X1 U10110 ( .A1(n8710), .A2(n9264), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8669), .ZN(n8670) );
  AOI21_X1 U10111 ( .B1(n8713), .B2(n9230), .A(n8670), .ZN(n8671) );
  OAI21_X1 U10112 ( .B1(n8715), .B2(n9224), .A(n8671), .ZN(n8672) );
  AOI21_X1 U10113 ( .B1(n9380), .B2(n8717), .A(n8672), .ZN(n8673) );
  OAI21_X1 U10114 ( .B1(n8674), .B2(n8719), .A(n8673), .ZN(P1_U3233) );
  NOR2_X1 U10115 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7057), .ZN(n9723) );
  AOI21_X1 U10116 ( .B1(n8713), .B2(n9016), .A(n9723), .ZN(n8677) );
  OR2_X1 U10117 ( .A1(n8710), .A2(n8675), .ZN(n8676) );
  OAI211_X1 U10118 ( .C1(n8715), .C2(n8678), .A(n8677), .B(n8676), .ZN(n8683)
         );
  INV_X1 U10119 ( .A(n8679), .ZN(n8680) );
  AOI211_X1 U10120 ( .C1(n8681), .C2(n8603), .A(n8719), .B(n8680), .ZN(n8682)
         );
  AOI211_X1 U10121 ( .C1(n9431), .C2(n8692), .A(n8683), .B(n8682), .ZN(n8684)
         );
  INV_X1 U10122 ( .A(n8684), .ZN(P1_U3234) );
  NAND2_X1 U10123 ( .A1(n4549), .A2(n8685), .ZN(n8686) );
  XOR2_X1 U10124 ( .A(n8687), .B(n8686), .Z(n8694) );
  NOR2_X1 U10125 ( .A1(n8715), .A2(n9293), .ZN(n8691) );
  NAND2_X1 U10126 ( .A1(n8713), .A2(n9284), .ZN(n8688) );
  NAND2_X1 U10127 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9743) );
  OAI211_X1 U10128 ( .C1(n8710), .C2(n8689), .A(n8688), .B(n9743), .ZN(n8690)
         );
  AOI211_X1 U10129 ( .C1(n9404), .C2(n8692), .A(n8691), .B(n8690), .ZN(n8693)
         );
  OAI21_X1 U10130 ( .B1(n8694), .B2(n8719), .A(n8693), .ZN(P1_U3236) );
  NAND2_X1 U10131 ( .A1(n8696), .A2(n8695), .ZN(n8697) );
  XNOR2_X1 U10132 ( .A(n8698), .B(n8697), .ZN(n8703) );
  NOR2_X1 U10133 ( .A1(n8715), .A2(n9170), .ZN(n8701) );
  AOI22_X1 U10134 ( .A1(n9012), .A2(n8713), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8699) );
  OAI21_X1 U10135 ( .B1(n9195), .B2(n8710), .A(n8699), .ZN(n8700) );
  AOI211_X1 U10136 ( .C1(n9362), .C2(n8717), .A(n8701), .B(n8700), .ZN(n8702)
         );
  OAI21_X1 U10137 ( .B1(n8703), .B2(n8719), .A(n8702), .ZN(P1_U3238) );
  INV_X1 U10138 ( .A(n8704), .ZN(n8706) );
  NOR2_X1 U10139 ( .A1(n8706), .A2(n8705), .ZN(n8708) );
  XNOR2_X1 U10140 ( .A(n8708), .B(n8707), .ZN(n8720) );
  NOR2_X1 U10141 ( .A1(n8710), .A2(n8709), .ZN(n8711) );
  AOI211_X1 U10142 ( .C1(n8713), .C2(n9329), .A(n8712), .B(n8711), .ZN(n8714)
         );
  OAI21_X1 U10143 ( .B1(n8715), .B2(n9318), .A(n8714), .ZN(n8716) );
  AOI21_X1 U10144 ( .B1(n9419), .B2(n8717), .A(n8716), .ZN(n8718) );
  OAI21_X1 U10145 ( .B1(n8720), .B2(n8719), .A(n8718), .ZN(P1_U3239) );
  NAND2_X1 U10146 ( .A1(n8721), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8725) );
  INV_X1 U10147 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8722) );
  OR2_X1 U10148 ( .A1(n6273), .A2(n8722), .ZN(n8724) );
  INV_X1 U10149 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10275) );
  OR2_X1 U10150 ( .A1(n6274), .A2(n10275), .ZN(n8723) );
  AND3_X1 U10151 ( .A1(n8725), .A2(n8724), .A3(n8723), .ZN(n9132) );
  NAND2_X1 U10152 ( .A1(n8726), .A2(n4475), .ZN(n8728) );
  NAND2_X1 U10153 ( .A1(n8730), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U10154 ( .A1(n8729), .A2(n4475), .ZN(n8732) );
  NAND2_X1 U10155 ( .A1(n8730), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U10156 ( .A1(n9344), .A2(n7632), .ZN(n8987) );
  INV_X1 U10157 ( .A(n8987), .ZN(n8786) );
  INV_X1 U10158 ( .A(n8880), .ZN(n8733) );
  NAND2_X1 U10159 ( .A1(n8895), .A2(n8733), .ZN(n8734) );
  NAND3_X1 U10160 ( .A1(n9128), .A2(n8881), .A3(n8734), .ZN(n8781) );
  INV_X1 U10161 ( .A(n8893), .ZN(n8735) );
  NAND2_X1 U10162 ( .A1(n8877), .A2(n8735), .ZN(n8775) );
  NAND2_X1 U10163 ( .A1(n8931), .A2(n8736), .ZN(n8867) );
  AND2_X1 U10164 ( .A1(n8886), .A2(n8933), .ZN(n8737) );
  OR2_X1 U10165 ( .A1(n8867), .A2(n8737), .ZN(n8885) );
  NAND2_X1 U10166 ( .A1(n8816), .A2(n4478), .ZN(n8825) );
  NAND2_X1 U10167 ( .A1(n8738), .A2(n8812), .ZN(n8739) );
  NAND2_X1 U10168 ( .A1(n8739), .A2(n8815), .ZN(n8807) );
  NOR2_X1 U10169 ( .A1(n8825), .A2(n8807), .ZN(n8758) );
  NAND3_X1 U10170 ( .A1(n8888), .A2(n8758), .A3(n8863), .ZN(n8740) );
  OR3_X1 U10171 ( .A1(n8775), .A2(n8885), .A3(n8740), .ZN(n8741) );
  OR2_X1 U10172 ( .A1(n8781), .A2(n8741), .ZN(n8986) );
  INV_X1 U10173 ( .A(n8986), .ZN(n8784) );
  AND2_X1 U10174 ( .A1(n8848), .A2(n8844), .ZN(n8742) );
  NAND2_X1 U10175 ( .A1(n8849), .A2(n8742), .ZN(n8985) );
  INV_X1 U10176 ( .A(n8743), .ZN(n8744) );
  AND2_X1 U10177 ( .A1(n8829), .A2(n8744), .ZN(n8983) );
  INV_X1 U10178 ( .A(n8983), .ZN(n8757) );
  AOI21_X1 U10179 ( .B1(n9024), .B2(n9802), .A(n8992), .ZN(n8745) );
  NAND3_X1 U10180 ( .A1(n8747), .A2(n8746), .A3(n8745), .ZN(n8748) );
  NAND3_X1 U10181 ( .A1(n8749), .A2(n8971), .A3(n8748), .ZN(n8752) );
  AND2_X1 U10182 ( .A1(n8750), .A2(n8969), .ZN(n8978) );
  INV_X1 U10183 ( .A(n8972), .ZN(n8751) );
  AOI21_X1 U10184 ( .B1(n8752), .B2(n8978), .A(n8751), .ZN(n8755) );
  AND2_X1 U10185 ( .A1(n8753), .A2(n8800), .ZN(n8977) );
  INV_X1 U10186 ( .A(n8977), .ZN(n8754) );
  OAI211_X1 U10187 ( .C1(n8755), .C2(n8754), .A(n8801), .B(n8981), .ZN(n8756)
         );
  NOR4_X1 U10188 ( .A1(n8985), .A2(n4642), .A3(n8757), .A4(n8756), .ZN(n8783)
         );
  INV_X1 U10189 ( .A(n8892), .ZN(n8777) );
  INV_X1 U10190 ( .A(n8885), .ZN(n8771) );
  INV_X1 U10191 ( .A(n8985), .ZN(n8768) );
  AND2_X1 U10192 ( .A1(n8818), .A2(n8810), .ZN(n8805) );
  INV_X1 U10193 ( .A(n8758), .ZN(n8764) );
  INV_X1 U10194 ( .A(n8816), .ZN(n8759) );
  OR2_X1 U10195 ( .A1(n8760), .A2(n8759), .ZN(n8763) );
  OR2_X1 U10196 ( .A1(n8762), .A2(n8761), .ZN(n8827) );
  AND2_X1 U10197 ( .A1(n8763), .A2(n8827), .ZN(n8833) );
  OAI21_X1 U10198 ( .B1(n8805), .B2(n8764), .A(n8833), .ZN(n8765) );
  AOI21_X1 U10199 ( .B1(n8765), .B2(n8983), .A(n9324), .ZN(n8766) );
  OAI211_X1 U10200 ( .C1(n8766), .C2(n4642), .A(n8839), .B(n8845), .ZN(n8767)
         );
  NAND4_X1 U10201 ( .A1(n8771), .A2(n8768), .A3(n8863), .A4(n8767), .ZN(n8773)
         );
  AND2_X1 U10202 ( .A1(n8860), .A2(n8843), .ZN(n8850) );
  NAND2_X1 U10203 ( .A1(n8863), .A2(n8849), .ZN(n8856) );
  INV_X1 U10204 ( .A(n8861), .ZN(n8769) );
  NOR2_X1 U10205 ( .A1(n8934), .A2(n8769), .ZN(n8858) );
  OAI211_X1 U10206 ( .C1(n8850), .C2(n8856), .A(n8858), .B(n8886), .ZN(n8770)
         );
  NAND2_X1 U10207 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  NAND3_X1 U10208 ( .A1(n8773), .A2(n8772), .A3(n8932), .ZN(n8774) );
  AND2_X1 U10209 ( .A1(n8774), .A2(n8888), .ZN(n8776) );
  INV_X1 U10210 ( .A(n8775), .ZN(n8875) );
  OAI21_X1 U10211 ( .B1(n8777), .B2(n8776), .A(n8875), .ZN(n8778) );
  AND3_X1 U10212 ( .A1(n8895), .A2(n8779), .A3(n8778), .ZN(n8780) );
  OR2_X1 U10213 ( .A1(n8781), .A2(n8780), .ZN(n8782) );
  NAND3_X1 U10214 ( .A1(n8782), .A2(n8914), .A3(n8896), .ZN(n8989) );
  AOI21_X1 U10215 ( .B1(n8784), .B2(n8783), .A(n8989), .ZN(n8785) );
  AOI211_X1 U10216 ( .C1(n9132), .C2(n9340), .A(n8786), .B(n8785), .ZN(n8788)
         );
  OR2_X1 U10217 ( .A1(n9340), .A2(n9132), .ZN(n8918) );
  INV_X1 U10218 ( .A(n8918), .ZN(n8787) );
  NOR2_X1 U10219 ( .A1(n8788), .A2(n8787), .ZN(n8793) );
  NAND2_X1 U10220 ( .A1(n8789), .A2(n4475), .ZN(n8791) );
  NAND2_X1 U10221 ( .A1(n8730), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8790) );
  INV_X1 U10222 ( .A(n8917), .ZN(n9115) );
  AOI21_X1 U10223 ( .B1(n8793), .B2(n8962), .A(n8991), .ZN(n8794) );
  XNOR2_X1 U10224 ( .A(n8794), .B(n4473), .ZN(n9002) );
  NOR2_X1 U10225 ( .A1(n8795), .A2(n8992), .ZN(n8796) );
  INV_X1 U10226 ( .A(n8991), .ZN(n8923) );
  AND2_X1 U10227 ( .A1(n8796), .A2(n8923), .ZN(n9000) );
  INV_X1 U10228 ( .A(n8973), .ZN(n8797) );
  OR2_X1 U10229 ( .A1(n8798), .A2(n8797), .ZN(n8802) );
  AND2_X1 U10230 ( .A1(n8800), .A2(n8799), .ZN(n8975) );
  AOI21_X1 U10231 ( .B1(n8802), .B2(n8975), .A(n4764), .ZN(n8803) );
  INV_X1 U10232 ( .A(n8921), .ZN(n8901) );
  NAND2_X1 U10233 ( .A1(n8811), .A2(n8981), .ZN(n8806) );
  NAND2_X1 U10234 ( .A1(n8806), .A2(n8805), .ZN(n8809) );
  INV_X1 U10235 ( .A(n8807), .ZN(n8808) );
  NAND2_X1 U10236 ( .A1(n8809), .A2(n8808), .ZN(n8820) );
  OAI21_X1 U10237 ( .B1(n8811), .B2(n4762), .A(n8810), .ZN(n8814) );
  INV_X1 U10238 ( .A(n8812), .ZN(n8813) );
  NAND2_X1 U10239 ( .A1(n8814), .A2(n8813), .ZN(n8819) );
  NAND2_X1 U10240 ( .A1(n8816), .A2(n8815), .ZN(n8817) );
  AND2_X1 U10241 ( .A1(n8824), .A2(n8821), .ZN(n8822) );
  NAND2_X1 U10242 ( .A1(n8823), .A2(n8822), .ZN(n8834) );
  NAND2_X1 U10243 ( .A1(n8825), .A2(n8824), .ZN(n8826) );
  NAND3_X1 U10244 ( .A1(n8834), .A2(n8983), .A3(n8826), .ZN(n8832) );
  NAND2_X1 U10245 ( .A1(n8828), .A2(n8827), .ZN(n8830) );
  NAND2_X1 U10246 ( .A1(n8830), .A2(n8829), .ZN(n8831) );
  NAND2_X1 U10247 ( .A1(n8832), .A2(n8831), .ZN(n8837) );
  NAND2_X1 U10248 ( .A1(n8834), .A2(n8833), .ZN(n8835) );
  AOI21_X1 U10249 ( .B1(n8835), .B2(n8983), .A(n9324), .ZN(n8836) );
  INV_X1 U10250 ( .A(n8956), .ZN(n8841) );
  MUX2_X1 U10251 ( .A(n8839), .B(n8838), .S(n8901), .Z(n8840) );
  OAI211_X1 U10252 ( .C1(n8842), .C2(n9323), .A(n8841), .B(n8840), .ZN(n8847)
         );
  NAND2_X1 U10253 ( .A1(n8843), .A2(n8848), .ZN(n8955) );
  INV_X1 U10254 ( .A(n8955), .ZN(n9308) );
  MUX2_X1 U10255 ( .A(n8845), .B(n8844), .S(n8921), .Z(n8846) );
  NAND3_X1 U10256 ( .A1(n8847), .A2(n9308), .A3(n8846), .ZN(n8855) );
  NAND2_X1 U10257 ( .A1(n8849), .A2(n8848), .ZN(n8852) );
  INV_X1 U10258 ( .A(n8850), .ZN(n8851) );
  MUX2_X1 U10259 ( .A(n8852), .B(n8851), .S(n8921), .Z(n8853) );
  INV_X1 U10260 ( .A(n8853), .ZN(n8854) );
  NAND2_X1 U10261 ( .A1(n8855), .A2(n8854), .ZN(n8862) );
  INV_X1 U10262 ( .A(n8856), .ZN(n8857) );
  NAND2_X1 U10263 ( .A1(n8862), .A2(n8857), .ZN(n8859) );
  NAND2_X1 U10264 ( .A1(n8859), .A2(n8858), .ZN(n8866) );
  NAND3_X1 U10265 ( .A1(n8862), .A2(n8861), .A3(n8860), .ZN(n8864) );
  NAND3_X1 U10266 ( .A1(n8864), .A2(n7616), .A3(n8863), .ZN(n8865) );
  INV_X1 U10267 ( .A(n8934), .ZN(n9236) );
  NAND3_X1 U10268 ( .A1(n8884), .A2(n8886), .A3(n9236), .ZN(n8870) );
  INV_X1 U10269 ( .A(n8867), .ZN(n8869) );
  NAND2_X1 U10270 ( .A1(n9190), .A2(n8932), .ZN(n8868) );
  AOI21_X1 U10271 ( .B1(n8870), .B2(n8869), .A(n8868), .ZN(n8874) );
  INV_X1 U10272 ( .A(n8888), .ZN(n8873) );
  INV_X1 U10273 ( .A(n8871), .ZN(n8872) );
  NOR2_X1 U10274 ( .A1(n8872), .A2(n8893), .ZN(n8889) );
  OAI21_X1 U10275 ( .B1(n8874), .B2(n8873), .A(n8889), .ZN(n8876) );
  NAND2_X1 U10276 ( .A1(n8876), .A2(n8875), .ZN(n8883) );
  NAND2_X1 U10277 ( .A1(n8894), .A2(n8880), .ZN(n9164) );
  MUX2_X1 U10278 ( .A(n9161), .B(n8877), .S(n8921), .Z(n8878) );
  INV_X1 U10279 ( .A(n8878), .ZN(n8879) );
  NOR2_X1 U10280 ( .A1(n9164), .A2(n8879), .ZN(n8898) );
  NAND4_X1 U10281 ( .A1(n9128), .A2(n8901), .A3(n8881), .A4(n8880), .ZN(n8882)
         );
  AOI21_X1 U10282 ( .B1(n8883), .B2(n8898), .A(n8882), .ZN(n8912) );
  INV_X1 U10283 ( .A(n8884), .ZN(n8887) );
  AOI21_X1 U10284 ( .B1(n8887), .B2(n8886), .A(n8885), .ZN(n8890) );
  OAI211_X1 U10285 ( .C1(n8890), .C2(n4645), .A(n8889), .B(n8888), .ZN(n8891)
         );
  OAI211_X1 U10286 ( .C1(n8893), .C2(n8892), .A(n8891), .B(n9161), .ZN(n8899)
         );
  NAND4_X1 U10287 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8921), .ZN(n8897)
         );
  AOI21_X1 U10288 ( .B1(n8899), .B2(n8898), .A(n8897), .ZN(n8911) );
  NAND2_X1 U10289 ( .A1(n9166), .A2(n8921), .ZN(n8902) );
  INV_X1 U10290 ( .A(n8902), .ZN(n8900) );
  AOI22_X1 U10291 ( .A1(n9356), .A2(n8900), .B1(n9150), .B2(n8921), .ZN(n8909)
         );
  NAND2_X1 U10292 ( .A1(n9012), .A2(n8901), .ZN(n8903) );
  OAI22_X1 U10293 ( .A1(n9356), .A2(n8903), .B1(n9150), .B2(n8921), .ZN(n8907)
         );
  OAI21_X1 U10294 ( .B1(n9124), .B2(n8902), .A(n9356), .ZN(n8906) );
  NOR2_X1 U10295 ( .A1(n8903), .A2(n9150), .ZN(n8904) );
  OR2_X1 U10296 ( .A1(n9356), .A2(n8904), .ZN(n8905) );
  AOI22_X1 U10297 ( .A1(n9123), .A2(n8907), .B1(n8906), .B2(n8905), .ZN(n8908)
         );
  OAI211_X1 U10298 ( .C1(n9123), .C2(n8909), .A(n9130), .B(n8908), .ZN(n8910)
         );
  INV_X1 U10299 ( .A(n9132), .ZN(n9010) );
  NAND2_X1 U10300 ( .A1(n9010), .A2(n8917), .ZN(n8913) );
  NAND2_X1 U10301 ( .A1(n9340), .A2(n8913), .ZN(n8988) );
  MUX2_X1 U10302 ( .A(n8987), .B(n8914), .S(n8921), .Z(n8915) );
  NAND3_X1 U10303 ( .A1(n8916), .A2(n8988), .A3(n8915), .ZN(n8920) );
  NAND2_X1 U10304 ( .A1(n8918), .A2(n8917), .ZN(n8919) );
  NAND2_X1 U10305 ( .A1(n8919), .A2(n9336), .ZN(n8994) );
  MUX2_X1 U10306 ( .A(n8921), .B(n8920), .S(n8994), .Z(n8926) );
  INV_X1 U10307 ( .A(n8988), .ZN(n8922) );
  NAND3_X1 U10308 ( .A1(n8962), .A2(n8922), .A3(n8921), .ZN(n8924) );
  AND2_X1 U10309 ( .A1(n8924), .A2(n8923), .ZN(n8925) );
  NAND2_X1 U10310 ( .A1(n8926), .A2(n8925), .ZN(n8999) );
  INV_X1 U10311 ( .A(n8927), .ZN(n8966) );
  INV_X1 U10312 ( .A(n8928), .ZN(n8930) );
  NAND2_X1 U10313 ( .A1(n8932), .A2(n8931), .ZN(n9228) );
  NOR2_X1 U10314 ( .A1(n8934), .A2(n8933), .ZN(n9261) );
  INV_X1 U10315 ( .A(n9323), .ZN(n8953) );
  NOR2_X1 U10316 ( .A1(n6576), .A2(n8935), .ZN(n8938) );
  NAND4_X1 U10317 ( .A1(n8938), .A2(n4513), .A3(n8937), .A4(n8936), .ZN(n8942)
         );
  NOR4_X1 U10318 ( .A1(n8942), .A2(n8941), .A3(n8940), .A4(n8939), .ZN(n8946)
         );
  INV_X1 U10319 ( .A(n8943), .ZN(n8944) );
  NAND3_X1 U10320 ( .A1(n8946), .A2(n8945), .A3(n8944), .ZN(n8949) );
  NOR4_X1 U10321 ( .A1(n8949), .A2(n8948), .A3(n8947), .A4(n9503), .ZN(n8951)
         );
  NAND4_X1 U10322 ( .A1(n8953), .A2(n8952), .A3(n8951), .A4(n8950), .ZN(n8954)
         );
  NOR4_X1 U10323 ( .A1(n9286), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n8957)
         );
  NAND4_X1 U10324 ( .A1(n9246), .A2(n9261), .A3(n9275), .A4(n8957), .ZN(n8958)
         );
  OR4_X1 U10325 ( .A1(n9192), .A2(n9213), .A3(n9228), .A4(n8958), .ZN(n8959)
         );
  NOR4_X1 U10326 ( .A1(n9147), .A2(n9164), .A3(n9182), .A4(n8959), .ZN(n8960)
         );
  XNOR2_X1 U10327 ( .A(n9340), .B(n9132), .ZN(n8963) );
  INV_X1 U10328 ( .A(n8996), .ZN(n8965) );
  OAI21_X1 U10329 ( .B1(n8999), .B2(n8966), .A(n8965), .ZN(n8998) );
  INV_X1 U10330 ( .A(n8967), .ZN(n8970) );
  OAI21_X1 U10331 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n8974) );
  AOI22_X1 U10332 ( .A1(n8974), .A2(n8973), .B1(n8972), .B2(n8971), .ZN(n8976)
         );
  AOI21_X1 U10333 ( .B1(n8976), .B2(n8975), .A(n4764), .ZN(n8982) );
  NAND3_X1 U10334 ( .A1(n8979), .A2(n8978), .A3(n8977), .ZN(n8980) );
  NAND4_X1 U10335 ( .A1(n8983), .A2(n8982), .A3(n8981), .A4(n8980), .ZN(n8984)
         );
  NOR4_X1 U10336 ( .A1(n8986), .A2(n4642), .A3(n8985), .A4(n8984), .ZN(n8990)
         );
  OAI211_X1 U10337 ( .C1(n8990), .C2(n8989), .A(n8988), .B(n8987), .ZN(n8993)
         );
  AOI211_X1 U10338 ( .C1(n8994), .C2(n8993), .A(n8992), .B(n8991), .ZN(n8995)
         );
  NOR2_X1 U10339 ( .A1(n8996), .A2(n8995), .ZN(n8997) );
  INV_X1 U10340 ( .A(n9004), .ZN(n9009) );
  NAND2_X1 U10341 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  OAI211_X1 U10342 ( .C1(n9007), .C2(n9006), .A(P1_B_REG_SCAN_IN), .B(n9005), 
        .ZN(n9008) );
  MUX2_X1 U10343 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9010), .S(n9025), .Z(
        P1_U3585) );
  MUX2_X1 U10344 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9011), .S(n9025), .Z(
        P1_U3584) );
  MUX2_X1 U10345 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9124), .S(n9025), .Z(
        P1_U3583) );
  MUX2_X1 U10346 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9012), .S(n9025), .Z(
        P1_U3582) );
  MUX2_X1 U10347 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9184), .S(n9025), .Z(
        P1_U3581) );
  MUX2_X1 U10348 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9013), .S(n9025), .Z(
        P1_U3580) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9216), .S(n9025), .Z(
        P1_U3579) );
  MUX2_X1 U10350 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9230), .S(n9025), .Z(
        P1_U3578) );
  MUX2_X1 U10351 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9240), .S(n9025), .Z(
        P1_U3577) );
  MUX2_X1 U10352 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9231), .S(n9025), .Z(
        P1_U3576) );
  MUX2_X1 U10353 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9277), .S(n9025), .Z(
        P1_U3575) );
  MUX2_X1 U10354 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9284), .S(n9025), .Z(
        P1_U3574) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9276), .S(n9025), .Z(
        P1_U3573) );
  MUX2_X1 U10356 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9283), .S(n9025), .Z(
        P1_U3572) );
  MUX2_X1 U10357 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9329), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10358 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9014), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10359 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9328), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10360 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9015), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10361 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9016), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10362 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9505), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9017), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10364 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9506), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10365 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9018), .S(n9025), .Z(
        P1_U3563) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9019), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9020), .S(n9025), .Z(
        P1_U3561) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9021), .S(n9025), .Z(
        P1_U3560) );
  MUX2_X1 U10369 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9022), .S(n9025), .Z(
        P1_U3559) );
  MUX2_X1 U10370 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9023), .S(n9025), .Z(
        P1_U3558) );
  MUX2_X1 U10371 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9024), .S(n9025), .Z(
        P1_U3557) );
  MUX2_X1 U10372 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6570), .S(n9025), .Z(
        P1_U3556) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9026), .S(n9025), .Z(
        P1_U3555) );
  AOI22_X1 U10374 ( .A1(n9742), .A2(n9027), .B1(n9749), .B2(
        P1_ADDR_REG_7__SCAN_IN), .ZN(n9039) );
  OAI21_X1 U10375 ( .B1(n9030), .B2(n9029), .A(n9028), .ZN(n9032) );
  AOI21_X1 U10376 ( .B1(n9750), .B2(n9032), .A(n9031), .ZN(n9038) );
  OAI21_X1 U10377 ( .B1(n9035), .B2(n9034), .A(n9033), .ZN(n9036) );
  NAND2_X1 U10378 ( .A1(n9740), .A2(n9036), .ZN(n9037) );
  NAND3_X1 U10379 ( .A1(n9039), .A2(n9038), .A3(n9037), .ZN(P1_U3248) );
  OAI21_X1 U10380 ( .B1(n9042), .B2(n9041), .A(n9040), .ZN(n9043) );
  NAND2_X1 U10381 ( .A1(n9043), .A2(n9750), .ZN(n9053) );
  INV_X1 U10382 ( .A(n9044), .ZN(n9052) );
  AOI211_X1 U10383 ( .C1(n9047), .C2(n9046), .A(n9045), .B(n9713), .ZN(n9048)
         );
  AOI21_X1 U10384 ( .B1(n9742), .B2(n9049), .A(n9048), .ZN(n9051) );
  NAND2_X1 U10385 ( .A1(n9749), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n9050) );
  NAND4_X1 U10386 ( .A1(n9053), .A2(n9052), .A3(n9051), .A4(n9050), .ZN(
        P1_U3253) );
  OAI21_X1 U10387 ( .B1(n9056), .B2(n9055), .A(n9054), .ZN(n9057) );
  NAND2_X1 U10388 ( .A1(n9057), .A2(n9750), .ZN(n9066) );
  AOI211_X1 U10389 ( .C1(n9060), .C2(n9059), .A(n9058), .B(n9713), .ZN(n9061)
         );
  AOI21_X1 U10390 ( .B1(n9742), .B2(n9062), .A(n9061), .ZN(n9065) );
  NAND2_X1 U10391 ( .A1(n9749), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n9063) );
  NAND4_X1 U10392 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(
        P1_U3254) );
  NOR2_X1 U10393 ( .A1(n9067), .A2(n9074), .ZN(n9069) );
  NAND2_X1 U10394 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9091), .ZN(n9070) );
  OAI21_X1 U10395 ( .B1(n9091), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9070), .ZN(
        n9071) );
  AOI211_X1 U10396 ( .C1(n9072), .C2(n9071), .A(n9086), .B(n9713), .ZN(n9085)
         );
  NOR2_X1 U10397 ( .A1(n9074), .A2(n9073), .ZN(n9076) );
  NOR2_X1 U10398 ( .A1(n9076), .A2(n9075), .ZN(n9078) );
  XNOR2_X1 U10399 ( .A(n9091), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9077) );
  NOR2_X1 U10400 ( .A1(n9078), .A2(n9077), .ZN(n9090) );
  AOI211_X1 U10401 ( .C1(n9078), .C2(n9077), .A(n9090), .B(n9657), .ZN(n9084)
         );
  NAND2_X1 U10402 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n9080) );
  NAND2_X1 U10403 ( .A1(n9749), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9079) );
  OAI211_X1 U10404 ( .C1(n9082), .C2(n9081), .A(n9080), .B(n9079), .ZN(n9083)
         );
  OR3_X1 U10405 ( .A1(n9085), .A2(n9084), .A3(n9083), .ZN(P1_U3257) );
  NAND2_X1 U10406 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9105), .ZN(n9087) );
  OAI21_X1 U10407 ( .B1(n9105), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9087), .ZN(
        n9088) );
  AOI211_X1 U10408 ( .C1(n9089), .C2(n9088), .A(n9099), .B(n9713), .ZN(n9096)
         );
  AOI21_X1 U10409 ( .B1(n9091), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9090), .ZN(
        n9093) );
  XNOR2_X1 U10410 ( .A(n9105), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9092) );
  NOR2_X1 U10411 ( .A1(n9093), .A2(n9092), .ZN(n9104) );
  AOI211_X1 U10412 ( .C1(n9093), .C2(n9092), .A(n9104), .B(n9657), .ZN(n9095)
         );
  AND2_X1 U10413 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9094) );
  NOR3_X1 U10414 ( .A1(n9096), .A2(n9095), .A3(n9094), .ZN(n9098) );
  AOI22_X1 U10415 ( .A1(n9742), .A2(n9105), .B1(n9749), .B2(
        P1_ADDR_REG_17__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U10416 ( .A1(n9098), .A2(n9097), .ZN(P1_U3258) );
  AOI21_X1 U10417 ( .B1(n9105), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9099), .ZN(
        n9737) );
  OR2_X1 U10418 ( .A1(n9741), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U10419 ( .A1(n9741), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U10420 ( .A1(n9101), .A2(n9100), .ZN(n9738) );
  NOR2_X1 U10421 ( .A1(n9737), .A2(n9738), .ZN(n9736) );
  AOI21_X1 U10422 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9741), .A(n9736), .ZN(
        n9102) );
  XNOR2_X1 U10423 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9102), .ZN(n9109) );
  AOI22_X1 U10424 ( .A1(n9741), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n10262), 
        .B2(n9103), .ZN(n9748) );
  AOI21_X1 U10425 ( .B1(n9105), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9104), .ZN(
        n9747) );
  NAND2_X1 U10426 ( .A1(n9748), .A2(n9747), .ZN(n9746) );
  OAI21_X1 U10427 ( .B1(n9741), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9746), .ZN(
        n9106) );
  XNOR2_X1 U10428 ( .A(n9106), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9107) );
  AOI22_X1 U10429 ( .A1(n9109), .A2(n9740), .B1(n9750), .B2(n9107), .ZN(n9111)
         );
  INV_X1 U10430 ( .A(n9107), .ZN(n9110) );
  INV_X1 U10431 ( .A(n9340), .ZN(n9119) );
  XNOR2_X1 U10432 ( .A(n9336), .B(n4495), .ZN(n9338) );
  NAND2_X1 U10433 ( .A1(n9113), .A2(P1_B_REG_SCAN_IN), .ZN(n9114) );
  NAND2_X1 U10434 ( .A1(n9504), .A2(n9114), .ZN(n9131) );
  NOR2_X1 U10435 ( .A1(n9115), .A2(n9131), .ZN(n9339) );
  NAND2_X1 U10436 ( .A1(n9339), .A2(n9786), .ZN(n9120) );
  OAI21_X1 U10437 ( .B1(n9786), .B2(n9116), .A(n9120), .ZN(n9117) );
  AOI21_X1 U10438 ( .B1(n9336), .B2(n9516), .A(n9117), .ZN(n9118) );
  OAI21_X1 U10439 ( .B1(n9338), .B2(n9139), .A(n9118), .ZN(P1_U3261) );
  OAI21_X1 U10440 ( .B1(n9136), .B2(n9119), .A(n4495), .ZN(n9342) );
  OAI21_X1 U10441 ( .B1(n9786), .B2(n10275), .A(n9120), .ZN(n9121) );
  AOI21_X1 U10442 ( .B1(n9340), .B2(n9516), .A(n9121), .ZN(n9122) );
  OAI21_X1 U10443 ( .B1(n9342), .B2(n9139), .A(n9122), .ZN(P1_U3262) );
  NAND2_X1 U10444 ( .A1(n9350), .A2(n9124), .ZN(n9125) );
  NAND2_X1 U10445 ( .A1(n9126), .A2(n9125), .ZN(n9127) );
  XNOR2_X1 U10446 ( .A(n9127), .B(n9130), .ZN(n9343) );
  INV_X1 U10447 ( .A(n9343), .ZN(n9144) );
  OAI22_X1 U10448 ( .A1(n9150), .A2(n9773), .B1(n9132), .B2(n9131), .ZN(n9133)
         );
  OAI21_X1 U10449 ( .B1(n9135), .B2(n9790), .A(n9347), .ZN(n9142) );
  AOI21_X1 U10450 ( .B1(n9344), .B2(n9137), .A(n9136), .ZN(n9345) );
  INV_X1 U10451 ( .A(n9345), .ZN(n9140) );
  AOI22_X1 U10452 ( .A1(n9344), .A2(n9516), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9767), .ZN(n9138) );
  OAI21_X1 U10453 ( .B1(n9140), .B2(n9139), .A(n9138), .ZN(n9141) );
  AOI21_X1 U10454 ( .B1(n9142), .B2(n9786), .A(n9141), .ZN(n9143) );
  OAI21_X1 U10455 ( .B1(n9144), .B2(n9335), .A(n9143), .ZN(P1_U3355) );
  XOR2_X1 U10456 ( .A(n9147), .B(n9145), .Z(n9359) );
  NOR2_X1 U10457 ( .A1(n9146), .A2(n9321), .ZN(n9159) );
  AOI21_X1 U10458 ( .B1(n9148), .B2(n9147), .A(n9509), .ZN(n9153) );
  OAI22_X1 U10459 ( .A1(n9150), .A2(n9771), .B1(n9149), .B2(n9773), .ZN(n9151)
         );
  AOI21_X1 U10460 ( .B1(n9153), .B2(n9152), .A(n9151), .ZN(n9358) );
  INV_X1 U10461 ( .A(n9154), .ZN(n9155) );
  AOI211_X1 U10462 ( .C1(n9356), .C2(n9167), .A(n9830), .B(n9155), .ZN(n9355)
         );
  AOI22_X1 U10463 ( .A1(n9355), .A2(n4473), .B1(n9156), .B2(n9514), .ZN(n9157)
         );
  AOI21_X1 U10464 ( .B1(n9358), .B2(n9157), .A(n9767), .ZN(n9158) );
  AOI211_X1 U10465 ( .C1(n9767), .C2(P1_REG2_REG_27__SCAN_IN), .A(n9159), .B(
        n9158), .ZN(n9160) );
  OAI21_X1 U10466 ( .B1(n9359), .B2(n9335), .A(n9160), .ZN(P1_U3264) );
  XNOR2_X1 U10467 ( .A(n4540), .B(n9164), .ZN(n9364) );
  NAND2_X1 U10468 ( .A1(n9162), .A2(n9161), .ZN(n9163) );
  XOR2_X1 U10469 ( .A(n9164), .B(n9163), .Z(n9165) );
  OAI222_X1 U10470 ( .A1(n9771), .A2(n9166), .B1(n9773), .B2(n9195), .C1(n9509), .C2(n9165), .ZN(n9360) );
  INV_X1 U10471 ( .A(n9178), .ZN(n9169) );
  INV_X1 U10472 ( .A(n9167), .ZN(n9168) );
  AOI211_X1 U10473 ( .C1(n9362), .C2(n9169), .A(n9830), .B(n9168), .ZN(n9361)
         );
  NAND2_X1 U10474 ( .A1(n9361), .A2(n9521), .ZN(n9173) );
  INV_X1 U10475 ( .A(n9170), .ZN(n9171) );
  AOI22_X1 U10476 ( .A1(n9171), .A2(n9514), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9767), .ZN(n9172) );
  OAI211_X1 U10477 ( .C1(n9174), .C2(n9321), .A(n9173), .B(n9172), .ZN(n9175)
         );
  AOI21_X1 U10478 ( .B1(n9360), .B2(n9786), .A(n9175), .ZN(n9176) );
  OAI21_X1 U10479 ( .B1(n9364), .B2(n9335), .A(n9176), .ZN(P1_U3265) );
  XOR2_X1 U10480 ( .A(n9182), .B(n9177), .Z(n9369) );
  AOI21_X1 U10481 ( .B1(n9365), .B2(n4700), .A(n9178), .ZN(n9366) );
  AOI22_X1 U10482 ( .A1(n9179), .A2(n9514), .B1(n9767), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n9180) );
  OAI21_X1 U10483 ( .B1(n9181), .B2(n9321), .A(n9180), .ZN(n9187) );
  XNOR2_X1 U10484 ( .A(n9183), .B(n9182), .ZN(n9185) );
  AOI222_X1 U10485 ( .A1(n9776), .A2(n9185), .B1(n9184), .B2(n9504), .C1(n9216), .C2(n9507), .ZN(n9368) );
  NOR2_X1 U10486 ( .A1(n9368), .A2(n9767), .ZN(n9186) );
  AOI211_X1 U10487 ( .C1(n9366), .C2(n9333), .A(n9187), .B(n9186), .ZN(n9188)
         );
  OAI21_X1 U10488 ( .B1(n9369), .B2(n9335), .A(n9188), .ZN(P1_U3266) );
  XNOR2_X1 U10489 ( .A(n9189), .B(n9192), .ZN(n9374) );
  AOI22_X1 U10490 ( .A1(n9372), .A2(n9516), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9767), .ZN(n9202) );
  NAND2_X1 U10491 ( .A1(n9210), .A2(n9190), .ZN(n9191) );
  XOR2_X1 U10492 ( .A(n9192), .B(n9191), .Z(n9193) );
  OAI222_X1 U10493 ( .A1(n9771), .A2(n9195), .B1(n9773), .B2(n9194), .C1(n9193), .C2(n9509), .ZN(n9370) );
  AOI211_X1 U10494 ( .C1(n9372), .C2(n9204), .A(n9830), .B(n9196), .ZN(n9371)
         );
  INV_X1 U10495 ( .A(n9371), .ZN(n9199) );
  INV_X1 U10496 ( .A(n9197), .ZN(n9198) );
  OAI22_X1 U10497 ( .A1(n9199), .A2(n9785), .B1(n9198), .B2(n9790), .ZN(n9200)
         );
  OAI21_X1 U10498 ( .B1(n9370), .B2(n9200), .A(n9786), .ZN(n9201) );
  OAI211_X1 U10499 ( .C1(n9374), .C2(n9335), .A(n9202), .B(n9201), .ZN(
        P1_U3267) );
  XNOR2_X1 U10500 ( .A(n9203), .B(n9213), .ZN(n9379) );
  INV_X1 U10501 ( .A(n9204), .ZN(n9205) );
  AOI21_X1 U10502 ( .B1(n9375), .B2(n9221), .A(n9205), .ZN(n9376) );
  INV_X1 U10503 ( .A(n9206), .ZN(n9207) );
  AOI22_X1 U10504 ( .A1(n9767), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9207), .B2(
        n9514), .ZN(n9208) );
  OAI21_X1 U10505 ( .B1(n9209), .B2(n9321), .A(n9208), .ZN(n9218) );
  AND2_X1 U10506 ( .A1(n9240), .A2(n9507), .ZN(n9215) );
  INV_X1 U10507 ( .A(n9210), .ZN(n9211) );
  AOI211_X1 U10508 ( .C1(n9213), .C2(n9212), .A(n9509), .B(n9211), .ZN(n9214)
         );
  AOI211_X1 U10509 ( .C1(n9504), .C2(n9216), .A(n9215), .B(n9214), .ZN(n9378)
         );
  NOR2_X1 U10510 ( .A1(n9378), .A2(n9767), .ZN(n9217) );
  AOI211_X1 U10511 ( .C1(n9376), .C2(n9333), .A(n9218), .B(n9217), .ZN(n9219)
         );
  OAI21_X1 U10512 ( .B1(n9379), .B2(n9335), .A(n9219), .ZN(P1_U3268) );
  XOR2_X1 U10513 ( .A(n9228), .B(n9220), .Z(n9384) );
  INV_X1 U10514 ( .A(n9242), .ZN(n9223) );
  INV_X1 U10515 ( .A(n9221), .ZN(n9222) );
  AOI21_X1 U10516 ( .B1(n9380), .B2(n9223), .A(n9222), .ZN(n9381) );
  INV_X1 U10517 ( .A(n9224), .ZN(n9225) );
  AOI22_X1 U10518 ( .A1(n9767), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9225), .B2(
        n9514), .ZN(n9226) );
  OAI21_X1 U10519 ( .B1(n9227), .B2(n9321), .A(n9226), .ZN(n9234) );
  XOR2_X1 U10520 ( .A(n9229), .B(n9228), .Z(n9232) );
  AOI222_X1 U10521 ( .A1(n9776), .A2(n9232), .B1(n9231), .B2(n9507), .C1(n9230), .C2(n9504), .ZN(n9383) );
  NOR2_X1 U10522 ( .A1(n9383), .A2(n9767), .ZN(n9233) );
  AOI211_X1 U10523 ( .C1(n9381), .C2(n9333), .A(n9234), .B(n9233), .ZN(n9235)
         );
  OAI21_X1 U10524 ( .B1(n9384), .B2(n9335), .A(n9235), .ZN(P1_U3269) );
  AND2_X1 U10525 ( .A1(n9237), .A2(n9236), .ZN(n9239) );
  OAI21_X1 U10526 ( .B1(n9239), .B2(n9246), .A(n9238), .ZN(n9241) );
  AOI222_X1 U10527 ( .A1(n9776), .A2(n9241), .B1(n9277), .B2(n9507), .C1(n9240), .C2(n9504), .ZN(n9389) );
  INV_X1 U10528 ( .A(n9254), .ZN(n9243) );
  AOI211_X1 U10529 ( .C1(n9387), .C2(n9243), .A(n9830), .B(n9242), .ZN(n9386)
         );
  AOI22_X1 U10530 ( .A1(n9386), .A2(n4473), .B1(n9244), .B2(n9514), .ZN(n9245)
         );
  AND2_X1 U10531 ( .A1(n9389), .A2(n9245), .ZN(n9251) );
  INV_X1 U10532 ( .A(n9391), .ZN(n9248) );
  INV_X1 U10533 ( .A(n9335), .ZN(n9288) );
  NAND2_X1 U10534 ( .A1(n9247), .A2(n9246), .ZN(n9385) );
  NAND3_X1 U10535 ( .A1(n9248), .A2(n9288), .A3(n9385), .ZN(n9250) );
  AOI22_X1 U10536 ( .A1(n9387), .A2(n9516), .B1(n9767), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9249) );
  OAI211_X1 U10537 ( .C1(n9767), .C2(n9251), .A(n9250), .B(n9249), .ZN(
        P1_U3270) );
  XNOR2_X1 U10538 ( .A(n9253), .B(n9261), .ZN(n9396) );
  AOI211_X1 U10539 ( .C1(n9394), .C2(n9268), .A(n9830), .B(n9254), .ZN(n9393)
         );
  NOR2_X1 U10540 ( .A1(n9255), .A2(n9321), .ZN(n9259) );
  OAI22_X1 U10541 ( .A1(n9786), .A2(n9257), .B1(n9256), .B2(n9790), .ZN(n9258)
         );
  AOI211_X1 U10542 ( .C1(n9393), .C2(n9521), .A(n9259), .B(n9258), .ZN(n9266)
         );
  XOR2_X1 U10543 ( .A(n9261), .B(n9260), .Z(n9262) );
  OAI222_X1 U10544 ( .A1(n9771), .A2(n9264), .B1(n9773), .B2(n9263), .C1(n9262), .C2(n9509), .ZN(n9392) );
  NAND2_X1 U10545 ( .A1(n9392), .A2(n9786), .ZN(n9265) );
  OAI211_X1 U10546 ( .C1(n9396), .C2(n9335), .A(n9266), .B(n9265), .ZN(
        P1_U3271) );
  XOR2_X1 U10547 ( .A(n9267), .B(n9275), .Z(n9401) );
  INV_X1 U10548 ( .A(n9268), .ZN(n9269) );
  AOI211_X1 U10549 ( .C1(n9398), .C2(n9289), .A(n9830), .B(n9269), .ZN(n9397)
         );
  AOI22_X1 U10550 ( .A1(n9767), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9270), .B2(
        n9514), .ZN(n9271) );
  OAI21_X1 U10551 ( .B1(n9272), .B2(n9321), .A(n9271), .ZN(n9280) );
  OAI21_X1 U10552 ( .B1(n9275), .B2(n9274), .A(n9273), .ZN(n9278) );
  AOI222_X1 U10553 ( .A1(n9776), .A2(n9278), .B1(n9277), .B2(n9504), .C1(n9276), .C2(n9507), .ZN(n9400) );
  NOR2_X1 U10554 ( .A1(n9400), .A2(n9767), .ZN(n9279) );
  AOI211_X1 U10555 ( .C1(n9397), .C2(n9521), .A(n9280), .B(n9279), .ZN(n9281)
         );
  OAI21_X1 U10556 ( .B1(n9401), .B2(n9335), .A(n9281), .ZN(P1_U3272) );
  XNOR2_X1 U10557 ( .A(n9282), .B(n9286), .ZN(n9285) );
  AOI222_X1 U10558 ( .A1(n9776), .A2(n9285), .B1(n9284), .B2(n9504), .C1(n9283), .C2(n9507), .ZN(n9407) );
  OR2_X1 U10559 ( .A1(n9287), .A2(n9286), .ZN(n9403) );
  NAND3_X1 U10560 ( .A1(n9403), .A2(n9402), .A3(n9288), .ZN(n9298) );
  INV_X1 U10561 ( .A(n9300), .ZN(n9291) );
  INV_X1 U10562 ( .A(n9289), .ZN(n9290) );
  AOI21_X1 U10563 ( .B1(n9404), .B2(n9291), .A(n9290), .ZN(n9405) );
  NOR2_X1 U10564 ( .A1(n9292), .A2(n9321), .ZN(n9296) );
  OAI22_X1 U10565 ( .A1(n9786), .A2(n9294), .B1(n9293), .B2(n9790), .ZN(n9295)
         );
  AOI211_X1 U10566 ( .C1(n9405), .C2(n9333), .A(n9296), .B(n9295), .ZN(n9297)
         );
  OAI211_X1 U10567 ( .C1(n9767), .C2(n9407), .A(n9298), .B(n9297), .ZN(
        P1_U3273) );
  XNOR2_X1 U10568 ( .A(n9299), .B(n9308), .ZN(n9413) );
  AOI211_X1 U10569 ( .C1(n9411), .C2(n9301), .A(n9830), .B(n9300), .ZN(n9410)
         );
  NOR2_X1 U10570 ( .A1(n9302), .A2(n9321), .ZN(n9307) );
  OAI22_X1 U10571 ( .A1(n9786), .A2(n9304), .B1(n9303), .B2(n9790), .ZN(n9306)
         );
  AOI211_X1 U10572 ( .C1(n9410), .C2(n9521), .A(n9307), .B(n9306), .ZN(n9314)
         );
  XNOR2_X1 U10573 ( .A(n9309), .B(n9308), .ZN(n9310) );
  OAI222_X1 U10574 ( .A1(n9771), .A2(n9312), .B1(n9773), .B2(n9311), .C1(n9509), .C2(n9310), .ZN(n9409) );
  NAND2_X1 U10575 ( .A1(n9409), .A2(n9786), .ZN(n9313) );
  OAI211_X1 U10576 ( .C1(n9413), .C2(n9335), .A(n9314), .B(n9313), .ZN(
        P1_U3274) );
  XNOR2_X1 U10577 ( .A(n9315), .B(n9323), .ZN(n9423) );
  AOI21_X1 U10578 ( .B1(n9419), .B2(n9317), .A(n4701), .ZN(n9420) );
  INV_X1 U10579 ( .A(n9318), .ZN(n9319) );
  AOI22_X1 U10580 ( .A1(n9767), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9319), .B2(
        n9514), .ZN(n9320) );
  OAI21_X1 U10581 ( .B1(n9322), .B2(n9321), .A(n9320), .ZN(n9332) );
  INV_X1 U10582 ( .A(n7429), .ZN(n9325) );
  OAI21_X1 U10583 ( .B1(n9325), .B2(n9324), .A(n9323), .ZN(n9327) );
  NAND2_X1 U10584 ( .A1(n9327), .A2(n9326), .ZN(n9330) );
  AOI222_X1 U10585 ( .A1(n9776), .A2(n9330), .B1(n9329), .B2(n9504), .C1(n9328), .C2(n9507), .ZN(n9422) );
  NOR2_X1 U10586 ( .A1(n9422), .A2(n9767), .ZN(n9331) );
  AOI211_X1 U10587 ( .C1(n9420), .C2(n9333), .A(n9332), .B(n9331), .ZN(n9334)
         );
  OAI21_X1 U10588 ( .B1(n9335), .B2(n9423), .A(n9334), .ZN(P1_U3276) );
  AOI21_X1 U10589 ( .B1(n9336), .B2(n9524), .A(n9339), .ZN(n9337) );
  OAI21_X1 U10590 ( .B1(n9338), .B2(n9830), .A(n9337), .ZN(n9435) );
  MUX2_X1 U10591 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9435), .S(n9848), .Z(
        P1_U3554) );
  AOI21_X1 U10592 ( .B1(n9340), .B2(n9524), .A(n9339), .ZN(n9341) );
  OAI21_X1 U10593 ( .B1(n9342), .B2(n9830), .A(n9341), .ZN(n9436) );
  MUX2_X1 U10594 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9436), .S(n9848), .Z(
        P1_U3553) );
  INV_X1 U10595 ( .A(n9434), .ZN(n9824) );
  NAND2_X1 U10596 ( .A1(n9343), .A2(n9824), .ZN(n9349) );
  AOI22_X1 U10597 ( .A1(n9345), .A2(n9782), .B1(n9524), .B2(n9344), .ZN(n9346)
         );
  AND2_X1 U10598 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  NAND2_X1 U10599 ( .A1(n9349), .A2(n9348), .ZN(n9437) );
  MUX2_X1 U10600 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9437), .S(n9848), .Z(
        P1_U3552) );
  AOI22_X1 U10601 ( .A1(n9351), .A2(n9782), .B1(n9524), .B2(n9350), .ZN(n9352)
         );
  OAI211_X1 U10602 ( .C1(n9354), .C2(n9434), .A(n9353), .B(n9352), .ZN(n9438)
         );
  MUX2_X1 U10603 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9438), .S(n9848), .Z(
        P1_U3551) );
  AOI21_X1 U10604 ( .B1(n9524), .B2(n9356), .A(n9355), .ZN(n9357) );
  OAI211_X1 U10605 ( .C1(n9359), .C2(n9434), .A(n9358), .B(n9357), .ZN(n9439)
         );
  MUX2_X1 U10606 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9439), .S(n9848), .Z(
        P1_U3550) );
  AOI211_X1 U10607 ( .C1(n9524), .C2(n9362), .A(n9361), .B(n9360), .ZN(n9363)
         );
  OAI21_X1 U10608 ( .B1(n9364), .B2(n9434), .A(n9363), .ZN(n9440) );
  MUX2_X1 U10609 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9440), .S(n9848), .Z(
        P1_U3549) );
  AOI22_X1 U10610 ( .A1(n9366), .A2(n9782), .B1(n9524), .B2(n9365), .ZN(n9367)
         );
  OAI211_X1 U10611 ( .C1(n9369), .C2(n9434), .A(n9368), .B(n9367), .ZN(n9441)
         );
  MUX2_X1 U10612 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9441), .S(n9848), .Z(
        P1_U3548) );
  AOI211_X1 U10613 ( .C1(n9524), .C2(n9372), .A(n9371), .B(n9370), .ZN(n9373)
         );
  OAI21_X1 U10614 ( .B1(n9374), .B2(n9434), .A(n9373), .ZN(n9442) );
  MUX2_X1 U10615 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9442), .S(n9848), .Z(
        P1_U3547) );
  AOI22_X1 U10616 ( .A1(n9376), .A2(n9782), .B1(n9524), .B2(n9375), .ZN(n9377)
         );
  OAI211_X1 U10617 ( .C1(n9379), .C2(n9434), .A(n9378), .B(n9377), .ZN(n9443)
         );
  MUX2_X1 U10618 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9443), .S(n9848), .Z(
        P1_U3546) );
  AOI22_X1 U10619 ( .A1(n9381), .A2(n9782), .B1(n9524), .B2(n9380), .ZN(n9382)
         );
  OAI211_X1 U10620 ( .C1(n9384), .C2(n9434), .A(n9383), .B(n9382), .ZN(n9444)
         );
  MUX2_X1 U10621 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9444), .S(n9848), .Z(
        P1_U3545) );
  NAND2_X1 U10622 ( .A1(n9385), .A2(n9824), .ZN(n9390) );
  AOI21_X1 U10623 ( .B1(n9524), .B2(n9387), .A(n9386), .ZN(n9388) );
  OAI211_X1 U10624 ( .C1(n9391), .C2(n9390), .A(n9389), .B(n9388), .ZN(n9445)
         );
  MUX2_X1 U10625 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9445), .S(n9848), .Z(
        P1_U3544) );
  AOI211_X1 U10626 ( .C1(n9524), .C2(n9394), .A(n9393), .B(n9392), .ZN(n9395)
         );
  OAI21_X1 U10627 ( .B1(n9396), .B2(n9434), .A(n9395), .ZN(n9446) );
  MUX2_X1 U10628 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9446), .S(n9848), .Z(
        P1_U3543) );
  AOI21_X1 U10629 ( .B1(n9524), .B2(n9398), .A(n9397), .ZN(n9399) );
  OAI211_X1 U10630 ( .C1(n9401), .C2(n9434), .A(n9400), .B(n9399), .ZN(n9447)
         );
  MUX2_X1 U10631 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9447), .S(n9848), .Z(
        P1_U3542) );
  NAND3_X1 U10632 ( .A1(n9403), .A2(n9402), .A3(n9824), .ZN(n9408) );
  AOI22_X1 U10633 ( .A1(n9405), .A2(n9782), .B1(n9524), .B2(n9404), .ZN(n9406)
         );
  NAND3_X1 U10634 ( .A1(n9408), .A2(n9407), .A3(n9406), .ZN(n9448) );
  MUX2_X1 U10635 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9448), .S(n9848), .Z(
        P1_U3541) );
  AOI211_X1 U10636 ( .C1(n9524), .C2(n9411), .A(n9410), .B(n9409), .ZN(n9412)
         );
  OAI21_X1 U10637 ( .B1(n9413), .B2(n9434), .A(n9412), .ZN(n9449) );
  MUX2_X1 U10638 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9449), .S(n9848), .Z(
        P1_U3540) );
  AOI211_X1 U10639 ( .C1(n9524), .C2(n9416), .A(n9415), .B(n9414), .ZN(n9417)
         );
  OAI21_X1 U10640 ( .B1(n9418), .B2(n9434), .A(n9417), .ZN(n9450) );
  MUX2_X1 U10641 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9450), .S(n9848), .Z(
        P1_U3539) );
  AOI22_X1 U10642 ( .A1(n9420), .A2(n9782), .B1(n9524), .B2(n9419), .ZN(n9421)
         );
  OAI211_X1 U10643 ( .C1(n9423), .C2(n9434), .A(n9422), .B(n9421), .ZN(n9451)
         );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9451), .S(n9848), .Z(
        P1_U3538) );
  AOI211_X1 U10645 ( .C1(n9524), .C2(n9426), .A(n9425), .B(n9424), .ZN(n9427)
         );
  OAI21_X1 U10646 ( .B1(n9428), .B2(n9434), .A(n9427), .ZN(n9452) );
  MUX2_X1 U10647 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9452), .S(n9848), .Z(
        P1_U3537) );
  AOI211_X1 U10648 ( .C1(n9524), .C2(n9431), .A(n9430), .B(n9429), .ZN(n9432)
         );
  OAI21_X1 U10649 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9453) );
  MUX2_X1 U10650 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9453), .S(n9848), .Z(
        P1_U3534) );
  MUX2_X1 U10651 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9435), .S(n4474), .Z(
        P1_U3522) );
  MUX2_X1 U10652 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9436), .S(n4474), .Z(
        P1_U3521) );
  MUX2_X1 U10653 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9437), .S(n4474), .Z(
        P1_U3520) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9438), .S(n4474), .Z(
        P1_U3519) );
  MUX2_X1 U10655 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9439), .S(n4474), .Z(
        P1_U3518) );
  MUX2_X1 U10656 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9440), .S(n4474), .Z(
        P1_U3517) );
  MUX2_X1 U10657 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9441), .S(n4474), .Z(
        P1_U3516) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9442), .S(n4474), .Z(
        P1_U3515) );
  MUX2_X1 U10659 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9443), .S(n4474), .Z(
        P1_U3514) );
  MUX2_X1 U10660 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9444), .S(n4474), .Z(
        P1_U3513) );
  MUX2_X1 U10661 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9445), .S(n4474), .Z(
        P1_U3512) );
  MUX2_X1 U10662 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9446), .S(n4474), .Z(
        P1_U3511) );
  MUX2_X1 U10663 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9447), .S(n4474), .Z(
        P1_U3510) );
  MUX2_X1 U10664 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9448), .S(n4474), .Z(
        P1_U3508) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9449), .S(n4474), .Z(
        P1_U3505) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9450), .S(n4474), .Z(
        P1_U3502) );
  MUX2_X1 U10667 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9451), .S(n4474), .Z(
        P1_U3499) );
  MUX2_X1 U10668 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9452), .S(n4474), .Z(
        P1_U3496) );
  MUX2_X1 U10669 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9453), .S(n4474), .Z(
        P1_U3487) );
  MUX2_X1 U10670 ( .A(n9455), .B(P1_D_REG_0__SCAN_IN), .S(n9454), .Z(P1_U3440)
         );
  NOR4_X1 U10671 ( .A1(n9457), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9456), .ZN(n9458) );
  AOI21_X1 U10672 ( .B1(n9465), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9458), .ZN(
        n9459) );
  OAI21_X1 U10673 ( .B1(n9460), .B2(n9463), .A(n9459), .ZN(P1_U3322) );
  AOI22_X1 U10674 ( .A1(n9461), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9465), .ZN(n9462) );
  OAI21_X1 U10675 ( .B1(n9464), .B2(n9463), .A(n9462), .ZN(P1_U3323) );
  AOI22_X1 U10676 ( .A1(n9466), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9465), .ZN(n9467) );
  OAI21_X1 U10677 ( .B1(n9468), .B2(n9463), .A(n9467), .ZN(P1_U3324) );
  MUX2_X1 U10678 ( .A(n9469), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10679 ( .A(n9470), .ZN(n9471) );
  AOI21_X1 U10680 ( .B1(n9857), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n9471), .ZN(
        n9483) );
  AOI211_X1 U10681 ( .C1(n9474), .C2(n9473), .A(n9472), .B(n9854), .ZN(n9475)
         );
  AOI21_X1 U10682 ( .B1(n9477), .B2(n9476), .A(n9475), .ZN(n9482) );
  NOR2_X1 U10683 ( .A1(n5098), .A2(n5082), .ZN(n9480) );
  OAI211_X1 U10684 ( .C1(n9480), .C2(n9479), .A(n9850), .B(n9478), .ZN(n9481)
         );
  NAND3_X1 U10685 ( .A1(n9483), .A2(n9482), .A3(n9481), .ZN(P2_U3246) );
  AOI21_X1 U10686 ( .B1(n9486), .B2(n9485), .A(n9484), .ZN(n9487) );
  NAND2_X1 U10687 ( .A1(n9849), .A2(n9487), .ZN(n9491) );
  INV_X1 U10688 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9538) );
  OAI22_X1 U10689 ( .A1(n9488), .A2(n9538), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5145), .ZN(n9489) );
  INV_X1 U10690 ( .A(n9489), .ZN(n9490) );
  OAI211_X1 U10691 ( .C1(n9852), .C2(n9492), .A(n9491), .B(n9490), .ZN(n9493)
         );
  INV_X1 U10692 ( .A(n9493), .ZN(n9498) );
  OAI211_X1 U10693 ( .C1(n9496), .C2(n9495), .A(n9850), .B(n9494), .ZN(n9497)
         );
  NAND2_X1 U10694 ( .A1(n9498), .A2(n9497), .ZN(P2_U3247) );
  XNOR2_X1 U10695 ( .A(n9499), .B(n9503), .ZN(n9530) );
  NAND2_X1 U10696 ( .A1(n9501), .A2(n9500), .ZN(n9502) );
  XOR2_X1 U10697 ( .A(n9503), .B(n9502), .Z(n9510) );
  AOI22_X1 U10698 ( .A1(n9507), .A2(n9506), .B1(n9505), .B2(n9504), .ZN(n9508)
         );
  OAI21_X1 U10699 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9511) );
  AOI21_X1 U10700 ( .B1(n9530), .B2(n9512), .A(n9511), .ZN(n9527) );
  INV_X1 U10701 ( .A(n9513), .ZN(n9515) );
  AOI222_X1 U10702 ( .A1(n9517), .A2(n9516), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n9767), .C1(n9515), .C2(n9514), .ZN(n9523) );
  OAI211_X1 U10703 ( .C1(n9519), .C2(n9526), .A(n9782), .B(n9518), .ZN(n9525)
         );
  INV_X1 U10704 ( .A(n9525), .ZN(n9520) );
  AOI22_X1 U10705 ( .A1(n9530), .A2(n9768), .B1(n9521), .B2(n9520), .ZN(n9522)
         );
  OAI211_X1 U10706 ( .C1(n9767), .C2(n9527), .A(n9523), .B(n9522), .ZN(
        P1_U3281) );
  INV_X1 U10707 ( .A(n9524), .ZN(n9828) );
  OAI21_X1 U10708 ( .B1(n9526), .B2(n9828), .A(n9525), .ZN(n9529) );
  INV_X1 U10709 ( .A(n9527), .ZN(n9528) );
  AOI211_X1 U10710 ( .C1(n9835), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9532)
         );
  AOI22_X1 U10711 ( .A1(n4474), .A2(n9532), .B1(n6989), .B2(n9836), .ZN(
        P1_U3484) );
  AOI22_X1 U10712 ( .A1(n9848), .A2(n9532), .B1(n9531), .B2(n9845), .ZN(
        P1_U3533) );
  NOR2_X1 U10713 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9533) );
  AOI21_X1 U10714 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9533), .ZN(n10002) );
  NOR2_X1 U10715 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9534) );
  AOI21_X1 U10716 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9534), .ZN(n10005) );
  NOR2_X1 U10717 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9535) );
  AOI21_X1 U10718 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9535), .ZN(n10008) );
  NOR2_X1 U10719 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9536) );
  AOI21_X1 U10720 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9536), .ZN(n10011) );
  NOR2_X1 U10721 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9537) );
  AOI21_X1 U10722 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9537), .ZN(n10014) );
  NOR2_X1 U10723 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9545) );
  XNOR2_X1 U10724 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10416) );
  NAND2_X1 U10725 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n9543) );
  INV_X1 U10726 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U10727 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .B1(n10263), .B2(n10171), .ZN(n10414) );
  NAND2_X1 U10728 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9541) );
  AOI22_X1 U10729 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .B1(n10090), .B2(n9538), .ZN(n10412) );
  AOI21_X1 U10730 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9996) );
  INV_X1 U10731 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9539) );
  NAND3_X1 U10732 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9998) );
  OAI21_X1 U10733 ( .B1(n9996), .B2(n9539), .A(n9998), .ZN(n10411) );
  NAND2_X1 U10734 ( .A1(n10412), .A2(n10411), .ZN(n9540) );
  NAND2_X1 U10735 ( .A1(n9541), .A2(n9540), .ZN(n10413) );
  NAND2_X1 U10736 ( .A1(n10414), .A2(n10413), .ZN(n9542) );
  NAND2_X1 U10737 ( .A1(n9543), .A2(n9542), .ZN(n10415) );
  NOR2_X1 U10738 ( .A1(n10416), .A2(n10415), .ZN(n9544) );
  NOR2_X1 U10739 ( .A1(n9545), .A2(n9544), .ZN(n9546) );
  NOR2_X1 U10740 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9546), .ZN(n10400) );
  AND2_X1 U10741 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9546), .ZN(n10399) );
  NOR2_X1 U10742 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10399), .ZN(n9547) );
  NOR2_X1 U10743 ( .A1(n10400), .A2(n9547), .ZN(n9548) );
  NAND2_X1 U10744 ( .A1(n9548), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9550) );
  XOR2_X1 U10745 ( .A(n9548), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10398) );
  NAND2_X1 U10746 ( .A1(n10398), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U10747 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  NAND2_X1 U10748 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9551), .ZN(n9553) );
  XOR2_X1 U10749 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9551), .Z(n10410) );
  NAND2_X1 U10750 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10410), .ZN(n9552) );
  NAND2_X1 U10751 ( .A1(n9553), .A2(n9552), .ZN(n9554) );
  NAND2_X1 U10752 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9554), .ZN(n9556) );
  XOR2_X1 U10753 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9554), .Z(n10409) );
  NAND2_X1 U10754 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10409), .ZN(n9555) );
  NAND2_X1 U10755 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  AND2_X1 U10756 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9557), .ZN(n9558) );
  INV_X1 U10757 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10408) );
  XNOR2_X1 U10758 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9557), .ZN(n10407) );
  NAND2_X1 U10759 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9559) );
  OAI21_X1 U10760 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9559), .ZN(n10022) );
  NAND2_X1 U10761 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9560) );
  OAI21_X1 U10762 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9560), .ZN(n10019) );
  AOI21_X1 U10763 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10018), .ZN(n10017) );
  NOR2_X1 U10764 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n9561) );
  AOI21_X1 U10765 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9561), .ZN(n10016) );
  NAND2_X1 U10766 ( .A1(n10017), .A2(n10016), .ZN(n10015) );
  OAI21_X1 U10767 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10015), .ZN(n10013) );
  NAND2_X1 U10768 ( .A1(n10014), .A2(n10013), .ZN(n10012) );
  OAI21_X1 U10769 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10012), .ZN(n10010) );
  NAND2_X1 U10770 ( .A1(n10011), .A2(n10010), .ZN(n10009) );
  OAI21_X1 U10771 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10009), .ZN(n10007) );
  NAND2_X1 U10772 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  OAI21_X1 U10773 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10006), .ZN(n10004) );
  NAND2_X1 U10774 ( .A1(n10005), .A2(n10004), .ZN(n10003) );
  OAI21_X1 U10775 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10003), .ZN(n10001) );
  NAND2_X1 U10776 ( .A1(n10002), .A2(n10001), .ZN(n10000) );
  OAI21_X1 U10777 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10000), .ZN(n10403) );
  NOR2_X1 U10778 ( .A1(n10404), .A2(n10403), .ZN(n9562) );
  NAND2_X1 U10779 ( .A1(n10404), .A2(n10403), .ZN(n10402) );
  OAI21_X1 U10780 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9562), .A(n10402), .ZN(
        n9564) );
  XOR2_X1 U10781 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9563) );
  XNOR2_X1 U10782 ( .A(n9564), .B(n9563), .ZN(ADD_1071_U4) );
  INV_X1 U10783 ( .A(n9565), .ZN(n9583) );
  OAI21_X1 U10784 ( .B1(n9566), .B2(n9574), .A(n9567), .ZN(n9597) );
  INV_X1 U10785 ( .A(n9569), .ZN(n9570) );
  OAI211_X1 U10786 ( .C1(n4602), .C2(n9570), .A(n4491), .B(n9963), .ZN(n9594)
         );
  INV_X1 U10787 ( .A(n9571), .ZN(n9572) );
  OAI22_X1 U10788 ( .A1(n9594), .A2(n9573), .B1(n4602), .B2(n9572), .ZN(n9582)
         );
  XNOR2_X1 U10789 ( .A(n9575), .B(n9574), .ZN(n9577) );
  OAI222_X1 U10790 ( .A1(n9581), .A2(n9580), .B1(n9579), .B2(n9578), .C1(n9577), .C2(n9576), .ZN(n9595) );
  AOI211_X1 U10791 ( .C1(n9583), .C2(n9597), .A(n9582), .B(n9595), .ZN(n9592)
         );
  INV_X1 U10792 ( .A(n9584), .ZN(n9588) );
  INV_X1 U10793 ( .A(n9585), .ZN(n9587) );
  AOI22_X1 U10794 ( .A1(n9597), .A2(n9588), .B1(n9587), .B2(n9586), .ZN(n9589)
         );
  OAI221_X1 U10795 ( .B1(n9593), .B2(n9592), .C1(n9591), .C2(n9590), .A(n9589), 
        .ZN(P2_U3279) );
  OAI21_X1 U10796 ( .B1(n4602), .B2(n9971), .A(n9594), .ZN(n9596) );
  AOI211_X1 U10797 ( .C1(n9978), .C2(n9597), .A(n9596), .B(n9595), .ZN(n9622)
         );
  AOI22_X1 U10798 ( .A1(n9995), .A2(n9622), .B1(n7186), .B2(n9993), .ZN(
        P2_U3537) );
  INV_X1 U10799 ( .A(n9618), .ZN(n9959) );
  INV_X1 U10800 ( .A(n9598), .ZN(n9603) );
  OAI22_X1 U10801 ( .A1(n9600), .A2(n9973), .B1(n9599), .B2(n9971), .ZN(n9602)
         );
  AOI211_X1 U10802 ( .C1(n9959), .C2(n9603), .A(n9602), .B(n9601), .ZN(n9623)
         );
  AOI22_X1 U10803 ( .A1(n9995), .A2(n9623), .B1(n6962), .B2(n9993), .ZN(
        P2_U3536) );
  OAI22_X1 U10804 ( .A1(n9605), .A2(n9973), .B1(n9604), .B2(n9971), .ZN(n9607)
         );
  AOI211_X1 U10805 ( .C1(n9978), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9625)
         );
  AOI22_X1 U10806 ( .A1(n9995), .A2(n9625), .B1(n5462), .B2(n9993), .ZN(
        P2_U3535) );
  OAI22_X1 U10807 ( .A1(n9610), .A2(n9973), .B1(n4594), .B2(n9971), .ZN(n9612)
         );
  AOI211_X1 U10808 ( .C1(n9978), .C2(n9613), .A(n9612), .B(n9611), .ZN(n9626)
         );
  AOI22_X1 U10809 ( .A1(n9995), .A2(n9626), .B1(n9614), .B2(n9993), .ZN(
        P2_U3534) );
  AOI22_X1 U10810 ( .A1(n9616), .A2(n9963), .B1(n9962), .B2(n9615), .ZN(n9617)
         );
  OAI21_X1 U10811 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(n9620) );
  NOR2_X1 U10812 ( .A1(n9621), .A2(n9620), .ZN(n9627) );
  AOI22_X1 U10813 ( .A1(n9995), .A2(n9627), .B1(n5409), .B2(n9993), .ZN(
        P2_U3533) );
  AOI22_X1 U10814 ( .A1(n9979), .A2(n9622), .B1(n5505), .B2(n4579), .ZN(
        P2_U3502) );
  AOI22_X1 U10815 ( .A1(n9979), .A2(n9623), .B1(n5483), .B2(n4579), .ZN(
        P2_U3499) );
  INV_X1 U10816 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9624) );
  AOI22_X1 U10817 ( .A1(n9979), .A2(n9625), .B1(n9624), .B2(n4579), .ZN(
        P2_U3496) );
  AOI22_X1 U10818 ( .A1(n9979), .A2(n9626), .B1(n5431), .B2(n4579), .ZN(
        P2_U3493) );
  INV_X1 U10819 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U10820 ( .A1(n9979), .A2(n9627), .B1(n10278), .B2(n4579), .ZN(
        P2_U3490) );
  OAI22_X1 U10821 ( .A1(n9629), .A2(n9830), .B1(n9628), .B2(n9828), .ZN(n9630)
         );
  AOI21_X1 U10822 ( .B1(n9631), .B2(n9835), .A(n9630), .ZN(n9632) );
  AND2_X1 U10823 ( .A1(n9633), .A2(n9632), .ZN(n9641) );
  AOI22_X1 U10824 ( .A1(n9848), .A2(n9641), .B1(n5957), .B2(n9845), .ZN(
        P1_U3536) );
  INV_X1 U10825 ( .A(n9634), .ZN(n9636) );
  OAI21_X1 U10826 ( .B1(n9636), .B2(n9828), .A(n9635), .ZN(n9637) );
  AOI21_X1 U10827 ( .B1(n9638), .B2(n9835), .A(n9637), .ZN(n9639) );
  AND2_X1 U10828 ( .A1(n9640), .A2(n9639), .ZN(n9642) );
  AOI22_X1 U10829 ( .A1(n9848), .A2(n9642), .B1(n7070), .B2(n9845), .ZN(
        P1_U3535) );
  AOI22_X1 U10830 ( .A1(n4474), .A2(n9641), .B1(n7143), .B2(n9836), .ZN(
        P1_U3493) );
  AOI22_X1 U10831 ( .A1(n4474), .A2(n9642), .B1(n7074), .B2(n9836), .ZN(
        P1_U3490) );
  XNOR2_X1 U10832 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10833 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10834 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9656) );
  OAI21_X1 U10835 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(n9647) );
  AOI22_X1 U10836 ( .A1(n9740), .A2(n9647), .B1(n9742), .B2(n9646), .ZN(n9655)
         );
  OAI21_X1 U10837 ( .B1(n9650), .B2(n9649), .A(n9648), .ZN(n9653) );
  AOI211_X1 U10838 ( .C1(n9750), .C2(n9653), .A(n9652), .B(n9651), .ZN(n9654)
         );
  OAI211_X1 U10839 ( .C1(n9735), .C2(n9656), .A(n9655), .B(n9654), .ZN(
        P1_U3245) );
  AOI211_X1 U10840 ( .C1(n9660), .C2(n9659), .A(n9658), .B(n9657), .ZN(n9661)
         );
  AOI211_X1 U10841 ( .C1(n9742), .C2(n9663), .A(n9662), .B(n9661), .ZN(n9669)
         );
  OAI21_X1 U10842 ( .B1(n9666), .B2(n9665), .A(n9664), .ZN(n9667) );
  AOI22_X1 U10843 ( .A1(n9740), .A2(n9667), .B1(n9749), .B2(
        P1_ADDR_REG_5__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U10844 ( .A1(n9669), .A2(n9668), .ZN(P1_U3246) );
  OAI21_X1 U10845 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n9678) );
  AOI211_X1 U10846 ( .C1(n9675), .C2(n9674), .A(n9673), .B(n9713), .ZN(n9676)
         );
  AOI211_X1 U10847 ( .C1(n9750), .C2(n9678), .A(n9677), .B(n9676), .ZN(n9681)
         );
  AOI22_X1 U10848 ( .A1(n9742), .A2(n9679), .B1(n9749), .B2(
        P1_ADDR_REG_6__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U10849 ( .A1(n9681), .A2(n9680), .ZN(P1_U3247) );
  NAND2_X1 U10850 ( .A1(n9742), .A2(n9682), .ZN(n9691) );
  INV_X1 U10851 ( .A(n9683), .ZN(n9690) );
  NAND2_X1 U10852 ( .A1(n9685), .A2(n9684), .ZN(n9688) );
  INV_X1 U10853 ( .A(n9686), .ZN(n9687) );
  NAND3_X1 U10854 ( .A1(n9750), .A2(n9688), .A3(n9687), .ZN(n9689) );
  AND3_X1 U10855 ( .A1(n9691), .A2(n9690), .A3(n9689), .ZN(n9697) );
  OAI21_X1 U10856 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9695) );
  AOI22_X1 U10857 ( .A1(n9740), .A2(n9695), .B1(n9749), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U10858 ( .A1(n9697), .A2(n9696), .ZN(P1_U3249) );
  OAI21_X1 U10859 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9706) );
  AOI211_X1 U10860 ( .C1(n9703), .C2(n9702), .A(n9701), .B(n9713), .ZN(n9704)
         );
  AOI211_X1 U10861 ( .C1(n9750), .C2(n9706), .A(n9705), .B(n9704), .ZN(n9709)
         );
  AOI22_X1 U10862 ( .A1(n9742), .A2(n9707), .B1(n9749), .B2(
        P1_ADDR_REG_9__SCAN_IN), .ZN(n9708) );
  NAND2_X1 U10863 ( .A1(n9709), .A2(n9708), .ZN(P1_U3250) );
  OAI21_X1 U10864 ( .B1(n9712), .B2(n9711), .A(n9710), .ZN(n9719) );
  AOI211_X1 U10865 ( .C1(n9716), .C2(n9715), .A(n9714), .B(n9713), .ZN(n9717)
         );
  AOI211_X1 U10866 ( .C1(n9750), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9722)
         );
  AOI22_X1 U10867 ( .A1(n9742), .A2(n9720), .B1(n9749), .B2(
        P1_ADDR_REG_10__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U10868 ( .A1(n9722), .A2(n9721), .ZN(P1_U3251) );
  INV_X1 U10869 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10147) );
  AOI21_X1 U10870 ( .B1(n9742), .B2(n9724), .A(n9723), .ZN(n9734) );
  OAI21_X1 U10871 ( .B1(n9727), .B2(n9726), .A(n9725), .ZN(n9732) );
  OAI21_X1 U10872 ( .B1(n9730), .B2(n9729), .A(n9728), .ZN(n9731) );
  AOI22_X1 U10873 ( .A1(n9732), .A2(n9750), .B1(n9740), .B2(n9731), .ZN(n9733)
         );
  OAI211_X1 U10874 ( .C1(n9735), .C2(n10147), .A(n9734), .B(n9733), .ZN(
        P1_U3252) );
  AOI21_X1 U10875 ( .B1(n9738), .B2(n9737), .A(n9736), .ZN(n9739) );
  NAND2_X1 U10876 ( .A1(n9740), .A2(n9739), .ZN(n9745) );
  NAND2_X1 U10877 ( .A1(n9742), .A2(n9741), .ZN(n9744) );
  AND3_X1 U10878 ( .A1(n9745), .A2(n9744), .A3(n9743), .ZN(n9753) );
  OAI21_X1 U10879 ( .B1(n9748), .B2(n9747), .A(n9746), .ZN(n9751) );
  AOI22_X1 U10880 ( .A1(n9751), .A2(n9750), .B1(n9749), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U10881 ( .A1(n9753), .A2(n9752), .ZN(P1_U3259) );
  OAI22_X1 U10882 ( .A1(n9755), .A2(n9784), .B1(n9790), .B2(n9754), .ZN(n9756)
         );
  AOI21_X1 U10883 ( .B1(n9757), .B2(n4473), .A(n9756), .ZN(n9758) );
  OAI211_X1 U10884 ( .C1(n9761), .C2(n9760), .A(n9759), .B(n9758), .ZN(n9762)
         );
  INV_X1 U10885 ( .A(n9762), .ZN(n9763) );
  AOI22_X1 U10886 ( .A1(n9767), .A2(n6481), .B1(n9763), .B2(n9786), .ZN(
        P1_U3286) );
  NAND2_X1 U10887 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  XNOR2_X1 U10888 ( .A(n9766), .B(n4513), .ZN(n9780) );
  INV_X1 U10889 ( .A(n9780), .ZN(n9811) );
  AOI22_X1 U10890 ( .A1(n9811), .A2(n9768), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n9767), .ZN(n9789) );
  OAI21_X1 U10891 ( .B1(n4513), .B2(n9770), .A(n9769), .ZN(n9777) );
  OAI22_X1 U10892 ( .A1(n9774), .A2(n9773), .B1(n9772), .B2(n9771), .ZN(n9775)
         );
  AOI21_X1 U10893 ( .B1(n9777), .B2(n9776), .A(n9775), .ZN(n9778) );
  OAI21_X1 U10894 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(n9809) );
  OAI211_X1 U10895 ( .C1(n9783), .C2(n9808), .A(n9782), .B(n9781), .ZN(n9807)
         );
  OAI22_X1 U10896 ( .A1(n9807), .A2(n9785), .B1(n9808), .B2(n9784), .ZN(n9787)
         );
  OAI21_X1 U10897 ( .B1(n9809), .B2(n9787), .A(n9786), .ZN(n9788) );
  OAI211_X1 U10898 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9788), .ZN(
        P1_U3287) );
  INV_X1 U10899 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10258) );
  NOR2_X1 U10900 ( .A1(n9794), .A2(n10258), .ZN(P1_U3292) );
  AND2_X1 U10901 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10024), .ZN(P1_U3293) );
  INV_X1 U10902 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10087) );
  NOR2_X1 U10903 ( .A1(n9794), .A2(n10087), .ZN(P1_U3294) );
  AND2_X1 U10904 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10024), .ZN(P1_U3295) );
  INV_X1 U10905 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10303) );
  NOR2_X1 U10906 ( .A1(n9794), .A2(n10303), .ZN(P1_U3296) );
  AND2_X1 U10907 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10024), .ZN(P1_U3297) );
  AND2_X1 U10908 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10024), .ZN(P1_U3298) );
  INV_X1 U10909 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10282) );
  NOR2_X1 U10910 ( .A1(n9794), .A2(n10282), .ZN(P1_U3299) );
  AND2_X1 U10911 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10024), .ZN(P1_U3300) );
  AND2_X1 U10912 ( .A1(n10024), .A2(P1_D_REG_22__SCAN_IN), .ZN(P1_U3301) );
  AND2_X1 U10913 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10024), .ZN(P1_U3302) );
  AND2_X1 U10914 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10024), .ZN(P1_U3303) );
  INV_X1 U10915 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10295) );
  NOR2_X1 U10916 ( .A1(n9794), .A2(n10295), .ZN(P1_U3304) );
  AND2_X1 U10917 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10024), .ZN(P1_U3305) );
  AND2_X1 U10918 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10024), .ZN(P1_U3306) );
  AND2_X1 U10919 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10024), .ZN(P1_U3307) );
  AND2_X1 U10920 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10024), .ZN(P1_U3308) );
  AND2_X1 U10921 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10024), .ZN(P1_U3309) );
  AND2_X1 U10922 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10024), .ZN(P1_U3310) );
  AND2_X1 U10923 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10024), .ZN(P1_U3311) );
  AND2_X1 U10924 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10024), .ZN(P1_U3312) );
  INV_X1 U10925 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10163) );
  NOR2_X1 U10926 ( .A1(n9794), .A2(n10163), .ZN(P1_U3313) );
  AND2_X1 U10927 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10024), .ZN(P1_U3314) );
  AND2_X1 U10928 ( .A1(n10024), .A2(P1_D_REG_7__SCAN_IN), .ZN(P1_U3316) );
  AND2_X1 U10929 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10024), .ZN(P1_U3317) );
  AND2_X1 U10930 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10024), .ZN(P1_U3318) );
  AND2_X1 U10931 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10024), .ZN(P1_U3319) );
  AND2_X1 U10932 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10024), .ZN(P1_U3320) );
  AND2_X1 U10933 ( .A1(n10024), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3321) );
  INV_X1 U10934 ( .A(n9795), .ZN(n9800) );
  OAI21_X1 U10935 ( .B1(n9797), .B2(n9828), .A(n9796), .ZN(n9799) );
  AOI211_X1 U10936 ( .C1(n9835), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9838)
         );
  AOI22_X1 U10937 ( .A1(n4474), .A2(n9838), .B1(n6229), .B2(n9836), .ZN(
        P1_U3457) );
  INV_X1 U10938 ( .A(n9801), .ZN(n9806) );
  OAI22_X1 U10939 ( .A1(n9803), .A2(n9830), .B1(n9802), .B2(n9828), .ZN(n9805)
         );
  AOI211_X1 U10940 ( .C1(n9835), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9840)
         );
  AOI22_X1 U10941 ( .A1(n4474), .A2(n9840), .B1(n6272), .B2(n9836), .ZN(
        P1_U3460) );
  OAI21_X1 U10942 ( .B1(n9808), .B2(n9828), .A(n9807), .ZN(n9810) );
  AOI211_X1 U10943 ( .C1(n9835), .C2(n9811), .A(n9810), .B(n9809), .ZN(n9842)
         );
  INV_X1 U10944 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9812) );
  AOI22_X1 U10945 ( .A1(n4474), .A2(n9842), .B1(n9812), .B2(n9836), .ZN(
        P1_U3466) );
  OAI22_X1 U10946 ( .A1(n9814), .A2(n9830), .B1(n9813), .B2(n9828), .ZN(n9816)
         );
  AOI211_X1 U10947 ( .C1(n9835), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9843)
         );
  INV_X1 U10948 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U10949 ( .A1(n4474), .A2(n9843), .B1(n9818), .B2(n9836), .ZN(
        P1_U3472) );
  INV_X1 U10950 ( .A(n9819), .ZN(n9825) );
  OAI22_X1 U10951 ( .A1(n9821), .A2(n9830), .B1(n9820), .B2(n9828), .ZN(n9823)
         );
  AOI211_X1 U10952 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9844)
         );
  INV_X1 U10953 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9826) );
  AOI22_X1 U10954 ( .A1(n4474), .A2(n9844), .B1(n9826), .B2(n9836), .ZN(
        P1_U3478) );
  INV_X1 U10955 ( .A(n9827), .ZN(n9834) );
  OAI22_X1 U10956 ( .A1(n9831), .A2(n9830), .B1(n9829), .B2(n9828), .ZN(n9833)
         );
  AOI211_X1 U10957 ( .C1(n9835), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9847)
         );
  AOI22_X1 U10958 ( .A1(n4474), .A2(n9847), .B1(n6759), .B2(n9836), .ZN(
        P1_U3481) );
  AOI22_X1 U10959 ( .A1(n9848), .A2(n9838), .B1(n9837), .B2(n9845), .ZN(
        P1_U3524) );
  AOI22_X1 U10960 ( .A1(n9848), .A2(n9840), .B1(n9839), .B2(n9845), .ZN(
        P1_U3525) );
  INV_X1 U10961 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9841) );
  AOI22_X1 U10962 ( .A1(n9848), .A2(n9842), .B1(n9841), .B2(n9845), .ZN(
        P1_U3527) );
  AOI22_X1 U10963 ( .A1(n9848), .A2(n9843), .B1(n6645), .B2(n9845), .ZN(
        P1_U3529) );
  AOI22_X1 U10964 ( .A1(n9848), .A2(n9844), .B1(n6741), .B2(n9845), .ZN(
        P1_U3531) );
  INV_X1 U10965 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9846) );
  AOI22_X1 U10966 ( .A1(n9848), .A2(n9847), .B1(n9846), .B2(n9845), .ZN(
        P1_U3532) );
  AOI22_X1 U10967 ( .A1(n9850), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9849), .ZN(n9860) );
  NAND2_X1 U10968 ( .A1(n9851), .A2(n5082), .ZN(n9853) );
  OAI211_X1 U10969 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9854), .A(n9853), .B(
        n9852), .ZN(n9855) );
  INV_X1 U10970 ( .A(n9855), .ZN(n9859) );
  AOI21_X1 U10971 ( .B1(n9857), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n9856), .ZN(
        n9858) );
  OAI221_X1 U10972 ( .B1(n9861), .B2(n9860), .C1(n5098), .C2(n9859), .A(n9858), 
        .ZN(P2_U3245) );
  XNOR2_X1 U10973 ( .A(n9863), .B(n9862), .ZN(n9867) );
  AOI222_X1 U10974 ( .A1(n9868), .A2(n9867), .B1(n9866), .B2(n9865), .C1(n5855), .C2(n9864), .ZN(n9921) );
  NOR2_X1 U10975 ( .A1(n8436), .A2(n6109), .ZN(n9875) );
  XNOR2_X1 U10976 ( .A(n9870), .B(n9869), .ZN(n9920) );
  OAI22_X1 U10977 ( .A1(n9873), .A2(n9920), .B1(n9872), .B2(n9871), .ZN(n9874)
         );
  NOR2_X1 U10978 ( .A1(n9875), .A2(n9874), .ZN(n9880) );
  XNOR2_X1 U10979 ( .A(n9877), .B(n9876), .ZN(n9924) );
  NAND2_X1 U10980 ( .A1(n9878), .A2(n9924), .ZN(n9879) );
  OAI211_X1 U10981 ( .C1(n9919), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9882)
         );
  INV_X1 U10982 ( .A(n9882), .ZN(n9883) );
  OAI21_X1 U10983 ( .B1(n9884), .B2(n9921), .A(n9883), .ZN(P2_U3292) );
  AND2_X1 U10984 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9890), .ZN(P2_U3297) );
  AND2_X1 U10985 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9890), .ZN(P2_U3298) );
  AND2_X1 U10986 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9890), .ZN(P2_U3299) );
  AND2_X1 U10987 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9890), .ZN(P2_U3300) );
  AND2_X1 U10988 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9890), .ZN(P2_U3301) );
  AND2_X1 U10989 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9890), .ZN(P2_U3302) );
  AND2_X1 U10990 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9890), .ZN(P2_U3303) );
  AND2_X1 U10991 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9890), .ZN(P2_U3304) );
  INV_X1 U10992 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U10993 ( .A1(n9887), .A2(n10231), .ZN(P2_U3305) );
  AND2_X1 U10994 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9890), .ZN(P2_U3306) );
  INV_X1 U10995 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10089) );
  NOR2_X1 U10996 ( .A1(n9887), .A2(n10089), .ZN(P2_U3307) );
  INV_X1 U10997 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U10998 ( .A1(n9887), .A2(n10198), .ZN(P2_U3308) );
  AND2_X1 U10999 ( .A1(n9890), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3309) );
  AND2_X1 U11000 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9890), .ZN(P2_U3310) );
  AND2_X1 U11001 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9890), .ZN(P2_U3311) );
  AND2_X1 U11002 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9890), .ZN(P2_U3312) );
  AND2_X1 U11003 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9890), .ZN(P2_U3313) );
  INV_X1 U11004 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10227) );
  NOR2_X1 U11005 ( .A1(n9887), .A2(n10227), .ZN(P2_U3314) );
  AND2_X1 U11006 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9890), .ZN(P2_U3315) );
  AND2_X1 U11007 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9890), .ZN(P2_U3316) );
  AND2_X1 U11008 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9890), .ZN(P2_U3317) );
  AND2_X1 U11009 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9890), .ZN(P2_U3318) );
  AND2_X1 U11010 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9890), .ZN(P2_U3319) );
  AND2_X1 U11011 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9890), .ZN(P2_U3320) );
  INV_X1 U11012 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10276) );
  NOR2_X1 U11013 ( .A1(n9887), .A2(n10276), .ZN(P2_U3321) );
  INV_X1 U11014 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10216) );
  NOR2_X1 U11015 ( .A1(n9887), .A2(n10216), .ZN(P2_U3322) );
  AND2_X1 U11016 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9890), .ZN(P2_U3323) );
  AND2_X1 U11017 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9890), .ZN(P2_U3324) );
  INV_X1 U11018 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10306) );
  NOR2_X1 U11019 ( .A1(n9887), .A2(n10306), .ZN(P2_U3325) );
  AND2_X1 U11020 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9890), .ZN(P2_U3326) );
  AOI22_X1 U11021 ( .A1(n9892), .A2(n9889), .B1(n9888), .B2(n9890), .ZN(
        P2_U3437) );
  AOI22_X1 U11022 ( .A1(n9892), .A2(n9891), .B1(n10293), .B2(n9890), .ZN(
        P2_U3438) );
  INV_X1 U11023 ( .A(n9893), .ZN(n9898) );
  OAI22_X1 U11024 ( .A1(n9896), .A2(n9966), .B1(n9895), .B2(n9894), .ZN(n9897)
         );
  NOR2_X1 U11025 ( .A1(n9898), .A2(n9897), .ZN(n9981) );
  AOI22_X1 U11026 ( .A1(n9979), .A2(n9981), .B1(n5085), .B2(n4579), .ZN(
        P2_U3451) );
  NOR3_X1 U11027 ( .A1(n9900), .A2(n9899), .A3(n9973), .ZN(n9901) );
  AOI21_X1 U11028 ( .B1(n9962), .B2(n9902), .A(n9901), .ZN(n9903) );
  OAI211_X1 U11029 ( .C1(n9966), .C2(n9905), .A(n9904), .B(n9903), .ZN(n9906)
         );
  INV_X1 U11030 ( .A(n9906), .ZN(n9982) );
  AOI22_X1 U11031 ( .A1(n9979), .A2(n9982), .B1(n5124), .B2(n4579), .ZN(
        P2_U3454) );
  NOR2_X1 U11032 ( .A1(n9907), .A2(n9966), .ZN(n9911) );
  OAI22_X1 U11033 ( .A1(n9909), .A2(n9973), .B1(n9908), .B2(n9971), .ZN(n9910)
         );
  NOR3_X1 U11034 ( .A1(n9912), .A2(n9911), .A3(n9910), .ZN(n9983) );
  AOI22_X1 U11035 ( .A1(n9979), .A2(n9983), .B1(n5144), .B2(n4579), .ZN(
        P2_U3457) );
  INV_X1 U11036 ( .A(n9913), .ZN(n9918) );
  OAI22_X1 U11037 ( .A1(n9915), .A2(n9973), .B1(n9914), .B2(n9971), .ZN(n9917)
         );
  AOI211_X1 U11038 ( .C1(n9959), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9985)
         );
  AOI22_X1 U11039 ( .A1(n9979), .A2(n9985), .B1(n5153), .B2(n4579), .ZN(
        P2_U3460) );
  OAI22_X1 U11040 ( .A1(n9920), .A2(n9973), .B1(n9919), .B2(n9971), .ZN(n9923)
         );
  INV_X1 U11041 ( .A(n9921), .ZN(n9922) );
  AOI211_X1 U11042 ( .C1(n9978), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9986)
         );
  INV_X1 U11043 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U11044 ( .A1(n9979), .A2(n9986), .B1(n9925), .B2(n4579), .ZN(
        P2_U3463) );
  AOI22_X1 U11045 ( .A1(n9927), .A2(n9963), .B1(n9962), .B2(n9926), .ZN(n9930)
         );
  OR2_X1 U11046 ( .A1(n9928), .A2(n9966), .ZN(n9929) );
  AND3_X1 U11047 ( .A1(n9931), .A2(n9930), .A3(n9929), .ZN(n9987) );
  INV_X1 U11048 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U11049 ( .A1(n9979), .A2(n9987), .B1(n9932), .B2(n4579), .ZN(
        P2_U3469) );
  AOI22_X1 U11050 ( .A1(n9934), .A2(n9963), .B1(n9962), .B2(n9933), .ZN(n9935)
         );
  OAI211_X1 U11051 ( .C1(n9966), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9938)
         );
  INV_X1 U11052 ( .A(n9938), .ZN(n9988) );
  INV_X1 U11053 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9939) );
  AOI22_X1 U11054 ( .A1(n9979), .A2(n9988), .B1(n9939), .B2(n4579), .ZN(
        P2_U3472) );
  INV_X1 U11055 ( .A(n9940), .ZN(n9945) );
  OAI22_X1 U11056 ( .A1(n9942), .A2(n9973), .B1(n9941), .B2(n9971), .ZN(n9944)
         );
  AOI211_X1 U11057 ( .C1(n9959), .C2(n9945), .A(n9944), .B(n9943), .ZN(n9989)
         );
  INV_X1 U11058 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9946) );
  AOI22_X1 U11059 ( .A1(n9979), .A2(n9989), .B1(n9946), .B2(n4579), .ZN(
        P2_U3475) );
  INV_X1 U11060 ( .A(n9947), .ZN(n9952) );
  OAI22_X1 U11061 ( .A1(n9949), .A2(n9973), .B1(n9948), .B2(n9971), .ZN(n9951)
         );
  AOI211_X1 U11062 ( .C1(n9959), .C2(n9952), .A(n9951), .B(n9950), .ZN(n9990)
         );
  AOI22_X1 U11063 ( .A1(n9979), .A2(n9990), .B1(n5311), .B2(n4579), .ZN(
        P2_U3478) );
  INV_X1 U11064 ( .A(n9953), .ZN(n9958) );
  OAI22_X1 U11065 ( .A1(n9955), .A2(n9973), .B1(n9954), .B2(n9971), .ZN(n9957)
         );
  AOI211_X1 U11066 ( .C1(n9959), .C2(n9958), .A(n9957), .B(n9956), .ZN(n9991)
         );
  INV_X1 U11067 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U11068 ( .A1(n9979), .A2(n9991), .B1(n9960), .B2(n4579), .ZN(
        P2_U3481) );
  AOI22_X1 U11069 ( .A1(n9964), .A2(n9963), .B1(n9962), .B2(n9961), .ZN(n9965)
         );
  OAI21_X1 U11070 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(n9968) );
  NOR2_X1 U11071 ( .A1(n9969), .A2(n9968), .ZN(n9992) );
  INV_X1 U11072 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11073 ( .A1(n9979), .A2(n9992), .B1(n9970), .B2(n4579), .ZN(
        P2_U3484) );
  OAI22_X1 U11074 ( .A1(n9974), .A2(n9973), .B1(n9972), .B2(n9971), .ZN(n9976)
         );
  AOI211_X1 U11075 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9994)
         );
  AOI22_X1 U11076 ( .A1(n9979), .A2(n9994), .B1(n5384), .B2(n4579), .ZN(
        P2_U3487) );
  INV_X1 U11077 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U11078 ( .A1(n9995), .A2(n9981), .B1(n9980), .B2(n9993), .ZN(
        P2_U3520) );
  AOI22_X1 U11079 ( .A1(n9995), .A2(n9982), .B1(n6080), .B2(n9993), .ZN(
        P2_U3521) );
  AOI22_X1 U11080 ( .A1(n9995), .A2(n9983), .B1(n6081), .B2(n9993), .ZN(
        P2_U3522) );
  INV_X1 U11081 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U11082 ( .A1(n9995), .A2(n9985), .B1(n9984), .B2(n9993), .ZN(
        P2_U3523) );
  AOI22_X1 U11083 ( .A1(n9995), .A2(n9986), .B1(n6079), .B2(n9993), .ZN(
        P2_U3524) );
  AOI22_X1 U11084 ( .A1(n9995), .A2(n9987), .B1(n6089), .B2(n9993), .ZN(
        P2_U3526) );
  AOI22_X1 U11085 ( .A1(n9995), .A2(n9988), .B1(n5253), .B2(n9993), .ZN(
        P2_U3527) );
  AOI22_X1 U11086 ( .A1(n9995), .A2(n9989), .B1(n6093), .B2(n9993), .ZN(
        P2_U3528) );
  AOI22_X1 U11087 ( .A1(n9995), .A2(n9990), .B1(n6094), .B2(n9993), .ZN(
        P2_U3529) );
  AOI22_X1 U11088 ( .A1(n9995), .A2(n9991), .B1(n6123), .B2(n9993), .ZN(
        P2_U3530) );
  AOI22_X1 U11089 ( .A1(n9995), .A2(n9992), .B1(n6288), .B2(n9993), .ZN(
        P2_U3531) );
  AOI22_X1 U11090 ( .A1(n9995), .A2(n9994), .B1(n6307), .B2(n9993), .ZN(
        P2_U3532) );
  INV_X1 U11091 ( .A(n9996), .ZN(n9997) );
  NAND2_X1 U11092 ( .A1(n9998), .A2(n9997), .ZN(n9999) );
  XNOR2_X1 U11093 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9999), .ZN(ADD_1071_U5) );
  XOR2_X1 U11094 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11095 ( .B1(n10002), .B2(n10001), .A(n10000), .ZN(ADD_1071_U56) );
  OAI21_X1 U11096 ( .B1(n10005), .B2(n10004), .A(n10003), .ZN(ADD_1071_U57) );
  OAI21_X1 U11097 ( .B1(n10008), .B2(n10007), .A(n10006), .ZN(ADD_1071_U58) );
  OAI21_X1 U11098 ( .B1(n10011), .B2(n10010), .A(n10009), .ZN(ADD_1071_U59) );
  OAI21_X1 U11099 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(ADD_1071_U60) );
  OAI21_X1 U11100 ( .B1(n10017), .B2(n10016), .A(n10015), .ZN(ADD_1071_U61) );
  AOI21_X1 U11101 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(ADD_1071_U62) );
  AOI21_X1 U11102 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(ADD_1071_U63) );
  NAND2_X1 U11103 ( .A1(n10024), .A2(P1_D_REG_8__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U11104 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput234), .B1(
        P1_REG3_REG_11__SCAN_IN), .B2(keyinput203), .ZN(n10025) );
  OAI221_X1 U11105 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput234), .C1(
        P1_REG3_REG_11__SCAN_IN), .C2(keyinput203), .A(n10025), .ZN(n10032) );
  AOI22_X1 U11106 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(keyinput169), .B1(SI_9_), 
        .B2(keyinput221), .ZN(n10026) );
  OAI221_X1 U11107 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(keyinput169), .C1(SI_9_), 
        .C2(keyinput221), .A(n10026), .ZN(n10031) );
  AOI22_X1 U11108 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput200), .B1(
        P1_REG0_REG_22__SCAN_IN), .B2(keyinput142), .ZN(n10027) );
  OAI221_X1 U11109 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput200), .C1(
        P1_REG0_REG_22__SCAN_IN), .C2(keyinput142), .A(n10027), .ZN(n10030) );
  AOI22_X1 U11110 ( .A1(SI_29_), .A2(keyinput152), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput151), .ZN(n10028) );
  OAI221_X1 U11111 ( .B1(SI_29_), .B2(keyinput152), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput151), .A(n10028), .ZN(n10029)
         );
  NOR4_X1 U11112 ( .A1(n10032), .A2(n10031), .A3(n10030), .A4(n10029), .ZN(
        n10060) );
  AOI22_X1 U11113 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(keyinput189), .B1(SI_23_), 
        .B2(keyinput136), .ZN(n10033) );
  OAI221_X1 U11114 ( .B1(P2_IR_REG_17__SCAN_IN), .B2(keyinput189), .C1(SI_23_), 
        .C2(keyinput136), .A(n10033), .ZN(n10040) );
  AOI22_X1 U11115 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(keyinput179), .B1(
        P1_D_REG_22__SCAN_IN), .B2(keyinput137), .ZN(n10034) );
  OAI221_X1 U11116 ( .B1(P2_IR_REG_13__SCAN_IN), .B2(keyinput179), .C1(
        P1_D_REG_22__SCAN_IN), .C2(keyinput137), .A(n10034), .ZN(n10039) );
  AOI22_X1 U11117 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(keyinput155), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput232), .ZN(n10035) );
  OAI221_X1 U11118 ( .B1(P1_DATAO_REG_2__SCAN_IN), .B2(keyinput155), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput232), .A(n10035), .ZN(n10038) );
  AOI22_X1 U11119 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(keyinput229), .B1(SI_26_), .B2(keyinput223), .ZN(n10036) );
  OAI221_X1 U11120 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(keyinput229), .C1(
        SI_26_), .C2(keyinput223), .A(n10036), .ZN(n10037) );
  NOR4_X1 U11121 ( .A1(n10040), .A2(n10039), .A3(n10038), .A4(n10037), .ZN(
        n10059) );
  AOI22_X1 U11122 ( .A1(P1_REG1_REG_29__SCAN_IN), .A2(keyinput196), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput197), .ZN(n10041) );
  OAI221_X1 U11123 ( .B1(P1_REG1_REG_29__SCAN_IN), .B2(keyinput196), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput197), .A(n10041), .ZN(n10048)
         );
  AOI22_X1 U11124 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(keyinput177), .B1(
        P1_D_REG_7__SCAN_IN), .B2(keyinput168), .ZN(n10042) );
  OAI221_X1 U11125 ( .B1(P2_REG0_REG_14__SCAN_IN), .B2(keyinput177), .C1(
        P1_D_REG_7__SCAN_IN), .C2(keyinput168), .A(n10042), .ZN(n10047) );
  AOI22_X1 U11126 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput134), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(keyinput244), .ZN(n10043) );
  OAI221_X1 U11127 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput134), .C1(
        P1_DATAO_REG_0__SCAN_IN), .C2(keyinput244), .A(n10043), .ZN(n10046) );
  AOI22_X1 U11128 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput224), .B1(
        P2_REG1_REG_13__SCAN_IN), .B2(keyinput170), .ZN(n10044) );
  OAI221_X1 U11129 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput224), .C1(
        P2_REG1_REG_13__SCAN_IN), .C2(keyinput170), .A(n10044), .ZN(n10045) );
  NOR4_X1 U11130 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10058) );
  AOI22_X1 U11131 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput129), .B1(SI_12_), 
        .B2(keyinput199), .ZN(n10049) );
  OAI221_X1 U11132 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput129), .C1(SI_12_), .C2(keyinput199), .A(n10049), .ZN(n10056) );
  AOI22_X1 U11133 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(keyinput130), .B1(
        P2_D_REG_23__SCAN_IN), .B2(keyinput180), .ZN(n10050) );
  OAI221_X1 U11134 ( .B1(P2_REG0_REG_13__SCAN_IN), .B2(keyinput130), .C1(
        P2_D_REG_23__SCAN_IN), .C2(keyinput180), .A(n10050), .ZN(n10055) );
  AOI22_X1 U11135 ( .A1(SI_31_), .A2(keyinput191), .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput216), .ZN(n10051) );
  OAI221_X1 U11136 ( .B1(SI_31_), .B2(keyinput191), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput216), .A(n10051), .ZN(n10054) );
  AOI22_X1 U11137 ( .A1(P2_REG0_REG_12__SCAN_IN), .A2(keyinput213), .B1(
        P2_REG2_REG_19__SCAN_IN), .B2(keyinput230), .ZN(n10052) );
  OAI221_X1 U11138 ( .B1(P2_REG0_REG_12__SCAN_IN), .B2(keyinput213), .C1(
        P2_REG2_REG_19__SCAN_IN), .C2(keyinput230), .A(n10052), .ZN(n10053) );
  NOR4_X1 U11139 ( .A1(n10056), .A2(n10055), .A3(n10054), .A4(n10053), .ZN(
        n10057) );
  NAND4_X1 U11140 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10196) );
  AOI22_X1 U11141 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(keyinput233), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput160), .ZN(n10061) );
  OAI221_X1 U11142 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(keyinput233), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput160), .A(n10061), .ZN(n10068) );
  AOI22_X1 U11143 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(keyinput254), .B1(
        P1_REG3_REG_23__SCAN_IN), .B2(keyinput210), .ZN(n10062) );
  OAI221_X1 U11144 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(keyinput254), .C1(
        P1_REG3_REG_23__SCAN_IN), .C2(keyinput210), .A(n10062), .ZN(n10067) );
  AOI22_X1 U11145 ( .A1(P1_REG0_REG_21__SCAN_IN), .A2(keyinput193), .B1(SI_15_), .B2(keyinput128), .ZN(n10063) );
  OAI221_X1 U11146 ( .B1(P1_REG0_REG_21__SCAN_IN), .B2(keyinput193), .C1(
        SI_15_), .C2(keyinput128), .A(n10063), .ZN(n10066) );
  AOI22_X1 U11147 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(keyinput173), .B1(
        P1_REG1_REG_26__SCAN_IN), .B2(keyinput240), .ZN(n10064) );
  OAI221_X1 U11148 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(keyinput173), .C1(
        P1_REG1_REG_26__SCAN_IN), .C2(keyinput240), .A(n10064), .ZN(n10065) );
  NOR4_X1 U11149 ( .A1(n10068), .A2(n10067), .A3(n10066), .A4(n10065), .ZN(
        n10099) );
  AOI22_X1 U11150 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(keyinput236), .B1(
        P1_D_REG_24__SCAN_IN), .B2(keyinput141), .ZN(n10069) );
  OAI221_X1 U11151 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(keyinput236), .C1(
        P1_D_REG_24__SCAN_IN), .C2(keyinput141), .A(n10069), .ZN(n10076) );
  AOI22_X1 U11152 ( .A1(P2_D_REG_6__SCAN_IN), .A2(keyinput249), .B1(
        P1_REG1_REG_28__SCAN_IN), .B2(keyinput198), .ZN(n10070) );
  OAI221_X1 U11153 ( .B1(P2_D_REG_6__SCAN_IN), .B2(keyinput249), .C1(
        P1_REG1_REG_28__SCAN_IN), .C2(keyinput198), .A(n10070), .ZN(n10075) );
  AOI22_X1 U11154 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(keyinput220), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput188), .ZN(n10071) );
  OAI221_X1 U11155 ( .B1(P2_IR_REG_8__SCAN_IN), .B2(keyinput220), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput188), .A(n10071), .ZN(n10074) );
  AOI22_X1 U11156 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(keyinput143), .B1(
        P2_IR_REG_22__SCAN_IN), .B2(keyinput157), .ZN(n10072) );
  OAI221_X1 U11157 ( .B1(P2_REG0_REG_9__SCAN_IN), .B2(keyinput143), .C1(
        P2_IR_REG_22__SCAN_IN), .C2(keyinput157), .A(n10072), .ZN(n10073) );
  NOR4_X1 U11158 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10098) );
  AOI22_X1 U11159 ( .A1(P2_REG0_REG_17__SCAN_IN), .A2(keyinput187), .B1(
        P2_D_REG_19__SCAN_IN), .B2(keyinput255), .ZN(n10077) );
  OAI221_X1 U11160 ( .B1(P2_REG0_REG_17__SCAN_IN), .B2(keyinput187), .C1(
        P2_D_REG_19__SCAN_IN), .C2(keyinput255), .A(n10077), .ZN(n10084) );
  AOI22_X1 U11161 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput243), .B1(SI_8_), 
        .B2(keyinput165), .ZN(n10078) );
  OAI221_X1 U11162 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput243), .C1(SI_8_), .C2(keyinput165), .A(n10078), .ZN(n10083) );
  AOI22_X1 U11163 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(keyinput252), .B1(
        P1_REG0_REG_30__SCAN_IN), .B2(keyinput147), .ZN(n10079) );
  OAI221_X1 U11164 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(keyinput252), .C1(
        P1_REG0_REG_30__SCAN_IN), .C2(keyinput147), .A(n10079), .ZN(n10082) );
  AOI22_X1 U11165 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput194), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput195), .ZN(n10080) );
  OAI221_X1 U11166 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput194), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput195), .A(n10080), .ZN(n10081)
         );
  NOR4_X1 U11167 ( .A1(n10084), .A2(n10083), .A3(n10082), .A4(n10081), .ZN(
        n10097) );
  AOI22_X1 U11168 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput138), .B1(
        P1_STATE_REG_SCAN_IN), .B2(keyinput139), .ZN(n10085) );
  OAI221_X1 U11169 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput138), .C1(
        P1_STATE_REG_SCAN_IN), .C2(keyinput139), .A(n10085), .ZN(n10095) );
  AOI22_X1 U11170 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput185), .B1(n10087), 
        .B2(keyinput246), .ZN(n10086) );
  OAI221_X1 U11171 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput185), .C1(n10087), 
        .C2(keyinput246), .A(n10086), .ZN(n10094) );
  AOI22_X1 U11172 ( .A1(n10090), .A2(keyinput182), .B1(n10089), .B2(
        keyinput209), .ZN(n10088) );
  OAI221_X1 U11173 ( .B1(n10090), .B2(keyinput182), .C1(n10089), .C2(
        keyinput209), .A(n10088), .ZN(n10093) );
  AOI22_X1 U11174 ( .A1(n10306), .A2(keyinput239), .B1(keyinput135), .B2(
        n10290), .ZN(n10091) );
  OAI221_X1 U11175 ( .B1(n10306), .B2(keyinput239), .C1(n10290), .C2(
        keyinput135), .A(n10091), .ZN(n10092) );
  NOR4_X1 U11176 ( .A1(n10095), .A2(n10094), .A3(n10093), .A4(n10092), .ZN(
        n10096) );
  NAND4_X1 U11177 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n10195) );
  AOI22_X1 U11178 ( .A1(n10102), .A2(keyinput201), .B1(n10101), .B2(
        keyinput241), .ZN(n10100) );
  OAI221_X1 U11179 ( .B1(n10102), .B2(keyinput201), .C1(n10101), .C2(
        keyinput241), .A(n10100), .ZN(n10109) );
  INV_X1 U11180 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U11181 ( .A1(n10242), .A2(keyinput250), .B1(n10218), .B2(
        keyinput211), .ZN(n10103) );
  OAI221_X1 U11182 ( .B1(n10242), .B2(keyinput250), .C1(n10218), .C2(
        keyinput211), .A(n10103), .ZN(n10108) );
  AOI22_X1 U11183 ( .A1(n10202), .A2(keyinput161), .B1(n6645), .B2(keyinput133), .ZN(n10104) );
  OAI221_X1 U11184 ( .B1(n10202), .B2(keyinput161), .C1(n6645), .C2(
        keyinput133), .A(n10104), .ZN(n10107) );
  AOI22_X1 U11185 ( .A1(n10263), .A2(keyinput167), .B1(n10275), .B2(
        keyinput251), .ZN(n10105) );
  OAI221_X1 U11186 ( .B1(n10263), .B2(keyinput167), .C1(n10275), .C2(
        keyinput251), .A(n10105), .ZN(n10106) );
  NOR4_X1 U11187 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n10145) );
  AOI22_X1 U11188 ( .A1(n10303), .A2(keyinput140), .B1(keyinput245), .B2(n6183), .ZN(n10110) );
  OAI221_X1 U11189 ( .B1(n10303), .B2(keyinput140), .C1(n6183), .C2(
        keyinput245), .A(n10110), .ZN(n10119) );
  AOI22_X1 U11190 ( .A1(n5153), .A2(keyinput131), .B1(n10295), .B2(keyinput176), .ZN(n10111) );
  OAI221_X1 U11191 ( .B1(n5153), .B2(keyinput131), .C1(n10295), .C2(
        keyinput176), .A(n10111), .ZN(n10118) );
  INV_X1 U11192 ( .A(SI_21_), .ZN(n10113) );
  INV_X1 U11193 ( .A(SI_7_), .ZN(n10302) );
  AOI22_X1 U11194 ( .A1(n10113), .A2(keyinput154), .B1(keyinput190), .B2(
        n10302), .ZN(n10112) );
  OAI221_X1 U11195 ( .B1(n10113), .B2(keyinput154), .C1(n10302), .C2(
        keyinput190), .A(n10112), .ZN(n10117) );
  XOR2_X1 U11196 ( .A(n5820), .B(keyinput184), .Z(n10115) );
  XNOR2_X1 U11197 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput248), .ZN(n10114) );
  NAND2_X1 U11198 ( .A1(n10115), .A2(n10114), .ZN(n10116) );
  NOR4_X1 U11199 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n10144) );
  AOI22_X1 U11200 ( .A1(n10121), .A2(keyinput146), .B1(keyinput204), .B2(
        n10276), .ZN(n10120) );
  OAI221_X1 U11201 ( .B1(n10121), .B2(keyinput146), .C1(n10276), .C2(
        keyinput204), .A(n10120), .ZN(n10129) );
  AOI22_X1 U11202 ( .A1(n6902), .A2(keyinput227), .B1(n10243), .B2(keyinput226), .ZN(n10122) );
  OAI221_X1 U11203 ( .B1(n6902), .B2(keyinput227), .C1(n10243), .C2(
        keyinput226), .A(n10122), .ZN(n10128) );
  XOR2_X1 U11204 ( .A(n8590), .B(keyinput217), .Z(n10126) );
  XNOR2_X1 U11205 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput132), .ZN(n10125) );
  XNOR2_X1 U11206 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput164), .ZN(n10124) );
  XNOR2_X1 U11207 ( .A(P2_REG1_REG_27__SCAN_IN), .B(keyinput145), .ZN(n10123)
         );
  NAND4_X1 U11208 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n10127) );
  NOR3_X1 U11209 ( .A1(n10129), .A2(n10128), .A3(n10127), .ZN(n10143) );
  AOI22_X1 U11210 ( .A1(n10245), .A2(keyinput144), .B1(n10288), .B2(
        keyinput174), .ZN(n10130) );
  OAI221_X1 U11211 ( .B1(n10245), .B2(keyinput144), .C1(n10288), .C2(
        keyinput174), .A(n10130), .ZN(n10133) );
  XNOR2_X1 U11212 ( .A(n10293), .B(keyinput186), .ZN(n10132) );
  XOR2_X1 U11213 ( .A(SI_0_), .B(keyinput231), .Z(n10131) );
  OR3_X1 U11214 ( .A1(n10133), .A2(n10132), .A3(n10131), .ZN(n10141) );
  AOI22_X1 U11215 ( .A1(n10135), .A2(keyinput166), .B1(keyinput212), .B2(
        n10262), .ZN(n10134) );
  OAI221_X1 U11216 ( .B1(n10135), .B2(keyinput166), .C1(n10262), .C2(
        keyinput212), .A(n10134), .ZN(n10140) );
  AOI22_X1 U11217 ( .A1(n10138), .A2(keyinput225), .B1(keyinput178), .B2(
        n10137), .ZN(n10136) );
  OAI221_X1 U11218 ( .B1(n10138), .B2(keyinput225), .C1(n10137), .C2(
        keyinput178), .A(n10136), .ZN(n10139) );
  NOR3_X1 U11219 ( .A1(n10141), .A2(n10140), .A3(n10139), .ZN(n10142) );
  NAND4_X1 U11220 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10194) );
  AOI22_X1 U11221 ( .A1(n10201), .A2(keyinput159), .B1(keyinput208), .B2(
        n10147), .ZN(n10146) );
  OAI221_X1 U11222 ( .B1(n10201), .B2(keyinput159), .C1(n10147), .C2(
        keyinput208), .A(n10146), .ZN(n10156) );
  AOI22_X1 U11223 ( .A1(n10149), .A2(keyinput162), .B1(n10225), .B2(
        keyinput235), .ZN(n10148) );
  OAI221_X1 U11224 ( .B1(n10149), .B2(keyinput162), .C1(n10225), .C2(
        keyinput235), .A(n10148), .ZN(n10155) );
  INV_X1 U11225 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10272) );
  XNOR2_X1 U11226 ( .A(n10272), .B(keyinput149), .ZN(n10154) );
  XNOR2_X1 U11227 ( .A(P2_REG1_REG_23__SCAN_IN), .B(keyinput181), .ZN(n10152)
         );
  XNOR2_X1 U11228 ( .A(SI_1_), .B(keyinput238), .ZN(n10151) );
  XNOR2_X1 U11229 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput207), .ZN(n10150) );
  NAND3_X1 U11230 ( .A1(n10152), .A2(n10151), .A3(n10150), .ZN(n10153) );
  NOR4_X1 U11231 ( .A1(n10156), .A2(n10155), .A3(n10154), .A4(n10153), .ZN(
        n10192) );
  AOI22_X1 U11232 ( .A1(n5378), .A2(keyinput150), .B1(n10158), .B2(keyinput206), .ZN(n10157) );
  OAI221_X1 U11233 ( .B1(n5378), .B2(keyinput150), .C1(n10158), .C2(
        keyinput206), .A(n10157), .ZN(n10167) );
  INV_X1 U11234 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U11235 ( .A1(n10160), .A2(keyinput183), .B1(n10281), .B2(
        keyinput253), .ZN(n10159) );
  OAI221_X1 U11236 ( .B1(n10160), .B2(keyinput183), .C1(n10281), .C2(
        keyinput253), .A(n10159), .ZN(n10166) );
  AOI22_X1 U11237 ( .A1(n10240), .A2(keyinput215), .B1(keyinput219), .B2(n5611), .ZN(n10161) );
  OAI221_X1 U11238 ( .B1(n10240), .B2(keyinput215), .C1(n5611), .C2(
        keyinput219), .A(n10161), .ZN(n10165) );
  AOI22_X1 U11239 ( .A1(n10163), .A2(keyinput172), .B1(keyinput242), .B2(
        n10233), .ZN(n10162) );
  OAI221_X1 U11240 ( .B1(n10163), .B2(keyinput172), .C1(n10233), .C2(
        keyinput242), .A(n10162), .ZN(n10164) );
  NOR4_X1 U11241 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10191) );
  AOI22_X1 U11242 ( .A1(n10258), .A2(keyinput214), .B1(keyinput171), .B2(
        n10169), .ZN(n10168) );
  OAI221_X1 U11243 ( .B1(n10258), .B2(keyinput214), .C1(n10169), .C2(
        keyinput171), .A(n10168), .ZN(n10177) );
  AOI22_X1 U11244 ( .A1(n10171), .A2(keyinput237), .B1(keyinput192), .B2(
        n10408), .ZN(n10170) );
  OAI221_X1 U11245 ( .B1(n10171), .B2(keyinput237), .C1(n10408), .C2(
        keyinput192), .A(n10170), .ZN(n10176) );
  AOI22_X1 U11246 ( .A1(n10287), .A2(keyinput148), .B1(keyinput228), .B2(n6105), .ZN(n10172) );
  OAI221_X1 U11247 ( .B1(n10287), .B2(keyinput148), .C1(n6105), .C2(
        keyinput228), .A(n10172), .ZN(n10175) );
  INV_X1 U11248 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U11249 ( .A1(n10257), .A2(keyinput205), .B1(n10198), .B2(
        keyinput175), .ZN(n10173) );
  OAI221_X1 U11250 ( .B1(n10257), .B2(keyinput205), .C1(n10198), .C2(
        keyinput175), .A(n10173), .ZN(n10174) );
  NOR4_X1 U11251 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10190) );
  AOI22_X1 U11252 ( .A1(n10179), .A2(keyinput156), .B1(keyinput158), .B2(n6337), .ZN(n10178) );
  OAI221_X1 U11253 ( .B1(n10179), .B2(keyinput156), .C1(n6337), .C2(
        keyinput158), .A(n10178), .ZN(n10188) );
  INV_X1 U11254 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U11255 ( .A1(n10181), .A2(keyinput247), .B1(n10265), .B2(
        keyinput163), .ZN(n10180) );
  OAI221_X1 U11256 ( .B1(n10181), .B2(keyinput247), .C1(n10265), .C2(
        keyinput163), .A(n10180), .ZN(n10187) );
  AOI22_X1 U11257 ( .A1(n5144), .A2(keyinput153), .B1(n10227), .B2(keyinput202), .ZN(n10182) );
  OAI221_X1 U11258 ( .B1(n5144), .B2(keyinput153), .C1(n10227), .C2(
        keyinput202), .A(n10182), .ZN(n10186) );
  INV_X1 U11259 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U11260 ( .A1(n10228), .A2(keyinput222), .B1(keyinput218), .B2(
        n10184), .ZN(n10183) );
  OAI221_X1 U11261 ( .B1(n10228), .B2(keyinput222), .C1(n10184), .C2(
        keyinput218), .A(n10183), .ZN(n10185) );
  NOR4_X1 U11262 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10189) );
  NAND4_X1 U11263 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10193) );
  NOR4_X1 U11264 ( .A1(n10196), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(
        n10395) );
  AOI22_X1 U11265 ( .A1(n10199), .A2(keyinput24), .B1(n10198), .B2(keyinput47), 
        .ZN(n10197) );
  OAI221_X1 U11266 ( .B1(n10199), .B2(keyinput24), .C1(n10198), .C2(keyinput47), .A(n10197), .ZN(n10209) );
  AOI22_X1 U11267 ( .A1(n10202), .A2(keyinput33), .B1(n10201), .B2(keyinput31), 
        .ZN(n10200) );
  OAI221_X1 U11268 ( .B1(n10202), .B2(keyinput33), .C1(n10201), .C2(keyinput31), .A(n10200), .ZN(n10208) );
  AOI22_X1 U11269 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput6), .B1(SI_31_), 
        .B2(keyinput63), .ZN(n10203) );
  OAI221_X1 U11270 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput6), .C1(SI_31_), 
        .C2(keyinput63), .A(n10203), .ZN(n10207) );
  XOR2_X1 U11271 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput92), .Z(n10205) );
  XNOR2_X1 U11272 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput27), .ZN(n10204)
         );
  NAND2_X1 U11273 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  NOR4_X1 U11274 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10255) );
  AOI22_X1 U11275 ( .A1(n5145), .A2(keyinput32), .B1(n8047), .B2(keyinput66), 
        .ZN(n10210) );
  OAI221_X1 U11276 ( .B1(n5145), .B2(keyinput32), .C1(n8047), .C2(keyinput66), 
        .A(n10210), .ZN(n10223) );
  AOI22_X1 U11277 ( .A1(n10213), .A2(keyinput95), .B1(keyinput106), .B2(n10212), .ZN(n10211) );
  OAI221_X1 U11278 ( .B1(n10213), .B2(keyinput95), .C1(n10212), .C2(
        keyinput106), .A(n10211), .ZN(n10222) );
  INV_X1 U11279 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U11280 ( .A1(n10216), .A2(keyinput121), .B1(n10215), .B2(keyinput70), .ZN(n10214) );
  OAI221_X1 U11281 ( .B1(n10216), .B2(keyinput121), .C1(n10215), .C2(
        keyinput70), .A(n10214), .ZN(n10221) );
  AOI22_X1 U11282 ( .A1(n10219), .A2(keyinput14), .B1(n10218), .B2(keyinput83), 
        .ZN(n10217) );
  OAI221_X1 U11283 ( .B1(n10219), .B2(keyinput14), .C1(n10218), .C2(keyinput83), .A(n10217), .ZN(n10220) );
  NOR4_X1 U11284 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10254) );
  AOI22_X1 U11285 ( .A1(n6645), .A2(keyinput5), .B1(n10225), .B2(keyinput107), 
        .ZN(n10224) );
  OAI221_X1 U11286 ( .B1(n6645), .B2(keyinput5), .C1(n10225), .C2(keyinput107), 
        .A(n10224), .ZN(n10238) );
  AOI22_X1 U11287 ( .A1(n10228), .A2(keyinput94), .B1(keyinput74), .B2(n10227), 
        .ZN(n10226) );
  OAI221_X1 U11288 ( .B1(n10228), .B2(keyinput94), .C1(n10227), .C2(keyinput74), .A(n10226), .ZN(n10237) );
  AOI22_X1 U11289 ( .A1(n10231), .A2(keyinput52), .B1(keyinput102), .B2(n10230), .ZN(n10229) );
  OAI221_X1 U11290 ( .B1(n10231), .B2(keyinput52), .C1(n10230), .C2(
        keyinput102), .A(n10229), .ZN(n10236) );
  AOI22_X1 U11291 ( .A1(n10234), .A2(keyinput69), .B1(keyinput114), .B2(n10233), .ZN(n10232) );
  OAI221_X1 U11292 ( .B1(n10234), .B2(keyinput69), .C1(n10233), .C2(
        keyinput114), .A(n10232), .ZN(n10235) );
  NOR4_X1 U11293 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10253) );
  AOI22_X1 U11294 ( .A1(n5820), .A2(keyinput56), .B1(keyinput87), .B2(n10240), 
        .ZN(n10239) );
  OAI221_X1 U11295 ( .B1(n5820), .B2(keyinput56), .C1(n10240), .C2(keyinput87), 
        .A(n10239), .ZN(n10251) );
  AOI22_X1 U11296 ( .A1(n10243), .A2(keyinput98), .B1(keyinput122), .B2(n10242), .ZN(n10241) );
  OAI221_X1 U11297 ( .B1(n10243), .B2(keyinput98), .C1(n10242), .C2(
        keyinput122), .A(n10241), .ZN(n10250) );
  AOI22_X1 U11298 ( .A1(n5378), .A2(keyinput22), .B1(keyinput16), .B2(n10245), 
        .ZN(n10244) );
  OAI221_X1 U11299 ( .B1(n5378), .B2(keyinput22), .C1(n10245), .C2(keyinput16), 
        .A(n10244), .ZN(n10249) );
  XOR2_X1 U11300 ( .A(n5611), .B(keyinput91), .Z(n10247) );
  XNOR2_X1 U11301 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput120), .ZN(n10246) );
  NAND2_X1 U11302 ( .A1(n10247), .A2(n10246), .ZN(n10248) );
  NOR4_X1 U11303 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10252) );
  NAND4_X1 U11304 ( .A1(n10255), .A2(n10254), .A3(n10253), .A4(n10252), .ZN(
        n10394) );
  AOI22_X1 U11305 ( .A1(n10258), .A2(keyinput86), .B1(keyinput77), .B2(n10257), 
        .ZN(n10256) );
  OAI221_X1 U11306 ( .B1(n10258), .B2(keyinput86), .C1(n10257), .C2(keyinput77), .A(n10256), .ZN(n10270) );
  AOI22_X1 U11307 ( .A1(n6902), .A2(keyinput99), .B1(keyinput53), .B2(n10260), 
        .ZN(n10259) );
  OAI221_X1 U11308 ( .B1(n6902), .B2(keyinput99), .C1(n10260), .C2(keyinput53), 
        .A(n10259), .ZN(n10269) );
  AOI22_X1 U11309 ( .A1(n10263), .A2(keyinput39), .B1(n10262), .B2(keyinput84), 
        .ZN(n10261) );
  OAI221_X1 U11310 ( .B1(n10263), .B2(keyinput39), .C1(n10262), .C2(keyinput84), .A(n10261), .ZN(n10268) );
  INV_X1 U11311 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U11312 ( .A1(n10266), .A2(keyinput105), .B1(n10265), .B2(keyinput35), .ZN(n10264) );
  OAI221_X1 U11313 ( .B1(n10266), .B2(keyinput105), .C1(n10265), .C2(
        keyinput35), .A(n10264), .ZN(n10267) );
  NOR4_X1 U11314 ( .A1(n10270), .A2(n10269), .A3(n10268), .A4(n10267), .ZN(
        n10392) );
  AOI22_X1 U11315 ( .A1(n10273), .A2(keyinput115), .B1(n10272), .B2(keyinput21), .ZN(n10271) );
  OAI221_X1 U11316 ( .B1(n10273), .B2(keyinput115), .C1(n10272), .C2(
        keyinput21), .A(n10271), .ZN(n10316) );
  OAI22_X1 U11317 ( .A1(n10276), .A2(keyinput76), .B1(n10275), .B2(keyinput123), .ZN(n10274) );
  AOI221_X1 U11318 ( .B1(n10276), .B2(keyinput76), .C1(keyinput123), .C2(
        n10275), .A(n10274), .ZN(n10285) );
  OAI22_X1 U11319 ( .A1(n10279), .A2(keyinput10), .B1(n10278), .B2(keyinput2), 
        .ZN(n10277) );
  AOI221_X1 U11320 ( .B1(n10279), .B2(keyinput10), .C1(keyinput2), .C2(n10278), 
        .A(n10277), .ZN(n10284) );
  OAI22_X1 U11321 ( .A1(n10282), .A2(keyinput13), .B1(n10281), .B2(keyinput125), .ZN(n10280) );
  AOI221_X1 U11322 ( .B1(n10282), .B2(keyinput13), .C1(keyinput125), .C2(
        n10281), .A(n10280), .ZN(n10283) );
  NAND3_X1 U11323 ( .A1(n10285), .A2(n10284), .A3(n10283), .ZN(n10315) );
  OAI22_X1 U11324 ( .A1(n10288), .A2(keyinput46), .B1(n10287), .B2(keyinput20), 
        .ZN(n10286) );
  AOI221_X1 U11325 ( .B1(n10288), .B2(keyinput46), .C1(keyinput20), .C2(n10287), .A(n10286), .ZN(n10299) );
  OAI22_X1 U11326 ( .A1(n10291), .A2(keyinput57), .B1(n10290), .B2(keyinput7), 
        .ZN(n10289) );
  AOI221_X1 U11327 ( .B1(n10291), .B2(keyinput57), .C1(keyinput7), .C2(n10290), 
        .A(n10289), .ZN(n10298) );
  OAI22_X1 U11328 ( .A1(n6998), .A2(keyinput41), .B1(n10293), .B2(keyinput58), 
        .ZN(n10292) );
  AOI221_X1 U11329 ( .B1(n6998), .B2(keyinput41), .C1(keyinput58), .C2(n10293), 
        .A(n10292), .ZN(n10297) );
  OAI22_X1 U11330 ( .A1(n10295), .A2(keyinput48), .B1(n5153), .B2(keyinput3), 
        .ZN(n10294) );
  AOI221_X1 U11331 ( .B1(n10295), .B2(keyinput48), .C1(keyinput3), .C2(n5153), 
        .A(n10294), .ZN(n10296) );
  NAND4_X1 U11332 ( .A1(n10299), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10314) );
  OAI22_X1 U11333 ( .A1(n7057), .A2(keyinput75), .B1(n6137), .B2(keyinput72), 
        .ZN(n10300) );
  AOI221_X1 U11334 ( .B1(n7057), .B2(keyinput75), .C1(keyinput72), .C2(n6137), 
        .A(n10300), .ZN(n10312) );
  OAI22_X1 U11335 ( .A1(n10303), .A2(keyinput12), .B1(n10302), .B2(keyinput62), 
        .ZN(n10301) );
  AOI221_X1 U11336 ( .B1(n10303), .B2(keyinput12), .C1(keyinput62), .C2(n10302), .A(n10301), .ZN(n10311) );
  OAI22_X1 U11337 ( .A1(n10306), .A2(keyinput111), .B1(n10305), .B2(keyinput88), .ZN(n10304) );
  AOI221_X1 U11338 ( .B1(n10306), .B2(keyinput111), .C1(keyinput88), .C2(
        n10305), .A(n10304), .ZN(n10310) );
  XOR2_X1 U11339 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput79), .Z(n10308) );
  XNOR2_X1 U11340 ( .A(keyinput15), .B(n5311), .ZN(n10307) );
  NOR2_X1 U11341 ( .A1(n10308), .A2(n10307), .ZN(n10309) );
  NAND4_X1 U11342 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n10309), .ZN(
        n10313) );
  NOR4_X1 U11343 ( .A1(n10316), .A2(n10315), .A3(n10314), .A4(n10313), .ZN(
        n10391) );
  OAI22_X1 U11344 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(keyinput101), .B1(
        keyinput30), .B2(P1_REG0_REG_3__SCAN_IN), .ZN(n10317) );
  AOI221_X1 U11345 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(keyinput101), .C1(
        P1_REG0_REG_3__SCAN_IN), .C2(keyinput30), .A(n10317), .ZN(n10324) );
  OAI22_X1 U11346 ( .A1(P2_REG0_REG_12__SCAN_IN), .A2(keyinput85), .B1(
        keyinput19), .B2(P1_REG0_REG_30__SCAN_IN), .ZN(n10318) );
  AOI221_X1 U11347 ( .B1(P2_REG0_REG_12__SCAN_IN), .B2(keyinput85), .C1(
        P1_REG0_REG_30__SCAN_IN), .C2(keyinput19), .A(n10318), .ZN(n10323) );
  OAI22_X1 U11348 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput60), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(keyinput1), .ZN(n10319) );
  AOI221_X1 U11349 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput60), .C1(keyinput1), 
        .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10319), .ZN(n10322) );
  OAI22_X1 U11350 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput104), .B1(
        keyinput119), .B2(P2_ADDR_REG_17__SCAN_IN), .ZN(n10320) );
  AOI221_X1 U11351 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput104), .C1(
        P2_ADDR_REG_17__SCAN_IN), .C2(keyinput119), .A(n10320), .ZN(n10321) );
  NAND4_X1 U11352 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10352) );
  OAI22_X1 U11353 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput36), .B1(keyinput54), .B2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10325) );
  AOI221_X1 U11354 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput36), .C1(
        P1_ADDR_REG_2__SCAN_IN), .C2(keyinput54), .A(n10325), .ZN(n10332) );
  OAI22_X1 U11355 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(keyinput108), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(keyinput80), .ZN(n10326) );
  AOI221_X1 U11356 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(keyinput108), .C1(
        keyinput80), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10326), .ZN(n10331) );
  OAI22_X1 U11357 ( .A1(P2_REG0_REG_17__SCAN_IN), .A2(keyinput59), .B1(
        P2_REG1_REG_13__SCAN_IN), .B2(keyinput42), .ZN(n10327) );
  AOI221_X1 U11358 ( .B1(P2_REG0_REG_17__SCAN_IN), .B2(keyinput59), .C1(
        keyinput42), .C2(P2_REG1_REG_13__SCAN_IN), .A(n10327), .ZN(n10330) );
  OAI22_X1 U11359 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(keyinput113), .B1(
        P1_REG1_REG_31__SCAN_IN), .B2(keyinput55), .ZN(n10328) );
  AOI221_X1 U11360 ( .B1(P1_DATAO_REG_22__SCAN_IN), .B2(keyinput113), .C1(
        keyinput55), .C2(P1_REG1_REG_31__SCAN_IN), .A(n10328), .ZN(n10329) );
  NAND4_X1 U11361 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10351) );
  OAI22_X1 U11362 ( .A1(SI_23_), .A2(keyinput8), .B1(SI_0_), .B2(keyinput103), 
        .ZN(n10333) );
  AOI221_X1 U11363 ( .B1(SI_23_), .B2(keyinput8), .C1(keyinput103), .C2(SI_0_), 
        .A(n10333), .ZN(n10340) );
  OAI22_X1 U11364 ( .A1(P1_D_REG_10__SCAN_IN), .A2(keyinput44), .B1(SI_21_), 
        .B2(keyinput26), .ZN(n10334) );
  AOI221_X1 U11365 ( .B1(P1_D_REG_10__SCAN_IN), .B2(keyinput44), .C1(
        keyinput26), .C2(SI_21_), .A(n10334), .ZN(n10339) );
  OAI22_X1 U11366 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(keyinput38), .B1(
        P2_REG0_REG_2__SCAN_IN), .B2(keyinput25), .ZN(n10335) );
  AOI221_X1 U11367 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(keyinput38), .C1(
        keyinput25), .C2(P2_REG0_REG_2__SCAN_IN), .A(n10335), .ZN(n10338) );
  OAI22_X1 U11368 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(keyinput28), .B1(
        keyinput117), .B2(P1_REG2_REG_0__SCAN_IN), .ZN(n10336) );
  AOI221_X1 U11369 ( .B1(P1_DATAO_REG_4__SCAN_IN), .B2(keyinput28), .C1(
        P1_REG2_REG_0__SCAN_IN), .C2(keyinput117), .A(n10336), .ZN(n10337) );
  NAND4_X1 U11370 ( .A1(n10340), .A2(n10339), .A3(n10338), .A4(n10337), .ZN(
        n10350) );
  OAI22_X1 U11371 ( .A1(P1_D_REG_22__SCAN_IN), .A2(keyinput9), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput73), .ZN(n10341) );
  AOI221_X1 U11372 ( .B1(P1_D_REG_22__SCAN_IN), .B2(keyinput9), .C1(keyinput73), .C2(P2_REG3_REG_10__SCAN_IN), .A(n10341), .ZN(n10348) );
  OAI22_X1 U11373 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(keyinput17), .B1(
        P2_REG2_REG_2__SCAN_IN), .B2(keyinput100), .ZN(n10342) );
  AOI221_X1 U11374 ( .B1(P2_REG1_REG_27__SCAN_IN), .B2(keyinput17), .C1(
        keyinput100), .C2(P2_REG2_REG_2__SCAN_IN), .A(n10342), .ZN(n10347) );
  OAI22_X1 U11375 ( .A1(P1_D_REG_29__SCAN_IN), .A2(keyinput118), .B1(
        keyinput82), .B2(P1_REG3_REG_23__SCAN_IN), .ZN(n10343) );
  AOI221_X1 U11376 ( .B1(P1_D_REG_29__SCAN_IN), .B2(keyinput118), .C1(
        P1_REG3_REG_23__SCAN_IN), .C2(keyinput82), .A(n10343), .ZN(n10346) );
  OAI22_X1 U11377 ( .A1(P1_REG0_REG_28__SCAN_IN), .A2(keyinput50), .B1(
        P1_REG0_REG_15__SCAN_IN), .B2(keyinput34), .ZN(n10344) );
  AOI221_X1 U11378 ( .B1(P1_REG0_REG_28__SCAN_IN), .B2(keyinput50), .C1(
        keyinput34), .C2(P1_REG0_REG_15__SCAN_IN), .A(n10344), .ZN(n10345) );
  NAND4_X1 U11379 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10349) );
  NOR4_X1 U11380 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        n10390) );
  OAI22_X1 U11381 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(keyinput29), .B1(
        P2_IR_REG_17__SCAN_IN), .B2(keyinput61), .ZN(n10353) );
  AOI221_X1 U11382 ( .B1(P2_IR_REG_22__SCAN_IN), .B2(keyinput29), .C1(
        keyinput61), .C2(P2_IR_REG_17__SCAN_IN), .A(n10353), .ZN(n10360) );
  OAI22_X1 U11383 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(keyinput112), .B1(
        keyinput124), .B2(P2_ADDR_REG_0__SCAN_IN), .ZN(n10354) );
  AOI221_X1 U11384 ( .B1(P1_REG1_REG_26__SCAN_IN), .B2(keyinput112), .C1(
        P2_ADDR_REG_0__SCAN_IN), .C2(keyinput124), .A(n10354), .ZN(n10359) );
  OAI22_X1 U11385 ( .A1(P1_D_REG_7__SCAN_IN), .A2(keyinput40), .B1(SI_15_), 
        .B2(keyinput0), .ZN(n10355) );
  AOI221_X1 U11386 ( .B1(P1_D_REG_7__SCAN_IN), .B2(keyinput40), .C1(keyinput0), 
        .C2(SI_15_), .A(n10355), .ZN(n10358) );
  OAI22_X1 U11387 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput116), .B1(
        keyinput126), .B2(P1_ADDR_REG_14__SCAN_IN), .ZN(n10356) );
  AOI221_X1 U11388 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput116), .C1(
        P1_ADDR_REG_14__SCAN_IN), .C2(keyinput126), .A(n10356), .ZN(n10357) );
  NAND4_X1 U11389 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10388) );
  OAI22_X1 U11390 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(keyinput97), .B1(
        keyinput18), .B2(P1_REG0_REG_14__SCAN_IN), .ZN(n10361) );
  AOI221_X1 U11391 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(keyinput97), .C1(
        P1_REG0_REG_14__SCAN_IN), .C2(keyinput18), .A(n10361), .ZN(n10368) );
  OAI22_X1 U11392 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput96), .B1(
        P2_ADDR_REG_2__SCAN_IN), .B2(keyinput45), .ZN(n10362) );
  AOI221_X1 U11393 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput96), .C1(
        keyinput45), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10362), .ZN(n10367) );
  OAI22_X1 U11394 ( .A1(SI_19_), .A2(keyinput78), .B1(keyinput109), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n10363) );
  AOI221_X1 U11395 ( .B1(SI_19_), .B2(keyinput78), .C1(P2_ADDR_REG_3__SCAN_IN), 
        .C2(keyinput109), .A(n10363), .ZN(n10366) );
  OAI22_X1 U11396 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput23), .B1(SI_1_), 
        .B2(keyinput110), .ZN(n10364) );
  AOI221_X1 U11397 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput23), .C1(
        keyinput110), .C2(SI_1_), .A(n10364), .ZN(n10365) );
  NAND4_X1 U11398 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10387) );
  OAI22_X1 U11399 ( .A1(SI_9_), .A2(keyinput93), .B1(P1_REG1_REG_29__SCAN_IN), 
        .B2(keyinput68), .ZN(n10369) );
  AOI221_X1 U11400 ( .B1(SI_9_), .B2(keyinput93), .C1(keyinput68), .C2(
        P1_REG1_REG_29__SCAN_IN), .A(n10369), .ZN(n10376) );
  OAI22_X1 U11401 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput67), .B1(
        keyinput90), .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n10370) );
  AOI221_X1 U11402 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput67), .C1(
        P1_DATAO_REG_29__SCAN_IN), .C2(keyinput90), .A(n10370), .ZN(n10375) );
  OAI22_X1 U11403 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(keyinput49), .B1(
        keyinput64), .B2(P1_ADDR_REG_9__SCAN_IN), .ZN(n10371) );
  AOI221_X1 U11404 ( .B1(P2_REG0_REG_14__SCAN_IN), .B2(keyinput49), .C1(
        P1_ADDR_REG_9__SCAN_IN), .C2(keyinput64), .A(n10371), .ZN(n10374) );
  OAI22_X1 U11405 ( .A1(P2_D_REG_19__SCAN_IN), .A2(keyinput127), .B1(
        keyinput43), .B2(P2_REG0_REG_25__SCAN_IN), .ZN(n10372) );
  AOI221_X1 U11406 ( .B1(P2_D_REG_19__SCAN_IN), .B2(keyinput127), .C1(
        P2_REG0_REG_25__SCAN_IN), .C2(keyinput43), .A(n10372), .ZN(n10373) );
  NAND4_X1 U11407 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10386) );
  OAI22_X1 U11408 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput4), .B1(keyinput51), .B2(P2_IR_REG_13__SCAN_IN), .ZN(n10377) );
  AOI221_X1 U11409 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput4), .C1(
        P2_IR_REG_13__SCAN_IN), .C2(keyinput51), .A(n10377), .ZN(n10384) );
  OAI22_X1 U11410 ( .A1(SI_12_), .A2(keyinput71), .B1(keyinput37), .B2(SI_8_), 
        .ZN(n10378) );
  AOI221_X1 U11411 ( .B1(SI_12_), .B2(keyinput71), .C1(SI_8_), .C2(keyinput37), 
        .A(n10378), .ZN(n10383) );
  OAI22_X1 U11412 ( .A1(P1_STATE_REG_SCAN_IN), .A2(keyinput11), .B1(
        P1_REG3_REG_21__SCAN_IN), .B2(keyinput89), .ZN(n10379) );
  AOI221_X1 U11413 ( .B1(P1_STATE_REG_SCAN_IN), .B2(keyinput11), .C1(
        keyinput89), .C2(P1_REG3_REG_21__SCAN_IN), .A(n10379), .ZN(n10382) );
  OAI22_X1 U11414 ( .A1(P1_REG0_REG_21__SCAN_IN), .A2(keyinput65), .B1(
        P2_D_REG_21__SCAN_IN), .B2(keyinput81), .ZN(n10380) );
  AOI221_X1 U11415 ( .B1(P1_REG0_REG_21__SCAN_IN), .B2(keyinput65), .C1(
        keyinput81), .C2(P2_D_REG_21__SCAN_IN), .A(n10380), .ZN(n10381) );
  NAND4_X1 U11416 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10385) );
  NOR4_X1 U11417 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10389) );
  NAND4_X1 U11418 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10393) );
  NOR3_X1 U11419 ( .A1(n10395), .A2(n10394), .A3(n10393), .ZN(n10396) );
  XNOR2_X1 U11420 ( .A(n10397), .B(n10396), .ZN(P1_U3315) );
  XOR2_X1 U11421 ( .A(n10398), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11422 ( .A1(n10400), .A2(n10399), .ZN(n10401) );
  XOR2_X1 U11423 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10401), .Z(ADD_1071_U51) );
  OAI21_X1 U11424 ( .B1(n10404), .B2(n10403), .A(n10402), .ZN(n10405) );
  XNOR2_X1 U11425 ( .A(n10405), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11426 ( .B1(n10408), .B2(n10407), .A(n10406), .ZN(ADD_1071_U47) );
  XOR2_X1 U11427 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10409), .Z(ADD_1071_U48) );
  XOR2_X1 U11428 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10410), .Z(ADD_1071_U49) );
  XOR2_X1 U11429 ( .A(n10412), .B(n10411), .Z(ADD_1071_U54) );
  XOR2_X1 U11430 ( .A(n10414), .B(n10413), .Z(ADD_1071_U53) );
  XNOR2_X1 U11431 ( .A(n10416), .B(n10415), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4991 ( .A(n7473), .Z(n8730) );
  INV_X2 U6518 ( .A(n9767), .ZN(n9786) );
endmodule

