

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5054, n5055, n5056, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070;

  NOR3_X1 U5119 ( .A1(n9340), .A2(n9528), .A3(n9534), .ZN(n8085) );
  NOR2_X2 U5120 ( .A1(n10464), .A2(n10329), .ZN(n10307) );
  NAND2_X1 U5121 ( .A1(n8109), .A2(n8108), .ZN(n10500) );
  CLKBUF_X3 U5122 ( .A(n6600), .Z(n9080) );
  CLKBUF_X2 U5123 ( .A(n5901), .Z(n8013) );
  INV_X1 U5124 ( .A(n10178), .ZN(n10728) );
  INV_X1 U5125 ( .A(n5839), .ZN(n6133) );
  INV_X1 U5126 ( .A(n8850), .ZN(n8840) );
  AND2_X1 U5127 ( .A1(n7349), .A2(n6584), .ZN(n9083) );
  INV_X1 U5128 ( .A(n8927), .ZN(n8940) );
  INV_X1 U5129 ( .A(n5858), .ZN(n8685) );
  XNOR2_X1 U5130 ( .A(n9523), .B(n9308), .ZN(n9290) );
  OR2_X1 U5131 ( .A1(n9554), .A2(n9402), .ZN(n9381) );
  INV_X1 U5132 ( .A(n6013), .ZN(n6470) );
  INV_X2 U5133 ( .A(n9083), .ZN(n9076) );
  INV_X1 U5134 ( .A(n6813), .ZN(n10762) );
  AND3_X1 U5135 ( .A1(n5853), .A2(n5852), .A3(n5851), .ZN(n6659) );
  INV_X1 U5137 ( .A(n9290), .ZN(n8880) );
  OAI211_X1 U5138 ( .C1(n7005), .C2(n6912), .A(n6911), .B(n6910), .ZN(n10784)
         );
  CLKBUF_X2 U5139 ( .A(n6469), .Z(n8492) );
  NAND2_X1 U5140 ( .A1(n8568), .A2(n8567), .ZN(n10381) );
  NAND4_X1 U5141 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n9224)
         );
  BUF_X1 U5142 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n10662) );
  INV_X1 U5143 ( .A(n8675), .ZN(n10708) );
  OR3_X2 U5144 ( .A1(n9340), .A2(n5476), .A3(n5475), .ZN(n5054) );
  INV_X1 U5145 ( .A(n9225), .ZN(n6656) );
  INV_X1 U5146 ( .A(n5811), .ZN(n5804) );
  NAND4_X4 U5147 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .ZN(n9175)
         );
  AOI22_X2 U5148 ( .A1(n10104), .A2(n10105), .B1(n9069), .B2(n9068), .ZN(
        n10200) );
  OAI22_X2 U5149 ( .A1(n10132), .A2(n10133), .B1(n9063), .B2(n9062), .ZN(
        n10104) );
  OAI222_X1 U5150 ( .A1(n9112), .A2(P2_U3152), .B1(n10053), .B2(n10531), .C1(
        n9111), .C2(n9110), .ZN(P2_U3328) );
  OR2_X4 U5151 ( .A1(n9112), .A2(n5772), .ZN(n5839) );
  CLKBUF_X1 U5152 ( .A(n5988), .Z(n5055) );
  XNOR2_X1 U5153 ( .A(n5192), .B(n5809), .ZN(n5988) );
  NAND2_X2 U5154 ( .A1(n8158), .A2(n8157), .ZN(n10479) );
  NAND2_X2 U5155 ( .A1(n10050), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U5156 ( .A1(n10200), .A2(n10199), .ZN(n10198) );
  NAND2_X1 U5157 ( .A1(n9366), .A2(n8057), .ZN(n9365) );
  OR2_X1 U5158 ( .A1(n9528), .A2(n9521), .ZN(n5475) );
  NAND2_X1 U5159 ( .A1(n8997), .A2(n8996), .ZN(n10152) );
  AND2_X1 U5160 ( .A1(n8025), .A2(n9352), .ZN(n9353) );
  OAI21_X1 U5161 ( .B1(n7532), .B2(n7531), .A(n7530), .ZN(n7698) );
  NAND2_X1 U5162 ( .A1(n7281), .A2(n7280), .ZN(n7285) );
  NAND2_X1 U5163 ( .A1(n7130), .A2(n7131), .ZN(n7281) );
  NAND2_X1 U5164 ( .A1(n8121), .A2(n8120), .ZN(n10494) );
  NAND2_X1 U5165 ( .A1(n6919), .A2(n6918), .ZN(n7018) );
  NAND2_X1 U5166 ( .A1(n7642), .A2(n7641), .ZN(n10020) );
  NAND2_X1 U5167 ( .A1(n7372), .A2(n7568), .ZN(n10889) );
  MUX2_X1 U5168 ( .A(n8511), .B(n8510), .S(n8613), .Z(n8512) );
  NAND2_X1 U5169 ( .A1(n6966), .A2(n5520), .ZN(n5522) );
  NAND2_X1 U5170 ( .A1(n7603), .A2(n7602), .ZN(n10976) );
  NAND2_X1 U5171 ( .A1(n7705), .A2(n7704), .ZN(n10968) );
  NAND2_X2 U5172 ( .A1(n6889), .A2(n10935), .ZN(n10946) );
  AND3_X1 U5173 ( .A1(n5818), .A2(n5817), .A3(n5816), .ZN(n7111) );
  NAND2_X1 U5174 ( .A1(n5469), .A2(n6881), .ZN(n7094) );
  NAND2_X1 U5175 ( .A1(n6481), .A2(n10786), .ZN(n10223) );
  NAND2_X1 U5176 ( .A1(n5321), .A2(n5318), .ZN(n9170) );
  NAND2_X1 U5177 ( .A1(n6815), .A2(n6814), .ZN(n11035) );
  INV_X1 U5178 ( .A(n10235), .ZN(n10778) );
  INV_X2 U5179 ( .A(n5877), .ZN(n8941) );
  NAND4_X1 U5181 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n10235)
         );
  AND3_X1 U5182 ( .A1(n5876), .A2(n5875), .A3(n5874), .ZN(n10754) );
  NAND3_X1 U5183 ( .A1(n5838), .A2(n5621), .A3(n5620), .ZN(n9225) );
  AND2_X4 U5184 ( .A1(n6563), .A2(n6584), .ZN(n7122) );
  NAND4_X1 U5185 ( .A1(n6576), .A2(n6575), .A3(n6574), .A4(n6573), .ZN(n10731)
         );
  INV_X1 U5186 ( .A(n6465), .ZN(n8619) );
  INV_X1 U5187 ( .A(n6659), .ZN(n6655) );
  NAND4_X1 U5188 ( .A1(n6018), .A2(n6017), .A3(n6015), .A4(n6016), .ZN(n6803)
         );
  INV_X1 U5189 ( .A(n6804), .ZN(n5056) );
  NAND3_X1 U5190 ( .A1(n5861), .A2(n5860), .A3(n5859), .ZN(n6529) );
  INV_X4 U5191 ( .A(n6134), .ZN(n8093) );
  AND2_X1 U5192 ( .A1(n5755), .A2(n5754), .ZN(n8618) );
  INV_X2 U5195 ( .A(n5928), .ZN(n8693) );
  NAND2_X1 U5196 ( .A1(n6577), .A2(n7833), .ZN(n7005) );
  CLKBUF_X1 U5197 ( .A(n6478), .Z(n10789) );
  INV_X2 U5198 ( .A(n5833), .ZN(n5856) );
  AND2_X1 U5199 ( .A1(n6124), .A2(n6128), .ZN(n5722) );
  AOI21_X1 U5200 ( .B1(n5805), .B2(n5434), .A(n5108), .ZN(n5433) );
  XNOR2_X1 U5201 ( .A(n6019), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8675) );
  AND2_X1 U5202 ( .A1(n6019), .A2(n5750), .ZN(n5753) );
  INV_X1 U5203 ( .A(n6011), .ZN(n10530) );
  NAND2_X2 U5204 ( .A1(n5988), .A2(n5971), .ZN(n5833) );
  XNOR2_X1 U5205 ( .A(n6009), .B(n9973), .ZN(n6013) );
  XNOR2_X1 U5206 ( .A(n5691), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6011) );
  CLKBUF_X1 U5207 ( .A(n5971), .Z(n9104) );
  NAND2_X1 U5208 ( .A1(n5749), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U5209 ( .A1(n10523), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5691) );
  NOR2_X1 U5210 ( .A1(n6490), .A2(n5747), .ZN(n6844) );
  CLKBUF_X1 U5211 ( .A(n5804), .Z(n5153) );
  AND2_X1 U5212 ( .A1(n5734), .A2(n5536), .ZN(n5765) );
  OR2_X1 U5213 ( .A1(n5372), .A2(n5072), .ZN(n10523) );
  NAND2_X2 U5214 ( .A1(n7833), .A2(P1_U3084), .ZN(n10532) );
  NAND2_X2 U5215 ( .A1(n8483), .A2(P1_U3084), .ZN(n10528) );
  NAND2_X1 U5216 ( .A1(n5617), .A2(n5618), .ZN(n5811) );
  AND2_X1 U5217 ( .A1(n5177), .A2(n5662), .ZN(n5659) );
  NAND2_X1 U5218 ( .A1(n5663), .A2(n5569), .ZN(n5570) );
  INV_X2 U5219 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9956) );
  INV_X1 U5220 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9734) );
  NOR2_X1 U5221 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5706) );
  NOR2_X1 U5222 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5707) );
  INV_X1 U5223 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9954) );
  NOR2_X1 U5224 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5703) );
  INV_X1 U5225 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9729) );
  NOR2_X1 U5226 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6036) );
  INV_X4 U5227 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5228 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5178) );
  NOR2_X1 U5229 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6792) );
  NOR2_X1 U5230 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5729) );
  INV_X4 U5231 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U5232 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5728) );
  NOR2_X1 U5233 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5727) );
  INV_X1 U5234 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6484) );
  INV_X1 U5235 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6284) );
  AOI21_X2 U5236 ( .B1(n5676), .B2(n5119), .A(n5339), .ZN(n10132) );
  XNOR2_X2 U5237 ( .A(n5855), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10661) );
  NAND2_X1 U5238 ( .A1(n8600), .A2(n5100), .ZN(n8602) );
  NOR2_X1 U5239 ( .A1(n5607), .A2(n5432), .ZN(n5431) );
  INV_X1 U5240 ( .A(n5433), .ZN(n5432) );
  NAND2_X1 U5241 ( .A1(n6107), .A2(n9808), .ZN(n6139) );
  OR2_X1 U5242 ( .A1(n9554), .A2(n9216), .ZN(n8811) );
  OR2_X1 U5243 ( .A1(n10005), .A2(n9186), .ZN(n8789) );
  NAND2_X1 U5244 ( .A1(n10020), .A2(n9502), .ZN(n5333) );
  BUF_X1 U5245 ( .A(n6011), .Z(n6471) );
  INV_X1 U5246 ( .A(n7821), .ZN(n5551) );
  INV_X1 U5247 ( .A(n5550), .ZN(n5549) );
  OAI21_X1 U5248 ( .B1(n8652), .B2(n5551), .A(n8653), .ZN(n5550) );
  NAND2_X1 U5249 ( .A1(n8471), .A2(n8470), .ZN(n8478) );
  AOI21_X1 U5250 ( .B1(n5586), .B2(n5059), .A(n5091), .ZN(n5585) );
  INV_X1 U5251 ( .A(n5415), .ZN(n5414) );
  OAI21_X1 U5252 ( .B1(n5416), .B2(n5586), .A(n8974), .ZN(n5415) );
  INV_X1 U5253 ( .A(n8708), .ZN(n8887) );
  NOR2_X1 U5254 ( .A1(n8363), .A2(n7094), .ZN(n7095) );
  AND2_X1 U5255 ( .A1(n5661), .A2(n5112), .ZN(n5177) );
  NOR2_X1 U5256 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  AND2_X2 U5257 ( .A1(n6471), .A2(n6470), .ZN(n8254) );
  AND2_X1 U5259 ( .A1(n6471), .A2(n6013), .ZN(n6571) );
  NOR2_X1 U5260 ( .A1(n5250), .A2(n9303), .ZN(n5249) );
  NOR2_X1 U5261 ( .A1(n8880), .A2(n5076), .ZN(n5250) );
  NOR2_X1 U5262 ( .A1(n7793), .A2(n5461), .ZN(n5460) );
  INV_X1 U5263 ( .A(n7728), .ZN(n5461) );
  INV_X1 U5264 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6786) );
  INV_X1 U5265 ( .A(n6276), .ZN(n5612) );
  NAND2_X1 U5266 ( .A1(n6371), .A2(n9589), .ZN(n6489) );
  INV_X1 U5267 ( .A(n6110), .ZN(n5608) );
  INV_X1 U5268 ( .A(n7928), .ZN(n5410) );
  AND2_X1 U5269 ( .A1(n5957), .A2(n5937), .ZN(n5595) );
  AOI21_X1 U5270 ( .B1(n5247), .B2(n5242), .A(n9514), .ZN(n5241) );
  INV_X1 U5271 ( .A(n5249), .ZN(n5242) );
  OR2_X1 U5272 ( .A1(n9528), .A2(n9202), .ZN(n8836) );
  OR2_X1 U5273 ( .A1(n9549), .A2(n9160), .ZN(n8817) );
  INV_X1 U5274 ( .A(n8801), .ZN(n5316) );
  AOI21_X1 U5275 ( .B1(n5314), .B2(n5639), .A(n5632), .ZN(n5313) );
  NAND2_X1 U5276 ( .A1(n5635), .A2(n5636), .ZN(n5632) );
  OR2_X1 U5277 ( .A1(n9993), .A2(n8346), .ZN(n8804) );
  AND2_X1 U5278 ( .A1(n9998), .A2(n9394), .ZN(n8801) );
  NAND2_X1 U5279 ( .A1(n5642), .A2(n9416), .ZN(n5639) );
  OR2_X1 U5280 ( .A1(n10015), .A2(n9447), .ZN(n8781) );
  OR2_X1 U5281 ( .A1(n10023), .A2(n8969), .ZN(n8706) );
  INV_X1 U5282 ( .A(n7420), .ZN(n7418) );
  AND2_X1 U5283 ( .A1(n5809), .A2(n5807), .ZN(n5762) );
  NAND2_X1 U5284 ( .A1(n8498), .A2(n5439), .ZN(n5438) );
  AND2_X1 U5285 ( .A1(n10444), .A2(n9094), .ZN(n8466) );
  NOR2_X1 U5286 ( .A1(n8665), .A2(n5482), .ZN(n5481) );
  OR2_X1 U5287 ( .A1(n10449), .A2(n10295), .ZN(n8629) );
  NAND2_X1 U5288 ( .A1(n10454), .A2(n10107), .ZN(n10285) );
  INV_X1 U5289 ( .A(n8656), .ZN(n7851) );
  NAND2_X1 U5290 ( .A1(n8619), .A2(n6461), .ZN(n7350) );
  NAND2_X1 U5291 ( .A1(n7973), .A2(n7972), .ZN(n8468) );
  NAND2_X1 U5292 ( .A1(n8081), .A2(n8080), .ZN(n7973) );
  AND2_X1 U5293 ( .A1(n7964), .A2(n7836), .ZN(n7958) );
  OAI21_X1 U5294 ( .B1(n5460), .B2(n5137), .A(n7840), .ZN(n5457) );
  OAI21_X1 U5295 ( .B1(n7578), .B2(n7577), .A(n7576), .ZN(n7727) );
  AND2_X1 U5296 ( .A1(n7728), .A2(n7582), .ZN(n7726) );
  NAND2_X1 U5297 ( .A1(n9729), .A2(n5746), .ZN(n5747) );
  OAI21_X1 U5298 ( .B1(n5603), .B2(n7184), .A(n5601), .ZN(n7264) );
  AOI21_X1 U5299 ( .B1(n7185), .B2(n5602), .A(n5131), .ZN(n5601) );
  INV_X1 U5300 ( .A(n6978), .ZN(n5602) );
  XNOR2_X1 U5301 ( .A(n6275), .B(n9800), .ZN(n6274) );
  AOI21_X1 U5302 ( .B1(n8340), .B2(n5421), .A(n5122), .ZN(n5420) );
  NAND2_X1 U5303 ( .A1(n5193), .A2(n8340), .ZN(n5419) );
  INV_X1 U5304 ( .A(n8338), .ZN(n5193) );
  NAND2_X1 U5305 ( .A1(n7878), .A2(n5592), .ZN(n7884) );
  NOR2_X1 U5306 ( .A1(n5107), .A2(n5593), .ZN(n5592) );
  INV_X1 U5307 ( .A(n7877), .ZN(n5593) );
  AOI21_X1 U5308 ( .B1(n5414), .B2(n5416), .A(n5130), .ZN(n5413) );
  INV_X1 U5309 ( .A(n8889), .ZN(n8859) );
  NOR2_X1 U5310 ( .A1(n5187), .A2(n5186), .ZN(n8856) );
  AND2_X1 U5311 ( .A1(n8851), .A2(n8852), .ZN(n5186) );
  AOI21_X1 U5312 ( .B1(n5189), .B2(n5068), .A(n5188), .ZN(n5187) );
  NAND2_X1 U5313 ( .A1(n8846), .A2(n8845), .ZN(n9303) );
  OR2_X1 U5314 ( .A1(n9375), .A2(n9160), .ZN(n5696) );
  AND2_X1 U5315 ( .A1(n5251), .A2(n8811), .ZN(n9366) );
  OAI21_X1 U5316 ( .B1(n9417), .B2(n5511), .A(n5082), .ZN(n5251) );
  INV_X1 U5317 ( .A(n5512), .ZN(n5511) );
  INV_X1 U5318 ( .A(n8055), .ZN(n5516) );
  AOI21_X1 U5319 ( .B1(n5642), .B2(n5641), .A(n5111), .ZN(n5640) );
  NAND2_X1 U5320 ( .A1(n5322), .A2(n5324), .ZN(n9453) );
  AOI21_X1 U5321 ( .B1(n5326), .B2(n5325), .A(n9462), .ZN(n5324) );
  INV_X1 U5322 ( .A(n5328), .ZN(n5325) );
  OR2_X1 U5323 ( .A1(n10023), .A2(n9218), .ZN(n5334) );
  NAND2_X1 U5324 ( .A1(n7684), .A2(n8752), .ZN(n10922) );
  OR2_X1 U5325 ( .A1(n10878), .A2(n7461), .ZN(n8748) );
  INV_X1 U5326 ( .A(n6838), .ZN(n5469) );
  INV_X1 U5327 ( .A(n9486), .ZN(n10923) );
  AND2_X1 U5328 ( .A1(n9104), .A2(n5996), .ZN(n9501) );
  OR2_X1 U5329 ( .A1(n11011), .A2(n5819), .ZN(n8927) );
  NAND2_X2 U5330 ( .A1(n5833), .A2(n8483), .ZN(n5928) );
  AND2_X1 U5331 ( .A1(n8700), .A2(n8854), .ZN(n9486) );
  AND2_X1 U5332 ( .A1(n5979), .A2(n10649), .ZN(n10543) );
  XNOR2_X1 U5333 ( .A(n5766), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5772) );
  OR2_X1 U5334 ( .A1(n5765), .A2(n6287), .ZN(n5766) );
  INV_X1 U5335 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5809) );
  AND4_X1 U5336 ( .A1(n5779), .A2(n5778), .A3(n5733), .A4(n5781), .ZN(n5662)
         );
  INV_X1 U5337 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5726) );
  NOR2_X1 U5338 ( .A1(n10098), .A2(n5681), .ZN(n5680) );
  INV_X1 U5339 ( .A(n10141), .ZN(n5681) );
  AND2_X1 U5340 ( .A1(n10208), .A2(n10114), .ZN(n5688) );
  NOR2_X1 U5341 ( .A1(n7303), .A2(n5669), .ZN(n5670) );
  NAND2_X1 U5342 ( .A1(n5683), .A2(n5679), .ZN(n5678) );
  AOI21_X1 U5343 ( .B1(n10789), .B2(n8616), .A(n8621), .ZN(n8617) );
  NAND2_X1 U5344 ( .A1(n6465), .A2(n10359), .ZN(n7349) );
  INV_X1 U5345 ( .A(n6571), .ZN(n6629) );
  INV_X1 U5346 ( .A(n8254), .ZN(n8209) );
  NOR2_X1 U5347 ( .A1(n8603), .A2(n8466), .ZN(n8665) );
  AOI21_X1 U5348 ( .B1(n9091), .B2(n8254), .A(n8253), .ZN(n10058) );
  INV_X1 U5349 ( .A(n5566), .ZN(n8255) );
  OAI21_X1 U5350 ( .B1(n8217), .B2(n5563), .A(n5560), .ZN(n5566) );
  AOI21_X1 U5351 ( .B1(n10277), .B2(n5561), .A(n5106), .ZN(n5560) );
  NAND2_X1 U5352 ( .A1(n10277), .A2(n5567), .ZN(n5563) );
  NOR2_X1 U5353 ( .A1(n8230), .A2(n5565), .ZN(n5564) );
  INV_X1 U5354 ( .A(n8216), .ZN(n5565) );
  NAND2_X1 U5355 ( .A1(n10454), .A2(n10318), .ZN(n5567) );
  OAI21_X1 U5356 ( .B1(n10365), .B2(n5222), .A(n5220), .ZN(n10306) );
  INV_X1 U5357 ( .A(n5223), .ZN(n5222) );
  AOI21_X1 U5358 ( .B1(n5223), .B2(n5221), .A(n5105), .ZN(n5220) );
  AND2_X1 U5359 ( .A1(n5062), .A2(n5118), .ZN(n5223) );
  AOI21_X1 U5360 ( .B1(n5578), .B2(n10373), .A(n5087), .ZN(n5576) );
  AND2_X1 U5361 ( .A1(n8446), .A2(n8571), .ZN(n10355) );
  INV_X1 U5362 ( .A(n10365), .ZN(n5582) );
  NOR2_X1 U5363 ( .A1(n5558), .A2(n5557), .ZN(n5556) );
  INV_X1 U5364 ( .A(n8106), .ZN(n5558) );
  INV_X1 U5365 ( .A(n8100), .ZN(n5557) );
  NAND2_X1 U5366 ( .A1(n7752), .A2(n5549), .ZN(n5548) );
  OAI21_X1 U5367 ( .B1(n7737), .B2(n8424), .A(n8435), .ZN(n10957) );
  OR2_X1 U5368 ( .A1(n6498), .A2(n8675), .ZN(n11043) );
  INV_X2 U5369 ( .A(n7005), .ZN(n8487) );
  NAND2_X1 U5371 ( .A1(n5258), .A2(n5744), .ZN(n5372) );
  AND2_X1 U5372 ( .A1(n5744), .A2(n9972), .ZN(n5256) );
  NAND2_X1 U5373 ( .A1(n5427), .A2(n5425), .ZN(n6785) );
  INV_X1 U5374 ( .A(n5426), .ZN(n5425) );
  NAND2_X1 U5375 ( .A1(n5799), .A2(n5798), .ZN(n5911) );
  CLKBUF_X1 U5376 ( .A(n5811), .Z(n8483) );
  NAND2_X1 U5377 ( .A1(n5972), .A2(n5996), .ZN(n9466) );
  NAND2_X1 U5378 ( .A1(n5166), .A2(n8850), .ZN(n5165) );
  NAND2_X1 U5379 ( .A1(n8707), .A2(n5167), .ZN(n5166) );
  OR2_X1 U5380 ( .A1(n8709), .A2(n8708), .ZN(n5167) );
  NAND2_X1 U5381 ( .A1(n8711), .A2(n8840), .ZN(n5164) );
  NAND2_X1 U5382 ( .A1(n5174), .A2(n8775), .ZN(n5169) );
  NOR2_X1 U5383 ( .A1(n5098), .A2(n5176), .ZN(n5174) );
  NAND2_X1 U5384 ( .A1(n5083), .A2(n5173), .ZN(n5172) );
  NOR2_X1 U5385 ( .A1(n5175), .A2(n5176), .ZN(n5173) );
  MUX2_X1 U5386 ( .A(n8574), .B(n8573), .S(n8613), .Z(n8575) );
  NOR2_X1 U5387 ( .A1(n5162), .A2(n5161), .ZN(n5160) );
  AND2_X1 U5388 ( .A1(n8814), .A2(n5090), .ZN(n5161) );
  AND2_X1 U5389 ( .A1(n5455), .A2(n7390), .ZN(n5454) );
  NAND2_X1 U5390 ( .A1(n7263), .A2(n7265), .ZN(n5455) );
  OAI21_X1 U5391 ( .B1(n6771), .B2(n6770), .A(n6773), .ZN(n6775) );
  INV_X1 U5392 ( .A(n6769), .ZN(n6770) );
  AOI21_X1 U5393 ( .B1(n5447), .B2(n5610), .A(n5446), .ZN(n5445) );
  INV_X1 U5394 ( .A(n5700), .ZN(n5446) );
  INV_X1 U5395 ( .A(n5448), .ZN(n5447) );
  NAND2_X1 U5396 ( .A1(n6279), .A2(n9799), .ZN(n6370) );
  INV_X1 U5397 ( .A(P2_RD_REG_SCAN_IN), .ZN(n9611) );
  NAND2_X1 U5398 ( .A1(n8939), .A2(n5216), .ZN(n5215) );
  INV_X1 U5399 ( .A(n8846), .ZN(n5248) );
  NOR2_X1 U5400 ( .A1(n5501), .A2(n9445), .ZN(n5500) );
  NOR2_X1 U5401 ( .A1(n9462), .A2(n5502), .ZN(n5501) );
  INV_X1 U5402 ( .A(n8053), .ZN(n5502) );
  OR2_X1 U5403 ( .A1(n10020), .A2(n9465), .ZN(n8776) );
  NAND2_X1 U5404 ( .A1(n7616), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7630) );
  INV_X1 U5405 ( .A(n7617), .ZN(n7616) );
  AND2_X1 U5406 ( .A1(n10994), .A2(n5474), .ZN(n5473) );
  OR2_X1 U5407 ( .A1(n9175), .A2(n10754), .ZN(n8718) );
  NAND2_X1 U5408 ( .A1(n6656), .A2(n6655), .ZN(n8713) );
  NAND2_X1 U5409 ( .A1(n8709), .A2(n6661), .ZN(n8710) );
  NOR2_X1 U5410 ( .A1(n10939), .A2(n10976), .ZN(n5474) );
  NAND2_X1 U5411 ( .A1(n5737), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5740) );
  INV_X1 U5412 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5778) );
  XNOR2_X1 U5413 ( .A(n6585), .B(n9076), .ZN(n6670) );
  NAND2_X1 U5414 ( .A1(n6583), .A2(n6582), .ZN(n6585) );
  NAND2_X1 U5415 ( .A1(n9052), .A2(n9053), .ZN(n5683) );
  INV_X1 U5416 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5714) );
  OR2_X1 U5417 ( .A1(n10464), .A2(n8265), .ZN(n8586) );
  OR2_X1 U5418 ( .A1(n10474), .A2(n10082), .ZN(n8580) );
  NAND2_X1 U5419 ( .A1(n10474), .A2(n10082), .ZN(n8577) );
  NAND2_X1 U5420 ( .A1(n10402), .A2(n5272), .ZN(n5271) );
  INV_X1 U5421 ( .A(n8559), .ZN(n5272) );
  INV_X1 U5422 ( .A(n5487), .ZN(n5268) );
  AOI21_X1 U5423 ( .B1(n5488), .B2(n5490), .A(n5066), .ZN(n5487) );
  OR2_X1 U5424 ( .A1(n10500), .A2(n10400), .ZN(n8559) );
  OR2_X1 U5425 ( .A1(n11061), .A2(n10214), .ZN(n8555) );
  OR2_X1 U5426 ( .A1(n10224), .A2(n10068), .ZN(n8551) );
  OR2_X1 U5427 ( .A1(n10074), .A2(n10156), .ZN(n8544) );
  NOR2_X1 U5428 ( .A1(n10968), .A2(n10984), .ZN(n5391) );
  AND2_X1 U5429 ( .A1(n8432), .A2(n5286), .ZN(n5285) );
  INV_X1 U5430 ( .A(n8521), .ZN(n5286) );
  OAI21_X1 U5431 ( .B1(n10800), .B2(n5110), .A(n5544), .ZN(n5543) );
  AOI21_X1 U5432 ( .B1(n8645), .B2(n5545), .A(n5695), .ZN(n5544) );
  NAND2_X1 U5433 ( .A1(n10823), .A2(n10848), .ZN(n8506) );
  NAND2_X1 U5434 ( .A1(n8404), .A2(n7203), .ZN(n5277) );
  NAND2_X1 U5435 ( .A1(n8414), .A2(n8505), .ZN(n7200) );
  XNOR2_X1 U5436 ( .A(n10731), .B(n10749), .ZN(n6819) );
  AND2_X1 U5437 ( .A1(n6577), .A2(n8483), .ZN(n6609) );
  OAI21_X1 U5438 ( .B1(n7005), .B2(n6594), .A(n5492), .ZN(n5376) );
  OR2_X1 U5439 ( .A1(n6577), .A2(n5491), .ZN(n5492) );
  NAND2_X1 U5440 ( .A1(n6609), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6593) );
  AND2_X1 U5441 ( .A1(n5713), .A2(n5568), .ZN(n5258) );
  AND2_X1 U5442 ( .A1(n5663), .A2(n5370), .ZN(n5568) );
  NOR2_X1 U5443 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5370) );
  INV_X1 U5444 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9743) );
  INV_X1 U5445 ( .A(n7792), .ZN(n5458) );
  NAND2_X1 U5446 ( .A1(n5459), .A2(n7792), .ZN(n7963) );
  OAI21_X1 U5447 ( .B1(n5426), .B2(SI_15_), .A(n5427), .ZN(n6849) );
  AND2_X1 U5448 ( .A1(n6850), .A2(n6790), .ZN(n6848) );
  NOR2_X1 U5449 ( .A1(n6277), .A2(n5615), .ZN(n5614) );
  INV_X1 U5450 ( .A(n6210), .ZN(n5615) );
  INV_X1 U5451 ( .A(n6274), .ZN(n6277) );
  NAND2_X1 U5452 ( .A1(n5430), .A2(n5428), .ZN(n6190) );
  AND2_X1 U5453 ( .A1(n5429), .A2(n5604), .ZN(n5428) );
  AOI21_X1 U5454 ( .B1(n6101), .B2(n5606), .A(n5605), .ZN(n5604) );
  NAND2_X1 U5455 ( .A1(n6103), .A2(n6102), .ZN(n5609) );
  OAI21_X1 U5456 ( .B1(n5803), .B2(n5435), .A(n5433), .ZN(n6103) );
  INV_X1 U5457 ( .A(n5214), .ZN(n5213) );
  OAI22_X1 U5458 ( .A1(n9114), .A2(n5215), .B1(n8939), .B2(n5216), .ZN(n5214)
         );
  OR2_X1 U5459 ( .A1(n8938), .A2(n5215), .ZN(n5212) );
  INV_X1 U5460 ( .A(n6514), .ZN(n5400) );
  XNOR2_X1 U5461 ( .A(n8357), .B(n5196), .ZN(n5402) );
  INV_X1 U5462 ( .A(n5917), .ZN(n5196) );
  NAND2_X1 U5463 ( .A1(n5401), .A2(n5897), .ZN(n9166) );
  NAND2_X1 U5464 ( .A1(n7147), .A2(n7146), .ZN(n7178) );
  NAND2_X1 U5465 ( .A1(n7070), .A2(n7069), .ZN(n7147) );
  NAND2_X1 U5466 ( .A1(n5405), .A2(n5093), .ZN(n9181) );
  INV_X1 U5467 ( .A(n9184), .ZN(n5404) );
  NAND2_X1 U5468 ( .A1(n9181), .A2(n8333), .ZN(n8338) );
  AND2_X1 U5469 ( .A1(n10543), .A2(n5960), .ZN(n6877) );
  AND3_X1 U5470 ( .A1(n8033), .A2(n8032), .A3(n8031), .ZN(n9203) );
  NAND2_X1 U5471 ( .A1(n8687), .A2(n8686), .ZN(n9521) );
  AND2_X1 U5472 ( .A1(n8067), .A2(n8089), .ZN(n8907) );
  OR2_X1 U5473 ( .A1(n9540), .A2(n9203), .ZN(n9323) );
  OR2_X1 U5474 ( .A1(n9543), .A2(n8024), .ZN(n9333) );
  AND2_X1 U5475 ( .A1(n9333), .A2(n8816), .ZN(n9357) );
  INV_X1 U5476 ( .A(n5313), .ZN(n5312) );
  AOI21_X1 U5477 ( .B1(n5313), .B2(n5315), .A(n5071), .ZN(n5311) );
  AOI21_X1 U5478 ( .B1(n5515), .B2(n5519), .A(n5513), .ZN(n5512) );
  INV_X1 U5479 ( .A(n8804), .ZN(n5513) );
  AND2_X1 U5480 ( .A1(n5317), .A2(n5314), .ZN(n9399) );
  NAND2_X1 U5481 ( .A1(n9399), .A2(n9398), .ZN(n9397) );
  INV_X1 U5482 ( .A(n9417), .ZN(n5518) );
  NOR2_X1 U5483 ( .A1(n8798), .A2(n8801), .ZN(n9416) );
  NAND2_X1 U5484 ( .A1(n5638), .A2(n9416), .ZN(n5637) );
  INV_X1 U5485 ( .A(n5640), .ZN(n5638) );
  OR2_X1 U5486 ( .A1(n9438), .A2(n5639), .ZN(n5317) );
  OR2_X1 U5487 ( .A1(n7652), .A2(n9855), .ZN(n7911) );
  AND2_X1 U5488 ( .A1(n9497), .A2(n5333), .ZN(n5328) );
  INV_X1 U5489 ( .A(n5329), .ZN(n5327) );
  NOR2_X1 U5490 ( .A1(n9472), .A2(n5330), .ZN(n5329) );
  INV_X1 U5491 ( .A(n5334), .ZN(n5330) );
  NAND2_X1 U5492 ( .A1(n5332), .A2(n9497), .ZN(n5331) );
  NAND2_X1 U5493 ( .A1(n8050), .A2(n8049), .ZN(n9498) );
  NAND2_X1 U5494 ( .A1(n5655), .A2(n7995), .ZN(n5654) );
  INV_X1 U5495 ( .A(n5657), .ZN(n5655) );
  NOR2_X1 U5496 ( .A1(n8874), .A2(n5658), .ZN(n5657) );
  INV_X1 U5497 ( .A(n5701), .ZN(n5658) );
  AND2_X1 U5498 ( .A1(n7769), .A2(n7768), .ZN(n7771) );
  INV_X1 U5499 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5781) );
  OAI21_X1 U5500 ( .B1(n6796), .B2(n5208), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5782) );
  NAND2_X1 U5501 ( .A1(n5209), .A2(n5778), .ZN(n5208) );
  NAND2_X1 U5502 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n5209) );
  AND2_X1 U5503 ( .A1(n7450), .A2(n8748), .ZN(n5530) );
  AND4_X1 U5504 ( .A1(n7167), .A2(n7166), .A3(n7165), .A4(n7164), .ZN(n8386)
         );
  NAND2_X1 U5505 ( .A1(n10869), .A2(n7416), .ZN(n7420) );
  NAND2_X1 U5506 ( .A1(n5600), .A2(n5599), .ZN(n7425) );
  NAND2_X1 U5507 ( .A1(n5820), .A2(n8895), .ZN(n5600) );
  OAI21_X1 U5508 ( .B1(n8893), .B2(n8708), .A(n8704), .ZN(n5599) );
  NAND2_X1 U5509 ( .A1(n8866), .A2(n5234), .ZN(n5233) );
  INV_X1 U5510 ( .A(n7112), .ZN(n5648) );
  AND2_X1 U5511 ( .A1(n5523), .A2(n5521), .ZN(n5235) );
  AND2_X1 U5512 ( .A1(n8744), .A2(n8742), .ZN(n8866) );
  OR2_X1 U5513 ( .A1(n9221), .A2(n7111), .ZN(n8737) );
  INV_X1 U5514 ( .A(n5524), .ZN(n5523) );
  OAI21_X1 U5515 ( .B1(n8734), .B2(n5525), .A(n7090), .ZN(n5524) );
  NAND2_X1 U5516 ( .A1(n5527), .A2(n8730), .ZN(n5525) );
  NOR2_X1 U5517 ( .A1(n5526), .A2(n8734), .ZN(n5520) );
  INV_X1 U5518 ( .A(n8730), .ZN(n5526) );
  NOR2_X1 U5519 ( .A1(n9170), .A2(n5471), .ZN(n5470) );
  AND2_X1 U5520 ( .A1(n9227), .A2(n6521), .ZN(n6532) );
  OR2_X1 U5521 ( .A1(n6652), .A2(n8887), .ZN(n6869) );
  INV_X1 U5522 ( .A(n9501), .ZN(n9468) );
  NAND2_X1 U5523 ( .A1(n8000), .A2(n7999), .ZN(n9554) );
  NAND2_X1 U5524 ( .A1(n7998), .A2(n7997), .ZN(n9998) );
  AND2_X1 U5525 ( .A1(n7055), .A2(n7054), .ZN(n10872) );
  AND3_X1 U5526 ( .A1(n5932), .A2(n5931), .A3(n5930), .ZN(n7086) );
  OR2_X1 U5527 ( .A1(n5928), .A2(n6083), .ZN(n5932) );
  NAND2_X1 U5528 ( .A1(n6880), .A2(n5942), .ZN(n10925) );
  NAND2_X1 U5529 ( .A1(n5254), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5191) );
  INV_X1 U5530 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5661) );
  INV_X1 U5531 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5779) );
  INV_X1 U5532 ( .A(n5734), .ZN(n6796) );
  INV_X1 U5533 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6791) );
  OR2_X1 U5534 ( .A1(n10140), .A2(n10143), .ZN(n5682) );
  NAND2_X1 U5535 ( .A1(n7303), .A2(n5669), .ZN(n5668) );
  NAND2_X1 U5536 ( .A1(n6600), .A2(n6803), .ZN(n6030) );
  AND2_X1 U5537 ( .A1(n5358), .A2(n5361), .ZN(n6031) );
  NOR2_X1 U5538 ( .A1(n5359), .A2(n5362), .ZN(n5358) );
  NOR2_X1 U5539 ( .A1(n6563), .A2(n10584), .ZN(n5362) );
  NOR2_X1 U5540 ( .A1(n5121), .A2(n5690), .ZN(n5689) );
  INV_X1 U5541 ( .A(n9027), .ZN(n5690) );
  NOR2_X1 U5542 ( .A1(n5354), .A2(n5351), .ZN(n5350) );
  INV_X1 U5543 ( .A(n9034), .ZN(n5351) );
  INV_X1 U5544 ( .A(n5355), .ZN(n5354) );
  AND2_X1 U5545 ( .A1(n10088), .A2(n5356), .ZN(n5355) );
  NAND2_X1 U5546 ( .A1(n10183), .A2(n10188), .ZN(n5356) );
  NOR2_X1 U5547 ( .A1(n10183), .A2(n10188), .ZN(n5357) );
  INV_X1 U5548 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7712) );
  INV_X1 U5549 ( .A(n10165), .ZN(n5675) );
  NAND2_X1 U5550 ( .A1(n6757), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8149) );
  INV_X1 U5551 ( .A(n8123), .ZN(n6757) );
  NAND2_X1 U5552 ( .A1(n9035), .A2(n9034), .ZN(n10184) );
  OR2_X1 U5553 ( .A1(n8222), .A2(n8221), .ZN(n8235) );
  NAND2_X1 U5554 ( .A1(n5436), .A2(n5099), .ZN(n8615) );
  NAND4_X1 U5555 ( .A1(n6475), .A2(n6474), .A3(n6473), .A4(n6472), .ZN(n6804)
         );
  OR2_X1 U5556 ( .A1(n8496), .A2(n6010), .ZN(n6018) );
  NOR2_X1 U5557 ( .A1(n10444), .A2(n8309), .ZN(n10273) );
  AOI21_X1 U5558 ( .B1(n5481), .B2(n5484), .A(n5067), .ZN(n5479) );
  INV_X1 U5559 ( .A(n5481), .ZN(n5480) );
  AND2_X1 U5560 ( .A1(n8250), .A2(n8249), .ZN(n9091) );
  NAND2_X1 U5561 ( .A1(n8268), .A2(n5483), .ZN(n8313) );
  AND2_X1 U5562 ( .A1(n8594), .A2(n10285), .ZN(n10296) );
  OR2_X1 U5563 ( .A1(n10469), .A2(n10337), .ZN(n10329) );
  AND2_X1 U5564 ( .A1(n8586), .A2(n8587), .ZN(n8660) );
  AND2_X1 U5565 ( .A1(n8453), .A2(n8419), .ZN(n10326) );
  INV_X1 U5566 ( .A(n5573), .ZN(n5572) );
  OAI21_X1 U5567 ( .B1(n5575), .B2(n5574), .A(n5583), .ZN(n5573) );
  NAND2_X1 U5568 ( .A1(n5577), .A2(n5077), .ZN(n5574) );
  AND2_X1 U5569 ( .A1(n8580), .A2(n8577), .ZN(n10345) );
  INV_X1 U5570 ( .A(n5584), .ZN(n5579) );
  OR2_X1 U5571 ( .A1(n10484), .A2(n10394), .ZN(n5584) );
  INV_X1 U5572 ( .A(n5489), .ZN(n5488) );
  OAI21_X1 U5573 ( .B1(n8264), .B2(n5490), .A(n10373), .ZN(n5489) );
  INV_X1 U5574 ( .A(n5540), .ZN(n5539) );
  NAND2_X1 U5575 ( .A1(n10390), .A2(n8264), .ZN(n10391) );
  NAND2_X1 U5576 ( .A1(n10399), .A2(n10402), .ZN(n10390) );
  NAND2_X1 U5577 ( .A1(n5542), .A2(n5273), .ZN(n10405) );
  INV_X1 U5578 ( .A(n10403), .ZN(n5542) );
  NAND2_X1 U5579 ( .A1(n8262), .A2(n8559), .ZN(n10399) );
  AOI21_X1 U5580 ( .B1(n5555), .B2(n5554), .A(n10422), .ZN(n5553) );
  INV_X1 U5581 ( .A(n5556), .ZN(n5554) );
  OR2_X1 U5582 ( .A1(n11044), .A2(n11061), .ZN(n11045) );
  AOI21_X1 U5583 ( .B1(n5549), .B2(n5551), .A(n5103), .ZN(n5547) );
  NAND2_X1 U5584 ( .A1(n5548), .A2(n5064), .ZN(n8101) );
  AND2_X1 U5585 ( .A1(n8551), .A2(n8552), .ZN(n8656) );
  AND2_X1 U5586 ( .A1(n8537), .A2(n8436), .ZN(n7751) );
  INV_X1 U5587 ( .A(n5262), .ZN(n7855) );
  AOI21_X1 U5588 ( .B1(n10957), .B2(n8535), .A(n5265), .ZN(n5262) );
  AND2_X1 U5589 ( .A1(n10951), .A2(n7750), .ZN(n7752) );
  NAND2_X1 U5590 ( .A1(n5280), .A2(n5283), .ZN(n7737) );
  AOI21_X1 U5591 ( .B1(n8649), .B2(n8421), .A(n5284), .ZN(n5283) );
  INV_X1 U5592 ( .A(n8526), .ZN(n5284) );
  INV_X1 U5593 ( .A(n10232), .ZN(n7739) );
  NOR2_X1 U5594 ( .A1(n7568), .A2(n10907), .ZN(n10954) );
  AOI21_X1 U5595 ( .B1(n7342), .B2(n7341), .A(n7340), .ZN(n7347) );
  OR2_X1 U5596 ( .A1(n7371), .A2(n10887), .ZN(n7568) );
  NAND2_X1 U5597 ( .A1(n10845), .A2(n8428), .ZN(n5486) );
  OR2_X1 U5598 ( .A1(n10841), .A2(n7472), .ZN(n7371) );
  NAND2_X1 U5599 ( .A1(n7330), .A2(n8506), .ZN(n10845) );
  NAND2_X1 U5600 ( .A1(n7212), .A2(n7325), .ZN(n10844) );
  NAND2_X1 U5601 ( .A1(n8506), .A2(n10844), .ZN(n8645) );
  OR2_X1 U5602 ( .A1(n8501), .A2(n6497), .ZN(n10781) );
  NOR2_X1 U5603 ( .A1(n10727), .A2(n8406), .ZN(n6901) );
  NOR2_X1 U5604 ( .A1(n6803), .A2(n8297), .ZN(n8294) );
  INV_X1 U5605 ( .A(n10779), .ZN(n11040) );
  INV_X1 U5606 ( .A(n10781), .ZN(n11037) );
  NAND2_X1 U5607 ( .A1(n8218), .A2(n8487), .ZN(n8220) );
  AND2_X1 U5608 ( .A1(n7352), .A2(n7351), .ZN(n10851) );
  NOR2_X1 U5609 ( .A1(n6799), .A2(n6495), .ZN(n6503) );
  XNOR2_X1 U5610 ( .A(n8486), .B(n8485), .ZN(n10045) );
  INV_X1 U5611 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9973) );
  XNOR2_X1 U5612 ( .A(n7794), .B(n7790), .ZN(n8191) );
  XNOR2_X1 U5613 ( .A(n6022), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6478) );
  NOR2_X1 U5614 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5672) );
  NAND2_X1 U5615 ( .A1(n5444), .A2(n5610), .ZN(n6488) );
  OR2_X1 U5616 ( .A1(n6206), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U5617 ( .A1(n6211), .A2(n6210), .ZN(n6278) );
  INV_X1 U5618 ( .A(SI_5_), .ZN(n5800) );
  NAND2_X1 U5619 ( .A1(n5218), .A2(n5796), .ZN(n5894) );
  XNOR2_X1 U5620 ( .A(n5795), .B(n9602), .ZN(n5871) );
  OR2_X1 U5621 ( .A1(n5739), .A2(n7761), .ZN(n5979) );
  AND4_X1 U5622 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n7085)
         );
  NAND2_X1 U5623 ( .A1(n5419), .A2(n5420), .ZN(n8918) );
  NAND2_X1 U5624 ( .A1(n8010), .A2(n8009), .ZN(n9549) );
  AND4_X1 U5625 ( .A1(n7895), .A2(n7894), .A3(n7893), .A4(n7892), .ZN(n9467)
         );
  AND4_X1 U5626 ( .A1(n8008), .A2(n8007), .A3(n8006), .A4(n8005), .ZN(n9216)
         );
  NAND2_X1 U5627 ( .A1(n7987), .A2(n7986), .ZN(n9993) );
  NAND2_X1 U5628 ( .A1(n5204), .A2(n5095), .ZN(n7878) );
  OR2_X1 U5629 ( .A1(n8950), .A2(n5206), .ZN(n5205) );
  NAND2_X1 U5630 ( .A1(n7880), .A2(n7879), .ZN(n10015) );
  AND4_X1 U5631 ( .A1(n8017), .A2(n8016), .A3(n8015), .A4(n8014), .ZN(n9160)
         );
  INV_X1 U5632 ( .A(n6521), .ZN(n5464) );
  OAI21_X1 U5633 ( .B1(n5833), .B2(n5253), .A(n5252), .ZN(n6521) );
  NAND2_X1 U5634 ( .A1(n5833), .A2(n10054), .ZN(n5252) );
  NAND2_X1 U5635 ( .A1(n8338), .A2(n9137), .ZN(n8341) );
  NAND2_X1 U5636 ( .A1(n7235), .A2(n7234), .ZN(n8380) );
  AOI21_X1 U5637 ( .B1(n7070), .B2(n5200), .A(n5198), .ZN(n5197) );
  NAND2_X1 U5638 ( .A1(n5199), .A2(n7232), .ZN(n5198) );
  AND4_X1 U5639 ( .A1(n7917), .A2(n7916), .A3(n7915), .A4(n7914), .ZN(n9186)
         );
  NAND2_X1 U5640 ( .A1(n7902), .A2(n7901), .ZN(n10008) );
  INV_X1 U5641 ( .A(n9211), .ZN(n9171) );
  NAND2_X1 U5642 ( .A1(n7628), .A2(n7627), .ZN(n10023) );
  AOI21_X1 U5643 ( .B1(n8697), .B2(n8883), .A(n8701), .ZN(n8698) );
  NAND2_X1 U5644 ( .A1(n5237), .A2(n5236), .ZN(n8697) );
  XNOR2_X1 U5645 ( .A(n8856), .B(n8854), .ZN(n8855) );
  NAND2_X1 U5646 ( .A1(n8889), .A2(n8884), .ZN(n8893) );
  AND4_X1 U5647 ( .A1(n6161), .A2(n6160), .A3(n6159), .A4(n6158), .ZN(n7461)
         );
  INV_X1 U5648 ( .A(n5508), .ZN(n5507) );
  OR2_X1 U5649 ( .A1(n5839), .A2(n5986), .ZN(n5841) );
  OR2_X1 U5650 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  INV_X1 U5651 ( .A(n5534), .ZN(n5533) );
  OR2_X1 U5652 ( .A1(n9305), .A2(n9486), .ZN(n5535) );
  OAI22_X1 U5653 ( .A1(n9308), .A2(n9466), .B1(n9307), .B2(n9306), .ZN(n5534)
         );
  NAND2_X1 U5654 ( .A1(n5158), .A2(n5157), .ZN(n5156) );
  NAND2_X1 U5655 ( .A1(n9213), .A2(n9501), .ZN(n5157) );
  XNOR2_X1 U5656 ( .A(n8084), .B(n8880), .ZN(n9527) );
  NAND2_X1 U5657 ( .A1(n5628), .A2(n5626), .ZN(n8079) );
  NAND2_X1 U5658 ( .A1(n7930), .A2(n7929), .ZN(n10005) );
  NAND2_X1 U5659 ( .A1(n10946), .A2(n10938), .ZN(n9495) );
  INV_X1 U5660 ( .A(n9309), .ZN(n9507) );
  NAND2_X1 U5661 ( .A1(n10946), .A2(n10944), .ZN(n9509) );
  OR2_X1 U5662 ( .A1(n5928), .A2(n6594), .ZN(n5860) );
  NAND2_X1 U5663 ( .A1(n5808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U5664 ( .A1(n5734), .A2(n5465), .ZN(n5808) );
  AND2_X1 U5665 ( .A1(n5659), .A2(n5466), .ZN(n5465) );
  XNOR2_X1 U5666 ( .A(n5780), .B(n5779), .ZN(n8889) );
  NAND2_X1 U5667 ( .A1(n5783), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5780) );
  INV_X1 U5668 ( .A(n5819), .ZN(n8884) );
  NAND2_X1 U5669 ( .A1(n8231), .A2(n8487), .ZN(n8233) );
  AOI21_X1 U5670 ( .B1(n5063), .B2(n5670), .A(n5094), .ZN(n5665) );
  NAND2_X1 U5671 ( .A1(n5341), .A2(n5340), .ZN(n5339) );
  NAND2_X1 U5672 ( .A1(n5346), .A2(n5075), .ZN(n5341) );
  OR2_X1 U5673 ( .A1(n10281), .A2(n8209), .ZN(n8244) );
  NAND2_X1 U5674 ( .A1(n8215), .A2(n8214), .ZN(n10230) );
  OR2_X1 U5675 ( .A1(n8255), .A2(n8662), .ZN(n8256) );
  XNOR2_X1 U5676 ( .A(n5229), .B(n10296), .ZN(n10457) );
  NAND2_X1 U5677 ( .A1(n8217), .A2(n8216), .ZN(n5229) );
  NAND2_X1 U5678 ( .A1(n5165), .A2(n5164), .ZN(n8716) );
  OAI21_X1 U5679 ( .B1(n8534), .B2(n8533), .A(n5109), .ZN(n8540) );
  NOR2_X1 U5680 ( .A1(n5171), .A2(n8780), .ZN(n5170) );
  INV_X1 U5681 ( .A(n8778), .ZN(n5171) );
  AND2_X1 U5682 ( .A1(n8797), .A2(n8798), .ZN(n5183) );
  INV_X1 U5683 ( .A(n8814), .ZN(n5163) );
  INV_X1 U5684 ( .A(n8820), .ZN(n5162) );
  NAND2_X1 U5685 ( .A1(n8584), .A2(n8610), .ZN(n5151) );
  MUX2_X1 U5686 ( .A(n8594), .B(n10285), .S(n8610), .Z(n8595) );
  AOI21_X1 U5687 ( .B1(n8822), .B2(n8025), .A(n8821), .ZN(n8824) );
  INV_X1 U5688 ( .A(SI_12_), .ZN(n9799) );
  INV_X1 U5689 ( .A(SI_9_), .ZN(n9804) );
  INV_X1 U5690 ( .A(n8602), .ZN(n8606) );
  OR2_X1 U5691 ( .A1(n10459), .A2(n10294), .ZN(n8591) );
  INV_X1 U5692 ( .A(n7202), .ZN(n5545) );
  INV_X1 U5693 ( .A(n7265), .ZN(n5452) );
  INV_X1 U5694 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9733) );
  INV_X1 U5695 ( .A(SI_11_), .ZN(n9800) );
  INV_X1 U5696 ( .A(n6139), .ZN(n5605) );
  NAND2_X1 U5697 ( .A1(n5431), .A2(n5435), .ZN(n5429) );
  INV_X1 U5698 ( .A(n5802), .ZN(n5434) );
  INV_X1 U5699 ( .A(n5805), .ZN(n5435) );
  INV_X1 U5700 ( .A(n8943), .ZN(n5216) );
  AND2_X1 U5701 ( .A1(n8842), .A2(n8841), .ZN(n5190) );
  INV_X1 U5702 ( .A(n8853), .ZN(n5188) );
  OR2_X1 U5703 ( .A1(n9521), .A2(n8909), .ZN(n8846) );
  NAND2_X1 U5704 ( .A1(n8839), .A2(n9322), .ZN(n5476) );
  NAND2_X1 U5705 ( .A1(n5512), .A2(n5514), .ZN(n5510) );
  AND2_X1 U5706 ( .A1(n5656), .A2(n7768), .ZN(n5302) );
  AND2_X1 U5707 ( .A1(n7995), .A2(n7770), .ZN(n5656) );
  OR2_X1 U5708 ( .A1(n7162), .A2(n6170), .ZN(n7617) );
  OR2_X1 U5709 ( .A1(n10939), .A2(n8386), .ZN(n8760) );
  INV_X1 U5710 ( .A(n8737), .ZN(n5234) );
  INV_X1 U5711 ( .A(n8729), .ZN(n5527) );
  NOR2_X1 U5712 ( .A1(n9222), .A2(n7086), .ZN(n8734) );
  NAND2_X1 U5713 ( .A1(n9227), .A2(n5464), .ZN(n8858) );
  INV_X1 U5714 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5807) );
  INV_X1 U5715 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6117) );
  INV_X1 U5716 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6118) );
  INV_X1 U5717 ( .A(n9080), .ZN(n6027) );
  XNOR2_X1 U5718 ( .A(n6597), .B(n9083), .ZN(n6602) );
  NAND2_X1 U5719 ( .A1(n10078), .A2(n5345), .ZN(n5344) );
  INV_X1 U5720 ( .A(n5075), .ZN(n5345) );
  AND3_X1 U5721 ( .A1(n7369), .A2(n5363), .A3(n6563), .ZN(n5359) );
  NAND2_X1 U5722 ( .A1(n6908), .A2(n5686), .ZN(n5685) );
  AND2_X1 U5723 ( .A1(n7369), .A2(n6563), .ZN(n6600) );
  INV_X1 U5724 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9738) );
  NOR2_X1 U5725 ( .A1(n10449), .A2(n5380), .ZN(n5379) );
  INV_X1 U5726 ( .A(n5381), .ZN(n5380) );
  INV_X1 U5727 ( .A(n8601), .ZN(n5482) );
  NOR2_X1 U5728 ( .A1(n5564), .A2(n5562), .ZN(n5561) );
  INV_X1 U5729 ( .A(n5567), .ZN(n5562) );
  NAND2_X1 U5730 ( .A1(n9099), .A2(n10058), .ZN(n8601) );
  OR2_X1 U5731 ( .A1(n8248), .A2(n8247), .ZN(n8250) );
  OR2_X1 U5732 ( .A1(n10454), .A2(n10107), .ZN(n8594) );
  NOR2_X1 U5733 ( .A1(n10459), .A2(n10454), .ZN(n5381) );
  INV_X1 U5734 ( .A(n5079), .ZN(n5221) );
  INV_X1 U5735 ( .A(n5576), .ZN(n5575) );
  INV_X1 U5736 ( .A(n10479), .ZN(n5386) );
  OR2_X1 U5737 ( .A1(n10479), .A2(n8166), .ZN(n8446) );
  NOR2_X1 U5738 ( .A1(n10489), .A2(n10484), .ZN(n5387) );
  OAI21_X1 U5739 ( .B1(n5273), .B2(n5541), .A(n8142), .ZN(n5540) );
  INV_X1 U5740 ( .A(n5264), .ZN(n5263) );
  OAI21_X1 U5741 ( .B1(n5265), .B2(n8535), .A(n7854), .ZN(n5264) );
  NAND2_X1 U5742 ( .A1(n5266), .A2(n7751), .ZN(n5265) );
  NAND2_X1 U5743 ( .A1(n8438), .A2(n8535), .ZN(n5266) );
  NOR2_X1 U5744 ( .A1(n8522), .A2(n5282), .ZN(n5281) );
  INV_X1 U5745 ( .A(n5285), .ZN(n5282) );
  NAND2_X1 U5746 ( .A1(n10307), .A2(n5379), .ZN(n10279) );
  AND2_X1 U5747 ( .A1(n10954), .A2(n5065), .ZN(n7869) );
  AND2_X1 U5748 ( .A1(n6593), .A2(n8297), .ZN(n5374) );
  NAND2_X1 U5749 ( .A1(n7969), .A2(n7968), .ZN(n8081) );
  OAI21_X1 U5750 ( .B1(n7484), .B2(n7483), .A(n7482), .ZN(n7578) );
  OAI21_X1 U5751 ( .B1(n7264), .B2(n5453), .A(n5450), .ZN(n7484) );
  AOI21_X1 U5752 ( .B1(n5454), .B2(n5452), .A(n5451), .ZN(n5450) );
  INV_X1 U5753 ( .A(n5454), .ZN(n5453) );
  INV_X1 U5754 ( .A(n7392), .ZN(n5451) );
  AND2_X1 U5755 ( .A1(n7392), .A2(n7269), .ZN(n7390) );
  AND3_X1 U5756 ( .A1(n9956), .A2(n9734), .A3(n9733), .ZN(n6020) );
  NAND2_X1 U5757 ( .A1(n6851), .A2(n5073), .ZN(n5603) );
  NAND2_X1 U5758 ( .A1(n6849), .A2(n6848), .ZN(n6851) );
  INV_X1 U5759 ( .A(n6844), .ZN(n6852) );
  AND2_X1 U5760 ( .A1(n6775), .A2(n6774), .ZN(n5426) );
  NAND2_X1 U5761 ( .A1(n6777), .A2(n6776), .ZN(n5427) );
  INV_X1 U5762 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5745) );
  XNOR2_X1 U5763 ( .A(n6772), .B(n9588), .ZN(n6769) );
  NAND2_X1 U5764 ( .A1(n5443), .A2(n5441), .ZN(n6771) );
  AOI21_X1 U5765 ( .B1(n5445), .B2(n5611), .A(n5442), .ZN(n5441) );
  INV_X1 U5766 ( .A(n6489), .ZN(n5442) );
  NOR2_X1 U5767 ( .A1(n5080), .A2(n5449), .ZN(n5448) );
  INV_X1 U5768 ( .A(n5699), .ZN(n5449) );
  INV_X1 U5769 ( .A(SI_10_), .ZN(n6193) );
  NAND2_X1 U5770 ( .A1(n5911), .A2(n5910), .ZN(n5803) );
  INV_X1 U5771 ( .A(SI_4_), .ZN(n9812) );
  NAND2_X1 U5772 ( .A1(n5786), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U5773 ( .A1(n5787), .A2(n5619), .ZN(n5618) );
  INV_X1 U5774 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5619) );
  INV_X1 U5775 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5785) );
  NAND2_X1 U5776 ( .A1(n5963), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6156) );
  INV_X1 U5777 ( .A(n7146), .ZN(n5203) );
  NOR2_X1 U5778 ( .A1(n5418), .A2(n8916), .ZN(n5417) );
  INV_X1 U5779 ( .A(n5420), .ZN(n5418) );
  AOI21_X1 U5780 ( .B1(n5408), .B2(n5407), .A(n5139), .ZN(n5406) );
  INV_X1 U5781 ( .A(n7926), .ZN(n5407) );
  OR2_X1 U5782 ( .A1(n7927), .A2(n5409), .ZN(n5405) );
  AND2_X1 U5783 ( .A1(n5587), .A2(n8371), .ZN(n5586) );
  OR2_X1 U5784 ( .A1(n7605), .A2(n5059), .ZN(n5587) );
  NAND2_X1 U5785 ( .A1(n5200), .A2(n5203), .ZN(n5199) );
  AND2_X1 U5786 ( .A1(n5594), .A2(n5201), .ZN(n5200) );
  NAND2_X1 U5787 ( .A1(n7146), .A2(n5202), .ZN(n5201) );
  AND2_X1 U5788 ( .A1(n7158), .A2(n7151), .ZN(n5594) );
  INV_X1 U5789 ( .A(n7069), .ZN(n5202) );
  NAND2_X1 U5790 ( .A1(n7884), .A2(n7886), .ZN(n7927) );
  NAND2_X1 U5791 ( .A1(n5240), .A2(n5239), .ZN(n5238) );
  INV_X1 U5792 ( .A(n5241), .ZN(n5239) );
  INV_X1 U5793 ( .A(n5244), .ZN(n5240) );
  AOI22_X1 U5794 ( .A1(n5244), .A2(n5246), .B1(n5241), .B2(n5243), .ZN(n5236)
         );
  INV_X1 U5795 ( .A(n5247), .ZN(n5243) );
  AOI21_X1 U5796 ( .B1(n9124), .B2(n8095), .A(n7985), .ZN(n9202) );
  OR2_X1 U5797 ( .A1(n6401), .A2(n6313), .ZN(n6548) );
  AND2_X1 U5798 ( .A1(n6733), .A2(n6732), .ZN(n6995) );
  NAND2_X1 U5799 ( .A1(n5993), .A2(n5833), .ZN(n5985) );
  NAND2_X1 U5800 ( .A1(n9214), .A2(n9499), .ZN(n5158) );
  INV_X1 U5801 ( .A(n9292), .ZN(n5627) );
  INV_X1 U5802 ( .A(n9324), .ZN(n5631) );
  AOI21_X1 U5803 ( .B1(n9324), .B2(n5630), .A(n5129), .ZN(n5629) );
  INV_X1 U5804 ( .A(n8034), .ZN(n5630) );
  NAND2_X1 U5805 ( .A1(n8836), .A2(n8835), .ZN(n9292) );
  NOR2_X1 U5806 ( .A1(n9340), .A2(n9534), .ZN(n9318) );
  INV_X1 U5807 ( .A(n5299), .ZN(n5298) );
  OAI21_X1 U5808 ( .B1(n8058), .B2(n5300), .A(n9334), .ZN(n5299) );
  NAND2_X1 U5809 ( .A1(n9323), .A2(n8825), .ZN(n9334) );
  NOR2_X1 U5810 ( .A1(n8058), .A2(n8812), .ZN(n5616) );
  INV_X1 U5811 ( .A(n9334), .ZN(n9332) );
  NAND2_X1 U5812 ( .A1(n5301), .A2(n8058), .ZN(n9349) );
  INV_X1 U5813 ( .A(n7938), .ZN(n7937) );
  OR2_X1 U5814 ( .A1(n7988), .A2(n9845), .ZN(n8002) );
  AOI21_X1 U5815 ( .B1(n5500), .B2(n5502), .A(n5104), .ZN(n5498) );
  NAND2_X1 U5816 ( .A1(n9457), .A2(n9444), .ZN(n9439) );
  INV_X1 U5817 ( .A(n7645), .ZN(n7644) );
  NAND2_X1 U5818 ( .A1(n10929), .A2(n5070), .ZN(n9491) );
  NAND2_X1 U5819 ( .A1(n10929), .A2(n5473), .ZN(n7784) );
  NAND2_X1 U5820 ( .A1(n7780), .A2(n7779), .ZN(n8050) );
  AND2_X1 U5821 ( .A1(n8761), .A2(n8762), .ZN(n8872) );
  NAND2_X1 U5822 ( .A1(n10929), .A2(n10928), .ZN(n10926) );
  OAI21_X1 U5823 ( .B1(n7418), .B2(n5652), .A(n5650), .ZN(n10918) );
  AOI21_X1 U5824 ( .B1(n5651), .B2(n8868), .A(n5123), .ZN(n5650) );
  OAI21_X1 U5825 ( .B1(n6966), .B2(n5527), .A(n8730), .ZN(n7091) );
  NAND2_X1 U5826 ( .A1(n6956), .A2(n10754), .ZN(n6958) );
  NAND2_X1 U5827 ( .A1(n5255), .A2(n8713), .ZN(n6949) );
  NAND2_X1 U5828 ( .A1(n6535), .A2(n6887), .ZN(n5528) );
  AND2_X1 U5829 ( .A1(n6654), .A2(n6653), .ZN(n6657) );
  NAND2_X1 U5830 ( .A1(n8863), .A2(n8710), .ZN(n8707) );
  NAND2_X1 U5831 ( .A1(n6535), .A2(n6887), .ZN(n8863) );
  NAND2_X1 U5832 ( .A1(n6660), .A2(n6661), .ZN(n6534) );
  NAND2_X1 U5833 ( .A1(n6877), .A2(n6876), .ZN(n6889) );
  NAND2_X1 U5834 ( .A1(n8028), .A2(n8027), .ZN(n9540) );
  NAND2_X1 U5835 ( .A1(n8019), .A2(n8018), .ZN(n9543) );
  AND2_X1 U5836 ( .A1(n7464), .A2(n7463), .ZN(n7465) );
  INV_X1 U5837 ( .A(n11011), .ZN(n10927) );
  AND2_X1 U5838 ( .A1(n5659), .A2(n5537), .ZN(n5536) );
  AND2_X1 U5839 ( .A1(n5692), .A2(n5810), .ZN(n5537) );
  AND2_X1 U5840 ( .A1(n5467), .A2(n5807), .ZN(n5466) );
  NAND2_X1 U5841 ( .A1(n5084), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5777) );
  AND2_X1 U5842 ( .A1(n5662), .A2(n5661), .ZN(n5660) );
  INV_X1 U5843 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7313) );
  INV_X1 U5844 ( .A(n5668), .ZN(n5666) );
  OR2_X1 U5845 ( .A1(n8182), .A2(n8181), .ZN(n8195) );
  INV_X1 U5846 ( .A(n5343), .ZN(n5342) );
  OAI21_X1 U5847 ( .B1(n5060), .B2(n5344), .A(n10077), .ZN(n5343) );
  INV_X1 U5848 ( .A(n5347), .ZN(n5346) );
  OAI21_X1 U5849 ( .B1(n5060), .B2(n5075), .A(n5348), .ZN(n5347) );
  NAND2_X1 U5850 ( .A1(n5342), .A2(n5344), .ZN(n5340) );
  NAND2_X1 U5851 ( .A1(n6624), .A2(n6625), .ZN(n6674) );
  OR2_X1 U5852 ( .A1(n8170), .A2(n10167), .ZN(n8182) );
  INV_X1 U5853 ( .A(n5683), .ZN(n5677) );
  NAND2_X1 U5854 ( .A1(n10184), .A2(n10183), .ZN(n10187) );
  INV_X1 U5855 ( .A(n7022), .ZN(n7020) );
  OAI21_X1 U5856 ( .B1(n10152), .B2(n5364), .A(n5365), .ZN(n10208) );
  INV_X1 U5857 ( .A(n5366), .ZN(n5364) );
  AOI21_X1 U5858 ( .B1(n5367), .B2(n5366), .A(n5128), .ZN(n5365) );
  AOI22_X1 U5859 ( .A1(n9014), .A2(n9011), .B1(n9010), .B2(n10150), .ZN(n5366)
         );
  NOR2_X1 U5860 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5371) );
  INV_X1 U5861 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9967) );
  OR2_X1 U5862 ( .A1(n6144), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U5863 ( .A1(n8474), .A2(n8473), .ZN(n8609) );
  NAND2_X1 U5864 ( .A1(n10307), .A2(n5377), .ZN(n8309) );
  AND2_X1 U5865 ( .A1(n5379), .A2(n5378), .ZN(n5377) );
  NAND2_X1 U5866 ( .A1(n10307), .A2(n10314), .ZN(n10308) );
  INV_X1 U5867 ( .A(n8585), .ZN(n10317) );
  NAND2_X1 U5868 ( .A1(n10409), .A2(n5383), .ZN(n10337) );
  NOR2_X1 U5869 ( .A1(n5385), .A2(n10474), .ZN(n5383) );
  OR2_X1 U5870 ( .A1(n8149), .A2(n6758), .ZN(n8160) );
  NAND2_X1 U5871 ( .A1(n5269), .A2(n5267), .ZN(n10354) );
  AOI21_X1 U5872 ( .B1(n5270), .B2(n5273), .A(n5268), .ZN(n5267) );
  AND2_X1 U5873 ( .A1(n5488), .A2(n5271), .ZN(n5270) );
  NAND2_X1 U5874 ( .A1(n10409), .A2(n5387), .ZN(n10366) );
  NAND2_X1 U5875 ( .A1(n10409), .A2(n10388), .ZN(n10383) );
  AND2_X1 U5876 ( .A1(n10429), .A2(n10414), .ZN(n10409) );
  NAND2_X1 U5877 ( .A1(n6756), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8111) );
  INV_X1 U5878 ( .A(n7858), .ZN(n6756) );
  NOR2_X1 U5879 ( .A1(n11045), .A2(n10500), .ZN(n10429) );
  NAND2_X1 U5880 ( .A1(n10954), .A2(n5389), .ZN(n11044) );
  AND2_X1 U5881 ( .A1(n5065), .A2(n11024), .ZN(n5389) );
  INV_X1 U5882 ( .A(n6584), .ZN(n7369) );
  INV_X1 U5883 ( .A(n5259), .ZN(n8260) );
  AOI21_X1 U5884 ( .B1(n10957), .B2(n5263), .A(n5260), .ZN(n5259) );
  NAND2_X1 U5885 ( .A1(n5261), .A2(n8544), .ZN(n5260) );
  NAND2_X1 U5886 ( .A1(n5263), .A2(n5265), .ZN(n5261) );
  NAND2_X1 U5887 ( .A1(n6755), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U5888 ( .A1(n10954), .A2(n5391), .ZN(n7816) );
  NAND2_X1 U5889 ( .A1(n10954), .A2(n10955), .ZN(n10952) );
  INV_X1 U5890 ( .A(n7550), .ZN(n6754) );
  OR2_X1 U5891 ( .A1(n7314), .A2(n7313), .ZN(n7356) );
  NAND2_X1 U5892 ( .A1(n6753), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7550) );
  INV_X1 U5893 ( .A(n7356), .ZN(n6753) );
  NAND2_X1 U5894 ( .A1(n7354), .A2(n8649), .ZN(n7565) );
  NAND2_X1 U5895 ( .A1(n5287), .A2(n8514), .ZN(n7354) );
  NAND2_X1 U5896 ( .A1(n5486), .A2(n5285), .ZN(n5287) );
  NAND2_X1 U5897 ( .A1(n6182), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7289) );
  INV_X1 U5898 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7288) );
  NAND2_X1 U5899 ( .A1(n10838), .A2(n7328), .ZN(n7342) );
  AND2_X1 U5900 ( .A1(n10807), .A2(n10823), .ZN(n10842) );
  NOR2_X1 U5901 ( .A1(n10808), .A2(n10814), .ZN(n10807) );
  OR2_X1 U5902 ( .A1(n10770), .A2(n10774), .ZN(n7199) );
  OAI21_X1 U5903 ( .B1(n7205), .B2(n5277), .A(n8409), .ZN(n5275) );
  INV_X1 U5904 ( .A(n7200), .ZN(n10801) );
  NAND2_X1 U5905 ( .A1(n5373), .A2(n10728), .ZN(n10727) );
  INV_X1 U5906 ( .A(n8643), .ZN(n6816) );
  NAND2_X1 U5907 ( .A1(n8307), .A2(n8306), .ZN(n10444) );
  OR2_X1 U5908 ( .A1(n6498), .A2(n6461), .ZN(n11047) );
  XNOR2_X1 U5909 ( .A(n8478), .B(n8477), .ZN(n9109) );
  XNOR2_X1 U5910 ( .A(n8468), .B(n8467), .ZN(n8684) );
  XNOR2_X1 U5911 ( .A(n8081), .B(n8080), .ZN(n8392) );
  XNOR2_X1 U5912 ( .A(n7837), .B(n7958), .ZN(n8231) );
  NAND2_X1 U5913 ( .A1(n7832), .A2(n7831), .ZN(n7837) );
  OR2_X1 U5914 ( .A1(n7963), .A2(n7828), .ZN(n7832) );
  XNOR2_X1 U5915 ( .A(n5717), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U5916 ( .A1(n5716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5717) );
  XNOR2_X1 U5917 ( .A(n7843), .B(n7842), .ZN(n8218) );
  OAI21_X1 U5918 ( .B1(n7729), .B2(n5137), .A(n5456), .ZN(n7843) );
  INV_X1 U5919 ( .A(n5457), .ZN(n5456) );
  XNOR2_X1 U5920 ( .A(n5721), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U5921 ( .A1(n5720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5721) );
  OR2_X1 U5922 ( .A1(n5753), .A2(n5752), .ZN(n5755) );
  XNOR2_X1 U5923 ( .A(n7484), .B(n7480), .ZN(n8156) );
  NAND2_X1 U5924 ( .A1(n5613), .A2(n6276), .ZN(n6369) );
  NAND2_X1 U5925 ( .A1(n6211), .A2(n5614), .ZN(n5613) );
  NAND2_X1 U5926 ( .A1(n5609), .A2(n5606), .ZN(n6140) );
  NAND2_X1 U5927 ( .A1(n5609), .A2(n6105), .ZN(n6111) );
  NAND2_X1 U5928 ( .A1(n5792), .A2(n5791), .ZN(n5845) );
  OAI21_X1 U5929 ( .B1(n7833), .B2(n5424), .A(n5296), .ZN(n5423) );
  OR2_X1 U5930 ( .A1(n5811), .A2(n6592), .ZN(n5296) );
  NAND2_X1 U5931 ( .A1(n8365), .A2(n5937), .ZN(n5958) );
  NAND2_X1 U5932 ( .A1(n8938), .A2(n9114), .ZN(n9117) );
  OAI21_X1 U5933 ( .B1(n8380), .B2(n5416), .A(n5414), .ZN(n8982) );
  AND4_X1 U5934 ( .A1(n7636), .A2(n7635), .A3(n7634), .A4(n7633), .ZN(n8969)
         );
  NAND2_X1 U5935 ( .A1(n7178), .A2(n7151), .ZN(n7156) );
  OAI21_X1 U5936 ( .B1(n7070), .B2(n5203), .A(n5200), .ZN(n7233) );
  NAND2_X1 U5937 ( .A1(n5411), .A2(n7928), .ZN(n8328) );
  NAND2_X1 U5938 ( .A1(n7927), .A2(n7926), .ZN(n5411) );
  INV_X1 U5939 ( .A(n8945), .ZN(n5598) );
  NAND2_X1 U5940 ( .A1(n9214), .A2(n9189), .ZN(n5597) );
  AND2_X1 U5941 ( .A1(n5213), .A2(n9167), .ZN(n5211) );
  NOR2_X1 U5942 ( .A1(n9523), .A2(n9195), .ZN(n5393) );
  NAND2_X1 U5943 ( .A1(n5877), .A2(n5464), .ZN(n5834) );
  NAND2_X1 U5944 ( .A1(n8921), .A2(n8920), .ZN(n9145) );
  NAND2_X1 U5945 ( .A1(n9145), .A2(n9146), .ZN(n9197) );
  NAND2_X1 U5946 ( .A1(n5398), .A2(n5396), .ZN(n8967) );
  OR2_X1 U5947 ( .A1(n5897), .A2(n5399), .ZN(n5398) );
  INV_X1 U5948 ( .A(n5900), .ZN(n5399) );
  OR2_X1 U5949 ( .A1(n8963), .A2(n5195), .ZN(n5194) );
  INV_X1 U5950 ( .A(n5402), .ZN(n5195) );
  NAND2_X1 U5951 ( .A1(n7878), .A2(n7877), .ZN(n7885) );
  OR2_X1 U5952 ( .A1(n6678), .A2(n5928), .ZN(n5321) );
  AND2_X1 U5953 ( .A1(n5895), .A2(n5319), .ZN(n5318) );
  NAND2_X1 U5954 ( .A1(n5856), .A2(n5320), .ZN(n5319) );
  AND2_X1 U5955 ( .A1(n6069), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9188) );
  NAND2_X1 U5956 ( .A1(n5405), .A2(n5406), .ZN(n9183) );
  OAI21_X1 U5957 ( .B1(n8380), .B2(n5059), .A(n5586), .ZN(n8979) );
  NAND2_X1 U5958 ( .A1(n8380), .A2(n7605), .ZN(n8391) );
  INV_X1 U5959 ( .A(n5590), .ZN(n5589) );
  OAI21_X1 U5960 ( .B1(n9146), .B2(n5591), .A(n9194), .ZN(n5590) );
  AND4_X1 U5961 ( .A1(n7651), .A2(n7650), .A3(n7649), .A4(n7648), .ZN(n9465)
         );
  NAND2_X1 U5962 ( .A1(n5207), .A2(n8950), .ZN(n8956) );
  INV_X1 U5963 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9912) );
  AND4_X1 U5964 ( .A1(n6168), .A2(n6167), .A3(n6166), .A4(n6165), .ZN(n8372)
         );
  AND4_X1 U5965 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .ZN(n7448)
         );
  INV_X1 U5966 ( .A(P2_U3966), .ZN(n9226) );
  AND2_X1 U5967 ( .A1(n6400), .A2(n6399), .ZN(n6401) );
  AND2_X1 U5968 ( .A1(n6781), .A2(n6510), .ZN(n7613) );
  NAND2_X1 U5969 ( .A1(n5997), .A2(n5833), .ZN(n5998) );
  NAND2_X1 U5970 ( .A1(n8695), .A2(n8694), .ZN(n9510) );
  NAND2_X1 U5971 ( .A1(n9365), .A2(n8815), .ZN(n9358) );
  INV_X1 U5972 ( .A(n9543), .ZN(n8025) );
  AOI21_X1 U5973 ( .B1(n5311), .B2(n5312), .A(n8057), .ZN(n5309) );
  NAND2_X1 U5974 ( .A1(n5308), .A2(n5311), .ZN(n9370) );
  OR2_X1 U5975 ( .A1(n9438), .A2(n5312), .ZN(n5308) );
  NAND2_X1 U5976 ( .A1(n5509), .A2(n5512), .ZN(n9387) );
  NAND2_X1 U5977 ( .A1(n9417), .A2(n5515), .ZN(n5509) );
  NAND2_X1 U5978 ( .A1(n9397), .A2(n5636), .ZN(n9380) );
  NAND2_X1 U5979 ( .A1(n5517), .A2(n8055), .ZN(n9393) );
  NAND2_X1 U5980 ( .A1(n5518), .A2(n5058), .ZN(n5517) );
  OAI21_X1 U5981 ( .B1(n9438), .B2(n5643), .A(n5640), .ZN(n9412) );
  AND2_X1 U5982 ( .A1(n5644), .A2(n5086), .ZN(n9425) );
  NAND2_X1 U5983 ( .A1(n5644), .A2(n5642), .ZN(n9423) );
  NAND2_X1 U5984 ( .A1(n9438), .A2(n9445), .ZN(n5644) );
  NAND2_X1 U5985 ( .A1(n5499), .A2(n8053), .ZN(n9446) );
  NAND2_X1 U5986 ( .A1(n9463), .A2(n9462), .ZN(n5499) );
  NAND2_X1 U5987 ( .A1(n5323), .A2(n5326), .ZN(n9455) );
  NAND2_X1 U5988 ( .A1(n5332), .A2(n5328), .ZN(n5323) );
  NAND2_X1 U5989 ( .A1(n5331), .A2(n5334), .ZN(n9471) );
  NAND2_X1 U5990 ( .A1(n7777), .A2(n5701), .ZN(n7778) );
  NAND2_X1 U5991 ( .A1(n7771), .A2(n7770), .ZN(n7777) );
  OR2_X1 U5992 ( .A1(n5782), .A2(n5781), .ZN(n5784) );
  NAND2_X1 U5993 ( .A1(n7449), .A2(n8748), .ZN(n7452) );
  NAND2_X1 U5994 ( .A1(n7144), .A2(n7143), .ZN(n10878) );
  INV_X1 U5995 ( .A(n10872), .ZN(n7415) );
  AND2_X1 U5996 ( .A1(n5645), .A2(n5646), .ZN(n10869) );
  NOR2_X1 U5997 ( .A1(n8866), .A2(n5648), .ZN(n5647) );
  NAND2_X1 U5998 ( .A1(n7110), .A2(n8735), .ZN(n5649) );
  NAND2_X1 U5999 ( .A1(n5232), .A2(n8737), .ZN(n7421) );
  NAND2_X1 U6000 ( .A1(n5235), .A2(n5522), .ZN(n5232) );
  NAND2_X1 U6001 ( .A1(n5522), .A2(n5523), .ZN(n7101) );
  AND3_X1 U6002 ( .A1(n5915), .A2(n5914), .A3(n5913), .ZN(n6881) );
  NOR2_X1 U6003 ( .A1(n5464), .A2(n6538), .ZN(n6939) );
  NAND2_X1 U6004 ( .A1(n10543), .A2(n6870), .ZN(n10935) );
  AOI21_X1 U6005 ( .B1(n9495), .B2(n9309), .A(n5464), .ZN(n6893) );
  INV_X2 U6006 ( .A(n11017), .ZN(n11018) );
  NAND2_X1 U6007 ( .A1(n9522), .A2(n5306), .ZN(n10030) );
  NOR2_X1 U6008 ( .A1(n9519), .A2(n5307), .ZN(n5306) );
  OR2_X1 U6009 ( .A1(n9520), .A2(n5132), .ZN(n5307) );
  XNOR2_X1 U6010 ( .A(n5735), .B(P2_IR_REG_26__SCAN_IN), .ZN(n10540) );
  AND2_X1 U6011 ( .A1(n5981), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10649) );
  INV_X1 U6012 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n10046) );
  XNOR2_X1 U6013 ( .A(n5736), .B(P2_IR_REG_25__SCAN_IN), .ZN(n10541) );
  NAND2_X1 U6014 ( .A1(n5734), .A2(n5659), .ZN(n5761) );
  INV_X1 U6015 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7488) );
  XNOR2_X1 U6016 ( .A(n5422), .B(n5661), .ZN(n8708) );
  NAND2_X1 U6017 ( .A1(n5085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5422) );
  INV_X1 U6018 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7302) );
  INV_X1 U6019 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7192) );
  OAI21_X1 U6020 ( .B1(n6796), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6980) );
  INV_X1 U6021 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6487) );
  INV_X1 U6022 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6289) );
  INV_X1 U6023 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6201) );
  INV_X1 U6024 ( .A(n7212), .ZN(n10823) );
  INV_X1 U6025 ( .A(n5337), .ZN(n5336) );
  AND4_X1 U6026 ( .A1(n6607), .A2(n6608), .A3(n6606), .A4(n6605), .ZN(n6808)
         );
  INV_X1 U6027 ( .A(n10184), .ZN(n5352) );
  OR2_X1 U6028 ( .A1(n7285), .A2(n7284), .ZN(n7305) );
  NAND2_X1 U6029 ( .A1(n5682), .A2(n10141), .ZN(n10097) );
  NAND2_X1 U6030 ( .A1(n8193), .A2(n8192), .ZN(n10464) );
  NAND2_X1 U6031 ( .A1(n8191), .A2(n8487), .ZN(n8193) );
  NAND2_X1 U6032 ( .A1(n6674), .A2(n6673), .ZN(n6907) );
  OR2_X1 U6033 ( .A1(n7285), .A2(n5670), .ZN(n5667) );
  NAND2_X1 U6034 ( .A1(n7308), .A2(n7307), .ZN(n7472) );
  AOI21_X1 U6035 ( .B1(n5355), .B2(n5357), .A(n5127), .ZN(n5353) );
  AND2_X1 U6036 ( .A1(n5676), .A2(n5060), .ZN(n10164) );
  NAND2_X1 U6037 ( .A1(n5676), .A2(n5081), .ZN(n10166) );
  NAND2_X1 U6038 ( .A1(n7536), .A2(n7535), .ZN(n10907) );
  INV_X1 U6039 ( .A(n10126), .ZN(n10218) );
  OAI21_X1 U6040 ( .B1(n10184), .B2(n10183), .A(n10188), .ZN(n10087) );
  AND2_X1 U6041 ( .A1(n8235), .A2(n8223), .ZN(n10300) );
  NAND2_X1 U6042 ( .A1(n5702), .A2(n9014), .ZN(n5684) );
  NAND2_X1 U6043 ( .A1(n5754), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U6044 ( .A1(n8202), .A2(n8201), .ZN(n10327) );
  OR2_X1 U6045 ( .A1(n8209), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6574) );
  OR2_X1 U6046 ( .A1(n6629), .A2(n6572), .ZN(n6573) );
  CLKBUF_X1 U6047 ( .A(n6804), .Z(n10732) );
  OR2_X1 U6048 ( .A1(n6203), .A2(n6012), .ZN(n6017) );
  INV_X1 U6049 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5295) );
  INV_X1 U6050 ( .A(n8609), .ZN(n10442) );
  NOR2_X1 U6051 ( .A1(n8305), .A2(n8304), .ZN(n8308) );
  NOR2_X1 U6052 ( .A1(n5378), .A2(n10058), .ZN(n8304) );
  AND2_X1 U6053 ( .A1(n8323), .A2(n8322), .ZN(n10446) );
  NAND2_X1 U6054 ( .A1(n8272), .A2(n8271), .ZN(n8900) );
  OR2_X1 U6055 ( .A1(n8259), .A2(n10851), .ZN(n8272) );
  NAND2_X1 U6056 ( .A1(n5559), .A2(n5567), .ZN(n10278) );
  NAND2_X1 U6057 ( .A1(n8217), .A2(n5564), .ZN(n5559) );
  AOI21_X1 U6058 ( .B1(n10448), .B2(n10291), .A(n10290), .ZN(n5290) );
  AND2_X1 U6059 ( .A1(n5293), .A2(n5292), .ZN(n10451) );
  AOI22_X1 U6060 ( .A1(n10288), .A2(n11037), .B1(n11040), .B2(n10318), .ZN(
        n5292) );
  NAND2_X1 U6061 ( .A1(n10289), .A2(n11035), .ZN(n5293) );
  INV_X1 U6062 ( .A(n5227), .ZN(n10456) );
  OAI21_X1 U6063 ( .B1(n10457), .B2(n10851), .A(n5228), .ZN(n5227) );
  AOI21_X1 U6064 ( .B1(n10298), .B2(n11035), .A(n10297), .ZN(n5228) );
  NAND2_X1 U6065 ( .A1(n5224), .A2(n5062), .ZN(n8276) );
  NAND2_X1 U6066 ( .A1(n10365), .A2(n5079), .ZN(n5224) );
  NAND2_X1 U6067 ( .A1(n8180), .A2(n8179), .ZN(n10469) );
  OAI21_X1 U6068 ( .B1(n10365), .B2(n5088), .A(n5572), .ZN(n10323) );
  NAND2_X1 U6069 ( .A1(n5571), .A2(n5576), .ZN(n10336) );
  NAND2_X1 U6070 ( .A1(n10365), .A2(n5578), .ZN(n5571) );
  NAND2_X1 U6071 ( .A1(n5580), .A2(n5578), .ZN(n10351) );
  NAND2_X1 U6072 ( .A1(n5582), .A2(n5581), .ZN(n5580) );
  OAI21_X1 U6073 ( .B1(n10390), .B2(n5490), .A(n5488), .ZN(n10372) );
  NAND2_X1 U6074 ( .A1(n10391), .A2(n8567), .ZN(n10374) );
  NAND2_X1 U6075 ( .A1(n10405), .A2(n8131), .ZN(n10382) );
  NAND2_X1 U6076 ( .A1(n5552), .A2(n5555), .ZN(n10421) );
  NAND2_X1 U6077 ( .A1(n8101), .A2(n5556), .ZN(n5552) );
  NAND2_X1 U6078 ( .A1(n8105), .A2(n8104), .ZN(n11061) );
  NAND2_X1 U6079 ( .A1(n11032), .A2(n11033), .ZN(n11031) );
  NAND2_X1 U6080 ( .A1(n8101), .A2(n8100), .ZN(n11032) );
  NAND2_X1 U6081 ( .A1(n5548), .A2(n5547), .ZN(n7852) );
  NAND2_X1 U6082 ( .A1(n7850), .A2(n7849), .ZN(n10224) );
  NAND2_X1 U6083 ( .A1(n7822), .A2(n7821), .ZN(n7845) );
  OAI21_X1 U6084 ( .B1(n10957), .B2(n8438), .A(n8535), .ZN(n7740) );
  NAND2_X1 U6085 ( .A1(n7735), .A2(n7734), .ZN(n10984) );
  NAND2_X1 U6086 ( .A1(n7346), .A2(n7345), .ZN(n10887) );
  OR2_X1 U6087 ( .A1(n11043), .A2(n6480), .ZN(n10786) );
  NAND2_X1 U6088 ( .A1(n5486), .A2(n8432), .ZN(n7353) );
  NAND2_X1 U6089 ( .A1(n10798), .A2(n7202), .ZN(n7326) );
  NAND2_X1 U6090 ( .A1(n5279), .A2(n8404), .ZN(n10775) );
  OR2_X1 U6091 ( .A1(n7204), .A2(n7203), .ZN(n5279) );
  CLKBUF_X1 U6093 ( .A(n10178), .Z(n10740) );
  INV_X1 U6094 ( .A(n10430), .ZN(n11060) );
  INV_X1 U6095 ( .A(n10786), .ZN(n11059) );
  AND2_X2 U6096 ( .A1(n6503), .A2(n6496), .ZN(n11054) );
  AND2_X1 U6097 ( .A1(n6563), .A2(n6123), .ZN(n6479) );
  NAND2_X1 U6098 ( .A1(n5257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6009) );
  MUX2_X1 U6099 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5757), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5758) );
  INV_X1 U6100 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9679) );
  INV_X1 U6101 ( .A(n8618), .ZN(n8667) );
  INV_X1 U6102 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9684) );
  INV_X1 U6103 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9683) );
  INV_X1 U6104 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6846) );
  INV_X1 U6105 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9908) );
  INV_X1 U6106 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9916) );
  INV_X1 U6107 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6162) );
  XNOR2_X1 U6108 ( .A(n5894), .B(n5893), .ZN(n6678) );
  XNOR2_X1 U6109 ( .A(n5423), .B(n5857), .ZN(n6594) );
  NOR2_X1 U6110 ( .A1(n7517), .A2(n7516), .ZN(n10572) );
  NOR2_X1 U6111 ( .A1(n10570), .A2(n10569), .ZN(n7516) );
  NAND2_X1 U6112 ( .A1(n5394), .A2(n5392), .ZN(P2_U3222) );
  AOI21_X1 U6113 ( .B1(n8944), .B2(n5393), .A(n5596), .ZN(n5392) );
  NAND2_X1 U6114 ( .A1(n5395), .A2(n9523), .ZN(n5394) );
  NAND2_X1 U6115 ( .A1(n5598), .A2(n5597), .ZN(n5596) );
  OAI22_X1 U6116 ( .A1(n9198), .A2(n5463), .B1(n5464), .B2(n9195), .ZN(n6520)
         );
  NAND2_X1 U6117 ( .A1(n8341), .A2(n8340), .ZN(n8913) );
  NOR3_X1 U6118 ( .A1(n8892), .A2(n8891), .A3(n8890), .ZN(n8899) );
  NOR2_X1 U6119 ( .A1(n9526), .A2(n9426), .ZN(n8097) );
  NAND2_X1 U6120 ( .A1(n5532), .A2(n5531), .ZN(P2_U3549) );
  OR2_X1 U6121 ( .A1(n11018), .A2(n8092), .ZN(n5531) );
  NAND2_X1 U6122 ( .A1(n10030), .A2(n11018), .ZN(n5532) );
  NAND2_X1 U6123 ( .A1(n5305), .A2(n5303), .ZN(P2_U3517) );
  OR2_X1 U6124 ( .A1(n11001), .A2(n5304), .ZN(n5303) );
  NAND2_X1 U6125 ( .A1(n10030), .A2(n11001), .ZN(n5305) );
  INV_X1 U6126 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5304) );
  OAI21_X1 U6127 ( .B1(n10446), .B2(n11070), .A(n5493), .ZN(P1_U3355) );
  AOI21_X1 U6128 ( .B1(n10443), .B2(n10291), .A(n5494), .ZN(n5493) );
  OAI21_X1 U6129 ( .B1(n10447), .B2(n11064), .A(n5495), .ZN(n5494) );
  INV_X1 U6130 ( .A(n8324), .ZN(n5495) );
  NAND2_X1 U6131 ( .A1(n5291), .A2(n5288), .ZN(P1_U3264) );
  INV_X1 U6132 ( .A(n5289), .ZN(n5288) );
  OR2_X1 U6133 ( .A1(n10451), .A2(n11070), .ZN(n5291) );
  OAI21_X1 U6134 ( .B1(n10452), .B2(n11064), .A(n5290), .ZN(n5289) );
  OR2_X1 U6135 ( .A1(n9998), .A2(n9431), .ZN(n5058) );
  AND2_X1 U6136 ( .A1(n10207), .A2(n10208), .ZN(n10112) );
  INV_X1 U6137 ( .A(n7284), .ZN(n5669) );
  INV_X1 U6138 ( .A(n9445), .ZN(n5641) );
  INV_X1 U6139 ( .A(n5506), .ZN(n5901) );
  AND2_X1 U6140 ( .A1(n8373), .A2(n7607), .ZN(n5059) );
  AND2_X1 U6141 ( .A1(n8776), .A2(n8777), .ZN(n9472) );
  AND2_X1 U6142 ( .A1(n5081), .A2(n5675), .ZN(n5060) );
  XOR2_X1 U6143 ( .A(n9009), .B(n9083), .Z(n5061) );
  NAND2_X1 U6144 ( .A1(n5705), .A2(n5704), .ZN(n6082) );
  AND2_X1 U6145 ( .A1(n8629), .A2(n8597), .ZN(n10286) );
  AND2_X1 U6146 ( .A1(n5225), .A2(n8190), .ZN(n5062) );
  AND2_X1 U6147 ( .A1(n8706), .A2(n9483), .ZN(n8857) );
  INV_X1 U6148 ( .A(n10373), .ZN(n5581) );
  NOR2_X1 U6149 ( .A1(n7434), .A2(n5666), .ZN(n5063) );
  AND2_X1 U6150 ( .A1(n7851), .A2(n5547), .ZN(n5064) );
  INV_X1 U6151 ( .A(n8663), .ZN(n5439) );
  AND2_X1 U6152 ( .A1(n5391), .A2(n5390), .ZN(n5065) );
  AND2_X1 U6153 ( .A1(n10484), .A2(n10093), .ZN(n5066) );
  INV_X1 U6154 ( .A(n10318), .ZN(n10107) );
  NAND2_X1 U6155 ( .A1(n8229), .A2(n8228), .ZN(n10318) );
  AND2_X1 U6156 ( .A1(n8665), .A2(n5482), .ZN(n5067) );
  AND2_X1 U6157 ( .A1(n8849), .A2(n5101), .ZN(n5068) );
  NAND2_X1 U6158 ( .A1(n8169), .A2(n8168), .ZN(n10474) );
  OR2_X1 U6159 ( .A1(n10469), .A2(n10346), .ZN(n5069) );
  AND2_X1 U6160 ( .A1(n5473), .A2(n5472), .ZN(n5070) );
  NAND2_X1 U6161 ( .A1(n9385), .A2(n9216), .ZN(n5635) );
  AND2_X1 U6162 ( .A1(n5633), .A2(n5635), .ZN(n5071) );
  INV_X1 U6163 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U6164 ( .A1(n9972), .A2(n9973), .ZN(n5072) );
  AND2_X1 U6165 ( .A1(n6976), .A2(n6850), .ZN(n5073) );
  INV_X1 U6166 ( .A(n9137), .ZN(n5421) );
  AND2_X1 U6167 ( .A1(n8748), .A2(n8746), .ZN(n8868) );
  NAND2_X2 U6168 ( .A1(n8619), .A2(n10789), .ZN(n8613) );
  AND2_X1 U6169 ( .A1(n6965), .A2(n5623), .ZN(n5074) );
  INV_X1 U6170 ( .A(n5403), .ZN(n5401) );
  AND2_X1 U6171 ( .A1(n9055), .A2(n9056), .ZN(n5075) );
  AND2_X1 U6172 ( .A1(n5888), .A2(n5726), .ZN(n5812) );
  INV_X1 U6173 ( .A(n9528), .ZN(n9127) );
  NAND2_X1 U6174 ( .A1(n7978), .A2(n7977), .ZN(n9528) );
  NOR2_X1 U6175 ( .A1(n9523), .A2(n9308), .ZN(n5076) );
  NAND2_X1 U6176 ( .A1(n10474), .A2(n10356), .ZN(n5077) );
  NOR3_X1 U6177 ( .A1(n9340), .A2(n5476), .A3(n9528), .ZN(n5078) );
  AND2_X1 U6178 ( .A1(n5572), .A2(n5069), .ZN(n5079) );
  INV_X1 U6179 ( .A(n8775), .ZN(n5175) );
  OR2_X1 U6180 ( .A1(n6368), .A2(n5612), .ZN(n5080) );
  NAND2_X1 U6181 ( .A1(n9424), .A2(n5086), .ZN(n5643) );
  INV_X1 U6182 ( .A(n5058), .ZN(n5519) );
  INV_X1 U6183 ( .A(n6437), .ZN(n5320) );
  OR2_X1 U6184 ( .A1(n5680), .A2(n5677), .ZN(n5081) );
  AND2_X1 U6185 ( .A1(n9379), .A2(n5510), .ZN(n5082) );
  INV_X1 U6186 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5733) );
  AND3_X1 U6187 ( .A1(n8771), .A2(n8874), .A3(n8770), .ZN(n5083) );
  NAND2_X1 U6188 ( .A1(n5734), .A2(n5660), .ZN(n5084) );
  NAND2_X1 U6189 ( .A1(n5734), .A2(n5662), .ZN(n5085) );
  NAND2_X1 U6190 ( .A1(n5258), .A2(n5256), .ZN(n5257) );
  NAND2_X1 U6191 ( .A1(n9444), .A2(n9467), .ZN(n5086) );
  NAND2_X1 U6192 ( .A1(n9349), .A2(n8026), .ZN(n9331) );
  AND2_X1 U6193 ( .A1(n10113), .A2(n9027), .ZN(n10121) );
  AND2_X1 U6194 ( .A1(n10479), .A2(n10375), .ZN(n5087) );
  NAND2_X1 U6195 ( .A1(n5576), .A2(n5077), .ZN(n5088) );
  NOR2_X1 U6196 ( .A1(n10164), .A2(n5075), .ZN(n5089) );
  AND2_X1 U6197 ( .A1(n8809), .A2(n8850), .ZN(n5090) );
  NAND2_X1 U6198 ( .A1(n7975), .A2(n9112), .ZN(n5506) );
  NOR2_X1 U6199 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5846) );
  INV_X1 U6200 ( .A(n8297), .ZN(n5363) );
  AND2_X1 U6201 ( .A1(n5846), .A2(n5496), .ZN(n5888) );
  OAI21_X1 U6202 ( .B1(n5352), .B2(n5357), .A(n5355), .ZN(n10086) );
  AND2_X1 U6203 ( .A1(n8976), .A2(n7612), .ZN(n5091) );
  INV_X1 U6204 ( .A(n9369), .ZN(n8057) );
  NOR2_X1 U6205 ( .A1(n5723), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U6206 ( .A1(n10207), .A2(n5688), .ZN(n10113) );
  INV_X1 U6207 ( .A(n8704), .ZN(n8895) );
  XNOR2_X1 U6208 ( .A(n5777), .B(n5178), .ZN(n8704) );
  XNOR2_X1 U6209 ( .A(n9224), .B(n9170), .ZN(n8719) );
  AND2_X1 U6210 ( .A1(n8562), .A2(n8563), .ZN(n10402) );
  INV_X1 U6211 ( .A(n10402), .ZN(n5273) );
  AND2_X1 U6212 ( .A1(n8268), .A2(n8629), .ZN(n5092) );
  AND2_X1 U6213 ( .A1(n5406), .A2(n5404), .ZN(n5093) );
  NAND2_X1 U6214 ( .A1(n8205), .A2(n8204), .ZN(n10459) );
  NAND2_X1 U6215 ( .A1(n7225), .A2(n7224), .ZN(n10939) );
  INV_X1 U6216 ( .A(n5611), .ZN(n5610) );
  OAI21_X1 U6217 ( .B1(n5614), .B2(n5080), .A(n6370), .ZN(n5611) );
  AND2_X1 U6218 ( .A1(n7433), .A2(n7432), .ZN(n5094) );
  AND2_X1 U6219 ( .A1(n5205), .A2(n7660), .ZN(n5095) );
  INV_X1 U6220 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6287) );
  INV_X1 U6221 ( .A(n10754), .ZN(n5471) );
  NAND2_X1 U6222 ( .A1(n10307), .A2(n5381), .ZN(n5382) );
  AND2_X1 U6223 ( .A1(n10355), .A2(n10373), .ZN(n5096) );
  AND2_X1 U6224 ( .A1(n5580), .A2(n5584), .ZN(n5097) );
  INV_X1 U6225 ( .A(n5484), .ZN(n5483) );
  NAND2_X1 U6226 ( .A1(n8598), .A2(n8629), .ZN(n5484) );
  INV_X1 U6227 ( .A(n6881), .ZN(n8965) );
  INV_X1 U6228 ( .A(n5315), .ZN(n5314) );
  NAND2_X1 U6229 ( .A1(n5637), .A2(n5316), .ZN(n5315) );
  AND2_X1 U6230 ( .A1(n8857), .A2(n8774), .ZN(n5098) );
  OR2_X1 U6231 ( .A1(n8631), .A2(n8613), .ZN(n5099) );
  AND2_X1 U6232 ( .A1(n8598), .A2(n8599), .ZN(n5100) );
  AND2_X1 U6233 ( .A1(n8847), .A2(n8848), .ZN(n5101) );
  NAND2_X1 U6234 ( .A1(n8233), .A2(n8232), .ZN(n10449) );
  AND2_X1 U6235 ( .A1(n5682), .A2(n5680), .ZN(n5102) );
  OR2_X1 U6236 ( .A1(n9220), .A2(n10872), .ZN(n8744) );
  NOR2_X1 U6237 ( .A1(n10074), .A2(n10231), .ZN(n5103) );
  INV_X1 U6238 ( .A(n5607), .ZN(n5606) );
  NAND2_X1 U6239 ( .A1(n6105), .A2(n5608), .ZN(n5607) );
  NOR2_X1 U6240 ( .A1(n10008), .A2(n9467), .ZN(n5104) );
  NOR2_X1 U6241 ( .A1(n10464), .A2(n10327), .ZN(n5105) );
  NOR2_X1 U6242 ( .A1(n10449), .A2(n10229), .ZN(n5106) );
  AND3_X1 U6243 ( .A1(n5705), .A2(n5672), .A3(n5671), .ZN(n5744) );
  INV_X1 U6244 ( .A(n5636), .ZN(n5634) );
  OR2_X1 U6245 ( .A1(n9993), .A2(n9418), .ZN(n5636) );
  INV_X1 U6246 ( .A(n5385), .ZN(n5384) );
  NAND2_X1 U6247 ( .A1(n5387), .A2(n5386), .ZN(n5385) );
  AND2_X1 U6248 ( .A1(n7881), .A2(n7882), .ZN(n5107) );
  NAND2_X1 U6249 ( .A1(n5535), .A2(n5533), .ZN(n9519) );
  NAND2_X1 U6250 ( .A1(n8462), .A2(n8601), .ZN(n8662) );
  AND2_X1 U6251 ( .A1(n5806), .A2(SI_6_), .ZN(n5108) );
  AND2_X1 U6252 ( .A1(n8532), .A2(n8531), .ZN(n5109) );
  INV_X1 U6253 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9943) );
  XOR2_X1 U6254 ( .A(n9076), .B(n9057), .Z(n10078) );
  INV_X1 U6255 ( .A(n10078), .ZN(n5348) );
  INV_X1 U6256 ( .A(n8404), .ZN(n5278) );
  NAND2_X1 U6257 ( .A1(n8645), .A2(n7200), .ZN(n5110) );
  AND2_X1 U6258 ( .A1(n8781), .A2(n8780), .ZN(n9454) );
  NAND2_X1 U6259 ( .A1(n8689), .A2(n8688), .ZN(n9514) );
  NAND2_X1 U6260 ( .A1(n8220), .A2(n8219), .ZN(n10454) );
  AND2_X1 U6261 ( .A1(n8489), .A2(n8488), .ZN(n10439) );
  NOR2_X1 U6262 ( .A1(n7996), .A2(n9186), .ZN(n5111) );
  OAI21_X1 U6263 ( .B1(n9398), .B2(n5634), .A(n9386), .ZN(n5633) );
  INV_X1 U6264 ( .A(n5643), .ZN(n5642) );
  NAND2_X1 U6265 ( .A1(n8655), .A2(n8106), .ZN(n5555) );
  AND2_X1 U6266 ( .A1(n5371), .A2(n5714), .ZN(n5663) );
  AND3_X1 U6267 ( .A1(n5180), .A2(n5179), .A3(n5178), .ZN(n5112) );
  AND2_X1 U6268 ( .A1(n9114), .A2(n8943), .ZN(n5113) );
  AND2_X1 U6269 ( .A1(n5483), .A2(n8665), .ZN(n5114) );
  NAND2_X1 U6270 ( .A1(n8713), .A2(n8712), .ZN(n6708) );
  INV_X1 U6271 ( .A(n6708), .ZN(n5529) );
  INV_X1 U6272 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5467) );
  AND2_X1 U6273 ( .A1(n8432), .A2(n8520), .ZN(n10846) );
  AND2_X1 U6274 ( .A1(n5400), .A2(n5900), .ZN(n5115) );
  AND2_X1 U6275 ( .A1(n5233), .A2(n8744), .ZN(n5116) );
  NAND2_X1 U6276 ( .A1(n5327), .A2(n5333), .ZN(n5326) );
  INV_X1 U6277 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9972) );
  AND2_X1 U6278 ( .A1(n5555), .A2(n5064), .ZN(n5117) );
  INV_X1 U6279 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U6280 ( .A1(n10464), .A2(n10327), .ZN(n5118) );
  OR2_X1 U6281 ( .A1(n5346), .A2(n5342), .ZN(n5119) );
  INV_X1 U6282 ( .A(n8370), .ZN(n10994) );
  NAND2_X1 U6283 ( .A1(n7610), .A2(n7609), .ZN(n8370) );
  INV_X1 U6284 ( .A(n5409), .ZN(n5408) );
  OR2_X1 U6285 ( .A1(n8327), .A2(n5410), .ZN(n5409) );
  INV_X1 U6286 ( .A(n7639), .ZN(n5206) );
  NAND2_X1 U6287 ( .A1(n8246), .A2(n8245), .ZN(n9099) );
  INV_X1 U6288 ( .A(n9099), .ZN(n5378) );
  XNOR2_X1 U6289 ( .A(n10056), .B(n10055), .ZN(n5120) );
  NAND2_X1 U6290 ( .A1(n5310), .A2(n5309), .ZN(n9371) );
  INV_X1 U6291 ( .A(n10140), .ZN(n5679) );
  INV_X1 U6292 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5424) );
  OR2_X1 U6293 ( .A1(n8973), .A2(n9500), .ZN(n7995) );
  INV_X1 U6294 ( .A(n8567), .ZN(n5490) );
  INV_X1 U6295 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9744) );
  AND2_X1 U6296 ( .A1(n10123), .A2(n9032), .ZN(n5121) );
  NAND2_X1 U6297 ( .A1(n7752), .A2(n8652), .ZN(n7822) );
  INV_X1 U6298 ( .A(n5578), .ZN(n5577) );
  NOR2_X1 U6299 ( .A1(n10355), .A2(n5579), .ZN(n5578) );
  INV_X1 U6300 ( .A(n5515), .ZN(n5514) );
  NOR2_X1 U6301 ( .A1(n8056), .A2(n5516), .ZN(n5515) );
  AND2_X1 U6302 ( .A1(n8912), .A2(n8911), .ZN(n5122) );
  INV_X1 U6303 ( .A(n9322), .ZN(n9534) );
  AND2_X1 U6304 ( .A1(n8037), .A2(n8036), .ZN(n9322) );
  NAND2_X1 U6305 ( .A1(n8083), .A2(n8082), .ZN(n9523) );
  AND2_X1 U6306 ( .A1(n7679), .A2(n7678), .ZN(n5123) );
  NAND2_X1 U6307 ( .A1(n10409), .A2(n5384), .ZN(n5388) );
  INV_X1 U6308 ( .A(n5468), .ZN(n9432) );
  NOR2_X1 U6309 ( .A1(n9439), .A2(n10005), .ZN(n5468) );
  AND2_X1 U6310 ( .A1(n5317), .A2(n5637), .ZN(n5124) );
  AND2_X1 U6311 ( .A1(n7777), .A2(n5657), .ZN(n5125) );
  AND2_X1 U6312 ( .A1(n5331), .A2(n5329), .ZN(n5126) );
  NOR2_X1 U6313 ( .A1(n9043), .A2(n9042), .ZN(n5127) );
  NAND2_X1 U6314 ( .A1(n7418), .A2(n7417), .ZN(n7464) );
  XOR2_X1 U6315 ( .A(n9017), .B(n9076), .Z(n5128) );
  AND2_X1 U6316 ( .A1(n9322), .A2(n9121), .ZN(n5129) );
  AND2_X1 U6317 ( .A1(n7625), .A2(n7624), .ZN(n5130) );
  AND2_X1 U6318 ( .A1(n7187), .A2(SI_18_), .ZN(n5131) );
  INV_X1 U6319 ( .A(n5652), .ZN(n5651) );
  NAND2_X1 U6320 ( .A1(n8869), .A2(n7463), .ZN(n5652) );
  NAND2_X1 U6321 ( .A1(n8737), .A2(n8738), .ZN(n8735) );
  INV_X1 U6322 ( .A(n8735), .ZN(n5521) );
  AND2_X1 U6323 ( .A1(n9521), .A2(n10925), .ZN(n5132) );
  NOR2_X1 U6324 ( .A1(n8962), .A2(n5194), .ZN(n5133) );
  INV_X1 U6325 ( .A(n8131), .ZN(n5541) );
  AND2_X1 U6326 ( .A1(n5120), .A2(n9075), .ZN(n5134) );
  NAND2_X1 U6327 ( .A1(n5667), .A2(n5668), .ZN(n7435) );
  INV_X1 U6328 ( .A(n8026), .ZN(n5300) );
  AND2_X1 U6329 ( .A1(n7682), .A2(n7681), .ZN(n5135) );
  INV_X1 U6330 ( .A(n8926), .ZN(n5591) );
  NOR2_X1 U6331 ( .A1(n5673), .A2(n6082), .ZN(n5136) );
  INV_X1 U6332 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U6333 ( .A1(n7615), .A2(n7614), .ZN(n8973) );
  INV_X1 U6334 ( .A(n8973), .ZN(n5472) );
  NAND2_X1 U6335 ( .A1(n7464), .A2(n5651), .ZN(n7680) );
  XNOR2_X1 U6336 ( .A(n5751), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U6337 ( .A1(n7804), .A2(n7803), .ZN(n10074) );
  INV_X1 U6338 ( .A(n10074), .ZN(n5390) );
  OR2_X1 U6339 ( .A1(n5458), .A2(n7961), .ZN(n5137) );
  NOR2_X1 U6340 ( .A1(n9212), .A2(n8708), .ZN(n5138) );
  NAND2_X1 U6341 ( .A1(n7285), .A2(n7284), .ZN(n7304) );
  NAND2_X1 U6342 ( .A1(n5674), .A2(n7018), .ZN(n7019) );
  AND2_X1 U6343 ( .A1(n7932), .A2(n7931), .ZN(n5139) );
  NAND2_X1 U6344 ( .A1(n5744), .A2(n5713), .ZN(n5723) );
  NAND2_X1 U6345 ( .A1(n5649), .A2(n7112), .ZN(n7113) );
  AND2_X1 U6346 ( .A1(n10929), .A2(n5474), .ZN(n5140) );
  NOR2_X1 U6347 ( .A1(n6513), .A2(n6514), .ZN(n5403) );
  NAND2_X1 U6348 ( .A1(n5546), .A2(n7200), .ZN(n10798) );
  AND2_X1 U6349 ( .A1(n9003), .A2(n9004), .ZN(n10150) );
  INV_X1 U6350 ( .A(n10150), .ZN(n5368) );
  INV_X1 U6351 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5179) );
  INV_X1 U6352 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5180) );
  AND2_X1 U6353 ( .A1(n10917), .A2(n7681), .ZN(n5141) );
  AND2_X1 U6354 ( .A1(n5659), .A2(n5467), .ZN(n5142) );
  NAND2_X1 U6355 ( .A1(n5734), .A2(n5142), .ZN(n5143) );
  INV_X1 U6356 ( .A(n10226), .ZN(n10197) );
  INV_X1 U6357 ( .A(n9227), .ZN(n5463) );
  INV_X1 U6358 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U6359 ( .A1(n6532), .A2(n6534), .ZN(n6654) );
  NAND2_X1 U6360 ( .A1(n5375), .A2(n5374), .ZN(n10726) );
  INV_X1 U6361 ( .A(n10726), .ZN(n5373) );
  NAND2_X1 U6362 ( .A1(n6683), .A2(n6684), .ZN(n5144) );
  OR2_X1 U6363 ( .A1(n10618), .A2(n5295), .ZN(n5145) );
  AND2_X1 U6364 ( .A1(n5055), .A2(n5833), .ZN(n5146) );
  NAND2_X1 U6365 ( .A1(n8704), .A2(n8708), .ZN(n10713) );
  INV_X1 U6366 ( .A(n10713), .ZN(n5462) );
  AND2_X1 U6367 ( .A1(n6521), .A2(n5462), .ZN(n5147) );
  INV_X1 U6368 ( .A(n6591), .ZN(n5491) );
  INV_X1 U6369 ( .A(n10662), .ZN(n5253) );
  NAND2_X1 U6370 ( .A1(n5148), .A2(n5096), .ZN(n8576) );
  NAND2_X1 U6371 ( .A1(n8570), .A2(n8569), .ZN(n5148) );
  NAND2_X1 U6372 ( .A1(n5151), .A2(n5149), .ZN(n8589) );
  NAND2_X1 U6373 ( .A1(n5150), .A2(n8613), .ZN(n5149) );
  NAND2_X1 U6374 ( .A1(n8583), .A2(n8582), .ZN(n5150) );
  NAND2_X2 U6375 ( .A1(n5152), .A2(n5274), .ZN(n10802) );
  NAND2_X1 U6376 ( .A1(n5276), .A2(n7204), .ZN(n5152) );
  NAND2_X1 U6377 ( .A1(n5219), .A2(n5794), .ZN(n5294) );
  OAI211_X1 U6378 ( .C1(n8607), .C2(n8610), .A(n5440), .B(n5438), .ZN(n5437)
         );
  NAND2_X1 U6379 ( .A1(n5437), .A2(n8631), .ZN(n5436) );
  NAND2_X1 U6380 ( .A1(n5230), .A2(n8873), .ZN(n7780) );
  NAND2_X1 U6381 ( .A1(n5831), .A2(n6025), .ZN(n5790) );
  NAND2_X1 U6382 ( .A1(n5231), .A2(n8872), .ZN(n7762) );
  AND2_X2 U6383 ( .A1(n5154), .A2(n5116), .ZN(n7422) );
  NAND2_X1 U6384 ( .A1(n5235), .A2(n5155), .ZN(n5154) );
  AND2_X1 U6385 ( .A1(n5522), .A2(n8866), .ZN(n5155) );
  NAND2_X1 U6386 ( .A1(n5423), .A2(n5857), .ZN(n5792) );
  AOI21_X2 U6387 ( .B1(n8096), .B2(n10923), .A(n5156), .ZN(n9526) );
  NAND2_X1 U6388 ( .A1(n5159), .A2(n5160), .ZN(n8822) );
  OR2_X1 U6389 ( .A1(n8810), .A2(n5163), .ZN(n5159) );
  NAND2_X1 U6390 ( .A1(n5168), .A2(n8779), .ZN(n8785) );
  NAND3_X1 U6391 ( .A1(n5172), .A2(n5170), .A3(n5169), .ZN(n5168) );
  NAND3_X1 U6392 ( .A1(n5172), .A2(n8778), .A3(n5169), .ZN(n8783) );
  INV_X1 U6393 ( .A(n9472), .ZN(n5176) );
  NAND3_X1 U6394 ( .A1(n5185), .A2(n5184), .A3(n8797), .ZN(n8802) );
  OR2_X1 U6395 ( .A1(n8794), .A2(n8840), .ZN(n5184) );
  OR2_X1 U6396 ( .A1(n8793), .A2(n8850), .ZN(n5185) );
  NAND2_X1 U6397 ( .A1(n5181), .A2(n8800), .ZN(n5182) );
  NAND3_X1 U6398 ( .A1(n5184), .A2(n5185), .A3(n5183), .ZN(n5181) );
  AOI21_X1 U6399 ( .B1(n8803), .B2(n5182), .A(n9398), .ZN(n8806) );
  NAND3_X1 U6400 ( .A1(n8844), .A2(n8843), .A3(n5190), .ZN(n5189) );
  NAND2_X2 U6401 ( .A1(n5833), .A2(n7833), .ZN(n5858) );
  XNOR2_X1 U6402 ( .A(n5191), .B(n5810), .ZN(n5971) );
  INV_X1 U6403 ( .A(n5197), .ZN(n7235) );
  NAND2_X1 U6404 ( .A1(n5413), .A2(n5412), .ZN(n5207) );
  NAND3_X1 U6405 ( .A1(n5413), .A2(n5412), .A3(n7639), .ZN(n5204) );
  NAND3_X1 U6406 ( .A1(n5212), .A2(n5211), .A3(n5210), .ZN(n5217) );
  NAND2_X1 U6407 ( .A1(n8938), .A2(n5113), .ZN(n5210) );
  NAND3_X1 U6408 ( .A1(n5212), .A2(n5213), .A3(n5210), .ZN(n8944) );
  NAND2_X1 U6409 ( .A1(n5217), .A2(n9211), .ZN(n5395) );
  NAND2_X1 U6410 ( .A1(n5294), .A2(n5871), .ZN(n5218) );
  NAND2_X1 U6411 ( .A1(n5845), .A2(n5844), .ZN(n5219) );
  NAND3_X1 U6412 ( .A1(n5572), .A2(n5088), .A3(n5069), .ZN(n5225) );
  INV_X4 U6413 ( .A(n5811), .ZN(n7833) );
  NAND2_X1 U6414 ( .A1(n5548), .A2(n5117), .ZN(n5226) );
  NAND2_X1 U6415 ( .A1(n5226), .A2(n5553), .ZN(n10419) );
  NAND2_X1 U6416 ( .A1(n7762), .A2(n8762), .ZN(n5230) );
  NAND2_X1 U6417 ( .A1(n7686), .A2(n8758), .ZN(n5231) );
  NAND2_X1 U6418 ( .A1(n8683), .A2(n5238), .ZN(n5237) );
  AOI21_X1 U6419 ( .B1(n8683), .B2(n8880), .A(n5076), .ZN(n9304) );
  AOI21_X1 U6420 ( .B1(n5247), .B2(n5245), .A(n5138), .ZN(n5244) );
  NOR2_X1 U6421 ( .A1(n5249), .A2(n8702), .ZN(n5245) );
  NAND2_X1 U6422 ( .A1(n5247), .A2(n8849), .ZN(n5246) );
  AOI21_X2 U6423 ( .B1(n5249), .B2(n5076), .A(n5248), .ZN(n5247) );
  NAND2_X2 U6424 ( .A1(n8054), .A2(n8789), .ZN(n9417) );
  NAND3_X1 U6425 ( .A1(n5734), .A2(n5659), .A3(n5692), .ZN(n5254) );
  NAND3_X1 U6426 ( .A1(n5528), .A2(n8710), .A3(n5529), .ZN(n5255) );
  NAND3_X1 U6427 ( .A1(n7350), .A2(n7122), .A3(n6803), .ZN(n5361) );
  NAND2_X1 U6428 ( .A1(n8262), .A2(n5270), .ZN(n5269) );
  INV_X1 U6429 ( .A(n5275), .ZN(n5274) );
  NOR2_X1 U6430 ( .A1(n7205), .A2(n5278), .ZN(n5276) );
  NAND2_X1 U6431 ( .A1(n10802), .A2(n10801), .ZN(n7206) );
  NAND2_X1 U6432 ( .A1(n5486), .A2(n5281), .ZN(n5280) );
  XNOR2_X1 U6433 ( .A(n5294), .B(n5871), .ZN(n6581) );
  NAND2_X1 U6434 ( .A1(n5295), .A2(n5785), .ZN(n5787) );
  NAND3_X1 U6435 ( .A1(n10266), .A2(n10265), .A3(n5145), .ZN(P1_U3260) );
  MUX2_X1 U6436 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7833), .Z(n5795) );
  MUX2_X1 U6437 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7833), .Z(n5797) );
  MUX2_X1 U6438 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7833), .Z(n6104) );
  MUX2_X1 U6439 ( .A(n6784), .B(n9908), .S(n7833), .Z(n6776) );
  MUX2_X1 U6440 ( .A(n6786), .B(n6846), .S(n7833), .Z(n6788) );
  NAND2_X1 U6441 ( .A1(n9351), .A2(n8026), .ZN(n5297) );
  NAND2_X1 U6442 ( .A1(n5297), .A2(n5298), .ZN(n8035) );
  INV_X1 U6443 ( .A(n9351), .ZN(n5301) );
  NAND2_X1 U6444 ( .A1(n10917), .A2(n5135), .ZN(n7769) );
  NAND2_X1 U6445 ( .A1(n7769), .A2(n5302), .ZN(n5653) );
  NAND2_X1 U6446 ( .A1(n9438), .A2(n5311), .ZN(n5310) );
  INV_X1 U6447 ( .A(n9490), .ZN(n5332) );
  NAND2_X1 U6448 ( .A1(n9490), .A2(n5326), .ZN(n5322) );
  NAND2_X1 U6449 ( .A1(n10198), .A2(n9075), .ZN(n10057) );
  OAI211_X1 U6450 ( .C1(n10198), .C2(n5120), .A(n5336), .B(n5335), .ZN(n5338)
         );
  NAND2_X1 U6451 ( .A1(n10198), .A2(n5134), .ZN(n5335) );
  OAI21_X1 U6452 ( .B1(n5120), .B2(n9075), .A(n10197), .ZN(n5337) );
  NAND2_X1 U6453 ( .A1(n5338), .A2(n10062), .ZN(P1_U3212) );
  NAND2_X1 U6454 ( .A1(n9035), .A2(n5350), .ZN(n5349) );
  NAND2_X1 U6455 ( .A1(n5349), .A2(n5353), .ZN(n10143) );
  NAND2_X1 U6456 ( .A1(n7350), .A2(n7122), .ZN(n5360) );
  NAND2_X2 U6457 ( .A1(n5722), .A2(n6127), .ZN(n6563) );
  INV_X2 U6458 ( .A(n5360), .ZN(n9085) );
  INV_X1 U6459 ( .A(n10152), .ZN(n5369) );
  NOR2_X1 U6460 ( .A1(n9014), .A2(n9010), .ZN(n5367) );
  NAND2_X1 U6461 ( .A1(n10149), .A2(n9010), .ZN(n10065) );
  NAND2_X1 U6462 ( .A1(n5369), .A2(n5368), .ZN(n10149) );
  OR2_X1 U6463 ( .A1(n10152), .A2(n9011), .ZN(n5702) );
  NAND2_X1 U6464 ( .A1(n5372), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5757) );
  AND2_X2 U6465 ( .A1(n5375), .A2(n6593), .ZN(n10720) );
  INV_X1 U6466 ( .A(n5376), .ZN(n5375) );
  INV_X1 U6467 ( .A(n5382), .ZN(n10299) );
  INV_X1 U6468 ( .A(n5388), .ZN(n10358) );
  AOI21_X1 U6469 ( .B1(n5115), .B2(n5397), .A(n5402), .ZN(n5396) );
  INV_X1 U6470 ( .A(n6513), .ZN(n5397) );
  NAND2_X1 U6471 ( .A1(n5414), .A2(n8380), .ZN(n5412) );
  INV_X1 U6472 ( .A(n5585), .ZN(n5416) );
  NAND2_X1 U6473 ( .A1(n5419), .A2(n5417), .ZN(n5693) );
  AND2_X2 U6474 ( .A1(n5812), .A2(n5732), .ZN(n5734) );
  NAND2_X1 U6475 ( .A1(n5803), .A2(n5431), .ZN(n5430) );
  NAND2_X1 U6476 ( .A1(n5803), .A2(n5802), .ZN(n5927) );
  NAND3_X1 U6477 ( .A1(n8605), .A2(n8604), .A3(n8610), .ZN(n5440) );
  NAND2_X1 U6478 ( .A1(n6209), .A2(n5445), .ZN(n5443) );
  NAND2_X1 U6479 ( .A1(n6209), .A2(n5699), .ZN(n6211) );
  NAND2_X1 U6480 ( .A1(n6209), .A2(n5448), .ZN(n5444) );
  OAI21_X1 U6481 ( .B1(n7264), .B2(n7263), .A(n7265), .ZN(n7391) );
  NAND2_X1 U6482 ( .A1(n7729), .A2(n5460), .ZN(n5459) );
  NAND2_X1 U6483 ( .A1(n7729), .A2(n7728), .ZN(n7794) );
  NAND2_X1 U6484 ( .A1(n6192), .A2(n6191), .ZN(n6209) );
  NAND2_X1 U6485 ( .A1(n7727), .A2(n7726), .ZN(n7729) );
  NAND2_X1 U6486 ( .A1(n6820), .A2(n8401), .ZN(n7204) );
  NAND2_X1 U6487 ( .A1(n8294), .A2(n8643), .ZN(n5485) );
  NAND2_X1 U6488 ( .A1(n8261), .A2(n8551), .ZN(n11034) );
  NAND2_X1 U6489 ( .A1(n5477), .A2(n8555), .ZN(n10423) );
  NAND2_X1 U6490 ( .A1(n5719), .A2(n5714), .ZN(n5715) );
  INV_X1 U6491 ( .A(n6775), .ZN(n6777) );
  NAND2_X1 U6492 ( .A1(n10174), .A2(n6623), .ZN(n6624) );
  NAND2_X1 U6493 ( .A1(n7017), .A2(n7016), .ZN(n5674) );
  NAND2_X1 U6494 ( .A1(n6590), .A2(n6589), .ZN(n6603) );
  NAND2_X2 U6495 ( .A1(n8059), .A2(n9332), .ZN(n9337) );
  OAI22_X2 U6496 ( .A1(n8615), .A2(n8614), .B1(n8636), .B2(n8613), .ZN(n8621)
         );
  NAND2_X1 U6497 ( .A1(n5464), .A2(n6538), .ZN(n6937) );
  NAND2_X1 U6498 ( .A1(n5463), .A2(n6521), .ZN(n6887) );
  NOR2_X2 U6499 ( .A1(n9432), .A2(n9998), .ZN(n9401) );
  NOR2_X2 U6500 ( .A1(n9474), .A2(n10015), .ZN(n9457) );
  NAND2_X1 U6501 ( .A1(n5470), .A2(n6956), .ZN(n6838) );
  NAND2_X1 U6502 ( .A1(n10423), .A2(n10422), .ZN(n8262) );
  NAND2_X1 U6503 ( .A1(n11034), .A2(n8655), .ZN(n5477) );
  NAND2_X1 U6504 ( .A1(n8268), .A2(n5114), .ZN(n5478) );
  OAI211_X1 U6505 ( .C1(n8268), .C2(n5480), .A(n5478), .B(n5479), .ZN(n8314)
         );
  NAND2_X1 U6506 ( .A1(n5485), .A2(n6817), .ZN(n10730) );
  XNOR2_X2 U6507 ( .A(n10720), .B(n5056), .ZN(n8643) );
  INV_X2 U6508 ( .A(n6577), .ZN(n8133) );
  NAND2_X2 U6509 ( .A1(n6007), .A2(n6006), .ZN(n6577) );
  OAI21_X2 U6510 ( .B1(n5723), .B2(n5570), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5759) );
  NOR2_X1 U6511 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5496) );
  NAND2_X1 U6512 ( .A1(n9463), .A2(n5500), .ZN(n5497) );
  NAND2_X1 U6513 ( .A1(n5497), .A2(n5498), .ZN(n9429) );
  NAND2_X1 U6514 ( .A1(n5503), .A2(n5772), .ZN(n5882) );
  INV_X1 U6515 ( .A(n9112), .ZN(n5503) );
  OAI21_X1 U6516 ( .B1(n9112), .B2(n5505), .A(n5504), .ZN(n5508) );
  NAND3_X1 U6517 ( .A1(n7975), .A2(n9112), .A3(P2_REG0_REG_1__SCAN_IN), .ZN(
        n5504) );
  NAND2_X1 U6518 ( .A1(n5772), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5505) );
  NAND3_X2 U6519 ( .A1(n5841), .A2(n5840), .A3(n5507), .ZN(n6531) );
  NAND2_X1 U6520 ( .A1(n6949), .A2(n8860), .ZN(n6709) );
  NAND2_X1 U6521 ( .A1(n7449), .A2(n5530), .ZN(n7684) );
  NAND2_X2 U6522 ( .A1(n7422), .A2(n8868), .ZN(n7449) );
  NAND2_X1 U6523 ( .A1(n5538), .A2(n5539), .ZN(n8144) );
  NAND2_X1 U6524 ( .A1(n10403), .A2(n8131), .ZN(n5538) );
  INV_X1 U6525 ( .A(n10800), .ZN(n5546) );
  INV_X1 U6526 ( .A(n5543), .ZN(n10840) );
  OR2_X1 U6527 ( .A1(n10474), .A2(n10356), .ZN(n5583) );
  NAND3_X1 U6528 ( .A1(n8921), .A2(n8920), .A3(n8926), .ZN(n5588) );
  NAND2_X1 U6529 ( .A1(n5588), .A2(n5589), .ZN(n9113) );
  NAND2_X1 U6530 ( .A1(n8365), .A2(n5595), .ZN(n7068) );
  NAND2_X1 U6531 ( .A1(n7068), .A2(n7067), .ZN(n7070) );
  NAND2_X1 U6532 ( .A1(n5603), .A2(n6978), .ZN(n7186) );
  NAND2_X1 U6533 ( .A1(n6851), .A2(n6850), .ZN(n6979) );
  NAND2_X1 U6534 ( .A1(n9365), .A2(n5616), .ZN(n9335) );
  NAND3_X1 U6535 ( .A1(n5618), .A2(n5617), .A3(n5788), .ZN(n6025) );
  NAND2_X1 U6536 ( .A1(n5901), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5620) );
  INV_X1 U6537 ( .A(n5622), .ZN(n5621) );
  OAI22_X1 U6538 ( .A1(n5839), .A2(n5837), .B1(n6000), .B2(n5882), .ZN(n5622)
         );
  NAND3_X1 U6539 ( .A1(n6830), .A2(n6829), .A3(n8861), .ZN(n6965) );
  NAND2_X1 U6540 ( .A1(n6830), .A2(n6829), .ZN(n5624) );
  NAND2_X1 U6541 ( .A1(n5624), .A2(n8727), .ZN(n5623) );
  NAND2_X1 U6542 ( .A1(n5625), .A2(n5629), .ZN(n9294) );
  OR2_X1 U6543 ( .A1(n8035), .A2(n5631), .ZN(n5625) );
  AOI21_X1 U6544 ( .B1(n5629), .B2(n5631), .A(n5627), .ZN(n5626) );
  NAND2_X1 U6545 ( .A1(n8035), .A2(n5629), .ZN(n5628) );
  NAND2_X1 U6546 ( .A1(n8035), .A2(n8034), .ZN(n9317) );
  NAND3_X1 U6547 ( .A1(n7089), .A2(n7088), .A3(n5647), .ZN(n5645) );
  NAND2_X1 U6548 ( .A1(n5647), .A2(n5521), .ZN(n5646) );
  NAND2_X1 U6549 ( .A1(n7089), .A2(n7088), .ZN(n7110) );
  NAND2_X1 U6550 ( .A1(n5653), .A2(n5654), .ZN(n9490) );
  NAND2_X1 U6551 ( .A1(n7285), .A2(n5063), .ZN(n5664) );
  NAND2_X1 U6552 ( .A1(n5664), .A2(n5665), .ZN(n7532) );
  INV_X1 U6553 ( .A(n5673), .ZN(n5671) );
  NAND4_X1 U6554 ( .A1(n5708), .A2(n5706), .A3(n5707), .A4(n9936), .ZN(n5673)
         );
  NAND3_X1 U6555 ( .A1(n5674), .A2(n7018), .A3(n7020), .ZN(n7129) );
  OR2_X2 U6556 ( .A1(n10143), .A2(n5678), .ZN(n5676) );
  NAND3_X1 U6557 ( .A1(n10065), .A2(n5684), .A3(n5128), .ZN(n10210) );
  NAND2_X1 U6558 ( .A1(n5144), .A2(n6673), .ZN(n5686) );
  NAND2_X1 U6559 ( .A1(n5687), .A2(n5685), .ZN(n6916) );
  NAND3_X1 U6560 ( .A1(n6908), .A2(n6625), .A3(n6624), .ZN(n5687) );
  NAND2_X1 U6561 ( .A1(n10113), .A2(n5689), .ZN(n9035) );
  INV_X1 U6562 ( .A(n7927), .ZN(n7908) );
  NAND2_X1 U6563 ( .A1(n8314), .A2(n11035), .ZN(n8323) );
  INV_X1 U6564 ( .A(n8617), .ZN(n8674) );
  AOI21_X1 U6565 ( .B1(n8674), .B2(n8673), .A(n8672), .ZN(n8676) );
  OR2_X1 U6566 ( .A1(n7963), .A2(n7962), .ZN(n7969) );
  XNOR2_X1 U6567 ( .A(n7963), .B(n7961), .ZN(n8203) );
  MUX2_X1 U6568 ( .A(n10584), .B(n10533), .S(n6577), .Z(n8297) );
  NAND2_X1 U6569 ( .A1(n6471), .A2(n6470), .ZN(n6203) );
  INV_X1 U6570 ( .A(n5772), .ZN(n7975) );
  NAND2_X1 U6571 ( .A1(n8718), .A2(n8717), .ZN(n6950) );
  INV_X1 U6572 ( .A(n8496), .ZN(n8162) );
  OR2_X1 U6573 ( .A1(n8496), .A2(n6467), .ZN(n6475) );
  OR2_X1 U6574 ( .A1(n8496), .A2(n10738), .ZN(n6608) );
  INV_X2 U6575 ( .A(n6529), .ZN(n6538) );
  NAND2_X1 U6576 ( .A1(n6031), .A2(n6587), .ZN(n6589) );
  AND2_X1 U6577 ( .A1(n5762), .A2(n5467), .ZN(n5692) );
  OR2_X1 U6578 ( .A1(n6560), .A2(n6528), .ZN(n11019) );
  AND3_X1 U6579 ( .A1(n9096), .A2(n9095), .A3(n10197), .ZN(n5694) );
  AND2_X1 U6580 ( .A1(n7325), .A2(n10823), .ZN(n5695) );
  NAND2_X1 U6581 ( .A1(n6134), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5697) );
  AND2_X1 U6582 ( .A1(n6191), .A2(n6143), .ZN(n5698) );
  AND2_X1 U6583 ( .A1(n6210), .A2(n6196), .ZN(n5699) );
  INV_X1 U6584 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6106) );
  CLKBUF_X1 U6585 ( .A(n6076), .Z(n10053) );
  OR2_X1 U6586 ( .A1(n6822), .A2(n10789), .ZN(n11063) );
  AND2_X1 U6587 ( .A1(n6489), .A2(n6373), .ZN(n5700) );
  INV_X1 U6588 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6374) );
  OR2_X1 U6589 ( .A1(n10994), .A2(n8975), .ZN(n5701) );
  INV_X1 U6590 ( .A(n8002), .ZN(n7979) );
  INV_X1 U6591 ( .A(n9367), .ZN(n8024) );
  INV_X1 U6592 ( .A(n8869), .ZN(n7450) );
  INV_X1 U6593 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9936) );
  AND2_X1 U6594 ( .A1(n8696), .A2(n8848), .ZN(n8883) );
  NAND2_X1 U6595 ( .A1(n7979), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8011) );
  OR2_X1 U6596 ( .A1(n9540), .A2(n9360), .ZN(n8034) );
  OR2_X1 U6597 ( .A1(n7630), .A2(n7629), .ZN(n7645) );
  INV_X1 U6598 ( .A(n8868), .ZN(n7417) );
  NAND2_X1 U6599 ( .A1(n6599), .A2(n6598), .ZN(n8286) );
  NAND2_X1 U6600 ( .A1(n10210), .A2(n10212), .ZN(n10207) );
  INV_X1 U6601 ( .A(n8195), .ZN(n6760) );
  INV_X1 U6602 ( .A(n8160), .ZN(n6759) );
  INV_X1 U6603 ( .A(n7742), .ZN(n6755) );
  INV_X1 U6604 ( .A(n10424), .ZN(n10214) );
  INV_X1 U6605 ( .A(n7184), .ZN(n7185) );
  INV_X1 U6606 ( .A(SI_13_), .ZN(n9589) );
  INV_X1 U6607 ( .A(SI_8_), .ZN(n9808) );
  AND2_X1 U6608 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5769) );
  AND2_X1 U6609 ( .A1(n9174), .A2(n5896), .ZN(n5897) );
  OR2_X1 U6610 ( .A1(n7160), .A2(n7240), .ZN(n7162) );
  OR2_X1 U6611 ( .A1(n8011), .A2(n9620), .ZN(n8020) );
  NAND2_X1 U6612 ( .A1(n7937), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7988) );
  OR2_X1 U6613 ( .A1(n7911), .A2(n7910), .ZN(n7938) );
  NAND2_X1 U6614 ( .A1(n7644), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7652) );
  OR2_X1 U6615 ( .A1(n6156), .A2(n6149), .ZN(n7160) );
  OR2_X1 U6616 ( .A1(n6120), .A2(n6119), .ZN(n6146) );
  AND2_X1 U6617 ( .A1(n7541), .A2(n7542), .ZN(n7697) );
  NAND2_X1 U6618 ( .A1(n6761), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U6619 ( .A1(n6760), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8207) );
  OR2_X1 U6620 ( .A1(n7713), .A2(n7712), .ZN(n7742) );
  NAND2_X1 U6621 ( .A1(n6759), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8170) );
  OR2_X1 U6622 ( .A1(n8111), .A2(n8110), .ZN(n8123) );
  OR2_X1 U6623 ( .A1(n7808), .A2(n7807), .ZN(n7858) );
  NAND2_X1 U6624 ( .A1(n6754), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7713) );
  OR2_X1 U6625 ( .A1(n7289), .A2(n7288), .ZN(n7314) );
  NAND2_X1 U6626 ( .A1(n8468), .A2(n8467), .ZN(n8471) );
  INV_X1 U6627 ( .A(n5719), .ZN(n5720) );
  INV_X1 U6628 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5752) );
  INV_X1 U6629 ( .A(SI_17_), .ZN(n9579) );
  INV_X1 U6630 ( .A(SI_14_), .ZN(n9588) );
  NAND2_X1 U6631 ( .A1(n6194), .A2(n6193), .ZN(n6210) );
  INV_X1 U6632 ( .A(n9215), .ZN(n9121) );
  INV_X1 U6633 ( .A(n7157), .ZN(n7158) );
  INV_X1 U6634 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9855) );
  INV_X1 U6635 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7240) );
  OR2_X1 U6636 ( .A1(n9195), .A2(n8940), .ZN(n9198) );
  OR2_X1 U6637 ( .A1(n8020), .A2(n9854), .ZN(n8029) );
  NAND2_X1 U6638 ( .A1(n9112), .A2(n5772), .ZN(n5836) );
  AND2_X1 U6639 ( .A1(n8895), .A2(n8887), .ZN(n5996) );
  INV_X1 U6640 ( .A(n10925), .ZN(n11010) );
  NAND2_X1 U6641 ( .A1(n5740), .A2(n5179), .ZN(n5742) );
  XNOR2_X1 U6642 ( .A(n6670), .B(n6671), .ZN(n6625) );
  NAND2_X1 U6643 ( .A1(n6604), .A2(n8287), .ZN(n10175) );
  NAND2_X1 U6644 ( .A1(n6465), .A2(n8618), .ZN(n8501) );
  AOI21_X1 U6645 ( .B1(n8621), .B2(n8620), .A(n8635), .ZN(n8673) );
  INV_X1 U6646 ( .A(n10229), .ZN(n10295) );
  INV_X1 U6647 ( .A(n10233), .ZN(n7567) );
  NAND2_X1 U6648 ( .A1(n10795), .A2(n6460), .ZN(n10430) );
  AND2_X1 U6649 ( .A1(n10708), .A2(n10359), .ZN(n6461) );
  INV_X1 U6650 ( .A(n11047), .ZN(n10908) );
  OR2_X1 U6651 ( .A1(n8501), .A2(n6007), .ZN(n10779) );
  AND2_X1 U6652 ( .A1(n8412), .A2(n8409), .ZN(n10774) );
  OR2_X1 U6653 ( .A1(n6493), .A2(n6492), .ZN(n6799) );
  INV_X1 U6654 ( .A(n9188), .ZN(n9206) );
  NAND2_X1 U6655 ( .A1(n6519), .A2(n5834), .ZN(n6439) );
  INV_X1 U6656 ( .A(n9198), .ZN(n9128) );
  AND2_X1 U6657 ( .A1(n9208), .A2(n9499), .ZN(n9189) );
  AND2_X1 U6658 ( .A1(n6877), .A2(n5970), .ZN(n9208) );
  AND2_X1 U6659 ( .A1(n5956), .A2(n6877), .ZN(n9167) );
  AND2_X1 U6660 ( .A1(n8073), .A2(n8072), .ZN(n9308) );
  AND4_X1 U6661 ( .A1(n7994), .A2(n7993), .A3(n7992), .A4(n7991), .ZN(n8346)
         );
  AND4_X1 U6662 ( .A1(n6177), .A2(n6176), .A3(n6175), .A4(n6174), .ZN(n8975)
         );
  INV_X1 U6663 ( .A(n10674), .ZN(n9257) );
  OR2_X1 U6664 ( .A1(n6726), .A2(n6725), .ZN(n6988) );
  INV_X1 U6665 ( .A(n9278), .ZN(n10679) );
  AND2_X1 U6666 ( .A1(n7950), .A2(n9104), .ZN(n10660) );
  INV_X1 U6667 ( .A(n9466), .ZN(n9499) );
  INV_X1 U6668 ( .A(n8857), .ZN(n9497) );
  INV_X1 U6669 ( .A(n9495), .ZN(n9427) );
  INV_X1 U6670 ( .A(n9509), .ZN(n9400) );
  OR2_X1 U6671 ( .A1(n10648), .A2(n5941), .ZN(n6875) );
  INV_X1 U6672 ( .A(n11015), .ZN(n10992) );
  OR2_X1 U6673 ( .A1(n6527), .A2(n6526), .ZN(n6560) );
  NAND2_X1 U6674 ( .A1(n10540), .A2(n5940), .ZN(n10542) );
  NAND2_X1 U6675 ( .A1(n5742), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5738) );
  INV_X1 U6676 ( .A(n10221), .ZN(n10203) );
  OR2_X1 U6677 ( .A1(n8492), .A2(n6688), .ZN(n6696) );
  INV_X1 U6678 ( .A(n10618), .ZN(n10696) );
  OR2_X1 U6679 ( .A1(n6357), .A2(n6497), .ZN(n10692) );
  INV_X1 U6680 ( .A(n10692), .ZN(n10605) );
  INV_X1 U6681 ( .A(n11043), .ZN(n10953) );
  AND2_X1 U6682 ( .A1(n10851), .A2(n10911), .ZN(n10769) );
  OR2_X1 U6683 ( .A1(n8613), .A2(n8675), .ZN(n10911) );
  INV_X1 U6684 ( .A(n10769), .ZN(n11050) );
  OAI21_X1 U6685 ( .B1(n6455), .B2(P1_D_REG_0__SCAN_IN), .A(n6444), .ZN(n6800)
         );
  AND2_X1 U6686 ( .A1(n7583), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6123) );
  NOR2_X1 U6687 ( .A1(n10557), .A2(n7497), .ZN(n7498) );
  NOR2_X1 U6688 ( .A1(n10568), .A2(n10567), .ZN(n7514) );
  INV_X1 U6689 ( .A(n10649), .ZN(n5743) );
  NAND2_X1 U6690 ( .A1(n5974), .A2(n5962), .ZN(n9211) );
  INV_X1 U6691 ( .A(n10660), .ZN(n10670) );
  OR2_X1 U6692 ( .A1(n6889), .A2(n8927), .ZN(n9309) );
  INV_X1 U6693 ( .A(n10946), .ZN(n9504) );
  OR2_X1 U6694 ( .A1(n6560), .A2(n6875), .ZN(n11017) );
  NAND2_X1 U6695 ( .A1(n10543), .A2(n10542), .ZN(n10646) );
  XNOR2_X1 U6696 ( .A(n5738), .B(n5180), .ZN(n7761) );
  INV_X1 U6697 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6784) );
  INV_X1 U6698 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6148) );
  AND2_X1 U6699 ( .A1(n6569), .A2(n6568), .ZN(n10221) );
  OR2_X1 U6700 ( .A1(n6462), .A2(n6459), .ZN(n10226) );
  NAND2_X1 U6701 ( .A1(n8244), .A2(n8243), .ZN(n10229) );
  OR2_X1 U6702 ( .A1(n6357), .A2(n6007), .ZN(n10701) );
  OR2_X1 U6703 ( .A1(n10587), .A2(n10583), .ZN(n10693) );
  OR2_X1 U6704 ( .A1(P1_U3083), .A2(n6053), .ZN(n10618) );
  AND2_X1 U6705 ( .A1(n11042), .A2(n11041), .ZN(n11069) );
  NAND2_X1 U6706 ( .A1(n6822), .A2(n10786), .ZN(n10795) );
  NAND2_X1 U6707 ( .A1(n10795), .A2(n10794), .ZN(n11064) );
  INV_X1 U6708 ( .A(n11054), .ZN(n11052) );
  AND2_X1 U6709 ( .A1(n10893), .A2(n10892), .ZN(n10896) );
  INV_X1 U6710 ( .A(n11057), .ZN(n11055) );
  AND2_X2 U6711 ( .A1(n6503), .A2(n6800), .ZN(n11057) );
  NAND2_X1 U6712 ( .A1(n6479), .A2(n6455), .ZN(n10539) );
  AOI21_X1 U6713 ( .B1(n6457), .B2(n9979), .A(n6456), .ZN(n10522) );
  INV_X1 U6714 ( .A(n6478), .ZN(n10359) );
  INV_X1 U6715 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9695) );
  INV_X1 U6716 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6116) );
  NOR2_X1 U6717 ( .A1(n7515), .A2(n7514), .ZN(n10570) );
  NOR2_X1 U6718 ( .A1(n6563), .A2(n5725), .ZN(P1_U4006) );
  NAND2_X1 U6719 ( .A1(n6036), .A2(n5703), .ZN(n6084) );
  INV_X1 U6720 ( .A(n6084), .ZN(n5705) );
  NOR2_X1 U6721 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5708) );
  NOR2_X1 U6722 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5710) );
  NOR2_X1 U6723 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5709) );
  NAND4_X1 U6724 ( .A1(n5710), .A2(n5709), .A3(n9738), .A4(n5752), .ZN(n5712)
         );
  NAND4_X1 U6725 ( .A1(n9729), .A2(n9956), .A3(n9734), .A4(n9954), .ZN(n5711)
         );
  NOR2_X1 U6726 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  NAND2_X1 U6727 ( .A1(n5715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U6728 ( .A1(n5718), .A2(n9743), .ZN(n5716) );
  XNOR2_X1 U6729 ( .A(n5718), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U6730 ( .A1(n5723), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5724) );
  XNOR2_X1 U6731 ( .A(n5724), .B(n5569), .ZN(n7583) );
  INV_X1 U6732 ( .A(n6123), .ZN(n5725) );
  NAND4_X1 U6733 ( .A1(n6792), .A2(n5729), .A3(n5728), .A4(n5727), .ZN(n5731)
         );
  NAND4_X1 U6734 ( .A1(n6117), .A2(n6791), .A3(n6284), .A4(n6484), .ZN(n5730)
         );
  NAND2_X1 U6735 ( .A1(n5143), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U6736 ( .A1(n5761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U6737 ( .A1(n10540), .A2(n10541), .ZN(n5739) );
  NAND2_X1 U6738 ( .A1(n5777), .A2(n5178), .ZN(n5737) );
  OR2_X1 U6739 ( .A1(n5740), .A2(n5179), .ZN(n5741) );
  NAND2_X1 U6740 ( .A1(n5742), .A2(n5741), .ZN(n5981) );
  NOR2_X4 U6741 ( .A1(n5979), .A2(n5743), .ZN(P2_U3966) );
  NAND2_X1 U6742 ( .A1(n5744), .A2(n5745), .ZN(n6490) );
  AND2_X1 U6743 ( .A1(n9738), .A2(n6020), .ZN(n5748) );
  NAND2_X1 U6744 ( .A1(n6844), .A2(n5748), .ZN(n5749) );
  OR2_X1 U6745 ( .A1(n6374), .A2(n9954), .ZN(n5750) );
  NAND2_X1 U6746 ( .A1(n5753), .A2(n5752), .ZN(n5754) );
  NAND2_X1 U6747 ( .A1(n8501), .A2(n6563), .ZN(n5756) );
  NAND2_X1 U6748 ( .A1(n5756), .A2(n7583), .ZN(n6043) );
  NAND2_X2 U6749 ( .A1(n5257), .A2(n5758), .ZN(n6007) );
  XNOR2_X2 U6750 ( .A(n5759), .B(n9967), .ZN(n6006) );
  NAND2_X1 U6751 ( .A1(n6043), .A2(n6577), .ZN(n5760) );
  NAND2_X1 U6752 ( .A1(n5760), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U6753 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U6754 ( .A1(n5765), .A2(n5763), .ZN(n10050) );
  XNOR2_X2 U6755 ( .A(n5764), .B(n10046), .ZN(n9112) );
  NAND2_X1 U6756 ( .A1(n8013), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5776) );
  INV_X1 U6757 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7093) );
  OR2_X1 U6758 ( .A1(n5839), .A2(n7093), .ZN(n5775) );
  NAND2_X1 U6759 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5903) );
  INV_X1 U6760 ( .A(n5903), .ZN(n5767) );
  NAND2_X1 U6761 ( .A1(n5767), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5920) );
  INV_X1 U6762 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9871) );
  INV_X1 U6763 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5768) );
  OAI21_X1 U6764 ( .B1(n5920), .B2(n9871), .A(n5768), .ZN(n5771) );
  INV_X1 U6765 ( .A(n5920), .ZN(n5770) );
  NAND2_X1 U6766 ( .A1(n5770), .A2(n5769), .ZN(n5964) );
  NAND2_X1 U6767 ( .A1(n5771), .A2(n5964), .ZN(n7097) );
  OR2_X1 U6768 ( .A1(n8040), .A2(n7097), .ZN(n5774) );
  INV_X2 U6769 ( .A(n5836), .ZN(n6134) );
  INV_X1 U6770 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6310) );
  OR2_X1 U6771 ( .A1(n8093), .A2(n6310), .ZN(n5773) );
  NAND4_X1 U6772 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n9221)
         );
  NAND2_X1 U6773 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  AND2_X2 U6775 ( .A1(n5784), .A2(n5783), .ZN(n5819) );
  AND2_X1 U6776 ( .A1(n9221), .A2(n8927), .ZN(n5821) );
  NAND2_X1 U6777 ( .A1(n9611), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5786) );
  AND2_X1 U6778 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5788) );
  AND2_X1 U6779 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U6780 ( .A1(n5811), .A2(n5789), .ZN(n5831) );
  INV_X1 U6781 ( .A(SI_1_), .ZN(n9817) );
  XNOR2_X1 U6782 ( .A(n5790), .B(n9817), .ZN(n5857) );
  NAND2_X1 U6783 ( .A1(n5790), .A2(SI_1_), .ZN(n5791) );
  MUX2_X1 U6784 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5804), .Z(n5793) );
  INV_X1 U6785 ( .A(SI_2_), .ZN(n9818) );
  XNOR2_X1 U6786 ( .A(n5793), .B(n9818), .ZN(n5844) );
  NAND2_X1 U6787 ( .A1(n5793), .A2(SI_2_), .ZN(n5794) );
  INV_X1 U6788 ( .A(SI_3_), .ZN(n9602) );
  NAND2_X1 U6789 ( .A1(n5795), .A2(SI_3_), .ZN(n5796) );
  XNOR2_X1 U6790 ( .A(n5797), .B(n9812), .ZN(n5893) );
  NAND2_X1 U6791 ( .A1(n5894), .A2(n5893), .ZN(n5799) );
  NAND2_X1 U6792 ( .A1(n5797), .A2(SI_4_), .ZN(n5798) );
  MUX2_X1 U6793 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7833), .Z(n5801) );
  XNOR2_X1 U6794 ( .A(n5801), .B(n5800), .ZN(n5910) );
  NAND2_X1 U6795 ( .A1(n5801), .A2(SI_5_), .ZN(n5802) );
  MUX2_X1 U6796 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5804), .Z(n5806) );
  XNOR2_X1 U6797 ( .A(n5806), .B(SI_6_), .ZN(n5926) );
  INV_X1 U6798 ( .A(n5926), .ZN(n5805) );
  XNOR2_X1 U6799 ( .A(n6104), .B(SI_7_), .ZN(n6101) );
  XNOR2_X1 U6800 ( .A(n6103), .B(n6101), .ZN(n7119) );
  NAND2_X1 U6801 ( .A1(n7119), .A2(n8693), .ZN(n5818) );
  INV_X1 U6802 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U6803 ( .A1(n5812), .A2(n5813), .ZN(n6120) );
  NAND2_X1 U6804 ( .A1(n6120), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U6805 ( .A1(n5929), .A2(n6118), .ZN(n5814) );
  NAND2_X1 U6806 ( .A1(n5814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5815) );
  XNOR2_X1 U6807 ( .A(n5815), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U6808 ( .A1(n5856), .A2(n6319), .ZN(n5817) );
  NAND2_X1 U6809 ( .A1(n8685), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U6810 ( .A1(n8889), .A2(n8887), .ZN(n6879) );
  NAND2_X1 U6811 ( .A1(n6879), .A2(n8884), .ZN(n5820) );
  MUX2_X2 U6812 ( .A(n7425), .B(n8859), .S(n8887), .Z(n5877) );
  XNOR2_X1 U6813 ( .A(n7111), .B(n5877), .ZN(n7061) );
  NAND2_X1 U6814 ( .A1(n5821), .A2(n7061), .ZN(n7067) );
  INV_X1 U6815 ( .A(n7061), .ZN(n5823) );
  INV_X1 U6816 ( .A(n5821), .ZN(n5822) );
  NAND2_X1 U6817 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  NAND2_X1 U6818 ( .A1(n7067), .A2(n5824), .ZN(n5959) );
  NAND2_X1 U6819 ( .A1(n6133), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5828) );
  INV_X1 U6820 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6890) );
  OR2_X1 U6821 ( .A1(n5882), .A2(n6890), .ZN(n5827) );
  INV_X1 U6822 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5825) );
  OR2_X1 U6823 ( .A1(n5506), .A2(n5825), .ZN(n5826) );
  NAND4_X1 U6824 ( .A1(n5697), .A2(n5828), .A3(n5827), .A4(n5826), .ZN(n9227)
         );
  NAND2_X1 U6825 ( .A1(n8483), .A2(SI_0_), .ZN(n5830) );
  INV_X1 U6826 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U6827 ( .A1(n5830), .A2(n5829), .ZN(n5832) );
  AND2_X1 U6828 ( .A1(n5832), .A2(n5831), .ZN(n10054) );
  NAND2_X1 U6829 ( .A1(n6532), .A2(n8927), .ZN(n6519) );
  INV_X1 U6830 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5835) );
  OR2_X1 U6831 ( .A1(n5836), .A2(n5835), .ZN(n5838) );
  INV_X1 U6832 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5837) );
  INV_X1 U6833 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6000) );
  AND2_X1 U6834 ( .A1(n9225), .A2(n8927), .ZN(n5842) );
  INV_X1 U6835 ( .A(n5842), .ZN(n6063) );
  INV_X1 U6836 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5986) );
  INV_X1 U6837 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U6838 ( .A1(n6134), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5840) );
  AND2_X1 U6839 ( .A1(n6531), .A2(n8927), .ZN(n6059) );
  INV_X1 U6840 ( .A(n6059), .ZN(n6060) );
  NAND2_X1 U6841 ( .A1(n6063), .A2(n6060), .ZN(n5865) );
  OAI21_X1 U6842 ( .B1(n6439), .B2(n6059), .A(n5842), .ZN(n5854) );
  INV_X1 U6843 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5843) );
  OR2_X1 U6844 ( .A1(n5858), .A2(n5843), .ZN(n5853) );
  XNOR2_X1 U6845 ( .A(n5845), .B(n5844), .ZN(n6613) );
  OR2_X1 U6846 ( .A1(n5928), .A2(n6613), .ZN(n5852) );
  NOR2_X1 U6847 ( .A1(n5846), .A2(n6287), .ZN(n5847) );
  NAND2_X1 U6848 ( .A1(n5847), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5850) );
  INV_X1 U6849 ( .A(n5847), .ZN(n5849) );
  INV_X1 U6850 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U6851 ( .A1(n5849), .A2(n5848), .ZN(n5872) );
  AND2_X1 U6852 ( .A1(n5850), .A2(n5872), .ZN(n6296) );
  NAND2_X1 U6853 ( .A1(n5856), .A2(n6296), .ZN(n5851) );
  XNOR2_X1 U6854 ( .A(n6659), .B(n8941), .ZN(n6062) );
  NAND2_X1 U6855 ( .A1(n5854), .A2(n6062), .ZN(n5864) );
  NAND2_X1 U6856 ( .A1(n6439), .A2(n6059), .ZN(n5862) );
  NAND2_X1 U6857 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n10662), .ZN(n5855) );
  NAND2_X1 U6858 ( .A1(n5856), .A2(n10661), .ZN(n5861) );
  OR2_X1 U6859 ( .A1(n5858), .A2(n5424), .ZN(n5859) );
  XNOR2_X1 U6860 ( .A(n6538), .B(n8941), .ZN(n6061) );
  OAI211_X1 U6861 ( .C1(n6062), .C2(n6063), .A(n5862), .B(n6061), .ZN(n5863)
         );
  OAI211_X1 U6862 ( .C1(n6439), .C2(n5865), .A(n5864), .B(n5863), .ZN(n6513)
         );
  NAND2_X1 U6863 ( .A1(n6133), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5870) );
  INV_X1 U6864 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6297) );
  OR2_X1 U6865 ( .A1(n8093), .A2(n6297), .ZN(n5869) );
  INV_X1 U6866 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5866) );
  OR2_X1 U6867 ( .A1(n5506), .A2(n5866), .ZN(n5868) );
  OR2_X1 U6868 ( .A1(n5882), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5867) );
  AND2_X1 U6869 ( .A1(n9175), .A2(n8927), .ZN(n5878) );
  OR2_X1 U6870 ( .A1(n5928), .A2(n6581), .ZN(n5876) );
  INV_X1 U6871 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6075) );
  OR2_X1 U6872 ( .A1(n5858), .A2(n6075), .ZN(n5875) );
  NAND2_X1 U6873 ( .A1(n5872), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5873) );
  XNOR2_X1 U6874 ( .A(n5873), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U6875 ( .A1(n5856), .A2(n6298), .ZN(n5874) );
  XNOR2_X1 U6876 ( .A(n10754), .B(n5877), .ZN(n5879) );
  NAND2_X1 U6877 ( .A1(n5878), .A2(n5879), .ZN(n5896) );
  INV_X1 U6878 ( .A(n5878), .ZN(n5880) );
  INV_X1 U6879 ( .A(n5879), .ZN(n9173) );
  NAND2_X1 U6880 ( .A1(n5880), .A2(n9173), .ZN(n5881) );
  NAND2_X1 U6881 ( .A1(n5896), .A2(n5881), .ZN(n6514) );
  NAND2_X1 U6882 ( .A1(n6133), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5887) );
  INV_X1 U6883 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6299) );
  OR2_X1 U6884 ( .A1(n8093), .A2(n6299), .ZN(n5886) );
  OAI21_X1 U6885 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n5903), .ZN(n9169) );
  OR2_X1 U6886 ( .A1(n5882), .A2(n9169), .ZN(n5885) );
  INV_X1 U6887 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5883) );
  OR2_X1 U6888 ( .A1(n5506), .A2(n5883), .ZN(n5884) );
  NAND2_X1 U6889 ( .A1(n9224), .A2(n8927), .ZN(n5899) );
  NOR2_X1 U6890 ( .A1(n5888), .A2(n6287), .ZN(n5889) );
  MUX2_X1 U6891 ( .A(n6287), .B(n5889), .S(P2_IR_REG_4__SCAN_IN), .Z(n5890) );
  INV_X1 U6892 ( .A(n5890), .ZN(n5892) );
  INV_X1 U6893 ( .A(n5812), .ZN(n5891) );
  NAND2_X1 U6894 ( .A1(n5892), .A2(n5891), .ZN(n6437) );
  INV_X1 U6895 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6078) );
  OR2_X1 U6896 ( .A1(n5858), .A2(n6078), .ZN(n5895) );
  XNOR2_X1 U6897 ( .A(n9170), .B(n8941), .ZN(n8961) );
  XNOR2_X1 U6898 ( .A(n5899), .B(n8961), .ZN(n9174) );
  INV_X1 U6899 ( .A(n8961), .ZN(n5898) );
  NAND2_X1 U6900 ( .A1(n5899), .A2(n5898), .ZN(n5900) );
  NAND2_X1 U6901 ( .A1(n8013), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5909) );
  INV_X1 U6902 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5902) );
  OR2_X1 U6903 ( .A1(n5839), .A2(n5902), .ZN(n5908) );
  INV_X1 U6904 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U6905 ( .A1(n5903), .A2(n9853), .ZN(n5904) );
  NAND2_X1 U6906 ( .A1(n5920), .A2(n5904), .ZN(n8960) );
  OR2_X1 U6907 ( .A1(n8040), .A2(n8960), .ZN(n5907) );
  INV_X1 U6908 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5905) );
  OR2_X1 U6909 ( .A1(n8093), .A2(n5905), .ZN(n5906) );
  NAND4_X1 U6910 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(n9223)
         );
  NAND2_X1 U6911 ( .A1(n9223), .A2(n8927), .ZN(n5917) );
  XNOR2_X1 U6912 ( .A(n5911), .B(n5910), .ZN(n6912) );
  OR2_X1 U6913 ( .A1(n5928), .A2(n6912), .ZN(n5915) );
  INV_X1 U6914 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6080) );
  OR2_X1 U6915 ( .A1(n5858), .A2(n6080), .ZN(n5914) );
  OR2_X1 U6916 ( .A1(n5812), .A2(n6287), .ZN(n5912) );
  XNOR2_X1 U6917 ( .A(n5912), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U6918 ( .A1(n5856), .A2(n6322), .ZN(n5913) );
  XNOR2_X1 U6919 ( .A(n6881), .B(n5877), .ZN(n8357) );
  INV_X1 U6920 ( .A(n8357), .ZN(n5916) );
  NAND2_X1 U6921 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  NAND2_X1 U6922 ( .A1(n8967), .A2(n5918), .ZN(n5933) );
  NAND2_X1 U6923 ( .A1(n8013), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5925) );
  INV_X1 U6924 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5919) );
  OR2_X1 U6925 ( .A1(n5839), .A2(n5919), .ZN(n5924) );
  XNOR2_X1 U6926 ( .A(n5920), .B(n9871), .ZN(n7045) );
  OR2_X1 U6927 ( .A1(n8040), .A2(n7045), .ZN(n5923) );
  INV_X1 U6928 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5921) );
  OR2_X1 U6929 ( .A1(n8093), .A2(n5921), .ZN(n5922) );
  OR2_X1 U6930 ( .A1(n7085), .A2(n8940), .ZN(n5936) );
  XNOR2_X1 U6931 ( .A(n5927), .B(n5926), .ZN(n7006) );
  INV_X1 U6932 ( .A(n7006), .ZN(n6083) );
  INV_X1 U6933 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6081) );
  OR2_X1 U6934 ( .A1(n5858), .A2(n6081), .ZN(n5931) );
  XNOR2_X1 U6935 ( .A(n5929), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U6936 ( .A1(n5856), .A2(n6320), .ZN(n5930) );
  XNOR2_X1 U6937 ( .A(n7086), .B(n5877), .ZN(n5934) );
  XNOR2_X1 U6938 ( .A(n5936), .B(n5934), .ZN(n8358) );
  NAND2_X1 U6939 ( .A1(n5933), .A2(n8358), .ZN(n8365) );
  INV_X1 U6940 ( .A(n5934), .ZN(n5935) );
  NAND2_X1 U6941 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  INV_X1 U6942 ( .A(n10540), .ZN(n7925) );
  AND2_X1 U6943 ( .A1(n7925), .A2(n7761), .ZN(n10648) );
  INV_X1 U6944 ( .A(n7761), .ZN(n5938) );
  INV_X1 U6945 ( .A(P2_B_REG_SCAN_IN), .ZN(n9280) );
  AOI22_X1 U6946 ( .A1(P2_B_REG_SCAN_IN), .A2(n7761), .B1(n5938), .B2(n9280), 
        .ZN(n5939) );
  OR2_X1 U6947 ( .A1(n10541), .A2(n5939), .ZN(n5940) );
  NOR2_X1 U6948 ( .A1(n10542), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5941) );
  OR2_X1 U6949 ( .A1(n10713), .A2(n8889), .ZN(n6880) );
  OR2_X1 U6950 ( .A1(n10713), .A2(n8884), .ZN(n5942) );
  OR2_X1 U6951 ( .A1(n10925), .A2(n5996), .ZN(n5943) );
  NOR2_X1 U6952 ( .A1(n6875), .A2(n5943), .ZN(n5956) );
  NOR4_X1 U6953 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5952) );
  NOR4_X1 U6954 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5951) );
  OR4_X1 U6955 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5949) );
  NOR4_X1 U6956 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5947) );
  NOR4_X1 U6957 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5946) );
  NOR4_X1 U6958 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5945) );
  NOR4_X1 U6959 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5944) );
  NAND4_X1 U6960 ( .A1(n5947), .A2(n5946), .A3(n5945), .A4(n5944), .ZN(n5948)
         );
  NOR4_X1 U6961 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n5949), .A4(n5948), .ZN(n5950) );
  AND3_X1 U6962 ( .A1(n5952), .A2(n5951), .A3(n5950), .ZN(n5953) );
  NOR2_X1 U6963 ( .A1(n5953), .A2(n10542), .ZN(n6527) );
  OR2_X1 U6964 ( .A1(n10542), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5955) );
  OR2_X1 U6965 ( .A1(n10540), .A2(n10541), .ZN(n5954) );
  NAND2_X1 U6966 ( .A1(n5955), .A2(n5954), .ZN(n6525) );
  NOR2_X1 U6967 ( .A1(n6527), .A2(n6525), .ZN(n5960) );
  INV_X1 U6968 ( .A(n5959), .ZN(n5957) );
  INV_X1 U6969 ( .A(n7068), .ZN(n7066) );
  AOI211_X1 U6970 ( .C1(n5959), .C2(n5958), .A(n9195), .B(n7066), .ZN(n5978)
         );
  INV_X1 U6971 ( .A(n5960), .ZN(n5961) );
  NAND3_X1 U6972 ( .A1(n8889), .A2(n5819), .A3(n8704), .ZN(n6652) );
  OAI21_X1 U6973 ( .B1(n6875), .B2(n5961), .A(n6869), .ZN(n5974) );
  AND2_X1 U6974 ( .A1(n10543), .A2(n10925), .ZN(n5962) );
  NOR2_X1 U6975 ( .A1(n7111), .A2(n9211), .ZN(n5977) );
  NAND2_X1 U6976 ( .A1(n8013), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5969) );
  INV_X1 U6977 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6330) );
  OR2_X1 U6978 ( .A1(n5839), .A2(n6330), .ZN(n5968) );
  INV_X1 U6979 ( .A(n5964), .ZN(n5963) );
  INV_X1 U6980 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9841) );
  NAND2_X1 U6981 ( .A1(n5964), .A2(n9841), .ZN(n5965) );
  NAND2_X1 U6982 ( .A1(n6156), .A2(n5965), .ZN(n7104) );
  OR2_X1 U6983 ( .A1(n8040), .A2(n7104), .ZN(n5967) );
  INV_X1 U6984 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6307) );
  OR2_X1 U6985 ( .A1(n8093), .A2(n6307), .ZN(n5966) );
  NAND4_X1 U6986 ( .A1(n5969), .A2(n5968), .A3(n5967), .A4(n5966), .ZN(n9220)
         );
  INV_X1 U6987 ( .A(n9220), .ZN(n7171) );
  NOR2_X1 U6988 ( .A1(n6875), .A2(n8893), .ZN(n5970) );
  NAND2_X1 U6989 ( .A1(n9208), .A2(n9501), .ZN(n9161) );
  OAI22_X1 U6990 ( .A1(n7171), .A2(n9161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5768), .ZN(n5976) );
  INV_X1 U6991 ( .A(n9104), .ZN(n5972) );
  INV_X1 U6992 ( .A(n9189), .ZN(n9159) );
  NAND2_X1 U6993 ( .A1(n8893), .A2(n5996), .ZN(n6874) );
  AND3_X1 U6994 ( .A1(n5979), .A2(n5981), .A3(n6874), .ZN(n5973) );
  NAND2_X1 U6995 ( .A1(n5974), .A2(n5973), .ZN(n6069) );
  OAI22_X1 U6996 ( .A1(n7085), .A2(n9159), .B1(n9206), .B2(n7097), .ZN(n5975)
         );
  OR4_X1 U6997 ( .A1(n5978), .A2(n5977), .A3(n5976), .A4(n5975), .ZN(P2_U3215)
         );
  INV_X1 U6998 ( .A(n5979), .ZN(n5980) );
  NAND2_X1 U6999 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5980), .ZN(n5984) );
  OR2_X1 U7000 ( .A1(n5981), .A2(P2_U3152), .ZN(n8898) );
  INV_X1 U7001 ( .A(n5996), .ZN(n5982) );
  NAND2_X1 U7002 ( .A1(n10543), .A2(n5982), .ZN(n5983) );
  NAND3_X1 U7003 ( .A1(n5984), .A2(n8898), .A3(n5983), .ZN(n5993) );
  NAND2_X1 U7004 ( .A1(n5985), .A2(n9226), .ZN(n7950) );
  INV_X1 U7005 ( .A(n6296), .ZN(n6074) );
  NOR2_X1 U7006 ( .A1(n10670), .A2(n6074), .ZN(n6005) );
  MUX2_X1 U7007 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n5986), .S(n10661), .Z(n10664) );
  NAND3_X1 U7008 ( .A1(n10662), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n10664), .ZN(
        n10663) );
  INV_X1 U7009 ( .A(n10663), .ZN(n5987) );
  AOI21_X1 U7010 ( .B1(n10661), .B2(P2_REG2_REG_1__SCAN_IN), .A(n5987), .ZN(
        n5991) );
  MUX2_X1 U7011 ( .A(n5837), .B(P2_REG2_REG_2__SCAN_IN), .S(n6296), .Z(n5990)
         );
  NOR2_X1 U7012 ( .A1(n5990), .A2(n5991), .ZN(n6292) );
  NOR2_X1 U7013 ( .A1(n9104), .A2(n5055), .ZN(n5989) );
  NAND2_X1 U7014 ( .A1(n7950), .A2(n5989), .ZN(n9278) );
  AOI211_X1 U7015 ( .C1(n5991), .C2(n5990), .A(n6292), .B(n9278), .ZN(n6004)
         );
  NAND2_X1 U7016 ( .A1(n10662), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10650) );
  INV_X1 U7017 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5992) );
  MUX2_X1 U7018 ( .A(n5992), .B(P2_REG1_REG_1__SCAN_IN), .S(n10661), .Z(n10651) );
  NOR2_X1 U7019 ( .A1(n10650), .A2(n10651), .ZN(n10652) );
  AOI21_X1 U7020 ( .B1(n10661), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10652), .ZN(
        n5995) );
  XNOR2_X1 U7021 ( .A(n6296), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n5994) );
  NOR2_X1 U7022 ( .A1(n5994), .A2(n5995), .ZN(n6295) );
  NAND2_X1 U7023 ( .A1(n5993), .A2(n5146), .ZN(n10658) );
  AOI211_X1 U7024 ( .C1(n5995), .C2(n5994), .A(n6295), .B(n10658), .ZN(n6003)
         );
  INV_X1 U7025 ( .A(n10543), .ZN(n8894) );
  NAND2_X1 U7026 ( .A1(n8894), .A2(n8898), .ZN(n5999) );
  NAND2_X1 U7027 ( .A1(n10543), .A2(n5996), .ZN(n5997) );
  AND2_X1 U7028 ( .A1(n5999), .A2(n5998), .ZN(n10674) );
  INV_X1 U7029 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6001) );
  OAI22_X1 U7030 ( .A1(n9257), .A2(n6001), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6000), .ZN(n6002) );
  OR4_X1 U7031 ( .A1(n6005), .A2(n6004), .A3(n6003), .A4(n6002), .ZN(P2_U3247)
         );
  INV_X1 U7032 ( .A(n6006), .ZN(n10583) );
  INV_X1 U7033 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6008) );
  AOI21_X1 U7034 ( .B1(n10583), .B2(n6008), .A(n6007), .ZN(n10582) );
  AND2_X1 U7035 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n10642) );
  NAND2_X4 U7036 ( .A1(n10530), .A2(n6470), .ZN(n8496) );
  INV_X1 U7037 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6010) );
  INV_X1 U7038 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7039 ( .A1(n6571), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7040 ( .A1(n10530), .A2(n6013), .ZN(n6469) );
  INV_X1 U7041 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6014) );
  OR2_X1 U7042 ( .A1(n6469), .A2(n6014), .ZN(n6015) );
  NAND2_X1 U7043 ( .A1(n6844), .A2(n6020), .ZN(n6021) );
  NAND2_X1 U7044 ( .A1(n6021), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6022) );
  NAND2_X2 U7045 ( .A1(n8618), .A2(n10708), .ZN(n6584) );
  INV_X1 U7046 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10584) );
  INV_X1 U7047 ( .A(SI_0_), .ZN(n6024) );
  INV_X1 U7048 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6023) );
  OAI21_X1 U7049 ( .B1(n8483), .B2(n6024), .A(n6023), .ZN(n6026) );
  NAND2_X1 U7050 ( .A1(n6026), .A2(n6025), .ZN(n10533) );
  INV_X1 U7051 ( .A(n6563), .ZN(n6028) );
  AOI22_X1 U7052 ( .A1(n5363), .A2(n7122), .B1(n6028), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7053 ( .A1(n6030), .A2(n6029), .ZN(n6587) );
  OAI21_X1 U7054 ( .B1(n6031), .B2(n6587), .A(n6589), .ZN(n6464) );
  INV_X1 U7055 ( .A(n6464), .ZN(n6032) );
  MUX2_X1 U7056 ( .A(n10642), .B(n6032), .S(n6006), .Z(n6033) );
  INV_X1 U7057 ( .A(n6007), .ZN(n6497) );
  NAND2_X1 U7058 ( .A1(n6033), .A2(n6497), .ZN(n6034) );
  OAI211_X1 U7059 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10582), .A(n6034), .B(
        P1_U4006), .ZN(n10703) );
  INV_X1 U7060 ( .A(n10703), .ZN(n6058) );
  AND2_X1 U7061 ( .A1(n6577), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7062 ( .A1(n6043), .A2(n6035), .ZN(n10587) );
  INV_X1 U7063 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10738) );
  OR2_X1 U7064 ( .A1(n6036), .A2(n6374), .ZN(n6091) );
  XNOR2_X1 U7065 ( .A(n6091), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6610) );
  MUX2_X1 U7066 ( .A(n10738), .B(P1_REG1_REG_2__SCAN_IN), .S(n6610), .Z(n6038)
         );
  INV_X1 U7067 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7068 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6037) );
  XNOR2_X1 U7069 ( .A(n6037), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6591) );
  MUX2_X1 U7070 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6467), .S(n6591), .Z(n10637)
         );
  AND2_X1 U7071 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n10638) );
  NAND2_X1 U7072 ( .A1(n10637), .A2(n10638), .ZN(n10635) );
  NAND2_X1 U7073 ( .A1(n6591), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6039) );
  NAND3_X1 U7074 ( .A1(n6038), .A2(n10635), .A3(n6039), .ZN(n6042) );
  MUX2_X1 U7075 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10738), .S(n6610), .Z(n6041)
         );
  NAND2_X1 U7076 ( .A1(n10635), .A2(n6039), .ZN(n6040) );
  NAND2_X1 U7077 ( .A1(n6041), .A2(n6040), .ZN(n6229) );
  NAND2_X1 U7078 ( .A1(n6042), .A2(n6229), .ZN(n6051) );
  NOR2_X1 U7079 ( .A1(n6006), .A2(P1_U3084), .ZN(n7838) );
  NAND2_X1 U7080 ( .A1(n6043), .A2(n7838), .ZN(n6357) );
  INV_X1 U7081 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6222) );
  MUX2_X1 U7082 ( .A(n6222), .B(P1_REG2_REG_2__SCAN_IN), .S(n6610), .Z(n6045)
         );
  INV_X1 U7083 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6044) );
  MUX2_X1 U7084 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6044), .S(n6591), .Z(n10641)
         );
  NAND2_X1 U7085 ( .A1(n10641), .A2(n10642), .ZN(n10639) );
  NAND2_X1 U7086 ( .A1(n6591), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6046) );
  NAND3_X1 U7087 ( .A1(n6045), .A2(n10639), .A3(n6046), .ZN(n6049) );
  MUX2_X1 U7088 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6222), .S(n6610), .Z(n6048)
         );
  NAND2_X1 U7089 ( .A1(n10639), .A2(n6046), .ZN(n6047) );
  NAND2_X1 U7090 ( .A1(n6048), .A2(n6047), .ZN(n6221) );
  NAND2_X1 U7091 ( .A1(n6049), .A2(n6221), .ZN(n6050) );
  OAI22_X1 U7092 ( .A1(n10693), .A2(n6051), .B1(n10701), .B2(n6050), .ZN(n6057) );
  INV_X1 U7093 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6055) );
  INV_X1 U7094 ( .A(n7583), .ZN(n6052) );
  NOR2_X1 U7095 ( .A1(n6563), .A2(n6052), .ZN(n6053) );
  AOI22_X1 U7096 ( .A1(n10605), .A2(n6610), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n6054) );
  OAI21_X1 U7097 ( .B1(n6055), .B2(n10618), .A(n6054), .ZN(n6056) );
  OR3_X1 U7098 ( .A1(n6058), .A2(n6057), .A3(n6056), .ZN(P1_U3243) );
  INV_X1 U7099 ( .A(n6061), .ZN(n6065) );
  XNOR2_X1 U7100 ( .A(n6065), .B(n6059), .ZN(n6440) );
  NOR2_X1 U7101 ( .A1(n6440), .A2(n6439), .ZN(n6438) );
  AOI21_X1 U7102 ( .B1(n6061), .B2(n6060), .A(n6438), .ZN(n6064) );
  XNOR2_X1 U7103 ( .A(n6063), .B(n6062), .ZN(n6066) );
  NOR3_X1 U7104 ( .A1(n6064), .A2(n6066), .A3(n9195), .ZN(n6073) );
  INV_X2 U7105 ( .A(n9167), .ZN(n9195) );
  AOI22_X1 U7106 ( .A1(n6065), .A2(n9167), .B1(n9128), .B2(n6531), .ZN(n6068)
         );
  INV_X1 U7107 ( .A(n6066), .ZN(n6067) );
  NOR3_X1 U7108 ( .A1(n6438), .A2(n6068), .A3(n6067), .ZN(n6072) );
  INV_X1 U7109 ( .A(n9175), .ZN(n6713) );
  OAI22_X1 U7110 ( .A1(n6713), .A2(n9161), .B1(n6659), .B2(n9211), .ZN(n6071)
         );
  NOR2_X1 U7111 ( .A1(n6069), .A2(P2_U3152), .ZN(n6524) );
  OAI22_X1 U7112 ( .A1(n6530), .A2(n9159), .B1(n6524), .B2(n6000), .ZN(n6070)
         );
  OR4_X1 U7113 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(P2_U3239)
         );
  NAND2_X1 U7114 ( .A1(n8483), .A2(P2_U3152), .ZN(n6076) );
  NAND2_X1 U7115 ( .A1(n5153), .A2(P2_U3152), .ZN(n9110) );
  OAI222_X1 U7116 ( .A1(P2_U3152), .A2(n6074), .B1(n10053), .B2(n6613), .C1(
        n9110), .C2(n5843), .ZN(P2_U3356) );
  INV_X1 U7117 ( .A(n9110), .ZN(n7799) );
  INV_X1 U7118 ( .A(n7799), .ZN(n10047) );
  INV_X1 U7119 ( .A(n6298), .ZN(n6422) );
  OAI222_X1 U7120 ( .A1(n10047), .A2(n6075), .B1(n10053), .B2(n6581), .C1(
        P2_U3152), .C2(n6422), .ZN(P2_U3355) );
  INV_X1 U7121 ( .A(n10661), .ZN(n6077) );
  OAI222_X1 U7122 ( .A1(n10047), .A2(n5424), .B1(n10053), .B2(n6594), .C1(
        P2_U3152), .C2(n6077), .ZN(P2_U3357) );
  OAI222_X1 U7123 ( .A1(n10047), .A2(n6078), .B1(n10053), .B2(n6678), .C1(
        P2_U3152), .C2(n6437), .ZN(P2_U3354) );
  INV_X1 U7124 ( .A(n6322), .ZN(n6079) );
  OAI222_X1 U7125 ( .A1(n10047), .A2(n6080), .B1(n10053), .B2(n6912), .C1(
        P2_U3152), .C2(n6079), .ZN(P2_U3353) );
  INV_X1 U7126 ( .A(n6320), .ZN(n6398) );
  OAI222_X1 U7127 ( .A1(n10047), .A2(n6081), .B1(n10053), .B2(n6083), .C1(
        P2_U3152), .C2(n6398), .ZN(P2_U3352) );
  INV_X1 U7128 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7010) );
  NOR2_X1 U7129 ( .A1(n6082), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6114) );
  OR2_X1 U7130 ( .A1(n6114), .A2(n6374), .ZN(n6095) );
  XNOR2_X1 U7131 ( .A(n6095), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7007) );
  INV_X1 U7132 ( .A(n7007), .ZN(n10593) );
  OAI222_X1 U7133 ( .A1(n10528), .A2(n7010), .B1(n10532), .B2(n6083), .C1(
        P1_U3084), .C2(n10593), .ZN(P1_U3347) );
  INV_X1 U7134 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7135 ( .A1(n6084), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6085) );
  XNOR2_X1 U7136 ( .A(n6085), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6675) );
  INV_X1 U7137 ( .A(n6675), .ZN(n10691) );
  OAI222_X1 U7138 ( .A1(n10528), .A2(n6086), .B1(n10532), .B2(n6678), .C1(
        P1_U3084), .C2(n10691), .ZN(P1_U3349) );
  INV_X1 U7139 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6087) );
  INV_X1 U7140 ( .A(n6610), .ZN(n6230) );
  OAI222_X1 U7141 ( .A1(n10528), .A2(n6087), .B1(n10532), .B2(n6613), .C1(
        P1_U3084), .C2(n6230), .ZN(P1_U3351) );
  INV_X1 U7142 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6592) );
  OAI222_X1 U7143 ( .A1(n10528), .A2(n6592), .B1(n10532), .B2(n6594), .C1(
        P1_U3084), .C2(n5491), .ZN(P1_U3352) );
  INV_X1 U7144 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7145 ( .A1(n6082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6088) );
  XNOR2_X1 U7146 ( .A(n6088), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6909) );
  INV_X1 U7147 ( .A(n6909), .ZN(n6224) );
  OAI222_X1 U7148 ( .A1(n10528), .A2(n6089), .B1(n10532), .B2(n6912), .C1(
        P1_U3084), .C2(n6224), .ZN(P1_U3348) );
  INV_X1 U7149 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7150 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  NAND2_X1 U7151 ( .A1(n6092), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6093) );
  XNOR2_X1 U7152 ( .A(n6093), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6578) );
  INV_X1 U7153 ( .A(n6578), .ZN(n10622) );
  INV_X1 U7154 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6132) );
  OAI222_X1 U7155 ( .A1(n10622), .A2(P1_U3084), .B1(n10532), .B2(n6581), .C1(
        n10528), .C2(n6132), .ZN(P1_U3350) );
  INV_X1 U7156 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6098) );
  INV_X1 U7157 ( .A(n7119), .ZN(n6099) );
  INV_X1 U7158 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7159 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7160 ( .A1(n6096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6097) );
  XNOR2_X1 U7161 ( .A(n6097), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7118) );
  INV_X1 U7162 ( .A(n7118), .ZN(n6248) );
  OAI222_X1 U7163 ( .A1(n10528), .A2(n6098), .B1(n10532), .B2(n6099), .C1(
        P1_U3084), .C2(n6248), .ZN(P1_U3346) );
  INV_X1 U7164 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6100) );
  INV_X1 U7165 ( .A(n6319), .ZN(n6387) );
  OAI222_X1 U7166 ( .A1(n10047), .A2(n6100), .B1(n10053), .B2(n6099), .C1(
        P2_U3152), .C2(n6387), .ZN(P2_U3351) );
  INV_X1 U7167 ( .A(n6101), .ZN(n6102) );
  NAND2_X1 U7168 ( .A1(n6104), .A2(SI_7_), .ZN(n6105) );
  MUX2_X1 U7169 ( .A(n6106), .B(n6116), .S(n5804), .Z(n6107) );
  INV_X1 U7170 ( .A(n6107), .ZN(n6108) );
  NAND2_X1 U7171 ( .A1(n6108), .A2(SI_8_), .ZN(n6109) );
  NAND2_X1 U7172 ( .A1(n6139), .A2(n6109), .ZN(n6110) );
  NAND2_X1 U7173 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NAND2_X1 U7174 ( .A1(n6140), .A2(n6112), .ZN(n7270) );
  INV_X1 U7175 ( .A(n7270), .ZN(n6122) );
  NOR2_X1 U7176 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6113) );
  NAND2_X1 U7177 ( .A1(n6114), .A2(n6113), .ZN(n6144) );
  NAND2_X1 U7178 ( .A1(n6144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6115) );
  XNOR2_X1 U7179 ( .A(n6115), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7271) );
  INV_X1 U7180 ( .A(n7271), .ZN(n6268) );
  OAI222_X1 U7181 ( .A1(n10528), .A2(n6116), .B1(n10532), .B2(n6122), .C1(
        P1_U3084), .C2(n6268), .ZN(P1_U3345) );
  NAND2_X1 U7182 ( .A1(n6118), .A2(n6117), .ZN(n6119) );
  NAND2_X1 U7183 ( .A1(n6146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6121) );
  XNOR2_X1 U7184 ( .A(n6121), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7053) );
  INV_X1 U7185 ( .A(n7053), .ZN(n6410) );
  OAI222_X1 U7186 ( .A1(P2_U3152), .A2(n6410), .B1(n10053), .B2(n6122), .C1(
        n9110), .C2(n6106), .ZN(P2_U3350) );
  NOR2_X1 U7187 ( .A1(n10674), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7188 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6130) );
  INV_X1 U7189 ( .A(n6124), .ZN(n7825) );
  NAND2_X1 U7190 ( .A1(n7825), .A2(P1_B_REG_SCAN_IN), .ZN(n6125) );
  MUX2_X1 U7191 ( .A(n6125), .B(P1_B_REG_SCAN_IN), .S(n6128), .Z(n6126) );
  NAND2_X1 U7192 ( .A1(n6126), .A2(n6127), .ZN(n6455) );
  INV_X1 U7193 ( .A(n10539), .ZN(n10538) );
  INV_X1 U7194 ( .A(n6127), .ZN(n7844) );
  INV_X1 U7195 ( .A(n6128), .ZN(n7731) );
  NAND2_X1 U7196 ( .A1(n7844), .A2(n7731), .ZN(n6444) );
  OAI21_X1 U7197 ( .B1(n10538), .B2(P1_D_REG_0__SCAN_IN), .A(n6444), .ZN(n6129) );
  OAI21_X1 U7198 ( .B1(n6479), .B2(n6130), .A(n6129), .ZN(P1_U3440) );
  NAND2_X1 U7199 ( .A1(n9175), .A2(P2_U3966), .ZN(n6131) );
  OAI21_X1 U7200 ( .B1(P2_U3966), .B2(n6132), .A(n6131), .ZN(P2_U3555) );
  NAND2_X1 U7201 ( .A1(n8013), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7202 ( .A1(n6133), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7203 ( .A1(n6134), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6135) );
  AND3_X1 U7204 ( .A1(n6137), .A2(n6136), .A3(n6135), .ZN(n9306) );
  NAND2_X1 U7205 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n9226), .ZN(n6138) );
  OAI21_X1 U7206 ( .B1(n9306), .B2(n9226), .A(n6138), .ZN(P2_U3582) );
  MUX2_X1 U7207 ( .A(n6148), .B(n6162), .S(n5153), .Z(n6141) );
  NAND2_X1 U7208 ( .A1(n6141), .A2(n9804), .ZN(n6191) );
  INV_X1 U7209 ( .A(n6141), .ZN(n6142) );
  NAND2_X1 U7210 ( .A1(n6142), .A2(SI_9_), .ZN(n6143) );
  XNOR2_X1 U7211 ( .A(n6190), .B(n5698), .ZN(n7306) );
  INV_X1 U7212 ( .A(n7306), .ZN(n6147) );
  NAND2_X1 U7213 ( .A1(n6206), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6145) );
  XNOR2_X1 U7214 ( .A(n6145), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10604) );
  INV_X1 U7215 ( .A(n10604), .ZN(n6338) );
  OAI222_X1 U7216 ( .A1(n10532), .A2(n6147), .B1(n6338), .B2(P1_U3084), .C1(
        n6162), .C2(n10528), .ZN(P1_U3344) );
  NOR2_X1 U7217 ( .A1(n6146), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6286) );
  OR2_X1 U7218 ( .A1(n6286), .A2(n6287), .ZN(n6197) );
  XNOR2_X1 U7219 ( .A(n6197), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7142) );
  INV_X1 U7220 ( .A(n7142), .ZN(n6544) );
  OAI222_X1 U7221 ( .A1(n10047), .A2(n6148), .B1(n10053), .B2(n6147), .C1(
        n6544), .C2(P2_U3152), .ZN(P2_U3349) );
  NAND2_X1 U7222 ( .A1(n8013), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6154) );
  INV_X1 U7223 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7455) );
  OR2_X1 U7224 ( .A1(n5839), .A2(n7455), .ZN(n6153) );
  INV_X1 U7225 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9645) );
  INV_X1 U7226 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9624) );
  OAI21_X1 U7227 ( .B1(n6156), .B2(n9645), .A(n9624), .ZN(n6150) );
  NAND2_X1 U7228 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n6149) );
  NAND2_X1 U7229 ( .A1(n6150), .A2(n7160), .ZN(n7454) );
  OR2_X1 U7230 ( .A1(n8040), .A2(n7454), .ZN(n6152) );
  INV_X1 U7231 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6547) );
  OR2_X1 U7232 ( .A1(n8093), .A2(n6547), .ZN(n6151) );
  MUX2_X1 U7233 ( .A(n9916), .B(n7448), .S(P2_U3966), .Z(n6155) );
  INV_X1 U7234 ( .A(n6155), .ZN(P2_U3562) );
  NAND2_X1 U7235 ( .A1(n8013), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6161) );
  INV_X1 U7236 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6331) );
  OR2_X1 U7237 ( .A1(n5839), .A2(n6331), .ZN(n6160) );
  XNOR2_X1 U7238 ( .A(n6156), .B(n9645), .ZN(n7426) );
  OR2_X1 U7239 ( .A1(n8040), .A2(n7426), .ZN(n6159) );
  INV_X1 U7240 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6157) );
  OR2_X1 U7241 ( .A1(n8093), .A2(n6157), .ZN(n6158) );
  MUX2_X1 U7242 ( .A(n6162), .B(n7461), .S(P2_U3966), .Z(n6163) );
  INV_X1 U7243 ( .A(n6163), .ZN(P2_U3561) );
  NAND2_X1 U7244 ( .A1(n8013), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6168) );
  INV_X1 U7245 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7689) );
  OR2_X1 U7246 ( .A1(n5839), .A2(n7689), .ZN(n6167) );
  INV_X1 U7247 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6172) );
  XNOR2_X1 U7248 ( .A(n7162), .B(n6172), .ZN(n8385) );
  OR2_X1 U7249 ( .A1(n8040), .A2(n8385), .ZN(n6166) );
  INV_X1 U7250 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6164) );
  OR2_X1 U7251 ( .A1(n8093), .A2(n6164), .ZN(n6165) );
  MUX2_X1 U7252 ( .A(n9695), .B(n8372), .S(P2_U3966), .Z(n6169) );
  INV_X1 U7253 ( .A(n6169), .ZN(P2_U3564) );
  NAND2_X1 U7254 ( .A1(n8013), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6177) );
  INV_X1 U7255 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10675) );
  OR2_X1 U7256 ( .A1(n5839), .A2(n10675), .ZN(n6176) );
  NAND2_X1 U7257 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n6170) );
  INV_X1 U7258 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6171) );
  OAI21_X1 U7259 ( .B1(n7162), .B2(n6172), .A(n6171), .ZN(n6173) );
  NAND2_X1 U7260 ( .A1(n7617), .A2(n6173), .ZN(n8367) );
  OR2_X1 U7261 ( .A1(n8040), .A2(n8367), .ZN(n6175) );
  INV_X1 U7262 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6997) );
  OR2_X1 U7263 ( .A1(n8093), .A2(n6997), .ZN(n6174) );
  MUX2_X1 U7264 ( .A(n9912), .B(n8975), .S(P2_U3966), .Z(n6178) );
  INV_X1 U7265 ( .A(n6178), .ZN(P2_U3565) );
  NAND2_X1 U7266 ( .A1(n8490), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6188) );
  INV_X1 U7267 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6179) );
  OR2_X1 U7268 ( .A1(n8496), .A2(n6179), .ZN(n6187) );
  NAND3_X1 U7269 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6925) );
  INV_X1 U7270 ( .A(n6925), .ZN(n6180) );
  NAND2_X1 U7271 ( .A1(n6180), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7024) );
  INV_X1 U7272 ( .A(n7024), .ZN(n6181) );
  NAND2_X1 U7273 ( .A1(n6181), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7026) );
  INV_X1 U7274 ( .A(n7026), .ZN(n6182) );
  INV_X1 U7275 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7276 ( .A1(n7026), .A2(n6266), .ZN(n6183) );
  NAND2_X1 U7277 ( .A1(n7289), .A2(n6183), .ZN(n10858) );
  OR2_X1 U7278 ( .A1(n6203), .A2(n10858), .ZN(n6186) );
  INV_X1 U7279 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6184) );
  OR2_X1 U7280 ( .A1(n8492), .A2(n6184), .ZN(n6185) );
  NAND4_X1 U7281 ( .A1(n6188), .A2(n6187), .A3(n6186), .A4(n6185), .ZN(n7327)
         );
  NAND2_X1 U7282 ( .A1(n7327), .A2(P1_U4006), .ZN(n6189) );
  OAI21_X1 U7283 ( .B1(P1_U4006), .B2(n6106), .A(n6189), .ZN(P1_U3563) );
  NAND2_X1 U7284 ( .A1(n6190), .A2(n5698), .ZN(n6192) );
  MUX2_X1 U7285 ( .A(n6201), .B(n9916), .S(n5153), .Z(n6194) );
  INV_X1 U7286 ( .A(n6194), .ZN(n6195) );
  NAND2_X1 U7287 ( .A1(n6195), .A2(SI_10_), .ZN(n6196) );
  XNOR2_X1 U7288 ( .A(n6209), .B(n5699), .ZN(n7343) );
  INV_X1 U7289 ( .A(n7343), .ZN(n6208) );
  NAND2_X1 U7290 ( .A1(n6197), .A2(n6284), .ZN(n6198) );
  NAND2_X1 U7291 ( .A1(n6198), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6199) );
  INV_X1 U7292 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7293 ( .A1(n6199), .A2(n6283), .ZN(n6217) );
  OR2_X1 U7294 ( .A1(n6199), .A2(n6283), .ZN(n6200) );
  NAND2_X1 U7295 ( .A1(n6217), .A2(n6200), .ZN(n7139) );
  OAI222_X1 U7296 ( .A1(n10047), .A2(n6201), .B1(n10053), .B2(n6208), .C1(
        n7139), .C2(P2_U3152), .ZN(P2_U3348) );
  NAND2_X1 U7297 ( .A1(n6571), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6607) );
  INV_X1 U7298 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6202) );
  OR2_X1 U7299 ( .A1(n6203), .A2(n6202), .ZN(n6606) );
  INV_X1 U7300 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6204) );
  OR2_X1 U7301 ( .A1(n6469), .A2(n6204), .ZN(n6605) );
  INV_X1 U7302 ( .A(n6808), .ZN(n8295) );
  NAND2_X1 U7303 ( .A1(n8295), .A2(P1_U4006), .ZN(n6205) );
  OAI21_X1 U7304 ( .B1(P1_U4006), .B2(n5843), .A(n6205), .ZN(P1_U3557) );
  NAND2_X1 U7305 ( .A1(n6207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6212) );
  XNOR2_X1 U7306 ( .A(n6212), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7344) );
  INV_X1 U7307 ( .A(n7344), .ZN(n6353) );
  OAI222_X1 U7308 ( .A1(n10528), .A2(n9916), .B1(n6353), .B2(P1_U3084), .C1(
        n10532), .C2(n6208), .ZN(P1_U3343) );
  MUX2_X1 U7309 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7833), .Z(n6275) );
  XNOR2_X1 U7310 ( .A(n6278), .B(n6274), .ZN(n7533) );
  INV_X1 U7311 ( .A(n7533), .ZN(n6219) );
  INV_X1 U7312 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U7313 ( .A1(n6212), .A2(n9720), .ZN(n6213) );
  NAND2_X1 U7314 ( .A1(n6213), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6215) );
  INV_X1 U7315 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6214) );
  XNOR2_X1 U7316 ( .A(n6215), .B(n6214), .ZN(n6361) );
  INV_X1 U7317 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6216) );
  OAI222_X1 U7318 ( .A1(n10532), .A2(n6219), .B1(n6361), .B2(P1_U3084), .C1(
        n6216), .C2(n10528), .ZN(P1_U3342) );
  INV_X1 U7319 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7320 ( .A1(n6217), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6218) );
  XNOR2_X1 U7321 ( .A(n6218), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7223) );
  INV_X1 U7322 ( .A(n7223), .ZN(n6729) );
  OAI222_X1 U7323 ( .A1(n10047), .A2(n6220), .B1(n6076), .B2(n6219), .C1(n6729), .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7324 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6223) );
  INV_X1 U7325 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6572) );
  OAI21_X1 U7326 ( .B1(n6222), .B2(n6230), .A(n6221), .ZN(n10626) );
  MUX2_X1 U7327 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6572), .S(n6578), .Z(n10625)
         );
  NAND2_X1 U7328 ( .A1(n10626), .A2(n10625), .ZN(n10624) );
  OAI21_X1 U7329 ( .B1(n6572), .B2(n10622), .A(n10624), .ZN(n10698) );
  MUX2_X1 U7330 ( .A(n6223), .B(P1_REG2_REG_4__SCAN_IN), .S(n6675), .Z(n10699)
         );
  NOR2_X1 U7331 ( .A1(n10698), .A2(n10699), .ZN(n10697) );
  AOI21_X1 U7332 ( .B1(n10691), .B2(n6223), .A(n10697), .ZN(n6226) );
  INV_X1 U7333 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U7334 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6224), .B1(n6909), .B2(
        n10797), .ZN(n6225) );
  NOR2_X1 U7335 ( .A1(n6226), .A2(n6225), .ZN(n6239) );
  AOI21_X1 U7336 ( .B1(n6226), .B2(n6225), .A(n6239), .ZN(n6236) );
  AND2_X1 U7337 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6933) );
  INV_X1 U7338 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6227) );
  NOR2_X1 U7339 ( .A1(n10618), .A2(n6227), .ZN(n6228) );
  AOI211_X1 U7340 ( .C1(n10605), .C2(n6909), .A(n6933), .B(n6228), .ZN(n6235)
         );
  INV_X1 U7341 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10766) );
  INV_X1 U7342 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6231) );
  OAI21_X1 U7343 ( .B1(n10738), .B2(n6230), .A(n6229), .ZN(n10629) );
  MUX2_X1 U7344 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6231), .S(n6578), .Z(n10628)
         );
  NAND2_X1 U7345 ( .A1(n10629), .A2(n10628), .ZN(n10627) );
  OAI21_X1 U7346 ( .B1(n6231), .B2(n10622), .A(n10627), .ZN(n10690) );
  AOI22_X1 U7347 ( .A1(n6675), .A2(n10766), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n10691), .ZN(n10689) );
  NOR2_X1 U7348 ( .A1(n10690), .A2(n10689), .ZN(n10688) );
  AOI21_X1 U7349 ( .B1(n10691), .B2(n10766), .A(n10688), .ZN(n6233) );
  INV_X1 U7350 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6689) );
  MUX2_X1 U7351 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6689), .S(n6909), .Z(n6232)
         );
  INV_X1 U7352 ( .A(n10693), .ZN(n10636) );
  NAND2_X1 U7353 ( .A1(n6233), .A2(n6232), .ZN(n6245) );
  OAI211_X1 U7354 ( .C1(n6233), .C2(n6232), .A(n10636), .B(n6245), .ZN(n6234)
         );
  OAI211_X1 U7355 ( .C1(n6236), .C2(n10701), .A(n6235), .B(n6234), .ZN(
        P1_U3246) );
  NAND2_X1 U7356 ( .A1(n7007), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6241) );
  INV_X1 U7357 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6237) );
  MUX2_X1 U7358 ( .A(n6237), .B(P1_REG2_REG_6__SCAN_IN), .S(n7007), .Z(n6238)
         );
  INV_X1 U7359 ( .A(n6238), .ZN(n10596) );
  NOR2_X1 U7360 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6909), .ZN(n6240) );
  NOR2_X1 U7361 ( .A1(n6240), .A2(n6239), .ZN(n10597) );
  NAND2_X1 U7362 ( .A1(n10596), .A2(n10597), .ZN(n10595) );
  NAND2_X1 U7363 ( .A1(n6241), .A2(n10595), .ZN(n6244) );
  INV_X1 U7364 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6242) );
  AOI22_X1 U7365 ( .A1(n7118), .A2(n6242), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6248), .ZN(n6243) );
  NOR2_X1 U7366 ( .A1(n6244), .A2(n6243), .ZN(n6256) );
  AOI21_X1 U7367 ( .B1(n6244), .B2(n6243), .A(n6256), .ZN(n6255) );
  AND2_X1 U7368 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U7369 ( .A1(n7007), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6247) );
  INV_X1 U7370 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6924) );
  MUX2_X1 U7371 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6924), .S(n7007), .Z(n10599)
         );
  NAND2_X1 U7372 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6909), .ZN(n6246) );
  NAND2_X1 U7373 ( .A1(n6246), .A2(n6245), .ZN(n10600) );
  NAND2_X1 U7374 ( .A1(n10599), .A2(n10600), .ZN(n10598) );
  NAND2_X1 U7375 ( .A1(n6247), .A2(n10598), .ZN(n6250) );
  INV_X1 U7376 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U7377 ( .A1(n7118), .A2(n10827), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n6248), .ZN(n6249) );
  NOR2_X1 U7378 ( .A1(n6250), .A2(n6249), .ZN(n6261) );
  AOI21_X1 U7379 ( .B1(n6250), .B2(n6249), .A(n6261), .ZN(n6252) );
  INV_X1 U7380 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6251) );
  OAI22_X1 U7381 ( .A1(n6252), .A2(n10693), .B1(n10618), .B2(n6251), .ZN(n6253) );
  AOI211_X1 U7382 ( .C1(n10605), .C2(n7118), .A(n7133), .B(n6253), .ZN(n6254)
         );
  OAI21_X1 U7383 ( .B1(n6255), .B2(n10701), .A(n6254), .ZN(P1_U3248) );
  NOR2_X1 U7384 ( .A1(n7118), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6257) );
  NOR2_X1 U7385 ( .A1(n6257), .A2(n6256), .ZN(n6260) );
  INV_X1 U7386 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6258) );
  AOI22_X1 U7387 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6268), .B1(n7271), .B2(
        n6258), .ZN(n6259) );
  NOR2_X1 U7388 ( .A1(n6260), .A2(n6259), .ZN(n6342) );
  AOI21_X1 U7389 ( .B1(n6260), .B2(n6259), .A(n6342), .ZN(n6273) );
  NOR2_X1 U7390 ( .A1(n7118), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6262) );
  NOR2_X1 U7391 ( .A1(n6262), .A2(n6261), .ZN(n6264) );
  AOI22_X1 U7392 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6268), .B1(n7271), .B2(
        n6179), .ZN(n6263) );
  NOR2_X1 U7393 ( .A1(n6264), .A2(n6263), .ZN(n6337) );
  AOI21_X1 U7394 ( .B1(n6264), .B2(n6263), .A(n6337), .ZN(n6265) );
  NOR2_X1 U7395 ( .A1(n6265), .A2(n10693), .ZN(n6271) );
  NOR2_X1 U7396 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6266), .ZN(n7296) );
  INV_X1 U7397 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6267) );
  NOR2_X1 U7398 ( .A1(n10618), .A2(n6267), .ZN(n6270) );
  NOR2_X1 U7399 ( .A1(n10692), .A2(n6268), .ZN(n6269) );
  NOR4_X1 U7400 ( .A1(n6271), .A2(n7296), .A3(n6270), .A4(n6269), .ZN(n6272)
         );
  OAI21_X1 U7401 ( .B1(n6273), .B2(n10701), .A(n6272), .ZN(P1_U3249) );
  NAND2_X1 U7402 ( .A1(n6275), .A2(SI_11_), .ZN(n6276) );
  MUX2_X1 U7403 ( .A(n6289), .B(n9695), .S(n5153), .Z(n6279) );
  INV_X1 U7404 ( .A(n6279), .ZN(n6280) );
  NAND2_X1 U7405 ( .A1(n6280), .A2(SI_12_), .ZN(n6281) );
  NAND2_X1 U7406 ( .A1(n6370), .A2(n6281), .ZN(n6368) );
  XNOR2_X1 U7407 ( .A(n6369), .B(n6368), .ZN(n7702) );
  INV_X1 U7408 ( .A(n7702), .ZN(n6291) );
  INV_X1 U7409 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6282) );
  AND3_X1 U7410 ( .A1(n6284), .A2(n6283), .A3(n6282), .ZN(n6285) );
  AND2_X1 U7411 ( .A1(n6286), .A2(n6285), .ZN(n6485) );
  OR2_X1 U7412 ( .A1(n6485), .A2(n6287), .ZN(n6288) );
  XNOR2_X1 U7413 ( .A(n6288), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7601) );
  INV_X1 U7414 ( .A(n7601), .ZN(n6996) );
  OAI222_X1 U7415 ( .A1(n10047), .A2(n6289), .B1(n6076), .B2(n6291), .C1(
        P2_U3152), .C2(n6996), .ZN(P2_U3346) );
  OR2_X1 U7416 ( .A1(n5136), .A2(n6374), .ZN(n6290) );
  XNOR2_X1 U7417 ( .A(n6290), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7703) );
  INV_X1 U7418 ( .A(n7703), .ZN(n6644) );
  OAI222_X1 U7419 ( .A1(n10528), .A2(n9695), .B1(n10532), .B2(n6291), .C1(
        P1_U3084), .C2(n6644), .ZN(P1_U3341) );
  MUX2_X1 U7420 ( .A(n5902), .B(P2_REG2_REG_5__SCAN_IN), .S(n6322), .Z(n6323)
         );
  INV_X1 U7421 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7076) );
  AOI21_X1 U7422 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n6296), .A(n6292), .ZN(
        n6418) );
  INV_X1 U7423 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6955) );
  MUX2_X1 U7424 ( .A(n6955), .B(P2_REG2_REG_3__SCAN_IN), .S(n6298), .Z(n6417)
         );
  NOR2_X1 U7425 ( .A1(n6418), .A2(n6417), .ZN(n6434) );
  NOR2_X1 U7426 ( .A1(n6422), .A2(n6955), .ZN(n6429) );
  MUX2_X1 U7427 ( .A(n7076), .B(P2_REG2_REG_4__SCAN_IN), .S(n6437), .Z(n6293)
         );
  OAI21_X1 U7428 ( .B1(n6434), .B2(n6429), .A(n6293), .ZN(n6432) );
  OAI21_X1 U7429 ( .B1(n7076), .B2(n6437), .A(n6432), .ZN(n6325) );
  XOR2_X1 U7430 ( .A(n6323), .B(n6325), .Z(n6306) );
  INV_X1 U7431 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7432 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8958) );
  OAI21_X1 U7433 ( .B1(n9257), .B2(n6294), .A(n8958), .ZN(n6304) );
  AOI21_X1 U7434 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n6296), .A(n6295), .ZN(
        n6414) );
  MUX2_X1 U7435 ( .A(n6297), .B(P2_REG1_REG_3__SCAN_IN), .S(n6298), .Z(n6413)
         );
  NOR2_X1 U7436 ( .A1(n6414), .A2(n6413), .ZN(n6412) );
  AOI21_X1 U7437 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n6298), .A(n6412), .ZN(
        n6426) );
  MUX2_X1 U7438 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6299), .S(n6437), .Z(n6425)
         );
  NOR2_X1 U7439 ( .A1(n6426), .A2(n6425), .ZN(n6424) );
  AOI21_X1 U7440 ( .B1(n5320), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6424), .ZN(
        n6302) );
  NAND2_X1 U7441 ( .A1(n6322), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6300) );
  OAI21_X1 U7442 ( .B1(n6322), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6300), .ZN(
        n6301) );
  NOR2_X1 U7443 ( .A1(n6302), .A2(n6301), .ZN(n6308) );
  AOI211_X1 U7444 ( .C1(n6302), .C2(n6301), .A(n10658), .B(n6308), .ZN(n6303)
         );
  AOI211_X1 U7445 ( .C1(n10660), .C2(n6322), .A(n6304), .B(n6303), .ZN(n6305)
         );
  OAI21_X1 U7446 ( .B1(n9278), .B2(n6306), .A(n6305), .ZN(P2_U3250) );
  XNOR2_X1 U7447 ( .A(n7053), .B(n6307), .ZN(n6400) );
  NAND2_X1 U7448 ( .A1(n6319), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6312) );
  AOI21_X1 U7449 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n6322), .A(n6308), .ZN(
        n6390) );
  NAND2_X1 U7450 ( .A1(n6320), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6309) );
  OAI21_X1 U7451 ( .B1(n6320), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6309), .ZN(
        n6389) );
  NOR2_X1 U7452 ( .A1(n6390), .A2(n6389), .ZN(n6388) );
  AOI21_X1 U7453 ( .B1(n6320), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6388), .ZN(
        n6379) );
  MUX2_X1 U7454 ( .A(n6310), .B(P2_REG1_REG_7__SCAN_IN), .S(n6319), .Z(n6378)
         );
  NOR2_X1 U7455 ( .A1(n6379), .A2(n6378), .ZN(n6377) );
  INV_X1 U7456 ( .A(n6377), .ZN(n6311) );
  NAND2_X1 U7457 ( .A1(n6312), .A2(n6311), .ZN(n6399) );
  AND2_X1 U7458 ( .A1(n7053), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7459 ( .A1(n7142), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6550) );
  OAI21_X1 U7460 ( .B1(n7142), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6550), .ZN(
        n6314) );
  INV_X1 U7461 ( .A(n6314), .ZN(n6315) );
  XNOR2_X1 U7462 ( .A(n6548), .B(n6315), .ZN(n6317) );
  NAND2_X1 U7463 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7176) );
  NAND2_X1 U7464 ( .A1(n10674), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6316) );
  OAI211_X1 U7465 ( .C1(n10658), .C2(n6317), .A(n7176), .B(n6316), .ZN(n6318)
         );
  AOI21_X1 U7466 ( .B1(n7142), .B2(n10660), .A(n6318), .ZN(n6335) );
  MUX2_X1 U7467 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6330), .S(n7053), .Z(n6407)
         );
  NAND2_X1 U7468 ( .A1(n6319), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6329) );
  MUX2_X1 U7469 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7093), .S(n6319), .Z(n6383)
         );
  NAND2_X1 U7470 ( .A1(n6320), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6328) );
  MUX2_X1 U7471 ( .A(n5919), .B(P2_REG2_REG_6__SCAN_IN), .S(n6320), .Z(n6321)
         );
  INV_X1 U7472 ( .A(n6321), .ZN(n6394) );
  NAND2_X1 U7473 ( .A1(n6322), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6327) );
  INV_X1 U7474 ( .A(n6323), .ZN(n6324) );
  NAND2_X1 U7475 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  NAND2_X1 U7476 ( .A1(n6327), .A2(n6326), .ZN(n6395) );
  NAND2_X1 U7477 ( .A1(n6394), .A2(n6395), .ZN(n6393) );
  NAND2_X1 U7478 ( .A1(n6328), .A2(n6393), .ZN(n6384) );
  NAND2_X1 U7479 ( .A1(n6383), .A2(n6384), .ZN(n6382) );
  NAND2_X1 U7480 ( .A1(n6329), .A2(n6382), .ZN(n6406) );
  NAND2_X1 U7481 ( .A1(n6407), .A2(n6406), .ZN(n6405) );
  OAI21_X1 U7482 ( .B1(n6330), .B2(n6410), .A(n6405), .ZN(n6333) );
  MUX2_X1 U7483 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6331), .S(n7142), .Z(n6332)
         );
  NAND2_X1 U7484 ( .A1(n6332), .A2(n6333), .ZN(n6543) );
  OAI211_X1 U7485 ( .C1(n6333), .C2(n6332), .A(n10679), .B(n6543), .ZN(n6334)
         );
  NAND2_X1 U7486 ( .A1(n6335), .A2(n6334), .ZN(P2_U3254) );
  INV_X1 U7487 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7479) );
  NOR2_X1 U7488 ( .A1(n7271), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6336) );
  NOR2_X1 U7489 ( .A1(n6337), .A2(n6336), .ZN(n10608) );
  MUX2_X1 U7490 ( .A(n7479), .B(P1_REG1_REG_9__SCAN_IN), .S(n10604), .Z(n10607) );
  NOR2_X1 U7491 ( .A1(n10608), .A2(n10607), .ZN(n10606) );
  AOI21_X1 U7492 ( .B1(n6338), .B2(n7479), .A(n10606), .ZN(n6340) );
  INV_X1 U7493 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U7494 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6353), .B1(n7344), .B2(
        n10894), .ZN(n6339) );
  NOR2_X1 U7495 ( .A1(n6340), .A2(n6339), .ZN(n6352) );
  AOI21_X1 U7496 ( .B1(n6340), .B2(n6339), .A(n6352), .ZN(n6351) );
  INV_X1 U7497 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U7498 ( .A1(n10604), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6343) );
  INV_X1 U7499 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7287) );
  MUX2_X1 U7500 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n7287), .S(n10604), .Z(n10611) );
  NOR2_X1 U7501 ( .A1(n7271), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6341) );
  NOR2_X1 U7502 ( .A1(n6342), .A2(n6341), .ZN(n10612) );
  NAND2_X1 U7503 ( .A1(n10611), .A2(n10612), .ZN(n10610) );
  NAND2_X1 U7504 ( .A1(n6343), .A2(n10610), .ZN(n6345) );
  INV_X1 U7505 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7373) );
  MUX2_X1 U7506 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7373), .S(n7344), .Z(n6344)
         );
  INV_X1 U7507 ( .A(n10701), .ZN(n10640) );
  NAND2_X1 U7508 ( .A1(n6344), .A2(n6345), .ZN(n6355) );
  OAI211_X1 U7509 ( .C1(n6345), .C2(n6344), .A(n10640), .B(n6355), .ZN(n6347)
         );
  NOR2_X1 U7510 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7313), .ZN(n7442) );
  AOI21_X1 U7511 ( .B1(n10605), .B2(n7344), .A(n7442), .ZN(n6346) );
  OAI211_X1 U7512 ( .C1(n10618), .C2(n6348), .A(n6347), .B(n6346), .ZN(n6349)
         );
  INV_X1 U7513 ( .A(n6349), .ZN(n6350) );
  OAI21_X1 U7514 ( .B1(n6351), .B2(n10693), .A(n6350), .ZN(P1_U3251) );
  AOI21_X1 U7515 ( .B1(n10894), .B2(n6353), .A(n6352), .ZN(n6638) );
  INV_X1 U7516 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10915) );
  NOR2_X1 U7517 ( .A1(n6361), .A2(n10915), .ZN(n6637) );
  AOI21_X1 U7518 ( .B1(n6361), .B2(n10915), .A(n6637), .ZN(n6354) );
  XNOR2_X1 U7519 ( .A(n6638), .B(n6354), .ZN(n6367) );
  AND2_X1 U7520 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7557) );
  NAND2_X1 U7521 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7344), .ZN(n6356) );
  NAND2_X1 U7522 ( .A1(n6356), .A2(n6355), .ZN(n6364) );
  AND2_X1 U7523 ( .A1(n6364), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6362) );
  INV_X1 U7524 ( .A(n6357), .ZN(n6358) );
  NAND2_X1 U7525 ( .A1(n6362), .A2(n6358), .ZN(n6359) );
  AOI21_X1 U7526 ( .B1(n6359), .B2(n10692), .A(n6361), .ZN(n6360) );
  AOI211_X1 U7527 ( .C1(n10696), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7557), .B(
        n6360), .ZN(n6366) );
  INV_X1 U7528 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7571) );
  NAND2_X1 U7529 ( .A1(n6361), .A2(n7571), .ZN(n6363) );
  INV_X1 U7530 ( .A(n6361), .ZN(n7534) );
  OAI22_X1 U7531 ( .A1(n6362), .A2(n7534), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n6364), .ZN(n6647) );
  OAI211_X1 U7532 ( .C1(n6364), .C2(n6363), .A(n6647), .B(n10640), .ZN(n6365)
         );
  OAI211_X1 U7533 ( .C1(n6367), .C2(n10693), .A(n6366), .B(n6365), .ZN(
        P1_U3252) );
  MUX2_X1 U7534 ( .A(n6487), .B(n9912), .S(n7833), .Z(n6371) );
  INV_X1 U7535 ( .A(n6371), .ZN(n6372) );
  NAND2_X1 U7536 ( .A1(n6372), .A2(SI_13_), .ZN(n6373) );
  XNOR2_X1 U7537 ( .A(n6488), .B(n5700), .ZN(n7732) );
  INV_X1 U7538 ( .A(n7732), .ZN(n6486) );
  OR2_X1 U7539 ( .A1(n5744), .A2(n6374), .ZN(n6375) );
  XNOR2_X1 U7540 ( .A(n6375), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7733) );
  INV_X1 U7541 ( .A(n10528), .ZN(n10525) );
  AOI22_X1 U7542 ( .A1(n7733), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10525), .ZN(n6376) );
  OAI21_X1 U7543 ( .B1(n6486), .B2(n10532), .A(n6376), .ZN(P1_U3340) );
  NOR2_X1 U7544 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5768), .ZN(n6381) );
  AOI211_X1 U7545 ( .C1(n6379), .C2(n6378), .A(n6377), .B(n10658), .ZN(n6380)
         );
  AOI211_X1 U7546 ( .C1(n10674), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6381), .B(
        n6380), .ZN(n6386) );
  OAI211_X1 U7547 ( .C1(n6384), .C2(n6383), .A(n10679), .B(n6382), .ZN(n6385)
         );
  OAI211_X1 U7548 ( .C1(n10670), .C2(n6387), .A(n6386), .B(n6385), .ZN(
        P2_U3252) );
  NAND2_X1 U7549 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8354) );
  INV_X1 U7550 ( .A(n8354), .ZN(n6392) );
  AOI211_X1 U7551 ( .C1(n6390), .C2(n6389), .A(n6388), .B(n10658), .ZN(n6391)
         );
  AOI211_X1 U7552 ( .C1(n10674), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6392), .B(
        n6391), .ZN(n6397) );
  OAI211_X1 U7553 ( .C1(n6395), .C2(n6394), .A(n10679), .B(n6393), .ZN(n6396)
         );
  OAI211_X1 U7554 ( .C1(n10670), .C2(n6398), .A(n6397), .B(n6396), .ZN(
        P2_U3251) );
  NOR2_X1 U7555 ( .A1(n9841), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7058) );
  INV_X1 U7556 ( .A(n6399), .ZN(n6403) );
  INV_X1 U7557 ( .A(n6400), .ZN(n6402) );
  AOI211_X1 U7558 ( .C1(n6403), .C2(n6402), .A(n6401), .B(n10658), .ZN(n6404)
         );
  AOI211_X1 U7559 ( .C1(n10674), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7058), .B(
        n6404), .ZN(n6409) );
  OAI211_X1 U7560 ( .C1(n6407), .C2(n6406), .A(n10679), .B(n6405), .ZN(n6408)
         );
  OAI211_X1 U7561 ( .C1(n10670), .C2(n6410), .A(n6409), .B(n6408), .ZN(
        P2_U3253) );
  INV_X1 U7562 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6411) );
  NOR2_X1 U7563 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6411), .ZN(n6416) );
  AOI211_X1 U7564 ( .C1(n6414), .C2(n6413), .A(n6412), .B(n10658), .ZN(n6415)
         );
  AOI211_X1 U7565 ( .C1(n10674), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6416), .B(
        n6415), .ZN(n6421) );
  AOI211_X1 U7566 ( .C1(n6418), .C2(n6417), .A(n6434), .B(n9278), .ZN(n6419)
         );
  INV_X1 U7567 ( .A(n6419), .ZN(n6420) );
  OAI211_X1 U7568 ( .C1(n10670), .C2(n6422), .A(n6421), .B(n6420), .ZN(
        P2_U3248) );
  INV_X1 U7569 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6423) );
  NOR2_X1 U7570 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6423), .ZN(n6428) );
  AOI211_X1 U7571 ( .C1(n6426), .C2(n6425), .A(n6424), .B(n10658), .ZN(n6427)
         );
  AOI211_X1 U7572 ( .C1(n10674), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6428), .B(
        n6427), .ZN(n6436) );
  MUX2_X1 U7573 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7076), .S(n6437), .Z(n6431)
         );
  INV_X1 U7574 ( .A(n6429), .ZN(n6430) );
  NAND2_X1 U7575 ( .A1(n6431), .A2(n6430), .ZN(n6433) );
  OAI211_X1 U7576 ( .C1(n6434), .C2(n6433), .A(n10679), .B(n6432), .ZN(n6435)
         );
  OAI211_X1 U7577 ( .C1(n10670), .C2(n6437), .A(n6436), .B(n6435), .ZN(
        P2_U3249) );
  AOI21_X1 U7578 ( .B1(n6440), .B2(n6439), .A(n6438), .ZN(n6443) );
  OAI22_X1 U7579 ( .A1(n5463), .A2(n9466), .B1(n6656), .B2(n9468), .ZN(n6536)
         );
  OAI22_X1 U7580 ( .A1(n6524), .A2(n6936), .B1(n6538), .B2(n9211), .ZN(n6441)
         );
  AOI21_X1 U7581 ( .B1(n6536), .B2(n9208), .A(n6441), .ZN(n6442) );
  OAI21_X1 U7582 ( .B1(n6443), .B2(n9195), .A(n6442), .ZN(P2_U3224) );
  NOR4_X1 U7583 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6453) );
  NOR4_X1 U7584 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6452) );
  OR4_X1 U7585 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6450) );
  NOR4_X1 U7586 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6448) );
  NOR4_X1 U7587 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6447) );
  NOR4_X1 U7588 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6446) );
  NOR4_X1 U7589 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6445) );
  NAND4_X1 U7590 ( .A1(n6448), .A2(n6447), .A3(n6446), .A4(n6445), .ZN(n6449)
         );
  NOR4_X1 U7591 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        n6450), .A4(n6449), .ZN(n6451) );
  AND3_X1 U7592 ( .A1(n6453), .A2(n6452), .A3(n6451), .ZN(n6454) );
  NOR2_X1 U7593 ( .A1(n6455), .A2(n6454), .ZN(n6492) );
  NOR2_X1 U7594 ( .A1(n6800), .A2(n6492), .ZN(n6458) );
  INV_X1 U7595 ( .A(n6455), .ZN(n6457) );
  INV_X1 U7596 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9979) );
  AND2_X1 U7597 ( .A1(n7844), .A2(n7825), .ZN(n6456) );
  AND2_X1 U7598 ( .A1(n6458), .A2(n10522), .ZN(n6477) );
  INV_X1 U7599 ( .A(n6477), .ZN(n6462) );
  NAND2_X1 U7600 ( .A1(n8619), .A2(n8667), .ZN(n6498) );
  NAND3_X1 U7601 ( .A1(n11047), .A2(n6479), .A3(n8501), .ZN(n6459) );
  OR2_X1 U7602 ( .A1(n6498), .A2(n10708), .ZN(n6823) );
  INV_X1 U7603 ( .A(n6823), .ZN(n6460) );
  NAND3_X1 U7604 ( .A1(n6462), .A2(n6479), .A3(n6460), .ZN(n6568) );
  OR2_X1 U7605 ( .A1(n8501), .A2(n6461), .ZN(n6564) );
  NAND2_X1 U7606 ( .A1(n6564), .A2(n6479), .ZN(n6493) );
  INV_X1 U7607 ( .A(n6493), .ZN(n6463) );
  NAND2_X1 U7608 ( .A1(n6462), .A2(n11047), .ZN(n6565) );
  NAND3_X1 U7609 ( .A1(n6568), .A2(n6463), .A3(n6565), .ZN(n10179) );
  AOI22_X1 U7610 ( .A1(n6464), .A2(n10197), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10179), .ZN(n6483) );
  OR2_X1 U7611 ( .A1(n7349), .A2(n6584), .ZN(n8678) );
  INV_X1 U7612 ( .A(n6479), .ZN(n10521) );
  NOR2_X1 U7613 ( .A1(n8678), .A2(n10521), .ZN(n6466) );
  AND2_X1 U7614 ( .A1(n6477), .A2(n6466), .ZN(n6627) );
  NAND2_X1 U7615 ( .A1(n6627), .A2(n6007), .ZN(n10215) );
  INV_X1 U7616 ( .A(n10215), .ZN(n10191) );
  INV_X1 U7617 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6468) );
  OR2_X1 U7618 ( .A1(n6469), .A2(n6468), .ZN(n6474) );
  NAND2_X1 U7619 ( .A1(n6571), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U7620 ( .A1(n8254), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6472) );
  NOR2_X1 U7621 ( .A1(n6823), .A2(n10521), .ZN(n6476) );
  NAND2_X1 U7622 ( .A1(n6477), .A2(n6476), .ZN(n6481) );
  NAND2_X1 U7623 ( .A1(n6479), .A2(n10789), .ZN(n6480) );
  AOI22_X1 U7624 ( .A1(n10191), .A2(n10732), .B1(n5363), .B2(n10223), .ZN(
        n6482) );
  NAND2_X1 U7625 ( .A1(n6483), .A2(n6482), .ZN(P1_U3230) );
  NAND2_X1 U7626 ( .A1(n6485), .A2(n6484), .ZN(n6794) );
  NAND2_X1 U7627 ( .A1(n6794), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6507) );
  XNOR2_X1 U7628 ( .A(n6507), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7608) );
  INV_X1 U7629 ( .A(n7608), .ZN(n10676) );
  OAI222_X1 U7630 ( .A1(n9110), .A2(n6487), .B1(n6076), .B2(n6486), .C1(n10676), .C2(P2_U3152), .ZN(P2_U3345) );
  MUX2_X1 U7631 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7833), .Z(n6772) );
  XNOR2_X1 U7632 ( .A(n6771), .B(n6769), .ZN(n7801) );
  INV_X1 U7633 ( .A(n7801), .ZN(n6511) );
  NAND2_X1 U7634 ( .A1(n6490), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6778) );
  XNOR2_X1 U7635 ( .A(n6778), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7802) );
  AOI22_X1 U7636 ( .A1(n7802), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10525), .ZN(n6491) );
  OAI21_X1 U7637 ( .B1(n6511), .B2(n10532), .A(n6491), .ZN(P1_U3339) );
  INV_X1 U7638 ( .A(n10522), .ZN(n6494) );
  OAI21_X1 U7639 ( .B1(n11043), .B2(n10359), .A(n6494), .ZN(n6495) );
  INV_X1 U7640 ( .A(n6800), .ZN(n6496) );
  AND2_X1 U7641 ( .A1(n6803), .A2(n8297), .ZN(n8395) );
  NOR2_X1 U7642 ( .A1(n8294), .A2(n8395), .ZN(n8641) );
  INV_X1 U7643 ( .A(n8678), .ZN(n6499) );
  INV_X1 U7644 ( .A(n6498), .ZN(n6501) );
  NOR3_X1 U7645 ( .A1(n8641), .A2(n6499), .A3(n6501), .ZN(n6500) );
  AOI21_X1 U7646 ( .B1(n11037), .B2(n10732), .A(n6500), .ZN(n10706) );
  NAND2_X1 U7647 ( .A1(n5363), .A2(n6501), .ZN(n10707) );
  NAND2_X1 U7648 ( .A1(n10706), .A2(n10707), .ZN(n6504) );
  NAND2_X1 U7649 ( .A1(n6504), .A2(n11054), .ZN(n6502) );
  OAI21_X1 U7650 ( .B1(n11054), .B2(n6010), .A(n6502), .ZN(P1_U3523) );
  NAND2_X1 U7651 ( .A1(n6504), .A2(n11057), .ZN(n6505) );
  OAI21_X1 U7652 ( .B1(n11057), .B2(n6014), .A(n6505), .ZN(P1_U3454) );
  INV_X1 U7653 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6512) );
  INV_X1 U7654 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U7655 ( .A1(n6507), .A2(n6506), .ZN(n6508) );
  NAND2_X1 U7656 ( .A1(n6508), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U7657 ( .A1(n6509), .A2(n6791), .ZN(n6781) );
  OR2_X1 U7658 ( .A1(n6509), .A2(n6791), .ZN(n6510) );
  INV_X1 U7659 ( .A(n7613), .ZN(n7245) );
  OAI222_X1 U7660 ( .A1(n10047), .A2(n6512), .B1(n10053), .B2(n6511), .C1(
        n7245), .C2(P2_U3152), .ZN(P2_U3344) );
  AOI211_X1 U7661 ( .C1(n6514), .C2(n6513), .A(n9195), .B(n5403), .ZN(n6518)
         );
  MUX2_X1 U7662 ( .A(n9206), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6516) );
  INV_X1 U7663 ( .A(n9161), .ZN(n9185) );
  AOI22_X1 U7664 ( .A1(n9224), .A2(n9185), .B1(n5471), .B2(n9171), .ZN(n6515)
         );
  OAI211_X1 U7665 ( .C1(n6656), .C2(n9159), .A(n6516), .B(n6515), .ZN(n6517)
         );
  OR2_X1 U7666 ( .A1(n6518), .A2(n6517), .ZN(P2_U3220) );
  NAND2_X1 U7667 ( .A1(n6520), .A2(n6519), .ZN(n6523) );
  AOI22_X1 U7668 ( .A1(n6531), .A2(n9185), .B1(n9171), .B2(n6521), .ZN(n6522)
         );
  OAI211_X1 U7669 ( .C1(n6524), .C2(n6890), .A(n6523), .B(n6522), .ZN(P2_U3234) );
  NAND4_X1 U7670 ( .A1(n10543), .A2(n6869), .A3(n6525), .A4(n6874), .ZN(n6526)
         );
  INV_X1 U7671 ( .A(n6875), .ZN(n6528) );
  INV_X2 U7672 ( .A(n11019), .ZN(n11001) );
  INV_X1 U7673 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U7674 ( .A1(n7425), .A2(n6652), .ZN(n11015) );
  INV_X1 U7675 ( .A(n6531), .ZN(n6530) );
  NAND2_X1 U7676 ( .A1(n6530), .A2(n6529), .ZN(n6661) );
  NAND2_X1 U7677 ( .A1(n6531), .A2(n6538), .ZN(n6660) );
  OAI21_X1 U7678 ( .B1(n6534), .B2(n6532), .A(n6654), .ZN(n6942) );
  INV_X1 U7679 ( .A(n6887), .ZN(n6533) );
  NAND2_X1 U7680 ( .A1(n8859), .A2(n8887), .ZN(n8700) );
  NAND2_X1 U7681 ( .A1(n8895), .A2(n5819), .ZN(n8854) );
  AOI21_X1 U7682 ( .B1(n6534), .B2(n6533), .A(n9486), .ZN(n6537) );
  INV_X1 U7683 ( .A(n6534), .ZN(n6535) );
  AOI21_X1 U7684 ( .B1(n6537), .B2(n8863), .A(n6536), .ZN(n6945) );
  NOR2_X1 U7685 ( .A1(n6939), .A2(n11011), .ZN(n6539) );
  AOI22_X1 U7686 ( .A1(n6539), .A2(n6937), .B1(n6529), .B2(n10925), .ZN(n6540)
         );
  OAI211_X1 U7687 ( .C1(n10992), .C2(n6942), .A(n6945), .B(n6540), .ZN(n6561)
         );
  NAND2_X1 U7688 ( .A1(n6561), .A2(n11001), .ZN(n6541) );
  OAI21_X1 U7689 ( .B1(n11001), .B2(n6542), .A(n6541), .ZN(P2_U3454) );
  INV_X1 U7690 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U7691 ( .A1(n7223), .A2(n10948), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n6729), .ZN(n6546) );
  MUX2_X1 U7692 ( .A(n7455), .B(P2_REG2_REG_10__SCAN_IN), .S(n7139), .Z(n9230)
         );
  OAI21_X1 U7693 ( .B1(n6544), .B2(n6331), .A(n6543), .ZN(n9229) );
  NAND2_X1 U7694 ( .A1(n9230), .A2(n9229), .ZN(n9228) );
  OAI21_X1 U7695 ( .B1(n7455), .B2(n7139), .A(n9228), .ZN(n6545) );
  NOR2_X1 U7696 ( .A1(n6545), .A2(n6546), .ZN(n6726) );
  AOI21_X1 U7697 ( .B1(n6546), .B2(n6545), .A(n6726), .ZN(n6559) );
  INV_X1 U7698 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7163) );
  MUX2_X1 U7699 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7163), .S(n7223), .Z(n6553)
         );
  MUX2_X1 U7700 ( .A(n6547), .B(P2_REG1_REG_10__SCAN_IN), .S(n7139), .Z(n9234)
         );
  INV_X1 U7701 ( .A(n6548), .ZN(n6551) );
  NOR2_X1 U7702 ( .A1(n7142), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6549) );
  AOI21_X1 U7703 ( .B1(n6551), .B2(n6550), .A(n6549), .ZN(n9235) );
  NAND2_X1 U7704 ( .A1(n9234), .A2(n9235), .ZN(n9233) );
  OAI21_X1 U7705 ( .B1(n7139), .B2(n6547), .A(n9233), .ZN(n6552) );
  NAND2_X1 U7706 ( .A1(n6553), .A2(n6552), .ZN(n6728) );
  OAI21_X1 U7707 ( .B1(n6553), .B2(n6552), .A(n6728), .ZN(n6556) );
  OR2_X1 U7708 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7240), .ZN(n6555) );
  NAND2_X1 U7709 ( .A1(n10674), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6554) );
  OAI211_X1 U7710 ( .C1(n10658), .C2(n6556), .A(n6555), .B(n6554), .ZN(n6557)
         );
  AOI21_X1 U7711 ( .B1(n7223), .B2(n10660), .A(n6557), .ZN(n6558) );
  OAI21_X1 U7712 ( .B1(n6559), .B2(n9278), .A(n6558), .ZN(P2_U3256) );
  NAND2_X1 U7713 ( .A1(n6561), .A2(n11018), .ZN(n6562) );
  OAI21_X1 U7714 ( .B1(n11018), .B2(n5992), .A(n6562), .ZN(P2_U3521) );
  AND3_X1 U7715 ( .A1(n6564), .A2(n6563), .A3(n7583), .ZN(n6566) );
  NAND2_X1 U7716 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  NAND2_X1 U7717 ( .A1(n6567), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6569) );
  NAND2_X1 U7718 ( .A1(n8162), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6576) );
  INV_X1 U7719 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6570) );
  OR2_X1 U7720 ( .A1(n8492), .A2(n6570), .ZN(n6575) );
  NAND2_X1 U7721 ( .A1(n10731), .A2(n9086), .ZN(n6583) );
  NAND2_X1 U7723 ( .A1(n6609), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U7724 ( .A1(n8133), .A2(n6578), .ZN(n6579) );
  NAND2_X1 U7725 ( .A1(n8406), .A2(n7122), .ZN(n6582) );
  AND2_X1 U7726 ( .A1(n8406), .A2(n9080), .ZN(n6586) );
  AOI21_X1 U7727 ( .B1(n10731), .B2(n9085), .A(n6586), .ZN(n6671) );
  INV_X1 U7728 ( .A(n6587), .ZN(n6588) );
  NAND2_X1 U7729 ( .A1(n6588), .A2(n9076), .ZN(n6590) );
  INV_X1 U7730 ( .A(n6603), .ZN(n6599) );
  NAND2_X1 U7731 ( .A1(n6804), .A2(n6600), .ZN(n6596) );
  NAND2_X1 U7732 ( .A1(n8300), .A2(n7122), .ZN(n6595) );
  NAND2_X1 U7733 ( .A1(n6596), .A2(n6595), .ZN(n6597) );
  INV_X1 U7734 ( .A(n6602), .ZN(n6598) );
  INV_X1 U7735 ( .A(n10720), .ZN(n8300) );
  AND2_X1 U7736 ( .A1(n8300), .A2(n9080), .ZN(n6601) );
  AOI21_X1 U7737 ( .B1(n10732), .B2(n9085), .A(n6601), .ZN(n8288) );
  NAND2_X1 U7738 ( .A1(n8286), .A2(n8288), .ZN(n6604) );
  NAND2_X1 U7739 ( .A1(n6603), .A2(n6602), .ZN(n8287) );
  NAND4_X1 U7740 ( .A1(n6608), .A2(n6607), .A3(n6606), .A4(n6605), .ZN(n6807)
         );
  NAND2_X1 U7741 ( .A1(n6807), .A2(n9086), .ZN(n6615) );
  NAND2_X1 U7742 ( .A1(n6609), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U7743 ( .A1(n8133), .A2(n6610), .ZN(n6611) );
  OAI211_X1 U7744 ( .C1(n7005), .C2(n6613), .A(n6612), .B(n6611), .ZN(n10178)
         );
  NAND2_X1 U7745 ( .A1(n10178), .A2(n7122), .ZN(n6614) );
  NAND2_X1 U7746 ( .A1(n6615), .A2(n6614), .ZN(n6616) );
  XNOR2_X1 U7747 ( .A(n6616), .B(n9083), .ZN(n6618) );
  AND2_X1 U7748 ( .A1(n10178), .A2(n9086), .ZN(n6617) );
  AOI21_X1 U7749 ( .B1(n6807), .B2(n9085), .A(n6617), .ZN(n6619) );
  NAND2_X1 U7750 ( .A1(n6618), .A2(n6619), .ZN(n6623) );
  INV_X1 U7751 ( .A(n6618), .ZN(n6621) );
  INV_X1 U7752 ( .A(n6619), .ZN(n6620) );
  NAND2_X1 U7753 ( .A1(n6621), .A2(n6620), .ZN(n6622) );
  AND2_X1 U7754 ( .A1(n6623), .A2(n6622), .ZN(n10176) );
  NAND2_X1 U7755 ( .A1(n10175), .A2(n10176), .ZN(n10174) );
  OAI21_X1 U7756 ( .B1(n6625), .B2(n6624), .A(n6674), .ZN(n6626) );
  NAND2_X1 U7757 ( .A1(n6626), .A2(n10197), .ZN(n6636) );
  INV_X1 U7758 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6899) );
  NOR2_X1 U7759 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6899), .ZN(n10619) );
  INV_X1 U7760 ( .A(n6627), .ZN(n6628) );
  OR2_X1 U7761 ( .A1(n6628), .A2(n6007), .ZN(n10126) );
  INV_X2 U7762 ( .A(n8492), .ZN(n8238) );
  NAND2_X1 U7763 ( .A1(n8238), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6633) );
  OR2_X1 U7764 ( .A1(n6629), .A2(n6223), .ZN(n6632) );
  OR2_X1 U7765 ( .A1(n8496), .A2(n10766), .ZN(n6631) );
  XNOR2_X1 U7766 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6824) );
  OR2_X1 U7767 ( .A1(n6203), .A2(n6824), .ZN(n6630) );
  OAI22_X1 U7768 ( .A1(n10126), .A2(n6808), .B1(n10778), .B2(n10215), .ZN(
        n6634) );
  AOI211_X1 U7769 ( .C1(n8406), .C2(n10223), .A(n10619), .B(n6634), .ZN(n6635)
         );
  OAI211_X1 U7770 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n10221), .A(n6636), .B(
        n6635), .ZN(P1_U3216) );
  OAI22_X1 U7771 ( .A1(n6638), .A2(n6637), .B1(n7534), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n6641) );
  INV_X1 U7772 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10963) );
  NOR2_X1 U7773 ( .A1(n6644), .A2(n10963), .ZN(n6639) );
  AOI21_X1 U7774 ( .B1(n10963), .B2(n6644), .A(n6639), .ZN(n6640) );
  NAND2_X1 U7775 ( .A1(n6640), .A2(n6641), .ZN(n6740) );
  OAI21_X1 U7776 ( .B1(n6641), .B2(n6640), .A(n6740), .ZN(n6642) );
  INV_X1 U7777 ( .A(n6642), .ZN(n6651) );
  INV_X1 U7778 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7549) );
  NOR2_X1 U7779 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7549), .ZN(n7721) );
  INV_X1 U7780 ( .A(n7721), .ZN(n6643) );
  OAI21_X1 U7781 ( .B1(n10692), .B2(n6644), .A(n6643), .ZN(n6649) );
  NAND2_X1 U7782 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7703), .ZN(n6645) );
  OAI21_X1 U7783 ( .B1(n7703), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6645), .ZN(
        n6646) );
  NOR2_X1 U7784 ( .A1(n6647), .A2(n6646), .ZN(n6745) );
  AOI211_X1 U7785 ( .C1(n6647), .C2(n6646), .A(n6745), .B(n10701), .ZN(n6648)
         );
  AOI211_X1 U7786 ( .C1(n10696), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6649), .B(
        n6648), .ZN(n6650) );
  OAI21_X1 U7787 ( .B1(n6651), .B2(n10693), .A(n6650), .ZN(P1_U3253) );
  INV_X1 U7788 ( .A(n6652), .ZN(n10884) );
  NAND2_X1 U7789 ( .A1(n6531), .A2(n6529), .ZN(n6653) );
  NAND2_X1 U7790 ( .A1(n9225), .A2(n6659), .ZN(n8712) );
  NAND2_X1 U7791 ( .A1(n6657), .A2(n6708), .ZN(n6703) );
  OAI21_X1 U7792 ( .B1(n6657), .B2(n6708), .A(n6703), .ZN(n7042) );
  AND2_X1 U7793 ( .A1(n6937), .A2(n6655), .ZN(n6658) );
  NOR2_X1 U7794 ( .A1(n6937), .A2(n6655), .ZN(n6956) );
  OR2_X1 U7795 ( .A1(n6658), .A2(n6956), .ZN(n7038) );
  OAI22_X1 U7796 ( .A1(n7038), .A2(n11011), .B1(n6659), .B2(n11010), .ZN(n6665) );
  NAND2_X1 U7797 ( .A1(n8858), .A2(n6660), .ZN(n8709) );
  XNOR2_X1 U7798 ( .A(n8707), .B(n5529), .ZN(n6664) );
  INV_X1 U7799 ( .A(n7425), .ZN(n6951) );
  NAND2_X1 U7800 ( .A1(n7042), .A2(n6951), .ZN(n6663) );
  AOI22_X1 U7801 ( .A1(n9499), .A2(n6531), .B1(n9175), .B2(n9501), .ZN(n6662)
         );
  OAI211_X1 U7802 ( .C1(n6664), .C2(n9486), .A(n6663), .B(n6662), .ZN(n7039)
         );
  AOI211_X1 U7803 ( .C1(n10884), .C2(n7042), .A(n6665), .B(n7039), .ZN(n6667)
         );
  OR2_X1 U7804 ( .A1(n6667), .A2(n11017), .ZN(n6666) );
  OAI21_X1 U7805 ( .B1(n11018), .B2(n5835), .A(n6666), .ZN(P2_U3522) );
  INV_X1 U7806 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6669) );
  OR2_X1 U7807 ( .A1(n6667), .A2(n11019), .ZN(n6668) );
  OAI21_X1 U7808 ( .B1(n11001), .B2(n6669), .A(n6668), .ZN(P2_U3457) );
  INV_X1 U7809 ( .A(n6670), .ZN(n6672) );
  NAND2_X1 U7810 ( .A1(n6672), .A2(n6671), .ZN(n6673) );
  NAND2_X1 U7811 ( .A1(n10235), .A2(n9080), .ZN(n6680) );
  INV_X2 U7812 ( .A(n7011), .ZN(n8472) );
  NAND2_X1 U7813 ( .A1(n8472), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U7814 ( .A1(n8133), .A2(n6675), .ZN(n6676) );
  OAI211_X1 U7815 ( .C1(n7005), .C2(n6678), .A(n6677), .B(n6676), .ZN(n6813)
         );
  NAND2_X1 U7816 ( .A1(n6813), .A2(n7122), .ZN(n6679) );
  NAND2_X1 U7817 ( .A1(n6680), .A2(n6679), .ZN(n6681) );
  XNOR2_X1 U7818 ( .A(n6681), .B(n9083), .ZN(n6683) );
  AND2_X1 U7819 ( .A1(n6813), .A2(n9080), .ZN(n6682) );
  AOI21_X1 U7820 ( .B1(n10235), .B2(n9085), .A(n6682), .ZN(n6684) );
  INV_X1 U7821 ( .A(n6683), .ZN(n6686) );
  INV_X1 U7822 ( .A(n6684), .ZN(n6685) );
  NAND2_X1 U7823 ( .A1(n6686), .A2(n6685), .ZN(n6908) );
  NAND2_X1 U7824 ( .A1(n5144), .A2(n6908), .ZN(n6687) );
  XNOR2_X1 U7825 ( .A(n6907), .B(n6687), .ZN(n6701) );
  INV_X1 U7826 ( .A(n6824), .ZN(n6699) );
  INV_X1 U7827 ( .A(n10223), .ZN(n10206) );
  INV_X1 U7828 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6688) );
  OR2_X1 U7829 ( .A1(n6629), .A2(n10797), .ZN(n6695) );
  OR2_X1 U7830 ( .A1(n8496), .A2(n6689), .ZN(n6694) );
  INV_X1 U7831 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U7832 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6690) );
  NAND2_X1 U7833 ( .A1(n6691), .A2(n6690), .ZN(n6692) );
  NAND2_X1 U7834 ( .A1(n6925), .A2(n6692), .ZN(n10785) );
  OR2_X1 U7835 ( .A1(n8209), .A2(n10785), .ZN(n6693) );
  NAND4_X1 U7836 ( .A1(n6696), .A2(n6695), .A3(n6694), .A4(n6693), .ZN(n10803)
         );
  AOI22_X1 U7837 ( .A1(n10191), .A2(n10803), .B1(n10218), .B2(n10731), .ZN(
        n6697) );
  NAND2_X1 U7838 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n10704) );
  OAI211_X1 U7839 ( .C1(n10762), .C2(n10206), .A(n6697), .B(n10704), .ZN(n6698) );
  AOI21_X1 U7840 ( .B1(n6699), .B2(n10203), .A(n6698), .ZN(n6700) );
  OAI21_X1 U7841 ( .B1(n6701), .B2(n10226), .A(n6700), .ZN(P1_U3228) );
  OR2_X1 U7842 ( .A1(n9225), .A2(n6655), .ZN(n6702) );
  NAND2_X1 U7843 ( .A1(n6703), .A2(n6702), .ZN(n6947) );
  NAND2_X1 U7844 ( .A1(n9175), .A2(n10754), .ZN(n8717) );
  NAND2_X1 U7845 ( .A1(n6947), .A2(n6950), .ZN(n6946) );
  OR2_X1 U7846 ( .A1(n9175), .A2(n5471), .ZN(n6704) );
  NAND2_X1 U7847 ( .A1(n6946), .A2(n6704), .ZN(n6706) );
  INV_X1 U7848 ( .A(n6706), .ZN(n6705) );
  NAND2_X1 U7849 ( .A1(n6705), .A2(n8862), .ZN(n6830) );
  NAND2_X1 U7850 ( .A1(n6706), .A2(n8719), .ZN(n6707) );
  NAND2_X1 U7851 ( .A1(n6830), .A2(n6707), .ZN(n7081) );
  INV_X1 U7852 ( .A(n6950), .ZN(n8860) );
  NAND2_X1 U7853 ( .A1(n6709), .A2(n8718), .ZN(n6710) );
  INV_X1 U7854 ( .A(n8719), .ZN(n8862) );
  AOI21_X1 U7855 ( .B1(n6710), .B2(n8862), .A(n9486), .ZN(n6715) );
  INV_X1 U7856 ( .A(n6710), .ZN(n6711) );
  NAND2_X1 U7857 ( .A1(n6711), .A2(n8719), .ZN(n6833) );
  INV_X1 U7858 ( .A(n9223), .ZN(n6712) );
  OAI22_X1 U7859 ( .A1(n6713), .A2(n9466), .B1(n6712), .B2(n9468), .ZN(n6714)
         );
  AOI21_X1 U7860 ( .B1(n6715), .B2(n6833), .A(n6714), .ZN(n7084) );
  NAND2_X1 U7861 ( .A1(n6958), .A2(n9170), .ZN(n6716) );
  AND2_X1 U7862 ( .A1(n6838), .A2(n6716), .ZN(n7078) );
  AOI22_X1 U7863 ( .A1(n7078), .A2(n10927), .B1(n9170), .B2(n10925), .ZN(n6717) );
  OAI211_X1 U7864 ( .C1(n10992), .C2(n7081), .A(n7084), .B(n6717), .ZN(n6719)
         );
  NAND2_X1 U7865 ( .A1(n6719), .A2(n11001), .ZN(n6718) );
  OAI21_X1 U7866 ( .B1(n11001), .B2(n5883), .A(n6718), .ZN(P2_U3463) );
  NAND2_X1 U7867 ( .A1(n6719), .A2(n11018), .ZN(n6720) );
  OAI21_X1 U7868 ( .B1(n11018), .B2(n6299), .A(n6720), .ZN(P2_U3524) );
  OR2_X1 U7869 ( .A1(n7223), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6724) );
  INV_X1 U7870 ( .A(n6724), .ZN(n6722) );
  MUX2_X1 U7871 ( .A(n7689), .B(P2_REG2_REG_12__SCAN_IN), .S(n7601), .Z(n6721)
         );
  OAI21_X1 U7872 ( .B1(n6726), .B2(n6722), .A(n6721), .ZN(n6727) );
  MUX2_X1 U7873 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7689), .S(n7601), .Z(n6723)
         );
  NAND2_X1 U7874 ( .A1(n6724), .A2(n6723), .ZN(n6725) );
  NAND3_X1 U7875 ( .A1(n6727), .A2(n10679), .A3(n6988), .ZN(n6738) );
  INV_X1 U7876 ( .A(n10658), .ZN(n10682) );
  MUX2_X1 U7877 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6164), .S(n7601), .Z(n6733)
         );
  OAI21_X1 U7878 ( .B1(n7163), .B2(n6729), .A(n6728), .ZN(n6730) );
  INV_X1 U7879 ( .A(n6730), .ZN(n6732) );
  INV_X1 U7880 ( .A(n6995), .ZN(n6731) );
  OAI21_X1 U7881 ( .B1(n6733), .B2(n6732), .A(n6731), .ZN(n6736) );
  INV_X1 U7882 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U7883 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8384) );
  OAI21_X1 U7884 ( .B1(n9257), .B2(n6734), .A(n8384), .ZN(n6735) );
  AOI21_X1 U7885 ( .B1(n10682), .B2(n6736), .A(n6735), .ZN(n6737) );
  OAI211_X1 U7886 ( .C1(n10670), .C2(n6996), .A(n6738), .B(n6737), .ZN(
        P2_U3257) );
  INV_X1 U7887 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10990) );
  INV_X1 U7888 ( .A(n7733), .ZN(n6744) );
  NOR2_X1 U7889 ( .A1(n6744), .A2(n10990), .ZN(n6739) );
  AOI21_X1 U7890 ( .B1(n10990), .B2(n6744), .A(n6739), .ZN(n6742) );
  OAI21_X1 U7891 ( .B1(n7703), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6740), .ZN(
        n6741) );
  NAND2_X1 U7892 ( .A1(n6742), .A2(n6741), .ZN(n6855) );
  OAI21_X1 U7893 ( .B1(n6742), .B2(n6741), .A(n6855), .ZN(n6751) );
  NAND2_X1 U7894 ( .A1(n10696), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U7895 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10155) );
  OAI211_X1 U7896 ( .C1(n10692), .C2(n6744), .A(n6743), .B(n10155), .ZN(n6750)
         );
  AOI21_X1 U7897 ( .B1(n7703), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6745), .ZN(
        n6748) );
  NAND2_X1 U7898 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7733), .ZN(n6746) );
  OAI21_X1 U7899 ( .B1(n7733), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6746), .ZN(
        n6747) );
  NOR2_X1 U7900 ( .A1(n6748), .A2(n6747), .ZN(n6861) );
  AOI211_X1 U7901 ( .C1(n6748), .C2(n6747), .A(n6861), .B(n10701), .ZN(n6749)
         );
  AOI211_X1 U7902 ( .C1(n10636), .C2(n6751), .A(n6750), .B(n6749), .ZN(n6752)
         );
  INV_X1 U7903 ( .A(n6752), .ZN(P1_U3254) );
  INV_X1 U7904 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7807) );
  INV_X1 U7905 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U7906 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6758) );
  INV_X1 U7907 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10167) );
  INV_X1 U7908 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8181) );
  INV_X1 U7909 ( .A(n8207), .ZN(n6761) );
  INV_X1 U7910 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8221) );
  INV_X1 U7911 ( .A(n8235), .ZN(n6762) );
  NAND2_X1 U7912 ( .A1(n6762), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8248) );
  INV_X1 U7913 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8247) );
  INV_X1 U7914 ( .A(n8250), .ZN(n8310) );
  INV_X1 U7915 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U7916 ( .A1(n8490), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6765) );
  INV_X1 U7917 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6763) );
  OR2_X1 U7918 ( .A1(n8492), .A2(n6763), .ZN(n6764) );
  OAI211_X1 U7919 ( .C1(n8496), .C2(n6766), .A(n6765), .B(n6764), .ZN(n6767)
         );
  AOI21_X1 U7920 ( .B1(n8310), .B2(n8254), .A(n6767), .ZN(n9094) );
  INV_X2 U7921 ( .A(P1_U4006), .ZN(n10236) );
  NAND2_X1 U7922 ( .A1(n10236), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6768) );
  OAI21_X1 U7923 ( .B1(n9094), .B2(n10236), .A(n6768), .ZN(P1_U3584) );
  NAND2_X1 U7924 ( .A1(n6772), .A2(SI_14_), .ZN(n6773) );
  INV_X1 U7925 ( .A(n6776), .ZN(n6774) );
  XNOR2_X1 U7926 ( .A(n6785), .B(SI_15_), .ZN(n7846) );
  INV_X1 U7927 ( .A(n7846), .ZN(n6783) );
  NAND2_X1 U7928 ( .A1(n6778), .A2(n9729), .ZN(n6779) );
  NAND2_X1 U7929 ( .A1(n6779), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6780) );
  XNOR2_X1 U7930 ( .A(n6780), .B(n5746), .ZN(n7847) );
  OAI222_X1 U7931 ( .A1(n10532), .A2(n6783), .B1(n7847), .B2(P1_U3084), .C1(
        n9908), .C2(n10528), .ZN(P1_U3338) );
  NAND2_X1 U7932 ( .A1(n6781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6782) );
  XNOR2_X1 U7933 ( .A(n6782), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7626) );
  INV_X1 U7934 ( .A(n7626), .ZN(n7385) );
  OAI222_X1 U7935 ( .A1(n10047), .A2(n6784), .B1(n6076), .B2(n6783), .C1(n7385), .C2(P2_U3152), .ZN(P2_U3343) );
  INV_X1 U7936 ( .A(SI_16_), .ZN(n6787) );
  NAND2_X1 U7937 ( .A1(n6788), .A2(n6787), .ZN(n6850) );
  INV_X1 U7938 ( .A(n6788), .ZN(n6789) );
  NAND2_X1 U7939 ( .A1(n6789), .A2(SI_16_), .ZN(n6790) );
  XNOR2_X1 U7940 ( .A(n6849), .B(n6848), .ZN(n8102) );
  INV_X1 U7941 ( .A(n8102), .ZN(n6847) );
  NAND2_X1 U7942 ( .A1(n6792), .A2(n6791), .ZN(n6793) );
  OAI21_X1 U7943 ( .B1(n6794), .B2(n6793), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6795) );
  MUX2_X1 U7944 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6795), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6797) );
  AND2_X1 U7945 ( .A1(n6797), .A2(n6796), .ZN(n7640) );
  AOI22_X1 U7946 ( .A1(n7640), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n7799), .ZN(n6798) );
  OAI21_X1 U7947 ( .B1(n6847), .B2(n10053), .A(n6798), .ZN(P2_U3342) );
  INV_X1 U7948 ( .A(n6799), .ZN(n6802) );
  AND2_X1 U7949 ( .A1(n10522), .A2(n6800), .ZN(n6801) );
  NAND2_X1 U7950 ( .A1(n6802), .A2(n6801), .ZN(n6822) );
  AND2_X1 U7951 ( .A1(n8678), .A2(n9076), .ZN(n10794) );
  NAND2_X1 U7952 ( .A1(n6803), .A2(n5363), .ZN(n8293) );
  NAND2_X1 U7953 ( .A1(n6816), .A2(n8293), .ZN(n6806) );
  NAND2_X1 U7954 ( .A1(n5056), .A2(n10720), .ZN(n6805) );
  NAND2_X1 U7955 ( .A1(n6806), .A2(n6805), .ZN(n10725) );
  NAND2_X1 U7956 ( .A1(n6808), .A2(n10178), .ZN(n8396) );
  NAND2_X1 U7957 ( .A1(n6807), .A2(n10728), .ZN(n8400) );
  NAND2_X1 U7958 ( .A1(n8396), .A2(n8400), .ZN(n10729) );
  NAND2_X1 U7959 ( .A1(n10725), .A2(n10729), .ZN(n6810) );
  NAND2_X1 U7960 ( .A1(n6808), .A2(n10728), .ZN(n6809) );
  NAND2_X1 U7961 ( .A1(n6810), .A2(n6809), .ZN(n6896) );
  INV_X1 U7962 ( .A(n8406), .ZN(n10749) );
  NAND2_X1 U7963 ( .A1(n6896), .A2(n6819), .ZN(n6812) );
  INV_X1 U7964 ( .A(n10731), .ZN(n8407) );
  NAND2_X1 U7965 ( .A1(n8407), .A2(n10749), .ZN(n6811) );
  NAND2_X1 U7966 ( .A1(n6812), .A2(n6811), .ZN(n7194) );
  NAND2_X1 U7967 ( .A1(n10778), .A2(n6813), .ZN(n8408) );
  NAND2_X1 U7968 ( .A1(n10235), .A2(n10762), .ZN(n8404) );
  NAND2_X1 U7969 ( .A1(n8408), .A2(n8404), .ZN(n7193) );
  INV_X1 U7970 ( .A(n7193), .ZN(n8640) );
  XNOR2_X1 U7971 ( .A(n7194), .B(n8640), .ZN(n10763) );
  OR2_X1 U7972 ( .A1(n8619), .A2(n10359), .ZN(n6815) );
  OR2_X1 U7973 ( .A1(n8667), .A2(n10708), .ZN(n6814) );
  NAND2_X1 U7974 ( .A1(n5056), .A2(n8300), .ZN(n6817) );
  INV_X1 U7975 ( .A(n10729), .ZN(n8642) );
  NAND2_X1 U7976 ( .A1(n10730), .A2(n8642), .ZN(n6818) );
  NAND2_X1 U7977 ( .A1(n6818), .A2(n8396), .ZN(n6897) );
  INV_X1 U7978 ( .A(n6819), .ZN(n8639) );
  NAND2_X1 U7979 ( .A1(n6897), .A2(n8639), .ZN(n6820) );
  NAND2_X1 U7980 ( .A1(n8407), .A2(n8406), .ZN(n8401) );
  XNOR2_X1 U7981 ( .A(n7204), .B(n8640), .ZN(n6821) );
  AOI222_X1 U7982 ( .A1(n11035), .A2(n6821), .B1(n10803), .B2(n11037), .C1(
        n10731), .C2(n11040), .ZN(n10761) );
  MUX2_X1 U7983 ( .A(n6223), .B(n10761), .S(n10795), .Z(n6828) );
  NAND2_X1 U7984 ( .A1(n6901), .A2(n10762), .ZN(n10771) );
  OAI211_X1 U7985 ( .C1(n6901), .C2(n10762), .A(n10771), .B(n10953), .ZN(
        n10760) );
  INV_X1 U7986 ( .A(n10760), .ZN(n6826) );
  INV_X1 U7987 ( .A(n11063), .ZN(n10291) );
  OAI22_X1 U7988 ( .A1(n10430), .A2(n10762), .B1(n10786), .B2(n6824), .ZN(
        n6825) );
  AOI21_X1 U7989 ( .B1(n6826), .B2(n10291), .A(n6825), .ZN(n6827) );
  OAI211_X1 U7990 ( .C1(n11064), .C2(n10763), .A(n6828), .B(n6827), .ZN(
        P1_U3287) );
  INV_X1 U7991 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U7992 ( .A1(n9224), .A2(n9170), .ZN(n6829) );
  OR2_X1 U7993 ( .A1(n9223), .A2(n6881), .ZN(n8730) );
  NAND2_X1 U7994 ( .A1(n9223), .A2(n6881), .ZN(n8729) );
  NAND2_X1 U7995 ( .A1(n8730), .A2(n8729), .ZN(n8861) );
  INV_X1 U7996 ( .A(n9170), .ZN(n6831) );
  NAND2_X1 U7997 ( .A1(n9224), .A2(n6831), .ZN(n6832) );
  NAND2_X1 U7998 ( .A1(n6833), .A2(n6832), .ZN(n6966) );
  XNOR2_X1 U7999 ( .A(n6966), .B(n8861), .ZN(n6836) );
  OR2_X1 U8000 ( .A1(n7085), .A2(n9468), .ZN(n6835) );
  NAND2_X1 U8001 ( .A1(n9224), .A2(n9499), .ZN(n6834) );
  NAND2_X1 U8002 ( .A1(n6835), .A2(n6834), .ZN(n8957) );
  AOI21_X1 U8003 ( .B1(n6836), .B2(n10923), .A(n8957), .ZN(n6873) );
  INV_X1 U8004 ( .A(n7094), .ZN(n6837) );
  AOI211_X1 U8005 ( .C1(n8965), .C2(n6838), .A(n11011), .B(n6837), .ZN(n6871)
         );
  AOI21_X1 U8006 ( .B1(n8965), .B2(n10925), .A(n6871), .ZN(n6839) );
  OAI211_X1 U8007 ( .C1(n5074), .C2(n10992), .A(n6873), .B(n6839), .ZN(n6842)
         );
  NAND2_X1 U8008 ( .A1(n6842), .A2(n11001), .ZN(n6840) );
  OAI21_X1 U8009 ( .B1(n11001), .B2(n6841), .A(n6840), .ZN(P2_U3466) );
  NAND2_X1 U8010 ( .A1(n6842), .A2(n11018), .ZN(n6843) );
  OAI21_X1 U8011 ( .B1(n11018), .B2(n5905), .A(n6843), .ZN(P2_U3525) );
  NAND2_X1 U8012 ( .A1(n6852), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6845) );
  XNOR2_X1 U8013 ( .A(n6845), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8103) );
  INV_X1 U8014 ( .A(n8103), .ZN(n7411) );
  OAI222_X1 U8015 ( .A1(n10532), .A2(n6847), .B1(n7411), .B2(P1_U3084), .C1(
        n6846), .C2(n10528), .ZN(P1_U3337) );
  MUX2_X1 U8016 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7833), .Z(n6977) );
  XNOR2_X1 U8017 ( .A(n6977), .B(n9579), .ZN(n6976) );
  XNOR2_X1 U8018 ( .A(n6979), .B(n6976), .ZN(n8107) );
  INV_X1 U8019 ( .A(n8107), .ZN(n6885) );
  OAI21_X1 U8020 ( .B1(n6852), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6982) );
  XNOR2_X1 U8021 ( .A(n6982), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U8022 ( .A1(n10246), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10525), .ZN(n6853) );
  OAI21_X1 U8023 ( .B1(n6885), .B2(n10532), .A(n6853), .ZN(P1_U3336) );
  INV_X1 U8024 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11006) );
  INV_X1 U8025 ( .A(n7802), .ZN(n6860) );
  NOR2_X1 U8026 ( .A1(n6860), .A2(n11006), .ZN(n6854) );
  AOI21_X1 U8027 ( .B1(n11006), .B2(n6860), .A(n6854), .ZN(n6857) );
  OAI21_X1 U8028 ( .B1(n7733), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6855), .ZN(
        n6856) );
  NAND2_X1 U8029 ( .A1(n6857), .A2(n6856), .ZN(n7215) );
  OAI21_X1 U8030 ( .B1(n6857), .B2(n6856), .A(n7215), .ZN(n6867) );
  NAND2_X1 U8031 ( .A1(n10696), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n6859) );
  INV_X1 U8032 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7741) );
  NOR2_X1 U8033 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7741), .ZN(n10070) );
  INV_X1 U8034 ( .A(n10070), .ZN(n6858) );
  OAI211_X1 U8035 ( .C1(n10692), .C2(n6860), .A(n6859), .B(n6858), .ZN(n6866)
         );
  AOI21_X1 U8036 ( .B1(n7733), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6861), .ZN(
        n6864) );
  NAND2_X1 U8037 ( .A1(n7802), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6862) );
  OAI21_X1 U8038 ( .B1(n7802), .B2(P1_REG2_REG_14__SCAN_IN), .A(n6862), .ZN(
        n6863) );
  NOR2_X1 U8039 ( .A1(n6864), .A2(n6863), .ZN(n7217) );
  AOI211_X1 U8040 ( .C1(n6864), .C2(n6863), .A(n7217), .B(n10701), .ZN(n6865)
         );
  AOI211_X1 U8041 ( .C1(n10636), .C2(n6867), .A(n6866), .B(n6865), .ZN(n6868)
         );
  INV_X1 U8042 ( .A(n6868), .ZN(P1_U3255) );
  INV_X1 U8043 ( .A(n6869), .ZN(n6870) );
  NAND2_X1 U8044 ( .A1(n6871), .A2(n8884), .ZN(n6872) );
  OAI211_X1 U8045 ( .C1(n10935), .C2(n8960), .A(n6873), .B(n6872), .ZN(n6878)
         );
  AND2_X1 U8046 ( .A1(n6875), .A2(n6874), .ZN(n6876) );
  MUX2_X1 U8047 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6878), .S(n10946), .Z(n6883)
         );
  OR2_X1 U8048 ( .A1(n6879), .A2(n8884), .ZN(n6948) );
  NAND2_X1 U8049 ( .A1(n7425), .A2(n6948), .ZN(n10944) );
  INV_X1 U8050 ( .A(n6880), .ZN(n10938) );
  OAI22_X1 U8051 ( .A1(n5074), .A2(n9509), .B1(n6881), .B2(n9495), .ZN(n6882)
         );
  OR2_X1 U8052 ( .A1(n6883), .A2(n6882), .ZN(P2_U3291) );
  INV_X1 U8053 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6886) );
  NAND2_X1 U8054 ( .A1(n6796), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6884) );
  XNOR2_X1 U8055 ( .A(n6884), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9244) );
  INV_X1 U8056 ( .A(n9244), .ZN(n9249) );
  OAI222_X1 U8057 ( .A1(n9110), .A2(n6886), .B1(n6076), .B2(n6885), .C1(n9249), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  AND2_X1 U8058 ( .A1(n6887), .A2(n8858), .ZN(n6888) );
  OAI22_X1 U8059 ( .A1(n6888), .A2(n9486), .B1(n6530), .B2(n9468), .ZN(n10714)
         );
  INV_X1 U8060 ( .A(n10714), .ZN(n6895) );
  INV_X1 U8061 ( .A(n10946), .ZN(n9426) );
  INV_X1 U8062 ( .A(n6888), .ZN(n10715) );
  INV_X1 U8063 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6891) );
  OAI22_X1 U8064 ( .A1(n10946), .A2(n6891), .B1(n6890), .B2(n10935), .ZN(n6892) );
  AOI211_X1 U8065 ( .C1(n10715), .C2(n9400), .A(n6893), .B(n6892), .ZN(n6894)
         );
  OAI21_X1 U8066 ( .B1(n6895), .B2(n9426), .A(n6894), .ZN(P2_U3296) );
  XNOR2_X1 U8067 ( .A(n6896), .B(n8639), .ZN(n10750) );
  XNOR2_X1 U8068 ( .A(n6897), .B(n8639), .ZN(n6898) );
  AOI222_X1 U8069 ( .A1(n11035), .A2(n6898), .B1(n8295), .B2(n11040), .C1(
        n10235), .C2(n11037), .ZN(n10748) );
  INV_X2 U8070 ( .A(n10795), .ZN(n11070) );
  OR2_X1 U8071 ( .A1(n10748), .A2(n11070), .ZN(n6906) );
  OAI22_X1 U8072 ( .A1(n10795), .A2(n6572), .B1(n10786), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U8073 ( .A1(n10727), .A2(n8406), .ZN(n6900) );
  NAND2_X1 U8074 ( .A1(n6900), .A2(n10953), .ZN(n6902) );
  OR2_X1 U8075 ( .A1(n6902), .A2(n6901), .ZN(n10747) );
  NOR2_X1 U8076 ( .A1(n10747), .A2(n11063), .ZN(n6903) );
  AOI211_X1 U8077 ( .C1(n11060), .C2(n8406), .A(n6904), .B(n6903), .ZN(n6905)
         );
  OAI211_X1 U8078 ( .C1(n11064), .C2(n10750), .A(n6906), .B(n6905), .ZN(
        P1_U3288) );
  NAND2_X1 U8079 ( .A1(n10803), .A2(n9080), .ZN(n6914) );
  NAND2_X1 U8080 ( .A1(n8472), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U8081 ( .A1(n8133), .A2(n6909), .ZN(n6910) );
  NAND2_X1 U8082 ( .A1(n10784), .A2(n7122), .ZN(n6913) );
  NAND2_X1 U8083 ( .A1(n6914), .A2(n6913), .ZN(n6915) );
  XNOR2_X1 U8084 ( .A(n6915), .B(n9083), .ZN(n6917) );
  NAND2_X1 U8085 ( .A1(n6916), .A2(n6917), .ZN(n7017) );
  INV_X1 U8086 ( .A(n6916), .ZN(n6919) );
  INV_X1 U8087 ( .A(n6917), .ZN(n6918) );
  NAND2_X1 U8088 ( .A1(n7017), .A2(n7018), .ZN(n6922) );
  NAND2_X1 U8089 ( .A1(n10803), .A2(n9085), .ZN(n6921) );
  NAND2_X1 U8090 ( .A1(n10784), .A2(n9080), .ZN(n6920) );
  NAND2_X1 U8091 ( .A1(n6921), .A2(n6920), .ZN(n7016) );
  XNOR2_X1 U8092 ( .A(n6922), .B(n7016), .ZN(n6923) );
  NAND2_X1 U8093 ( .A1(n6923), .A2(n10197), .ZN(n6935) );
  NAND2_X1 U8094 ( .A1(n8490), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6931) );
  OR2_X1 U8095 ( .A1(n8496), .A2(n6924), .ZN(n6930) );
  INV_X1 U8096 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7031) );
  NAND2_X1 U8097 ( .A1(n6925), .A2(n7031), .ZN(n6926) );
  NAND2_X1 U8098 ( .A1(n7024), .A2(n6926), .ZN(n10812) );
  OR2_X1 U8099 ( .A1(n6203), .A2(n10812), .ZN(n6929) );
  INV_X1 U8100 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6927) );
  OR2_X1 U8101 ( .A1(n8492), .A2(n6927), .ZN(n6928) );
  NAND4_X1 U8102 ( .A1(n6931), .A2(n6930), .A3(n6929), .A4(n6928), .ZN(n10234)
         );
  INV_X1 U8103 ( .A(n10234), .ZN(n10780) );
  OAI22_X1 U8104 ( .A1(n10126), .A2(n10778), .B1(n10780), .B2(n10215), .ZN(
        n6932) );
  AOI211_X1 U8105 ( .C1(n10784), .C2(n10223), .A(n6933), .B(n6932), .ZN(n6934)
         );
  OAI211_X1 U8106 ( .C1(n10221), .C2(n10785), .A(n6935), .B(n6934), .ZN(
        P1_U3225) );
  OAI22_X1 U8107 ( .A1(n10946), .A2(n5986), .B1(n6936), .B2(n10935), .ZN(n6941) );
  INV_X1 U8108 ( .A(n6937), .ZN(n6938) );
  NOR3_X1 U8109 ( .A1(n6939), .A2(n6938), .A3(n9309), .ZN(n6940) );
  AOI211_X1 U8110 ( .C1(n9427), .C2(n6529), .A(n6941), .B(n6940), .ZN(n6944)
         );
  OR2_X1 U8111 ( .A1(n6942), .A2(n9509), .ZN(n6943) );
  OAI211_X1 U8112 ( .C1(n6945), .C2(n9504), .A(n6944), .B(n6943), .ZN(P2_U3295) );
  OAI21_X1 U8113 ( .B1(n6947), .B2(n6950), .A(n6946), .ZN(n10758) );
  INV_X1 U8114 ( .A(n10758), .ZN(n6963) );
  OR2_X1 U8115 ( .A1(n9426), .A2(n6948), .ZN(n7431) );
  XNOR2_X1 U8116 ( .A(n6950), .B(n6949), .ZN(n6954) );
  AOI22_X1 U8117 ( .A1(n9499), .A2(n9225), .B1(n9224), .B2(n9501), .ZN(n6953)
         );
  NAND2_X1 U8118 ( .A1(n10758), .A2(n6951), .ZN(n6952) );
  OAI211_X1 U8119 ( .C1(n6954), .C2(n9486), .A(n6953), .B(n6952), .ZN(n10756)
         );
  NAND2_X1 U8120 ( .A1(n10756), .A2(n10946), .ZN(n6962) );
  OAI22_X1 U8121 ( .A1(n10946), .A2(n6955), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10935), .ZN(n6960) );
  OR2_X1 U8122 ( .A1(n6956), .A2(n10754), .ZN(n6957) );
  NAND2_X1 U8123 ( .A1(n6958), .A2(n6957), .ZN(n10755) );
  NOR2_X1 U8124 ( .A1(n10755), .A2(n9309), .ZN(n6959) );
  AOI211_X1 U8125 ( .C1(n9427), .C2(n5471), .A(n6960), .B(n6959), .ZN(n6961)
         );
  OAI211_X1 U8126 ( .C1(n6963), .C2(n7431), .A(n6962), .B(n6961), .ZN(P2_U3293) );
  OR2_X1 U8127 ( .A1(n9223), .A2(n8965), .ZN(n6964) );
  NAND2_X1 U8128 ( .A1(n6965), .A2(n6964), .ZN(n7087) );
  INV_X1 U8129 ( .A(n7085), .ZN(n9222) );
  NAND2_X1 U8130 ( .A1(n9222), .A2(n7086), .ZN(n7090) );
  INV_X1 U8131 ( .A(n7090), .ZN(n8733) );
  OR2_X1 U8132 ( .A1(n8734), .A2(n8733), .ZN(n6967) );
  XNOR2_X1 U8133 ( .A(n7087), .B(n6967), .ZN(n7051) );
  INV_X1 U8134 ( .A(n7086), .ZN(n8363) );
  XNOR2_X1 U8135 ( .A(n7094), .B(n8363), .ZN(n7047) );
  OAI22_X1 U8136 ( .A1(n7047), .A2(n11011), .B1(n7086), .B2(n11010), .ZN(n6971) );
  INV_X1 U8137 ( .A(n6967), .ZN(n8865) );
  XNOR2_X1 U8138 ( .A(n7091), .B(n8865), .ZN(n6968) );
  NAND2_X1 U8139 ( .A1(n6968), .A2(n10923), .ZN(n6970) );
  AOI22_X1 U8140 ( .A1(n9499), .A2(n9223), .B1(n9221), .B2(n9501), .ZN(n6969)
         );
  NAND2_X1 U8141 ( .A1(n6970), .A2(n6969), .ZN(n7048) );
  AOI211_X1 U8142 ( .C1(n11015), .C2(n7051), .A(n6971), .B(n7048), .ZN(n6973)
         );
  OR2_X1 U8143 ( .A1(n6973), .A2(n11017), .ZN(n6972) );
  OAI21_X1 U8144 ( .B1(n11018), .B2(n5921), .A(n6972), .ZN(P2_U3526) );
  INV_X1 U8145 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6975) );
  OR2_X1 U8146 ( .A1(n6973), .A2(n11019), .ZN(n6974) );
  OAI21_X1 U8147 ( .B1(n11001), .B2(n6975), .A(n6974), .ZN(P2_U3469) );
  NAND2_X1 U8148 ( .A1(n6977), .A2(SI_17_), .ZN(n6978) );
  MUX2_X1 U8149 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7833), .Z(n7187) );
  XNOR2_X1 U8150 ( .A(n7187), .B(SI_18_), .ZN(n7184) );
  XNOR2_X1 U8151 ( .A(n7186), .B(n7184), .ZN(n8119) );
  INV_X1 U8152 ( .A(n8119), .ZN(n6986) );
  XNOR2_X1 U8153 ( .A(n6980), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9262) );
  AOI22_X1 U8154 ( .A1(n9262), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7799), .ZN(n6981) );
  OAI21_X1 U8155 ( .B1(n6986), .B2(n10053), .A(n6981), .ZN(P2_U3340) );
  NAND2_X1 U8156 ( .A1(n6982), .A2(n9734), .ZN(n6983) );
  NAND2_X1 U8157 ( .A1(n6983), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6984) );
  XNOR2_X1 U8158 ( .A(n6984), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U8159 ( .A1(n10259), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10525), .ZN(n6985) );
  OAI21_X1 U8160 ( .B1(n6986), .B2(n10532), .A(n6985), .ZN(P1_U3335) );
  NAND2_X1 U8161 ( .A1(n7601), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6987) );
  NAND2_X1 U8162 ( .A1(n6988), .A2(n6987), .ZN(n10669) );
  INV_X1 U8163 ( .A(n10669), .ZN(n10677) );
  NOR2_X1 U8164 ( .A1(n10677), .A2(n10675), .ZN(n6989) );
  OAI22_X1 U8165 ( .A1(n6989), .A2(n7608), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10669), .ZN(n10680) );
  INV_X1 U8166 ( .A(n10680), .ZN(n6994) );
  INV_X1 U8167 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6990) );
  MUX2_X1 U8168 ( .A(n6990), .B(P2_REG2_REG_14__SCAN_IN), .S(n7613), .Z(n6993)
         );
  INV_X1 U8169 ( .A(n6993), .ZN(n6991) );
  NAND2_X1 U8170 ( .A1(n10680), .A2(n6991), .ZN(n7252) );
  INV_X1 U8171 ( .A(n7252), .ZN(n6992) );
  AOI21_X1 U8172 ( .B1(n6994), .B2(n6993), .A(n6992), .ZN(n7004) );
  INV_X1 U8173 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7001) );
  AOI21_X1 U8174 ( .B1(n6164), .B2(n6996), .A(n6995), .ZN(n10684) );
  MUX2_X1 U8175 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n6997), .S(n7608), .Z(n10683) );
  NAND2_X1 U8176 ( .A1(n10684), .A2(n10683), .ZN(n10681) );
  OAI21_X1 U8177 ( .B1(n6997), .B2(n10676), .A(n10681), .ZN(n6999) );
  INV_X1 U8178 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7619) );
  MUX2_X1 U8179 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7619), .S(n7613), .Z(n6998)
         );
  NAND2_X1 U8180 ( .A1(n6998), .A2(n6999), .ZN(n7244) );
  OAI211_X1 U8181 ( .C1(n6999), .C2(n6998), .A(n10682), .B(n7244), .ZN(n7000)
         );
  NAND2_X1 U8182 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8968) );
  OAI211_X1 U8183 ( .C1(n9257), .C2(n7001), .A(n7000), .B(n8968), .ZN(n7002)
         );
  AOI21_X1 U8184 ( .B1(n7613), .B2(n10660), .A(n7002), .ZN(n7003) );
  OAI21_X1 U8185 ( .B1(n7004), .B2(n9278), .A(n7003), .ZN(P2_U3259) );
  NAND2_X1 U8186 ( .A1(n10234), .A2(n9080), .ZN(n7013) );
  NAND2_X1 U8187 ( .A1(n8487), .A2(n7006), .ZN(n7009) );
  NAND2_X1 U8188 ( .A1(n8133), .A2(n7007), .ZN(n7008) );
  OAI211_X1 U8189 ( .C1(n7011), .C2(n7010), .A(n7009), .B(n7008), .ZN(n10814)
         );
  NAND2_X1 U8190 ( .A1(n10814), .A2(n7122), .ZN(n7012) );
  NAND2_X1 U8191 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  XNOR2_X1 U8192 ( .A(n7014), .B(n9083), .ZN(n7127) );
  AND2_X1 U8193 ( .A1(n10814), .A2(n9080), .ZN(n7015) );
  AOI21_X1 U8194 ( .B1(n10234), .B2(n9085), .A(n7015), .ZN(n7126) );
  XNOR2_X1 U8195 ( .A(n7127), .B(n7126), .ZN(n7022) );
  INV_X1 U8196 ( .A(n7129), .ZN(n7021) );
  AOI21_X1 U8197 ( .B1(n7022), .B2(n7019), .A(n7021), .ZN(n7036) );
  NAND2_X1 U8198 ( .A1(n8238), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7030) );
  OR2_X1 U8199 ( .A1(n8496), .A2(n10827), .ZN(n7029) );
  OR2_X1 U8200 ( .A1(n6629), .A2(n6242), .ZN(n7028) );
  INV_X1 U8201 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7023) );
  NAND2_X1 U8202 ( .A1(n7024), .A2(n7023), .ZN(n7025) );
  NAND2_X1 U8203 ( .A1(n7026), .A2(n7025), .ZN(n7208) );
  OR2_X1 U8204 ( .A1(n8209), .A2(n7208), .ZN(n7027) );
  NAND4_X1 U8205 ( .A1(n7030), .A2(n7029), .A3(n7028), .A4(n7027), .ZN(n10848)
         );
  INV_X1 U8206 ( .A(n10848), .ZN(n7325) );
  NOR2_X1 U8207 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7031), .ZN(n10590) );
  AOI21_X1 U8208 ( .B1(n10218), .B2(n10803), .A(n10590), .ZN(n7032) );
  OAI21_X1 U8209 ( .B1(n7325), .B2(n10215), .A(n7032), .ZN(n7034) );
  NOR2_X1 U8210 ( .A1(n10221), .A2(n10812), .ZN(n7033) );
  AOI211_X1 U8211 ( .C1(n10814), .C2(n10223), .A(n7034), .B(n7033), .ZN(n7035)
         );
  OAI21_X1 U8212 ( .B1(n7036), .B2(n10226), .A(n7035), .ZN(P1_U3237) );
  INV_X1 U8213 ( .A(n7431), .ZN(n7043) );
  INV_X1 U8214 ( .A(n10935), .ZN(n9492) );
  AOI22_X1 U8215 ( .A1(n9427), .A2(n6655), .B1(n9492), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7037) );
  OAI21_X1 U8216 ( .B1(n7038), .B2(n9309), .A(n7037), .ZN(n7041) );
  MUX2_X1 U8217 ( .A(n7039), .B(P2_REG2_REG_2__SCAN_IN), .S(n9426), .Z(n7040)
         );
  AOI211_X1 U8218 ( .C1(n7043), .C2(n7042), .A(n7041), .B(n7040), .ZN(n7044)
         );
  INV_X1 U8219 ( .A(n7044), .ZN(P2_U3294) );
  INV_X1 U8220 ( .A(n7045), .ZN(n8353) );
  AOI22_X1 U8221 ( .A1(n9427), .A2(n8363), .B1(n8353), .B2(n9492), .ZN(n7046)
         );
  OAI21_X1 U8222 ( .B1(n7047), .B2(n9309), .A(n7046), .ZN(n7050) );
  MUX2_X1 U8223 ( .A(n7048), .B(P2_REG2_REG_6__SCAN_IN), .S(n9426), .Z(n7049)
         );
  AOI211_X1 U8224 ( .C1(n9400), .C2(n7051), .A(n7050), .B(n7049), .ZN(n7052)
         );
  INV_X1 U8225 ( .A(n7052), .ZN(P2_U3290) );
  NAND2_X1 U8226 ( .A1(n7270), .A2(n8693), .ZN(n7055) );
  AOI22_X1 U8227 ( .A1(n8685), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5856), .B2(
        n7053), .ZN(n7054) );
  OR2_X1 U8228 ( .A1(n7461), .A2(n9468), .ZN(n7057) );
  NAND2_X1 U8229 ( .A1(n9221), .A2(n9499), .ZN(n7056) );
  AND2_X1 U8230 ( .A1(n7057), .A2(n7056), .ZN(n7102) );
  INV_X1 U8231 ( .A(n9208), .ZN(n9148) );
  INV_X1 U8232 ( .A(n7104), .ZN(n7059) );
  AOI21_X1 U8233 ( .B1(n9188), .B2(n7059), .A(n7058), .ZN(n7060) );
  OAI21_X1 U8234 ( .B1(n7102), .B2(n9148), .A(n7060), .ZN(n7074) );
  NAND3_X1 U8235 ( .A1(n7061), .A2(n9128), .A3(n9221), .ZN(n7072) );
  XNOR2_X1 U8236 ( .A(n10872), .B(n5877), .ZN(n7062) );
  AND2_X1 U8237 ( .A1(n9220), .A2(n8927), .ZN(n7063) );
  NAND2_X1 U8238 ( .A1(n7062), .A2(n7063), .ZN(n7145) );
  INV_X1 U8239 ( .A(n7062), .ZN(n7172) );
  INV_X1 U8240 ( .A(n7063), .ZN(n7064) );
  NAND2_X1 U8241 ( .A1(n7172), .A2(n7064), .ZN(n7065) );
  AND2_X1 U8242 ( .A1(n7145), .A2(n7065), .ZN(n7069) );
  OAI21_X1 U8243 ( .B1(n7066), .B2(n7069), .A(n9167), .ZN(n7071) );
  INV_X1 U8244 ( .A(n7147), .ZN(n7174) );
  AOI21_X1 U8245 ( .B1(n7072), .B2(n7071), .A(n7174), .ZN(n7073) );
  AOI211_X1 U8246 ( .C1(n9171), .C2(n7415), .A(n7074), .B(n7073), .ZN(n7075)
         );
  INV_X1 U8247 ( .A(n7075), .ZN(P2_U3223) );
  OAI22_X1 U8248 ( .A1(n10946), .A2(n7076), .B1(n9169), .B2(n10935), .ZN(n7077) );
  AOI21_X1 U8249 ( .B1(n9427), .B2(n9170), .A(n7077), .ZN(n7080) );
  NAND2_X1 U8250 ( .A1(n7078), .A2(n9507), .ZN(n7079) );
  OAI211_X1 U8251 ( .C1(n7081), .C2(n9509), .A(n7080), .B(n7079), .ZN(n7082)
         );
  INV_X1 U8252 ( .A(n7082), .ZN(n7083) );
  OAI21_X1 U8253 ( .B1(n7084), .B2(n9426), .A(n7083), .ZN(P2_U3292) );
  OAI21_X1 U8254 ( .B1(n7087), .B2(n7086), .A(n7085), .ZN(n7089) );
  NAND2_X1 U8255 ( .A1(n7087), .A2(n7086), .ZN(n7088) );
  NAND2_X1 U8256 ( .A1(n9221), .A2(n7111), .ZN(n8738) );
  XNOR2_X1 U8257 ( .A(n7110), .B(n5521), .ZN(n10834) );
  XNOR2_X1 U8258 ( .A(n7101), .B(n8735), .ZN(n7092) );
  AOI222_X1 U8259 ( .A1(n10923), .A2(n7092), .B1(n9220), .B2(n9501), .C1(n9222), .C2(n9499), .ZN(n10833) );
  MUX2_X1 U8260 ( .A(n7093), .B(n10833), .S(n10946), .Z(n7100) );
  OR2_X1 U8261 ( .A1(n7095), .A2(n7111), .ZN(n7096) );
  NAND2_X1 U8262 ( .A1(n7095), .A2(n7111), .ZN(n7105) );
  AND2_X1 U8263 ( .A1(n7096), .A2(n7105), .ZN(n10831) );
  OAI22_X1 U8264 ( .A1(n9495), .A2(n7111), .B1(n10935), .B2(n7097), .ZN(n7098)
         );
  AOI21_X1 U8265 ( .B1(n10831), .B2(n9507), .A(n7098), .ZN(n7099) );
  OAI211_X1 U8266 ( .C1(n10834), .C2(n9509), .A(n7100), .B(n7099), .ZN(
        P2_U3289) );
  NAND2_X1 U8267 ( .A1(n9220), .A2(n10872), .ZN(n8742) );
  XOR2_X1 U8268 ( .A(n8866), .B(n7421), .Z(n7103) );
  OAI21_X1 U8269 ( .B1(n7103), .B2(n9486), .A(n7102), .ZN(n10874) );
  INV_X1 U8270 ( .A(n10874), .ZN(n7116) );
  OAI22_X1 U8271 ( .A1(n10946), .A2(n6330), .B1(n7104), .B2(n10935), .ZN(n7109) );
  INV_X1 U8272 ( .A(n7105), .ZN(n7106) );
  OR2_X2 U8273 ( .A1(n7105), .A2(n7415), .ZN(n7456) );
  OAI211_X1 U8274 ( .C1(n7106), .C2(n10872), .A(n10927), .B(n7456), .ZN(n10870) );
  AND2_X1 U8275 ( .A1(n10946), .A2(n8884), .ZN(n9481) );
  INV_X1 U8276 ( .A(n9481), .ZN(n7107) );
  NOR2_X1 U8277 ( .A1(n10870), .A2(n7107), .ZN(n7108) );
  AOI211_X1 U8278 ( .C1(n9427), .C2(n7415), .A(n7109), .B(n7108), .ZN(n7115)
         );
  INV_X1 U8279 ( .A(n7111), .ZN(n10830) );
  OR2_X1 U8280 ( .A1(n9221), .A2(n10830), .ZN(n7112) );
  NAND2_X1 U8281 ( .A1(n7113), .A2(n8866), .ZN(n10868) );
  NAND3_X1 U8282 ( .A1(n10869), .A2(n10868), .A3(n9400), .ZN(n7114) );
  OAI211_X1 U8283 ( .C1(n7116), .C2(n9504), .A(n7115), .B(n7114), .ZN(P2_U3288) );
  AOI22_X1 U8284 ( .A1(n8472), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8133), .B2(
        n7118), .ZN(n7121) );
  NAND2_X1 U8285 ( .A1(n7119), .A2(n8487), .ZN(n7120) );
  NAND2_X1 U8286 ( .A1(n7121), .A2(n7120), .ZN(n7212) );
  NAND2_X1 U8287 ( .A1(n10848), .A2(n9080), .ZN(n7124) );
  NAND2_X1 U8288 ( .A1(n7212), .A2(n7122), .ZN(n7123) );
  NAND2_X1 U8289 ( .A1(n7124), .A2(n7123), .ZN(n7125) );
  XNOR2_X1 U8290 ( .A(n7125), .B(n9076), .ZN(n7277) );
  AOI22_X1 U8291 ( .A1(n10848), .A2(n9085), .B1(n7212), .B2(n9080), .ZN(n7278)
         );
  XNOR2_X1 U8292 ( .A(n7277), .B(n7278), .ZN(n7131) );
  NAND2_X1 U8293 ( .A1(n7127), .A2(n7126), .ZN(n7128) );
  NAND2_X1 U8294 ( .A1(n7129), .A2(n7128), .ZN(n7130) );
  OAI21_X1 U8295 ( .B1(n7131), .B2(n7130), .A(n7281), .ZN(n7132) );
  NAND2_X1 U8296 ( .A1(n7132), .A2(n10197), .ZN(n7138) );
  INV_X1 U8297 ( .A(n7208), .ZN(n7136) );
  INV_X1 U8298 ( .A(n7327), .ZN(n7332) );
  AOI21_X1 U8299 ( .B1(n10218), .B2(n10234), .A(n7133), .ZN(n7134) );
  OAI21_X1 U8300 ( .B1(n7332), .B2(n10215), .A(n7134), .ZN(n7135) );
  AOI21_X1 U8301 ( .B1(n7136), .B2(n10203), .A(n7135), .ZN(n7137) );
  OAI211_X1 U8302 ( .C1(n10823), .C2(n10206), .A(n7138), .B(n7137), .ZN(
        P1_U3211) );
  NAND2_X1 U8303 ( .A1(n7343), .A2(n8693), .ZN(n7141) );
  INV_X1 U8304 ( .A(n7139), .ZN(n9232) );
  AOI22_X1 U8305 ( .A1(n8685), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5856), .B2(
        n9232), .ZN(n7140) );
  NAND2_X1 U8306 ( .A1(n7141), .A2(n7140), .ZN(n7679) );
  INV_X1 U8307 ( .A(n7679), .ZN(n10898) );
  NAND2_X1 U8308 ( .A1(n7306), .A2(n8693), .ZN(n7144) );
  AOI22_X1 U8309 ( .A1(n8685), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5856), .B2(
        n7142), .ZN(n7143) );
  XNOR2_X1 U8310 ( .A(n10878), .B(n5877), .ZN(n7150) );
  NOR2_X1 U8311 ( .A1(n7461), .A2(n8940), .ZN(n7148) );
  XNOR2_X1 U8312 ( .A(n7150), .B(n7148), .ZN(n7182) );
  AND2_X1 U8313 ( .A1(n7182), .A2(n7145), .ZN(n7146) );
  INV_X1 U8314 ( .A(n7148), .ZN(n7149) );
  NAND2_X1 U8315 ( .A1(n7150), .A2(n7149), .ZN(n7151) );
  XNOR2_X1 U8316 ( .A(n7679), .B(n8941), .ZN(n7152) );
  NOR2_X1 U8317 ( .A1(n7448), .A2(n8940), .ZN(n7153) );
  NAND2_X1 U8318 ( .A1(n7152), .A2(n7153), .ZN(n7232) );
  INV_X1 U8319 ( .A(n7152), .ZN(n7231) );
  INV_X1 U8320 ( .A(n7153), .ZN(n7154) );
  NAND2_X1 U8321 ( .A1(n7231), .A2(n7154), .ZN(n7155) );
  NAND2_X1 U8322 ( .A1(n7232), .A2(n7155), .ZN(n7157) );
  AOI21_X1 U8323 ( .B1(n7156), .B2(n7157), .A(n9195), .ZN(n7159) );
  NAND2_X1 U8324 ( .A1(n7159), .A2(n7233), .ZN(n7170) );
  NAND2_X1 U8325 ( .A1(n8013), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7167) );
  OR2_X1 U8326 ( .A1(n5839), .A2(n10948), .ZN(n7166) );
  NAND2_X1 U8327 ( .A1(n7160), .A2(n7240), .ZN(n7161) );
  NAND2_X1 U8328 ( .A1(n7162), .A2(n7161), .ZN(n10934) );
  OR2_X1 U8329 ( .A1(n8040), .A2(n10934), .ZN(n7165) );
  OR2_X1 U8330 ( .A1(n8093), .A2(n7163), .ZN(n7164) );
  INV_X1 U8331 ( .A(n8386), .ZN(n9219) );
  AND2_X1 U8332 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9231) );
  OAI22_X1 U8333 ( .A1(n7461), .A2(n9159), .B1(n9206), .B2(n7454), .ZN(n7168)
         );
  AOI211_X1 U8334 ( .C1(n9185), .C2(n9219), .A(n9231), .B(n7168), .ZN(n7169)
         );
  OAI211_X1 U8335 ( .C1(n10898), .C2(n9211), .A(n7170), .B(n7169), .ZN(
        P2_U3219) );
  NOR3_X1 U8336 ( .A1(n7172), .A2(n7171), .A3(n9198), .ZN(n7173) );
  AOI21_X1 U8337 ( .B1(n7174), .B2(n9167), .A(n7173), .ZN(n7183) );
  INV_X1 U8338 ( .A(n7426), .ZN(n7175) );
  AOI22_X1 U8339 ( .A1(n9220), .A2(n9189), .B1(n9188), .B2(n7175), .ZN(n7177)
         );
  OAI211_X1 U8340 ( .C1(n7448), .C2(n9161), .A(n7177), .B(n7176), .ZN(n7180)
         );
  NOR2_X1 U8341 ( .A1(n7178), .A2(n9195), .ZN(n7179) );
  AOI211_X1 U8342 ( .C1(n9171), .C2(n10878), .A(n7180), .B(n7179), .ZN(n7181)
         );
  OAI21_X1 U8343 ( .B1(n7183), .B2(n7182), .A(n7181), .ZN(P2_U3233) );
  MUX2_X1 U8344 ( .A(n7192), .B(n9683), .S(n7833), .Z(n7189) );
  INV_X1 U8345 ( .A(SI_19_), .ZN(n7188) );
  NAND2_X1 U8346 ( .A1(n7189), .A2(n7188), .ZN(n7265) );
  INV_X1 U8347 ( .A(n7189), .ZN(n7190) );
  NAND2_X1 U8348 ( .A1(n7190), .A2(SI_19_), .ZN(n7191) );
  NAND2_X1 U8349 ( .A1(n7265), .A2(n7191), .ZN(n7263) );
  XNOR2_X1 U8350 ( .A(n7264), .B(n7263), .ZN(n8132) );
  INV_X1 U8351 ( .A(n8132), .ZN(n8394) );
  OAI222_X1 U8352 ( .A1(n9110), .A2(n7192), .B1(n6076), .B2(n8394), .C1(
        P2_U3152), .C2(n8884), .ZN(P2_U3339) );
  NAND2_X1 U8353 ( .A1(n7194), .A2(n7193), .ZN(n7196) );
  NAND2_X1 U8354 ( .A1(n10778), .A2(n10762), .ZN(n7195) );
  NAND2_X1 U8355 ( .A1(n7196), .A2(n7195), .ZN(n10770) );
  INV_X1 U8356 ( .A(n10803), .ZN(n7197) );
  NAND2_X1 U8357 ( .A1(n7197), .A2(n10784), .ZN(n8409) );
  INV_X1 U8358 ( .A(n10784), .ZN(n10773) );
  NAND2_X1 U8359 ( .A1(n10803), .A2(n10773), .ZN(n8412) );
  NAND2_X1 U8360 ( .A1(n10803), .A2(n10784), .ZN(n7198) );
  NAND2_X1 U8361 ( .A1(n7199), .A2(n7198), .ZN(n10800) );
  NAND2_X1 U8362 ( .A1(n10780), .A2(n10814), .ZN(n8505) );
  INV_X1 U8363 ( .A(n10814), .ZN(n7201) );
  NAND2_X1 U8364 ( .A1(n10234), .A2(n7201), .ZN(n8414) );
  NAND2_X1 U8365 ( .A1(n10780), .A2(n7201), .ZN(n7202) );
  XOR2_X1 U8366 ( .A(n7326), .B(n8645), .Z(n10824) );
  INV_X1 U8367 ( .A(n8408), .ZN(n7203) );
  INV_X1 U8368 ( .A(n8412), .ZN(n7205) );
  NAND2_X1 U8369 ( .A1(n7206), .A2(n8505), .ZN(n7330) );
  XOR2_X1 U8370 ( .A(n7330), .B(n8645), .Z(n7207) );
  AOI222_X1 U8371 ( .A1(n11035), .A2(n7207), .B1(n7327), .B2(n11037), .C1(
        n10234), .C2(n11040), .ZN(n10822) );
  OR2_X1 U8372 ( .A1(n10822), .A2(n11070), .ZN(n7214) );
  OAI22_X1 U8373 ( .A1(n10795), .A2(n6242), .B1(n7208), .B2(n10786), .ZN(n7211) );
  OR2_X1 U8374 ( .A1(n10771), .A2(n10784), .ZN(n10808) );
  INV_X1 U8375 ( .A(n10842), .ZN(n7209) );
  OAI211_X1 U8376 ( .C1(n10823), .C2(n10807), .A(n7209), .B(n10953), .ZN(
        n10821) );
  NOR2_X1 U8377 ( .A1(n10821), .A2(n11063), .ZN(n7210) );
  AOI211_X1 U8378 ( .C1(n11060), .C2(n7212), .A(n7211), .B(n7210), .ZN(n7213)
         );
  OAI211_X1 U8379 ( .C1(n11064), .C2(n10824), .A(n7214), .B(n7213), .ZN(
        P1_U3284) );
  OAI21_X1 U8380 ( .B1(n7802), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7215), .ZN(
        n7403) );
  XNOR2_X1 U8381 ( .A(n7847), .B(n7403), .ZN(n7216) );
  INV_X1 U8382 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11029) );
  NOR2_X1 U8383 ( .A1(n11029), .A2(n7216), .ZN(n7404) );
  AOI211_X1 U8384 ( .C1(n7216), .C2(n11029), .A(n7404), .B(n10693), .ZN(n7222)
         );
  INV_X1 U8385 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7868) );
  AOI21_X1 U8386 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7802), .A(n7217), .ZN(
        n7397) );
  XNOR2_X1 U8387 ( .A(n7847), .B(n7397), .ZN(n7218) );
  NOR2_X1 U8388 ( .A1(n7868), .A2(n7218), .ZN(n7398) );
  AOI211_X1 U8389 ( .C1(n7868), .C2(n7218), .A(n7398), .B(n10701), .ZN(n7221)
         );
  NAND2_X1 U8390 ( .A1(n10696), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7219) );
  NAND2_X1 U8391 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10213) );
  OAI211_X1 U8392 ( .C1(n10692), .C2(n7847), .A(n7219), .B(n10213), .ZN(n7220)
         );
  OR3_X1 U8393 ( .A1(n7222), .A2(n7221), .A3(n7220), .ZN(P1_U3256) );
  NAND2_X1 U8394 ( .A1(n7533), .A2(n8693), .ZN(n7225) );
  AOI22_X1 U8395 ( .A1(n8685), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5856), .B2(
        n7223), .ZN(n7224) );
  INV_X1 U8396 ( .A(n10939), .ZN(n10928) );
  XNOR2_X1 U8397 ( .A(n10939), .B(n8941), .ZN(n8378) );
  NOR2_X1 U8398 ( .A1(n8386), .A2(n8940), .ZN(n7226) );
  NAND2_X1 U8399 ( .A1(n8378), .A2(n7226), .ZN(n7604) );
  INV_X1 U8400 ( .A(n8378), .ZN(n7228) );
  INV_X1 U8401 ( .A(n7226), .ZN(n7227) );
  NAND2_X1 U8402 ( .A1(n7228), .A2(n7227), .ZN(n7229) );
  AND2_X1 U8403 ( .A1(n7604), .A2(n7229), .ZN(n7234) );
  INV_X1 U8404 ( .A(n7234), .ZN(n7230) );
  AOI21_X1 U8405 ( .B1(n7233), .B2(n7230), .A(n9195), .ZN(n7237) );
  NOR3_X1 U8406 ( .A1(n7231), .A2(n7448), .A3(n9198), .ZN(n7236) );
  OAI21_X1 U8407 ( .B1(n7237), .B2(n7236), .A(n8380), .ZN(n7243) );
  OR2_X1 U8408 ( .A1(n8372), .A2(n9468), .ZN(n7239) );
  OR2_X1 U8409 ( .A1(n7448), .A2(n9466), .ZN(n7238) );
  NAND2_X1 U8410 ( .A1(n7239), .A2(n7238), .ZN(n10936) );
  OAI22_X1 U8411 ( .A1(n9206), .A2(n10934), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7240), .ZN(n7241) );
  AOI21_X1 U8412 ( .B1(n10936), .B2(n9208), .A(n7241), .ZN(n7242) );
  OAI211_X1 U8413 ( .C1(n10928), .C2(n9211), .A(n7243), .B(n7242), .ZN(
        P2_U3238) );
  OAI21_X1 U8414 ( .B1(n7619), .B2(n7245), .A(n7244), .ZN(n7246) );
  NAND2_X1 U8415 ( .A1(n7626), .A2(n7246), .ZN(n7247) );
  XNOR2_X1 U8416 ( .A(n7385), .B(n7246), .ZN(n7382) );
  NAND2_X1 U8417 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7382), .ZN(n7381) );
  NAND2_X1 U8418 ( .A1(n7247), .A2(n7381), .ZN(n7249) );
  XNOR2_X1 U8419 ( .A(n7640), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7248) );
  NOR2_X1 U8420 ( .A1(n7248), .A2(n7249), .ZN(n7593) );
  AOI21_X1 U8421 ( .B1(n7249), .B2(n7248), .A(n7593), .ZN(n7262) );
  INV_X1 U8422 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9846) );
  NOR2_X1 U8423 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9846), .ZN(n7250) );
  AOI21_X1 U8424 ( .B1(n10674), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7250), .ZN(
        n7251) );
  INV_X1 U8425 ( .A(n7251), .ZN(n7260) );
  OAI21_X1 U8426 ( .B1(n7613), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7252), .ZN(
        n7253) );
  NAND2_X1 U8427 ( .A1(n7385), .A2(n7253), .ZN(n7254) );
  XNOR2_X1 U8428 ( .A(n7626), .B(n7253), .ZN(n7380) );
  INV_X1 U8429 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7379) );
  NAND2_X1 U8430 ( .A1(n7380), .A2(n7379), .ZN(n7378) );
  NAND2_X1 U8431 ( .A1(n7254), .A2(n7378), .ZN(n7258) );
  INV_X1 U8432 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7255) );
  MUX2_X1 U8433 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n7255), .S(n7640), .Z(n7256)
         );
  INV_X1 U8434 ( .A(n7256), .ZN(n7257) );
  NOR2_X1 U8435 ( .A1(n7258), .A2(n7257), .ZN(n7589) );
  AOI211_X1 U8436 ( .C1(n7258), .C2(n7257), .A(n7589), .B(n9278), .ZN(n7259)
         );
  AOI211_X1 U8437 ( .C1(n7640), .C2(n10660), .A(n7260), .B(n7259), .ZN(n7261)
         );
  OAI21_X1 U8438 ( .B1(n7262), .B2(n10658), .A(n7261), .ZN(P2_U3261) );
  MUX2_X1 U8439 ( .A(n7302), .B(n9684), .S(n7833), .Z(n7267) );
  INV_X1 U8440 ( .A(SI_20_), .ZN(n7266) );
  NAND2_X1 U8441 ( .A1(n7267), .A2(n7266), .ZN(n7392) );
  INV_X1 U8442 ( .A(n7267), .ZN(n7268) );
  NAND2_X1 U8443 ( .A1(n7268), .A2(SI_20_), .ZN(n7269) );
  XNOR2_X1 U8444 ( .A(n7391), .B(n7390), .ZN(n8145) );
  INV_X1 U8445 ( .A(n8145), .ZN(n7301) );
  OAI222_X1 U8446 ( .A1(n10532), .A2(n7301), .B1(P1_U3084), .B2(n10708), .C1(
        n9684), .C2(n10528), .ZN(P1_U3333) );
  NAND2_X1 U8447 ( .A1(n7270), .A2(n8487), .ZN(n7273) );
  AOI22_X1 U8448 ( .A1(n8472), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8133), .B2(
        n7271), .ZN(n7272) );
  NAND2_X1 U8449 ( .A1(n7273), .A2(n7272), .ZN(n10860) );
  NAND2_X1 U8450 ( .A1(n10860), .A2(n7122), .ZN(n7275) );
  NAND2_X1 U8451 ( .A1(n7327), .A2(n9080), .ZN(n7274) );
  NAND2_X1 U8452 ( .A1(n7275), .A2(n7274), .ZN(n7276) );
  XNOR2_X1 U8453 ( .A(n7276), .B(n9076), .ZN(n7303) );
  INV_X1 U8454 ( .A(n7277), .ZN(n7279) );
  NAND2_X1 U8455 ( .A1(n7279), .A2(n7278), .ZN(n7280) );
  NAND2_X1 U8456 ( .A1(n10860), .A2(n9080), .ZN(n7283) );
  NAND2_X1 U8457 ( .A1(n7327), .A2(n9085), .ZN(n7282) );
  AND2_X1 U8458 ( .A1(n7283), .A2(n7282), .ZN(n7284) );
  NAND2_X1 U8459 ( .A1(n7305), .A2(n7304), .ZN(n7286) );
  XOR2_X1 U8460 ( .A(n7303), .B(n7286), .Z(n7300) );
  NAND2_X1 U8461 ( .A1(n8238), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7294) );
  OR2_X1 U8462 ( .A1(n8496), .A2(n7479), .ZN(n7293) );
  OR2_X1 U8463 ( .A1(n6629), .A2(n7287), .ZN(n7292) );
  NAND2_X1 U8464 ( .A1(n7289), .A2(n7288), .ZN(n7290) );
  NAND2_X1 U8465 ( .A1(n7314), .A2(n7290), .ZN(n7335) );
  OR2_X1 U8466 ( .A1(n8209), .A2(n7335), .ZN(n7291) );
  NAND4_X1 U8467 ( .A1(n7294), .A2(n7293), .A3(n7292), .A4(n7291), .ZN(n10849)
         );
  INV_X1 U8468 ( .A(n10849), .ZN(n7329) );
  NOR2_X1 U8469 ( .A1(n10215), .A2(n7329), .ZN(n7295) );
  AOI211_X1 U8470 ( .C1(n10218), .C2(n10848), .A(n7296), .B(n7295), .ZN(n7297)
         );
  OAI21_X1 U8471 ( .B1(n10221), .B2(n10858), .A(n7297), .ZN(n7298) );
  AOI21_X1 U8472 ( .B1(n10860), .B2(n10223), .A(n7298), .ZN(n7299) );
  OAI21_X1 U8473 ( .B1(n7300), .B2(n10226), .A(n7299), .ZN(P1_U3219) );
  OAI222_X1 U8474 ( .A1(n9110), .A2(n7302), .B1(n6076), .B2(n7301), .C1(n8889), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NAND2_X1 U8475 ( .A1(n7306), .A2(n8487), .ZN(n7308) );
  AOI22_X1 U8476 ( .A1(n8472), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8133), .B2(
        n10604), .ZN(n7307) );
  NAND2_X1 U8477 ( .A1(n7472), .A2(n7122), .ZN(n7310) );
  NAND2_X1 U8478 ( .A1(n10849), .A2(n9080), .ZN(n7309) );
  NAND2_X1 U8479 ( .A1(n7310), .A2(n7309), .ZN(n7311) );
  XNOR2_X1 U8480 ( .A(n7311), .B(n9083), .ZN(n7433) );
  AND2_X1 U8481 ( .A1(n10849), .A2(n9085), .ZN(n7312) );
  AOI21_X1 U8482 ( .B1(n7472), .B2(n9080), .A(n7312), .ZN(n7432) );
  XNOR2_X1 U8483 ( .A(n7433), .B(n7432), .ZN(n7434) );
  XOR2_X1 U8484 ( .A(n7435), .B(n7434), .Z(n7324) );
  NAND2_X1 U8485 ( .A1(n8238), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7319) );
  OR2_X1 U8486 ( .A1(n6629), .A2(n7373), .ZN(n7318) );
  OR2_X1 U8487 ( .A1(n8496), .A2(n10894), .ZN(n7317) );
  NAND2_X1 U8488 ( .A1(n7314), .A2(n7313), .ZN(n7315) );
  NAND2_X1 U8489 ( .A1(n7356), .A2(n7315), .ZN(n7444) );
  OR2_X1 U8490 ( .A1(n6203), .A2(n7444), .ZN(n7316) );
  NAND4_X1 U8491 ( .A1(n7319), .A2(n7318), .A3(n7317), .A4(n7316), .ZN(n10233)
         );
  NAND2_X1 U8492 ( .A1(n10218), .A2(n7327), .ZN(n7320) );
  NAND2_X1 U8493 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10615) );
  OAI211_X1 U8494 ( .C1(n7567), .C2(n10215), .A(n7320), .B(n10615), .ZN(n7322)
         );
  NOR2_X1 U8495 ( .A1(n10221), .A2(n7335), .ZN(n7321) );
  AOI211_X1 U8496 ( .C1(n7472), .C2(n10223), .A(n7322), .B(n7321), .ZN(n7323)
         );
  OAI21_X1 U8497 ( .B1(n7324), .B2(n10226), .A(n7323), .ZN(P1_U3229) );
  INV_X1 U8498 ( .A(n10860), .ZN(n10843) );
  NAND2_X1 U8499 ( .A1(n10843), .A2(n7327), .ZN(n8432) );
  NAND2_X1 U8500 ( .A1(n7332), .A2(n10860), .ZN(n8520) );
  NAND2_X1 U8501 ( .A1(n10840), .A2(n10839), .ZN(n10838) );
  NAND2_X1 U8502 ( .A1(n10860), .A2(n7327), .ZN(n7328) );
  NOR2_X1 U8503 ( .A1(n7472), .A2(n7329), .ZN(n8521) );
  NAND2_X1 U8504 ( .A1(n7472), .A2(n7329), .ZN(n8514) );
  INV_X1 U8505 ( .A(n8514), .ZN(n8421) );
  OR2_X1 U8506 ( .A1(n8521), .A2(n8421), .ZN(n8646) );
  XNOR2_X1 U8507 ( .A(n7342), .B(n8646), .ZN(n7474) );
  INV_X1 U8508 ( .A(n11035), .ZN(n10777) );
  AND2_X1 U8509 ( .A1(n10844), .A2(n8520), .ZN(n8428) );
  XOR2_X1 U8510 ( .A(n8646), .B(n7353), .Z(n7331) );
  OAI222_X1 U8511 ( .A1(n10779), .A2(n7332), .B1(n10781), .B2(n7567), .C1(
        n10777), .C2(n7331), .ZN(n7470) );
  NAND2_X1 U8512 ( .A1(n7470), .A2(n10795), .ZN(n7339) );
  NAND2_X1 U8513 ( .A1(n10842), .A2(n10843), .ZN(n10841) );
  INV_X1 U8514 ( .A(n7371), .ZN(n7333) );
  AOI211_X1 U8515 ( .C1(n7472), .C2(n10841), .A(n11043), .B(n7333), .ZN(n7471)
         );
  INV_X1 U8516 ( .A(n7472), .ZN(n7334) );
  NOR2_X1 U8517 ( .A1(n7334), .A2(n10430), .ZN(n7337) );
  OAI22_X1 U8518 ( .A1(n10795), .A2(n7287), .B1(n7335), .B2(n10786), .ZN(n7336) );
  AOI211_X1 U8519 ( .C1(n7471), .C2(n10291), .A(n7337), .B(n7336), .ZN(n7338)
         );
  OAI211_X1 U8520 ( .C1(n7474), .C2(n11064), .A(n7339), .B(n7338), .ZN(
        P1_U3282) );
  OR2_X1 U8521 ( .A1(n7472), .A2(n10849), .ZN(n7341) );
  AND2_X1 U8522 ( .A1(n7472), .A2(n10849), .ZN(n7340) );
  NAND2_X1 U8523 ( .A1(n7343), .A2(n8487), .ZN(n7346) );
  AOI22_X1 U8524 ( .A1(n8472), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8133), .B2(
        n7344), .ZN(n7345) );
  OR2_X1 U8525 ( .A1(n10887), .A2(n7567), .ZN(n8525) );
  NAND2_X1 U8526 ( .A1(n10887), .A2(n7567), .ZN(n8526) );
  NAND2_X1 U8527 ( .A1(n8525), .A2(n8526), .ZN(n8522) );
  NAND2_X1 U8528 ( .A1(n7347), .A2(n8522), .ZN(n7563) );
  OR2_X1 U8529 ( .A1(n7347), .A2(n8522), .ZN(n7348) );
  NAND2_X1 U8530 ( .A1(n7563), .A2(n7348), .ZN(n10891) );
  OR2_X1 U8531 ( .A1(n7349), .A2(n7369), .ZN(n7352) );
  OR2_X1 U8532 ( .A1(n7350), .A2(n8667), .ZN(n7351) );
  INV_X1 U8533 ( .A(n10851), .ZN(n10913) );
  NAND2_X1 U8534 ( .A1(n10891), .A2(n10913), .ZN(n7368) );
  INV_X1 U8535 ( .A(n8522), .ZN(n8649) );
  OAI21_X1 U8536 ( .B1(n8649), .B2(n7354), .A(n7565), .ZN(n7366) );
  NAND2_X1 U8537 ( .A1(n10849), .A2(n11040), .ZN(n7364) );
  NAND2_X1 U8538 ( .A1(n8490), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7362) );
  OR2_X1 U8539 ( .A1(n8496), .A2(n10915), .ZN(n7361) );
  INV_X1 U8540 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U8541 ( .A1(n7356), .A2(n7355), .ZN(n7357) );
  NAND2_X1 U8542 ( .A1(n7550), .A2(n7357), .ZN(n7570) );
  OR2_X1 U8543 ( .A1(n8209), .A2(n7570), .ZN(n7360) );
  INV_X1 U8544 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7358) );
  OR2_X1 U8545 ( .A1(n8492), .A2(n7358), .ZN(n7359) );
  NAND4_X1 U8546 ( .A1(n7362), .A2(n7361), .A3(n7360), .A4(n7359), .ZN(n10958)
         );
  NAND2_X1 U8547 ( .A1(n10958), .A2(n11037), .ZN(n7363) );
  NAND2_X1 U8548 ( .A1(n7364), .A2(n7363), .ZN(n7365) );
  AOI21_X1 U8549 ( .B1(n7366), .B2(n11035), .A(n7365), .ZN(n7367) );
  AND2_X1 U8550 ( .A1(n7368), .A2(n7367), .ZN(n10893) );
  AND2_X1 U8551 ( .A1(n7369), .A2(n10789), .ZN(n7370) );
  NAND2_X1 U8552 ( .A1(n10795), .A2(n7370), .ZN(n10415) );
  INV_X1 U8553 ( .A(n10415), .ZN(n10863) );
  AOI21_X1 U8554 ( .B1(n7371), .B2(n10887), .A(n11043), .ZN(n7372) );
  OAI22_X1 U8555 ( .A1(n10795), .A2(n7373), .B1(n7444), .B2(n10786), .ZN(n7374) );
  AOI21_X1 U8556 ( .B1(n11060), .B2(n10887), .A(n7374), .ZN(n7375) );
  OAI21_X1 U8557 ( .B1(n10889), .B2(n11063), .A(n7375), .ZN(n7376) );
  AOI21_X1 U8558 ( .B1(n10891), .B2(n10863), .A(n7376), .ZN(n7377) );
  OAI21_X1 U8559 ( .B1(n10893), .B2(n11070), .A(n7377), .ZN(P1_U3281) );
  OAI21_X1 U8560 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7388) );
  INV_X1 U8561 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7384) );
  OAI211_X1 U8562 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n7382), .A(n10682), .B(
        n7381), .ZN(n7383) );
  NAND2_X1 U8563 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8947) );
  OAI211_X1 U8564 ( .C1(n9257), .C2(n7384), .A(n7383), .B(n8947), .ZN(n7387)
         );
  NOR2_X1 U8565 ( .A1(n10670), .A2(n7385), .ZN(n7386) );
  AOI211_X1 U8566 ( .C1(n10679), .C2(n7388), .A(n7387), .B(n7386), .ZN(n7389)
         );
  INV_X1 U8567 ( .A(n7389), .ZN(P2_U3260) );
  MUX2_X1 U8568 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5153), .Z(n7481) );
  INV_X1 U8569 ( .A(SI_21_), .ZN(n7393) );
  XNOR2_X1 U8570 ( .A(n7481), .B(n7393), .ZN(n7480) );
  INV_X1 U8571 ( .A(n8156), .ZN(n7395) );
  INV_X1 U8572 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7394) );
  OAI222_X1 U8573 ( .A1(n10532), .A2(n7395), .B1(P1_U3084), .B2(n8667), .C1(
        n7394), .C2(n10528), .ZN(P1_U3332) );
  INV_X1 U8574 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7396) );
  OAI222_X1 U8575 ( .A1(n9110), .A2(n7396), .B1(n6076), .B2(n7395), .C1(n8708), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NOR2_X1 U8576 ( .A1(n7397), .A2(n7847), .ZN(n7399) );
  NOR2_X1 U8577 ( .A1(n7399), .A2(n7398), .ZN(n7402) );
  NAND2_X1 U8578 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8103), .ZN(n7400) );
  OAI21_X1 U8579 ( .B1(n8103), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7400), .ZN(
        n7401) );
  NOR2_X1 U8580 ( .A1(n7402), .A2(n7401), .ZN(n7669) );
  AOI211_X1 U8581 ( .C1(n7402), .C2(n7401), .A(n7669), .B(n10701), .ZN(n7414)
         );
  NOR2_X1 U8582 ( .A1(n7847), .A2(n7403), .ZN(n7405) );
  NOR2_X1 U8583 ( .A1(n7405), .A2(n7404), .ZN(n7408) );
  INV_X1 U8584 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11053) );
  NOR2_X1 U8585 ( .A1(n8103), .A2(n11053), .ZN(n7406) );
  AOI21_X1 U8586 ( .B1(n8103), .B2(n11053), .A(n7406), .ZN(n7407) );
  NOR2_X1 U8587 ( .A1(n7408), .A2(n7407), .ZN(n7666) );
  AOI211_X1 U8588 ( .C1(n7408), .C2(n7407), .A(n7666), .B(n10693), .ZN(n7413)
         );
  NAND2_X1 U8589 ( .A1(n10696), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7410) );
  NAND2_X1 U8590 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n7409) );
  OAI211_X1 U8591 ( .C1(n7411), .C2(n10692), .A(n7410), .B(n7409), .ZN(n7412)
         );
  OR3_X1 U8592 ( .A1(n7414), .A2(n7413), .A3(n7412), .ZN(P1_U3257) );
  NAND2_X1 U8593 ( .A1(n10878), .A2(n7461), .ZN(n8746) );
  NAND2_X1 U8594 ( .A1(n9220), .A2(n7415), .ZN(n7416) );
  INV_X1 U8595 ( .A(n7464), .ZN(n7419) );
  AOI21_X1 U8596 ( .B1(n8868), .B2(n7420), .A(n7419), .ZN(n10877) );
  INV_X1 U8597 ( .A(n7448), .ZN(n7678) );
  AOI22_X1 U8598 ( .A1(n7678), .A2(n9501), .B1(n9499), .B2(n9220), .ZN(n7424)
         );
  OAI211_X1 U8599 ( .C1(n7422), .C2(n8868), .A(n7449), .B(n10923), .ZN(n7423)
         );
  OAI211_X1 U8600 ( .C1(n10877), .C2(n7425), .A(n7424), .B(n7423), .ZN(n10881)
         );
  NAND2_X1 U8601 ( .A1(n10881), .A2(n10946), .ZN(n7430) );
  OAI22_X1 U8602 ( .A1(n10946), .A2(n6331), .B1(n7426), .B2(n10935), .ZN(n7428) );
  XNOR2_X1 U8603 ( .A(n7456), .B(n10878), .ZN(n10880) );
  NOR2_X1 U8604 ( .A1(n10880), .A2(n9309), .ZN(n7427) );
  AOI211_X1 U8605 ( .C1(n9427), .C2(n10878), .A(n7428), .B(n7427), .ZN(n7429)
         );
  OAI211_X1 U8606 ( .C1(n10877), .C2(n7431), .A(n7430), .B(n7429), .ZN(
        P2_U3287) );
  NAND2_X1 U8607 ( .A1(n10887), .A2(n7122), .ZN(n7437) );
  NAND2_X1 U8608 ( .A1(n10233), .A2(n9080), .ZN(n7436) );
  NAND2_X1 U8609 ( .A1(n7437), .A2(n7436), .ZN(n7438) );
  XNOR2_X1 U8610 ( .A(n7438), .B(n9083), .ZN(n7531) );
  AND2_X1 U8611 ( .A1(n10233), .A2(n9085), .ZN(n7439) );
  AOI21_X1 U8612 ( .B1(n10887), .B2(n9080), .A(n7439), .ZN(n7530) );
  XNOR2_X1 U8613 ( .A(n7531), .B(n7530), .ZN(n7440) );
  XNOR2_X1 U8614 ( .A(n7532), .B(n7440), .ZN(n7447) );
  INV_X1 U8615 ( .A(n10958), .ZN(n7738) );
  NOR2_X1 U8616 ( .A1(n10215), .A2(n7738), .ZN(n7441) );
  AOI211_X1 U8617 ( .C1(n10218), .C2(n10849), .A(n7442), .B(n7441), .ZN(n7443)
         );
  OAI21_X1 U8618 ( .B1(n10221), .B2(n7444), .A(n7443), .ZN(n7445) );
  AOI21_X1 U8619 ( .B1(n10887), .B2(n10223), .A(n7445), .ZN(n7446) );
  OAI21_X1 U8620 ( .B1(n7447), .B2(n10226), .A(n7446), .ZN(P1_U3215) );
  OR2_X1 U8621 ( .A1(n7679), .A2(n7448), .ZN(n8753) );
  NAND2_X1 U8622 ( .A1(n7679), .A2(n7448), .ZN(n8752) );
  NAND2_X1 U8623 ( .A1(n8753), .A2(n8752), .ZN(n8869) );
  INV_X1 U8624 ( .A(n7684), .ZN(n7451) );
  AOI21_X1 U8625 ( .B1(n8869), .B2(n7452), .A(n7451), .ZN(n7453) );
  OAI222_X1 U8626 ( .A1(n9468), .A2(n8386), .B1(n9466), .B2(n7461), .C1(n9486), 
        .C2(n7453), .ZN(n10900) );
  INV_X1 U8627 ( .A(n10900), .ZN(n7469) );
  OAI22_X1 U8628 ( .A1(n10946), .A2(n7455), .B1(n7454), .B2(n10935), .ZN(n7460) );
  NOR2_X1 U8629 ( .A1(n7456), .A2(n10878), .ZN(n7457) );
  AND2_X2 U8630 ( .A1(n7457), .A2(n10898), .ZN(n10929) );
  NOR2_X1 U8631 ( .A1(n7457), .A2(n10898), .ZN(n7458) );
  OR2_X1 U8632 ( .A1(n10929), .A2(n7458), .ZN(n10899) );
  NOR2_X1 U8633 ( .A1(n10899), .A2(n9309), .ZN(n7459) );
  AOI211_X1 U8634 ( .C1(n9427), .C2(n7679), .A(n7460), .B(n7459), .ZN(n7468)
         );
  INV_X1 U8635 ( .A(n7461), .ZN(n7462) );
  OR2_X1 U8636 ( .A1(n10878), .A2(n7462), .ZN(n7463) );
  NOR2_X1 U8637 ( .A1(n7465), .A2(n8869), .ZN(n10897) );
  INV_X1 U8638 ( .A(n10897), .ZN(n7466) );
  NAND3_X1 U8639 ( .A1(n7466), .A2(n9400), .A3(n7680), .ZN(n7467) );
  OAI211_X1 U8640 ( .C1(n7469), .C2(n9504), .A(n7468), .B(n7467), .ZN(P2_U3286) );
  INV_X1 U8641 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7476) );
  AOI211_X1 U8642 ( .C1(n10908), .C2(n7472), .A(n7471), .B(n7470), .ZN(n7473)
         );
  OAI21_X1 U8643 ( .B1(n10769), .B2(n7474), .A(n7473), .ZN(n7477) );
  NAND2_X1 U8644 ( .A1(n7477), .A2(n11057), .ZN(n7475) );
  OAI21_X1 U8645 ( .B1(n11057), .B2(n7476), .A(n7475), .ZN(P1_U3481) );
  NAND2_X1 U8646 ( .A1(n7477), .A2(n11054), .ZN(n7478) );
  OAI21_X1 U8647 ( .B1(n11054), .B2(n7479), .A(n7478), .ZN(P1_U3532) );
  INV_X1 U8648 ( .A(n7480), .ZN(n7483) );
  NAND2_X1 U8649 ( .A1(n7481), .A2(SI_21_), .ZN(n7482) );
  MUX2_X1 U8650 ( .A(n7488), .B(n9679), .S(n7833), .Z(n7485) );
  INV_X1 U8651 ( .A(SI_22_), .ZN(n9784) );
  NAND2_X1 U8652 ( .A1(n7485), .A2(n9784), .ZN(n7576) );
  INV_X1 U8653 ( .A(n7485), .ZN(n7486) );
  NAND2_X1 U8654 ( .A1(n7486), .A2(SI_22_), .ZN(n7487) );
  NAND2_X1 U8655 ( .A1(n7576), .A2(n7487), .ZN(n7577) );
  XNOR2_X1 U8656 ( .A(n7578), .B(n7577), .ZN(n8167) );
  INV_X1 U8657 ( .A(n8167), .ZN(n7956) );
  OAI222_X1 U8658 ( .A1(n9110), .A2(n7488), .B1(n6076), .B2(n7956), .C1(
        P2_U3152), .C2(n8704), .ZN(P2_U3336) );
  NOR2_X1 U8659 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7525) );
  NOR2_X1 U8660 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7523) );
  NOR2_X1 U8661 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7521) );
  NOR2_X1 U8662 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7519) );
  NOR2_X1 U8663 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7517) );
  NOR2_X1 U8664 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7515) );
  NAND2_X1 U8665 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7513) );
  XOR2_X1 U8666 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10566) );
  NAND2_X1 U8667 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7511) );
  XOR2_X1 U8668 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10564) );
  NOR2_X1 U8669 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7495) );
  XNOR2_X1 U8670 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10555) );
  NAND2_X1 U8671 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7493) );
  XOR2_X1 U8672 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10553) );
  NAND2_X1 U8673 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7491) );
  XOR2_X1 U8674 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10551) );
  AOI21_X1 U8675 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10546) );
  INV_X1 U8676 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7489) );
  NAND3_X1 U8677 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10548) );
  OAI21_X1 U8678 ( .B1(n10546), .B2(n7489), .A(n10548), .ZN(n10550) );
  NAND2_X1 U8679 ( .A1(n10551), .A2(n10550), .ZN(n7490) );
  NAND2_X1 U8680 ( .A1(n7491), .A2(n7490), .ZN(n10552) );
  NAND2_X1 U8681 ( .A1(n10553), .A2(n10552), .ZN(n7492) );
  NAND2_X1 U8682 ( .A1(n7493), .A2(n7492), .ZN(n10554) );
  NOR2_X1 U8683 ( .A1(n10555), .A2(n10554), .ZN(n7494) );
  NOR2_X1 U8684 ( .A1(n7495), .A2(n7494), .ZN(n7496) );
  NOR2_X1 U8685 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7496), .ZN(n10557) );
  AND2_X1 U8686 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7496), .ZN(n10556) );
  NOR2_X1 U8687 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10556), .ZN(n7497) );
  NAND2_X1 U8688 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7498), .ZN(n7500) );
  XOR2_X1 U8689 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7498), .Z(n10559) );
  NAND2_X1 U8690 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10559), .ZN(n7499) );
  NAND2_X1 U8691 ( .A1(n7500), .A2(n7499), .ZN(n7501) );
  NAND2_X1 U8692 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7501), .ZN(n7503) );
  XOR2_X1 U8693 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7501), .Z(n10560) );
  NAND2_X1 U8694 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10560), .ZN(n7502) );
  NAND2_X1 U8695 ( .A1(n7503), .A2(n7502), .ZN(n7504) );
  NAND2_X1 U8696 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7504), .ZN(n7506) );
  XOR2_X1 U8697 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7504), .Z(n10561) );
  NAND2_X1 U8698 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10561), .ZN(n7505) );
  NAND2_X1 U8699 ( .A1(n7506), .A2(n7505), .ZN(n7507) );
  NAND2_X1 U8700 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7507), .ZN(n7509) );
  XOR2_X1 U8701 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7507), .Z(n10562) );
  NAND2_X1 U8702 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10562), .ZN(n7508) );
  NAND2_X1 U8703 ( .A1(n7509), .A2(n7508), .ZN(n10563) );
  NAND2_X1 U8704 ( .A1(n10564), .A2(n10563), .ZN(n7510) );
  NAND2_X1 U8705 ( .A1(n7511), .A2(n7510), .ZN(n10565) );
  NAND2_X1 U8706 ( .A1(n10566), .A2(n10565), .ZN(n7512) );
  NAND2_X1 U8707 ( .A1(n7513), .A2(n7512), .ZN(n10568) );
  XNOR2_X1 U8708 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10567) );
  XNOR2_X1 U8709 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10569) );
  XNOR2_X1 U8710 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10571) );
  NOR2_X1 U8711 ( .A1(n10572), .A2(n10571), .ZN(n7518) );
  NOR2_X1 U8712 ( .A1(n7519), .A2(n7518), .ZN(n10574) );
  XNOR2_X1 U8713 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10573) );
  NOR2_X1 U8714 ( .A1(n10574), .A2(n10573), .ZN(n7520) );
  NOR2_X1 U8715 ( .A1(n7521), .A2(n7520), .ZN(n10576) );
  XNOR2_X1 U8716 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10575) );
  NOR2_X1 U8717 ( .A1(n10576), .A2(n10575), .ZN(n7522) );
  NOR2_X1 U8718 ( .A1(n7523), .A2(n7522), .ZN(n10578) );
  XNOR2_X1 U8719 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10577) );
  NOR2_X1 U8720 ( .A1(n10578), .A2(n10577), .ZN(n7524) );
  NOR2_X1 U8721 ( .A1(n7525), .A2(n7524), .ZN(n7526) );
  AND2_X1 U8722 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7526), .ZN(n10579) );
  NOR2_X1 U8723 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10579), .ZN(n7527) );
  NOR2_X1 U8724 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7526), .ZN(n10580) );
  NOR2_X1 U8725 ( .A1(n7527), .A2(n10580), .ZN(n7529) );
  XNOR2_X1 U8726 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7528) );
  XNOR2_X1 U8727 ( .A(n7529), .B(n7528), .ZN(ADD_1071_U4) );
  NAND2_X1 U8728 ( .A1(n7532), .A2(n7531), .ZN(n7695) );
  NAND2_X1 U8729 ( .A1(n7698), .A2(n7695), .ZN(n7547) );
  NAND2_X1 U8730 ( .A1(n7533), .A2(n8487), .ZN(n7536) );
  AOI22_X1 U8731 ( .A1(n8472), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8133), .B2(
        n7534), .ZN(n7535) );
  NAND2_X1 U8732 ( .A1(n10907), .A2(n7122), .ZN(n7538) );
  NAND2_X1 U8733 ( .A1(n10958), .A2(n9080), .ZN(n7537) );
  NAND2_X1 U8734 ( .A1(n7538), .A2(n7537), .ZN(n7539) );
  XNOR2_X1 U8735 ( .A(n7539), .B(n9083), .ZN(n7541) );
  AND2_X1 U8736 ( .A1(n10958), .A2(n9085), .ZN(n7540) );
  AOI21_X1 U8737 ( .B1(n10907), .B2(n9080), .A(n7540), .ZN(n7542) );
  INV_X1 U8738 ( .A(n7697), .ZN(n7545) );
  INV_X1 U8739 ( .A(n7541), .ZN(n7544) );
  INV_X1 U8740 ( .A(n7542), .ZN(n7543) );
  NAND2_X1 U8741 ( .A1(n7544), .A2(n7543), .ZN(n7700) );
  NAND2_X1 U8742 ( .A1(n7545), .A2(n7700), .ZN(n7546) );
  XNOR2_X1 U8743 ( .A(n7547), .B(n7546), .ZN(n7561) );
  NAND2_X1 U8744 ( .A1(n8238), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7555) );
  OR2_X1 U8745 ( .A1(n8496), .A2(n10963), .ZN(n7554) );
  INV_X1 U8746 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7548) );
  OR2_X1 U8747 ( .A1(n6629), .A2(n7548), .ZN(n7553) );
  NAND2_X1 U8748 ( .A1(n7550), .A2(n7549), .ZN(n7551) );
  NAND2_X1 U8749 ( .A1(n7713), .A2(n7551), .ZN(n10966) );
  OR2_X1 U8750 ( .A1(n6203), .A2(n10966), .ZN(n7552) );
  NAND4_X1 U8751 ( .A1(n7555), .A2(n7554), .A3(n7553), .A4(n7552), .ZN(n10232)
         );
  NOR2_X1 U8752 ( .A1(n10215), .A2(n7739), .ZN(n7556) );
  AOI211_X1 U8753 ( .C1(n10218), .C2(n10233), .A(n7557), .B(n7556), .ZN(n7558)
         );
  OAI21_X1 U8754 ( .B1(n10221), .B2(n7570), .A(n7558), .ZN(n7559) );
  AOI21_X1 U8755 ( .B1(n10907), .B2(n10223), .A(n7559), .ZN(n7560) );
  OAI21_X1 U8756 ( .B1(n7561), .B2(n10226), .A(n7560), .ZN(P1_U3234) );
  OR2_X1 U8757 ( .A1(n10887), .A2(n10233), .ZN(n7562) );
  NAND2_X1 U8758 ( .A1(n7563), .A2(n7562), .ZN(n7749) );
  NOR2_X1 U8759 ( .A1(n10907), .A2(n10958), .ZN(n8528) );
  NAND2_X1 U8760 ( .A1(n10907), .A2(n10958), .ZN(n8529) );
  INV_X1 U8761 ( .A(n8529), .ZN(n7564) );
  OR2_X1 U8762 ( .A1(n8528), .A2(n7564), .ZN(n8648) );
  XNOR2_X1 U8763 ( .A(n7749), .B(n8648), .ZN(n10910) );
  XOR2_X1 U8764 ( .A(n8648), .B(n7737), .Z(n7566) );
  OAI222_X1 U8765 ( .A1(n10781), .A2(n7739), .B1(n10779), .B2(n7567), .C1(
        n10777), .C2(n7566), .ZN(n10905) );
  NAND2_X1 U8766 ( .A1(n10905), .A2(n10795), .ZN(n7575) );
  AOI211_X1 U8767 ( .C1(n10907), .C2(n7568), .A(n11043), .B(n10954), .ZN(
        n10906) );
  INV_X1 U8768 ( .A(n10907), .ZN(n7569) );
  NOR2_X1 U8769 ( .A1(n7569), .A2(n10430), .ZN(n7573) );
  OAI22_X1 U8770 ( .A1(n10795), .A2(n7571), .B1(n7570), .B2(n10786), .ZN(n7572) );
  AOI211_X1 U8771 ( .C1(n10906), .C2(n10291), .A(n7573), .B(n7572), .ZN(n7574)
         );
  OAI211_X1 U8772 ( .C1(n11064), .C2(n10910), .A(n7575), .B(n7574), .ZN(
        P1_U3280) );
  INV_X1 U8773 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7579) );
  INV_X1 U8774 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9893) );
  MUX2_X1 U8775 ( .A(n7579), .B(n9893), .S(n7833), .Z(n7580) );
  INV_X1 U8776 ( .A(SI_23_), .ZN(n9569) );
  NAND2_X1 U8777 ( .A1(n7580), .A2(n9569), .ZN(n7728) );
  INV_X1 U8778 ( .A(n7580), .ZN(n7581) );
  NAND2_X1 U8779 ( .A1(n7581), .A2(SI_23_), .ZN(n7582) );
  XNOR2_X1 U8780 ( .A(n7727), .B(n7726), .ZN(n8178) );
  INV_X1 U8781 ( .A(n8178), .ZN(n7586) );
  OR2_X1 U8782 ( .A1(n7583), .A2(P1_U3084), .ZN(n8681) );
  NAND2_X1 U8783 ( .A1(n10525), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7584) );
  OAI211_X1 U8784 ( .C1(n7586), .C2(n10532), .A(n8681), .B(n7584), .ZN(
        P1_U3330) );
  NAND2_X1 U8785 ( .A1(n7799), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7585) );
  OAI211_X1 U8786 ( .C1(n7586), .C2(n10053), .A(n8898), .B(n7585), .ZN(
        P2_U3335) );
  INV_X1 U8787 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7588) );
  NOR2_X1 U8788 ( .A1(n9244), .A2(n7588), .ZN(n7587) );
  AOI21_X1 U8789 ( .B1(n9244), .B2(n7588), .A(n7587), .ZN(n7591) );
  AOI21_X1 U8790 ( .B1(n7640), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7589), .ZN(
        n7590) );
  NOR2_X1 U8791 ( .A1(n7590), .A2(n7591), .ZN(n9243) );
  AOI211_X1 U8792 ( .C1(n7591), .C2(n7590), .A(n9243), .B(n9278), .ZN(n7600)
         );
  NOR2_X1 U8793 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9855), .ZN(n7592) );
  AOI21_X1 U8794 ( .B1(n10674), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7592), .ZN(
        n7598) );
  XNOR2_X1 U8795 ( .A(n9249), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7596) );
  INV_X1 U8796 ( .A(n7640), .ZN(n7594) );
  INV_X1 U8797 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7647) );
  AOI21_X1 U8798 ( .B1(n7594), .B2(n7647), .A(n7593), .ZN(n7595) );
  NAND2_X1 U8799 ( .A1(n7596), .A2(n7595), .ZN(n9248) );
  OAI211_X1 U8800 ( .C1(n7596), .C2(n7595), .A(n10682), .B(n9248), .ZN(n7597)
         );
  OAI211_X1 U8801 ( .C1(n10670), .C2(n9249), .A(n7598), .B(n7597), .ZN(n7599)
         );
  OR2_X1 U8802 ( .A1(n7600), .A2(n7599), .ZN(P2_U3262) );
  NAND2_X1 U8803 ( .A1(n7702), .A2(n8693), .ZN(n7603) );
  AOI22_X1 U8804 ( .A1(n8685), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5856), .B2(
        n7601), .ZN(n7602) );
  XNOR2_X1 U8805 ( .A(n10976), .B(n5877), .ZN(n8373) );
  NOR2_X1 U8806 ( .A1(n8372), .A2(n8940), .ZN(n7606) );
  XNOR2_X1 U8807 ( .A(n8373), .B(n7606), .ZN(n8381) );
  AND2_X1 U8808 ( .A1(n8381), .A2(n7604), .ZN(n7605) );
  INV_X1 U8809 ( .A(n7606), .ZN(n7607) );
  NAND2_X1 U8810 ( .A1(n7732), .A2(n8693), .ZN(n7610) );
  AOI22_X1 U8811 ( .A1(n8685), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5856), .B2(
        n7608), .ZN(n7609) );
  XNOR2_X1 U8812 ( .A(n8370), .B(n5877), .ZN(n8976) );
  NOR2_X1 U8813 ( .A1(n8975), .A2(n8940), .ZN(n7611) );
  XNOR2_X1 U8814 ( .A(n8976), .B(n7611), .ZN(n8371) );
  INV_X1 U8815 ( .A(n7611), .ZN(n7612) );
  NAND2_X1 U8816 ( .A1(n7801), .A2(n8693), .ZN(n7615) );
  AOI22_X1 U8817 ( .A1(n8685), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5856), .B2(
        n7613), .ZN(n7614) );
  XNOR2_X1 U8818 ( .A(n8973), .B(n8941), .ZN(n8949) );
  NAND2_X1 U8819 ( .A1(n8013), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7623) );
  OR2_X1 U8820 ( .A1(n5839), .A2(n6990), .ZN(n7622) );
  INV_X1 U8821 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9619) );
  NAND2_X1 U8822 ( .A1(n7617), .A2(n9619), .ZN(n7618) );
  NAND2_X1 U8823 ( .A1(n7630), .A2(n7618), .ZN(n8970) );
  OR2_X1 U8824 ( .A1(n8040), .A2(n8970), .ZN(n7621) );
  OR2_X1 U8825 ( .A1(n8093), .A2(n7619), .ZN(n7620) );
  NAND4_X1 U8826 ( .A1(n7623), .A2(n7622), .A3(n7621), .A4(n7620), .ZN(n9500)
         );
  NAND2_X1 U8827 ( .A1(n9500), .A2(n8927), .ZN(n7624) );
  XNOR2_X1 U8828 ( .A(n8949), .B(n7624), .ZN(n8974) );
  INV_X1 U8829 ( .A(n8949), .ZN(n7625) );
  NAND2_X1 U8830 ( .A1(n7846), .A2(n8693), .ZN(n7628) );
  AOI22_X1 U8831 ( .A1(n8685), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5856), .B2(
        n7626), .ZN(n7627) );
  XNOR2_X1 U8832 ( .A(n10023), .B(n5877), .ZN(n7661) );
  NAND2_X1 U8833 ( .A1(n8013), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7636) );
  OR2_X1 U8834 ( .A1(n5839), .A2(n7379), .ZN(n7635) );
  INV_X1 U8835 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U8836 ( .A1(n7630), .A2(n7629), .ZN(n7631) );
  NAND2_X1 U8837 ( .A1(n7645), .A2(n7631), .ZN(n8946) );
  OR2_X1 U8838 ( .A1(n8040), .A2(n8946), .ZN(n7634) );
  INV_X1 U8839 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7632) );
  OR2_X1 U8840 ( .A1(n8093), .A2(n7632), .ZN(n7633) );
  NOR2_X1 U8841 ( .A1(n8969), .A2(n8940), .ZN(n7637) );
  XNOR2_X1 U8842 ( .A(n7661), .B(n7637), .ZN(n8950) );
  INV_X1 U8843 ( .A(n7637), .ZN(n7638) );
  NAND2_X1 U8844 ( .A1(n7661), .A2(n7638), .ZN(n7639) );
  NAND2_X1 U8845 ( .A1(n8102), .A2(n8693), .ZN(n7642) );
  AOI22_X1 U8846 ( .A1(n8685), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5856), .B2(
        n7640), .ZN(n7641) );
  XNOR2_X1 U8847 ( .A(n10020), .B(n5877), .ZN(n7876) );
  NAND2_X1 U8848 ( .A1(n6133), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7651) );
  INV_X1 U8849 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7643) );
  OR2_X1 U8850 ( .A1(n5506), .A2(n7643), .ZN(n7650) );
  NAND2_X1 U8851 ( .A1(n7645), .A2(n9846), .ZN(n7646) );
  NAND2_X1 U8852 ( .A1(n7652), .A2(n7646), .ZN(n9478) );
  OR2_X1 U8853 ( .A1(n8040), .A2(n9478), .ZN(n7649) );
  OR2_X1 U8854 ( .A1(n8093), .A2(n7647), .ZN(n7648) );
  NOR2_X1 U8855 ( .A1(n9465), .A2(n8940), .ZN(n7874) );
  XNOR2_X1 U8856 ( .A(n7876), .B(n7874), .ZN(n7660) );
  INV_X1 U8857 ( .A(n8969), .ZN(n9218) );
  NAND2_X1 U8858 ( .A1(n8013), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7657) );
  OR2_X1 U8859 ( .A1(n5839), .A2(n7588), .ZN(n7656) );
  NAND2_X1 U8860 ( .A1(n7652), .A2(n9855), .ZN(n7653) );
  NAND2_X1 U8861 ( .A1(n7911), .A2(n7653), .ZN(n9459) );
  OR2_X1 U8862 ( .A1(n8040), .A2(n9459), .ZN(n7655) );
  INV_X1 U8863 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9250) );
  OR2_X1 U8864 ( .A1(n8093), .A2(n9250), .ZN(n7654) );
  NAND4_X1 U8865 ( .A1(n7657), .A2(n7656), .A3(n7655), .A4(n7654), .ZN(n9447)
         );
  AOI22_X1 U8866 ( .A1(n9218), .A2(n9499), .B1(n9501), .B2(n9447), .ZN(n9485)
         );
  NOR2_X1 U8867 ( .A1(n9485), .A2(n9148), .ZN(n7659) );
  OAI22_X1 U8868 ( .A1(n9206), .A2(n9478), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9846), .ZN(n7658) );
  AOI211_X1 U8869 ( .C1(n10020), .C2(n9171), .A(n7659), .B(n7658), .ZN(n7665)
         );
  INV_X1 U8870 ( .A(n7660), .ZN(n7663) );
  OAI22_X1 U8871 ( .A1(n7661), .A2(n9195), .B1(n8969), .B2(n9198), .ZN(n7662)
         );
  NAND3_X1 U8872 ( .A1(n8956), .A2(n7663), .A3(n7662), .ZN(n7664) );
  OAI211_X1 U8873 ( .C1(n7878), .C2(n9195), .A(n7665), .B(n7664), .ZN(P2_U3228) );
  AOI21_X1 U8874 ( .B1(n8103), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7666), .ZN(
        n7668) );
  XNOR2_X1 U8875 ( .A(n10246), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7667) );
  NOR2_X1 U8876 ( .A1(n7668), .A2(n7667), .ZN(n10238) );
  AOI211_X1 U8877 ( .C1(n7668), .C2(n7667), .A(n10238), .B(n10693), .ZN(n7677)
         );
  AOI21_X1 U8878 ( .B1(n8103), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7669), .ZN(
        n7672) );
  NAND2_X1 U8879 ( .A1(n10246), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7670) );
  OAI21_X1 U8880 ( .B1(n10246), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7670), .ZN(
        n7671) );
  NOR2_X1 U8881 ( .A1(n7672), .A2(n7671), .ZN(n10245) );
  AOI211_X1 U8882 ( .C1(n7672), .C2(n7671), .A(n10245), .B(n10701), .ZN(n7676)
         );
  INV_X1 U8883 ( .A(n10246), .ZN(n7674) );
  NAND2_X1 U8884 ( .A1(n10696), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U8885 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10125) );
  OAI211_X1 U8886 ( .C1(n7674), .C2(n10692), .A(n7673), .B(n10125), .ZN(n7675)
         );
  OR3_X1 U8887 ( .A1(n7677), .A2(n7676), .A3(n7675), .ZN(P1_U3258) );
  NAND2_X1 U8888 ( .A1(n10939), .A2(n8386), .ZN(n8758) );
  NAND2_X1 U8889 ( .A1(n8760), .A2(n8758), .ZN(n10920) );
  NAND2_X1 U8890 ( .A1(n10918), .A2(n10920), .ZN(n10917) );
  NAND2_X1 U8891 ( .A1(n10939), .A2(n9219), .ZN(n7681) );
  OR2_X1 U8892 ( .A1(n10976), .A2(n8372), .ZN(n8761) );
  NAND2_X1 U8893 ( .A1(n10976), .A2(n8372), .ZN(n8762) );
  INV_X1 U8894 ( .A(n8872), .ZN(n7682) );
  OAI21_X1 U8895 ( .B1(n5141), .B2(n7682), .A(n7769), .ZN(n10981) );
  INV_X1 U8896 ( .A(n10981), .ZN(n7694) );
  INV_X1 U8897 ( .A(n8758), .ZN(n7683) );
  NOR2_X1 U8898 ( .A1(n8872), .A2(n7683), .ZN(n7687) );
  NAND2_X1 U8899 ( .A1(n10922), .A2(n8760), .ZN(n7686) );
  INV_X1 U8900 ( .A(n7762), .ZN(n7685) );
  AOI21_X1 U8901 ( .B1(n7687), .B2(n7686), .A(n7685), .ZN(n7688) );
  OAI222_X1 U8902 ( .A1(n9468), .A2(n8975), .B1(n9466), .B2(n8386), .C1(n9486), 
        .C2(n7688), .ZN(n10979) );
  XNOR2_X1 U8903 ( .A(n10926), .B(n10976), .ZN(n10978) );
  OAI22_X1 U8904 ( .A1(n10946), .A2(n7689), .B1(n8385), .B2(n10935), .ZN(n7690) );
  AOI21_X1 U8905 ( .B1(n10976), .B2(n9427), .A(n7690), .ZN(n7691) );
  OAI21_X1 U8906 ( .B1(n10978), .B2(n9309), .A(n7691), .ZN(n7692) );
  AOI21_X1 U8907 ( .B1(n10979), .B2(n10946), .A(n7692), .ZN(n7693) );
  OAI21_X1 U8908 ( .B1(n7694), .B2(n9509), .A(n7693), .ZN(P2_U3284) );
  INV_X1 U8909 ( .A(n7695), .ZN(n7696) );
  NOR2_X1 U8910 ( .A1(n7697), .A2(n7696), .ZN(n7699) );
  NAND2_X1 U8911 ( .A1(n7699), .A2(n7698), .ZN(n7701) );
  NAND2_X1 U8912 ( .A1(n7701), .A2(n7700), .ZN(n8995) );
  NAND2_X1 U8913 ( .A1(n7702), .A2(n8487), .ZN(n7705) );
  AOI22_X1 U8914 ( .A1(n8472), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8133), .B2(
        n7703), .ZN(n7704) );
  NAND2_X1 U8915 ( .A1(n10968), .A2(n9086), .ZN(n7707) );
  NAND2_X1 U8916 ( .A1(n10232), .A2(n9085), .ZN(n7706) );
  NAND2_X1 U8917 ( .A1(n7707), .A2(n7706), .ZN(n8993) );
  NAND2_X1 U8918 ( .A1(n10968), .A2(n7122), .ZN(n7709) );
  NAND2_X1 U8919 ( .A1(n10232), .A2(n9086), .ZN(n7708) );
  NAND2_X1 U8920 ( .A1(n7709), .A2(n7708), .ZN(n7710) );
  XNOR2_X1 U8921 ( .A(n7710), .B(n9076), .ZN(n8994) );
  XOR2_X1 U8922 ( .A(n8993), .B(n8994), .Z(n7711) );
  XNOR2_X1 U8923 ( .A(n8995), .B(n7711), .ZN(n7725) );
  NAND2_X1 U8924 ( .A1(n8490), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7719) );
  OR2_X1 U8925 ( .A1(n8496), .A2(n10990), .ZN(n7718) );
  NAND2_X1 U8926 ( .A1(n7713), .A2(n7712), .ZN(n7714) );
  NAND2_X1 U8927 ( .A1(n7742), .A2(n7714), .ZN(n10160) );
  OR2_X1 U8928 ( .A1(n8209), .A2(n10160), .ZN(n7717) );
  INV_X1 U8929 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7715) );
  OR2_X1 U8930 ( .A1(n8492), .A2(n7715), .ZN(n7716) );
  NAND4_X1 U8931 ( .A1(n7719), .A2(n7718), .A3(n7717), .A4(n7716), .ZN(n10959)
         );
  INV_X1 U8932 ( .A(n10959), .ZN(n7736) );
  NOR2_X1 U8933 ( .A1(n10215), .A2(n7736), .ZN(n7720) );
  AOI211_X1 U8934 ( .C1(n10218), .C2(n10958), .A(n7721), .B(n7720), .ZN(n7722)
         );
  OAI21_X1 U8935 ( .B1(n10221), .B2(n10966), .A(n7722), .ZN(n7723) );
  AOI21_X1 U8936 ( .B1(n10968), .B2(n10223), .A(n7723), .ZN(n7724) );
  OAI21_X1 U8937 ( .B1(n7725), .B2(n10226), .A(n7724), .ZN(P1_U3222) );
  MUX2_X1 U8938 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7833), .Z(n7791) );
  INV_X1 U8939 ( .A(SI_24_), .ZN(n9568) );
  XNOR2_X1 U8940 ( .A(n7791), .B(n9568), .ZN(n7790) );
  INV_X1 U8941 ( .A(n8191), .ZN(n7760) );
  INV_X1 U8942 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7730) );
  OAI222_X1 U8943 ( .A1(n10532), .A2(n7760), .B1(P1_U3084), .B2(n7731), .C1(
        n7730), .C2(n10528), .ZN(P1_U3329) );
  NAND2_X1 U8944 ( .A1(n7732), .A2(n8487), .ZN(n7735) );
  AOI22_X1 U8945 ( .A1(n8472), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8133), .B2(
        n7733), .ZN(n7734) );
  OR2_X1 U8946 ( .A1(n10984), .A2(n7736), .ZN(n8537) );
  NAND2_X1 U8947 ( .A1(n10984), .A2(n7736), .ZN(n8436) );
  AND2_X1 U8948 ( .A1(n10907), .A2(n7738), .ZN(n8424) );
  OR2_X1 U8949 ( .A1(n10907), .A2(n7738), .ZN(n8435) );
  OR2_X1 U8950 ( .A1(n10968), .A2(n7739), .ZN(n8536) );
  INV_X1 U8951 ( .A(n8536), .ZN(n8438) );
  NAND2_X1 U8952 ( .A1(n10968), .A2(n7739), .ZN(n8535) );
  OAI21_X1 U8953 ( .B1(n7751), .B2(n7740), .A(n7855), .ZN(n7748) );
  NAND2_X1 U8954 ( .A1(n8238), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7747) );
  OR2_X1 U8955 ( .A1(n8496), .A2(n11006), .ZN(n7746) );
  NAND2_X1 U8956 ( .A1(n7742), .A2(n7741), .ZN(n7743) );
  NAND2_X1 U8957 ( .A1(n7808), .A2(n7743), .ZN(n10072) );
  OR2_X1 U8958 ( .A1(n6203), .A2(n10072), .ZN(n7745) );
  INV_X1 U8959 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7815) );
  OR2_X1 U8960 ( .A1(n6629), .A2(n7815), .ZN(n7744) );
  NAND4_X1 U8961 ( .A1(n7747), .A2(n7746), .A3(n7745), .A4(n7744), .ZN(n10231)
         );
  AOI222_X1 U8962 ( .A1(n11035), .A2(n7748), .B1(n10231), .B2(n11037), .C1(
        n10232), .C2(n11040), .ZN(n10986) );
  OAI21_X1 U8963 ( .B1(n7749), .B2(n8528), .A(n8529), .ZN(n10949) );
  NAND2_X1 U8964 ( .A1(n8536), .A2(n8535), .ZN(n10956) );
  NAND2_X1 U8965 ( .A1(n10949), .A2(n10956), .ZN(n10951) );
  NAND2_X1 U8966 ( .A1(n10968), .A2(n10232), .ZN(n7750) );
  INV_X1 U8967 ( .A(n7751), .ZN(n8652) );
  OAI21_X1 U8968 ( .B1(n7752), .B2(n8652), .A(n7822), .ZN(n10989) );
  INV_X1 U8969 ( .A(n11064), .ZN(n10971) );
  INV_X1 U8970 ( .A(n10968), .ZN(n10955) );
  AOI21_X1 U8971 ( .B1(n10952), .B2(n10984), .A(n11043), .ZN(n7753) );
  NAND2_X1 U8972 ( .A1(n7753), .A2(n7816), .ZN(n10985) );
  INV_X1 U8973 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7754) );
  OAI22_X1 U8974 ( .A1(n10795), .A2(n7754), .B1(n10160), .B2(n10786), .ZN(
        n7755) );
  AOI21_X1 U8975 ( .B1(n10984), .B2(n11060), .A(n7755), .ZN(n7756) );
  OAI21_X1 U8976 ( .B1(n10985), .B2(n11063), .A(n7756), .ZN(n7757) );
  AOI21_X1 U8977 ( .B1(n10989), .B2(n10971), .A(n7757), .ZN(n7758) );
  OAI21_X1 U8978 ( .B1(n10986), .B2(n11070), .A(n7758), .ZN(P1_U3278) );
  INV_X1 U8979 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7759) );
  OAI222_X1 U8980 ( .A1(P2_U3152), .A2(n7761), .B1(n10053), .B2(n7760), .C1(
        n7759), .C2(n9110), .ZN(P2_U3334) );
  INV_X1 U8981 ( .A(n9500), .ZN(n8366) );
  OR2_X1 U8982 ( .A1(n8370), .A2(n8975), .ZN(n8768) );
  NAND2_X1 U8983 ( .A1(n8370), .A2(n8975), .ZN(n8769) );
  NAND2_X1 U8984 ( .A1(n8768), .A2(n8769), .ZN(n7770) );
  INV_X1 U8985 ( .A(n7770), .ZN(n8873) );
  NAND3_X1 U8986 ( .A1(n7762), .A2(n7770), .A3(n8762), .ZN(n7763) );
  AND2_X1 U8987 ( .A1(n7780), .A2(n7763), .ZN(n7764) );
  OAI222_X1 U8988 ( .A1(n9468), .A2(n8366), .B1(n9466), .B2(n8372), .C1(n9486), 
        .C2(n7764), .ZN(n10996) );
  INV_X1 U8989 ( .A(n10996), .ZN(n7775) );
  OAI22_X1 U8990 ( .A1(n10946), .A2(n10675), .B1(n8367), .B2(n10935), .ZN(
        n7766) );
  OAI21_X1 U8991 ( .B1(n5140), .B2(n10994), .A(n7784), .ZN(n10995) );
  NOR2_X1 U8992 ( .A1(n10995), .A2(n9309), .ZN(n7765) );
  AOI211_X1 U8993 ( .C1(n9427), .C2(n8370), .A(n7766), .B(n7765), .ZN(n7774)
         );
  INV_X1 U8994 ( .A(n8372), .ZN(n7767) );
  OR2_X1 U8995 ( .A1(n10976), .A2(n7767), .ZN(n7768) );
  NOR2_X1 U8996 ( .A1(n7771), .A2(n7770), .ZN(n10993) );
  INV_X1 U8997 ( .A(n10993), .ZN(n7772) );
  NAND3_X1 U8998 ( .A1(n7772), .A2(n9400), .A3(n7777), .ZN(n7773) );
  OAI211_X1 U8999 ( .C1(n7775), .C2(n9504), .A(n7774), .B(n7773), .ZN(P2_U3283) );
  NAND2_X1 U9000 ( .A1(n8973), .A2(n9500), .ZN(n7776) );
  NAND2_X1 U9001 ( .A1(n7995), .A2(n7776), .ZN(n8874) );
  AOI21_X1 U9002 ( .B1(n8874), .B2(n7778), .A(n5125), .ZN(n11009) );
  AND2_X1 U9003 ( .A1(n7780), .A2(n8769), .ZN(n7781) );
  AND2_X1 U9004 ( .A1(n8874), .A2(n8769), .ZN(n7779) );
  OAI211_X1 U9005 ( .C1(n7781), .C2(n8874), .A(n8050), .B(n10923), .ZN(n7783)
         );
  OR2_X1 U9006 ( .A1(n8975), .A2(n9466), .ZN(n7782) );
  OAI211_X1 U9007 ( .C1(n8969), .C2(n9468), .A(n7783), .B(n7782), .ZN(n11014)
         );
  INV_X1 U9008 ( .A(n7784), .ZN(n7785) );
  OAI21_X1 U9009 ( .B1(n7785), .B2(n5472), .A(n9491), .ZN(n11012) );
  OAI22_X1 U9010 ( .A1(n10946), .A2(n6990), .B1(n8970), .B2(n10935), .ZN(n7786) );
  AOI21_X1 U9011 ( .B1(n8973), .B2(n9427), .A(n7786), .ZN(n7787) );
  OAI21_X1 U9012 ( .B1(n11012), .B2(n9309), .A(n7787), .ZN(n7788) );
  AOI21_X1 U9013 ( .B1(n11014), .B2(n10946), .A(n7788), .ZN(n7789) );
  OAI21_X1 U9014 ( .B1(n11009), .B2(n9509), .A(n7789), .ZN(P2_U3282) );
  INV_X1 U9015 ( .A(n7790), .ZN(n7793) );
  NAND2_X1 U9016 ( .A1(n7791), .A2(SI_24_), .ZN(n7792) );
  INV_X1 U9017 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7795) );
  INV_X1 U9018 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9892) );
  MUX2_X1 U9019 ( .A(n7795), .B(n9892), .S(n5153), .Z(n7796) );
  INV_X1 U9020 ( .A(SI_25_), .ZN(n9777) );
  NAND2_X1 U9021 ( .A1(n7796), .A2(n9777), .ZN(n7840) );
  INV_X1 U9022 ( .A(n7796), .ZN(n7797) );
  NAND2_X1 U9023 ( .A1(n7797), .A2(SI_25_), .ZN(n7798) );
  NAND2_X1 U9024 ( .A1(n7840), .A2(n7798), .ZN(n7961) );
  INV_X1 U9025 ( .A(n8203), .ZN(n7826) );
  AOI22_X1 U9026 ( .A1(n10541), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n7799), .ZN(n7800) );
  OAI21_X1 U9027 ( .B1(n7826), .B2(n10053), .A(n7800), .ZN(P2_U3333) );
  NAND2_X1 U9028 ( .A1(n7801), .A2(n8487), .ZN(n7804) );
  AOI22_X1 U9029 ( .A1(n8472), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8133), .B2(
        n7802), .ZN(n7803) );
  INV_X1 U9030 ( .A(n10231), .ZN(n10156) );
  NAND2_X1 U9031 ( .A1(n10074), .A2(n10156), .ZN(n8546) );
  NAND2_X1 U9032 ( .A1(n8544), .A2(n8546), .ZN(n8653) );
  NAND2_X1 U9033 ( .A1(n7855), .A2(n8436), .ZN(n7805) );
  XOR2_X1 U9034 ( .A(n8653), .B(n7805), .Z(n7814) );
  NAND2_X1 U9035 ( .A1(n8162), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7813) );
  INV_X1 U9036 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7806) );
  OR2_X1 U9037 ( .A1(n8492), .A2(n7806), .ZN(n7812) );
  NAND2_X1 U9038 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  NAND2_X1 U9039 ( .A1(n7858), .A2(n7809), .ZN(n10220) );
  OR2_X1 U9040 ( .A1(n8209), .A2(n10220), .ZN(n7811) );
  OR2_X1 U9041 ( .A1(n6629), .A2(n7868), .ZN(n7810) );
  NAND4_X1 U9042 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n11039)
         );
  AOI222_X1 U9043 ( .A1(n11035), .A2(n7814), .B1(n11039), .B2(n11037), .C1(
        n10959), .C2(n11040), .ZN(n11003) );
  OAI22_X1 U9044 ( .A1(n10795), .A2(n7815), .B1(n10072), .B2(n10786), .ZN(
        n7820) );
  INV_X1 U9045 ( .A(n7816), .ZN(n7818) );
  INV_X1 U9046 ( .A(n7869), .ZN(n7817) );
  OAI211_X1 U9047 ( .C1(n5390), .C2(n7818), .A(n7817), .B(n10953), .ZN(n11002)
         );
  NOR2_X1 U9048 ( .A1(n11002), .A2(n11063), .ZN(n7819) );
  AOI211_X1 U9049 ( .C1(n11060), .C2(n10074), .A(n7820), .B(n7819), .ZN(n7824)
         );
  OR2_X1 U9050 ( .A1(n10984), .A2(n10959), .ZN(n7821) );
  XNOR2_X1 U9051 ( .A(n7845), .B(n8653), .ZN(n11005) );
  NAND2_X1 U9052 ( .A1(n11005), .A2(n10971), .ZN(n7823) );
  OAI211_X1 U9053 ( .C1(n11003), .C2(n11070), .A(n7824), .B(n7823), .ZN(
        P1_U3277) );
  OAI222_X1 U9054 ( .A1(n10528), .A2(n9892), .B1(n10532), .B2(n7826), .C1(
        n7825), .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9055 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7923) );
  INV_X1 U9056 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9670) );
  MUX2_X1 U9057 ( .A(n7923), .B(n9670), .S(n7833), .Z(n7829) );
  INV_X1 U9058 ( .A(n7829), .ZN(n7827) );
  NAND2_X1 U9059 ( .A1(n7827), .A2(SI_26_), .ZN(n7957) );
  INV_X1 U9060 ( .A(n7957), .ZN(n7830) );
  OR2_X1 U9061 ( .A1(n7961), .A2(n7830), .ZN(n7828) );
  INV_X1 U9062 ( .A(SI_26_), .ZN(n9776) );
  NAND2_X1 U9063 ( .A1(n7829), .A2(n9776), .ZN(n7841) );
  AND2_X1 U9064 ( .A1(n7840), .A2(n7841), .ZN(n7965) );
  OR2_X1 U9065 ( .A1(n7830), .A2(n7965), .ZN(n7831) );
  INV_X1 U9066 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8326) );
  INV_X1 U9067 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9887) );
  MUX2_X1 U9068 ( .A(n8326), .B(n9887), .S(n7833), .Z(n7834) );
  INV_X1 U9069 ( .A(SI_27_), .ZN(n9772) );
  NAND2_X1 U9070 ( .A1(n7834), .A2(n9772), .ZN(n7964) );
  INV_X1 U9071 ( .A(n7834), .ZN(n7835) );
  NAND2_X1 U9072 ( .A1(n7835), .A2(SI_27_), .ZN(n7836) );
  INV_X1 U9073 ( .A(n8231), .ZN(n8325) );
  AOI21_X1 U9074 ( .B1(n10525), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7838), .ZN(
        n7839) );
  OAI21_X1 U9075 ( .B1(n8325), .B2(n10532), .A(n7839), .ZN(P1_U3326) );
  AND2_X1 U9076 ( .A1(n7841), .A2(n7957), .ZN(n7842) );
  INV_X1 U9077 ( .A(n8218), .ZN(n7924) );
  OAI222_X1 U9078 ( .A1(n10532), .A2(n7924), .B1(P1_U3084), .B2(n7844), .C1(
        n9670), .C2(n10528), .ZN(P1_U3327) );
  NAND2_X1 U9079 ( .A1(n7846), .A2(n8487), .ZN(n7850) );
  INV_X1 U9080 ( .A(n7847), .ZN(n7848) );
  AOI22_X1 U9081 ( .A1(n8472), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8133), .B2(
        n7848), .ZN(n7849) );
  INV_X1 U9082 ( .A(n11039), .ZN(n10068) );
  NAND2_X1 U9083 ( .A1(n10224), .A2(n10068), .ZN(n8552) );
  NAND2_X1 U9084 ( .A1(n7852), .A2(n8656), .ZN(n7853) );
  NAND2_X1 U9085 ( .A1(n8101), .A2(n7853), .ZN(n11022) );
  INV_X1 U9086 ( .A(n8436), .ZN(n8543) );
  NOR2_X1 U9087 ( .A1(n8653), .A2(n8543), .ZN(n7854) );
  XOR2_X1 U9088 ( .A(n8260), .B(n8656), .Z(n7866) );
  NAND2_X1 U9089 ( .A1(n8162), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7864) );
  INV_X1 U9090 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7856) );
  OR2_X1 U9091 ( .A1(n8492), .A2(n7856), .ZN(n7863) );
  INV_X1 U9092 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7857) );
  NAND2_X1 U9093 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U9094 ( .A1(n8111), .A2(n7859), .ZN(n10116) );
  OR2_X1 U9095 ( .A1(n6203), .A2(n10116), .ZN(n7862) );
  INV_X1 U9096 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7860) );
  OR2_X1 U9097 ( .A1(n6629), .A2(n7860), .ZN(n7861) );
  NAND4_X1 U9098 ( .A1(n7864), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n10424)
         );
  OAI22_X1 U9099 ( .A1(n10156), .A2(n10779), .B1(n10214), .B2(n10781), .ZN(
        n7865) );
  AOI21_X1 U9100 ( .B1(n7866), .B2(n11035), .A(n7865), .ZN(n7867) );
  OAI21_X1 U9101 ( .B1(n11022), .B2(n10851), .A(n7867), .ZN(n11025) );
  NAND2_X1 U9102 ( .A1(n11025), .A2(n10795), .ZN(n7873) );
  OAI22_X1 U9103 ( .A1(n10795), .A2(n7868), .B1(n10220), .B2(n10786), .ZN(
        n7871) );
  INV_X1 U9104 ( .A(n10224), .ZN(n11024) );
  OAI211_X1 U9105 ( .C1(n7869), .C2(n11024), .A(n11044), .B(n10953), .ZN(
        n11023) );
  NOR2_X1 U9106 ( .A1(n11023), .A2(n11063), .ZN(n7870) );
  AOI211_X1 U9107 ( .C1(n11060), .C2(n10224), .A(n7871), .B(n7870), .ZN(n7872)
         );
  OAI211_X1 U9108 ( .C1(n11022), .C2(n10415), .A(n7873), .B(n7872), .ZN(
        P1_U3276) );
  INV_X1 U9109 ( .A(n7874), .ZN(n7875) );
  NAND2_X1 U9110 ( .A1(n7876), .A2(n7875), .ZN(n7877) );
  NAND2_X1 U9111 ( .A1(n8107), .A2(n8693), .ZN(n7880) );
  AOI22_X1 U9112 ( .A1(n8685), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5856), .B2(
        n9244), .ZN(n7879) );
  XNOR2_X1 U9113 ( .A(n10015), .B(n5877), .ZN(n7881) );
  NAND2_X1 U9114 ( .A1(n9447), .A2(n8927), .ZN(n7882) );
  INV_X1 U9115 ( .A(n7881), .ZN(n7889) );
  INV_X1 U9116 ( .A(n7882), .ZN(n7883) );
  NAND2_X1 U9117 ( .A1(n7889), .A2(n7883), .ZN(n7886) );
  INV_X1 U9118 ( .A(n7884), .ZN(n7887) );
  AOI21_X1 U9119 ( .B1(n7887), .B2(n7886), .A(n7885), .ZN(n7888) );
  AOI21_X1 U9120 ( .B1(n7908), .B2(n7889), .A(n7888), .ZN(n7900) );
  OAI22_X1 U9121 ( .A1(n9465), .A2(n9159), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9855), .ZN(n7897) );
  NAND2_X1 U9122 ( .A1(n8013), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7895) );
  INV_X1 U9123 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7890) );
  OR2_X1 U9124 ( .A1(n5839), .A2(n7890), .ZN(n7894) );
  INV_X1 U9125 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9872) );
  XNOR2_X1 U9126 ( .A(n7911), .B(n9872), .ZN(n7918) );
  OR2_X1 U9127 ( .A1(n8040), .A2(n7918), .ZN(n7893) );
  INV_X1 U9128 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7891) );
  OR2_X1 U9129 ( .A1(n8093), .A2(n7891), .ZN(n7892) );
  OAI22_X1 U9130 ( .A1(n9467), .A2(n9161), .B1(n9206), .B2(n9459), .ZN(n7896)
         );
  AOI211_X1 U9131 ( .C1(n10015), .C2(n9171), .A(n7897), .B(n7896), .ZN(n7899)
         );
  NAND3_X1 U9132 ( .A1(n7908), .A2(n9128), .A3(n9447), .ZN(n7898) );
  OAI211_X1 U9133 ( .C1(n7900), .C2(n9195), .A(n7899), .B(n7898), .ZN(P2_U3230) );
  NAND2_X1 U9134 ( .A1(n8119), .A2(n8693), .ZN(n7902) );
  AOI22_X1 U9135 ( .A1(n8685), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5856), .B2(
        n9262), .ZN(n7901) );
  XNOR2_X1 U9136 ( .A(n10008), .B(n5877), .ZN(n7903) );
  OR2_X1 U9137 ( .A1(n9467), .A2(n8940), .ZN(n7904) );
  NAND2_X1 U9138 ( .A1(n7903), .A2(n7904), .ZN(n7926) );
  INV_X1 U9139 ( .A(n7903), .ZN(n7906) );
  INV_X1 U9140 ( .A(n7904), .ZN(n7905) );
  NAND2_X1 U9141 ( .A1(n7906), .A2(n7905), .ZN(n7928) );
  NAND2_X1 U9142 ( .A1(n7926), .A2(n7928), .ZN(n7907) );
  XNOR2_X1 U9143 ( .A(n7908), .B(n7907), .ZN(n7922) );
  NAND2_X1 U9144 ( .A1(n8013), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7917) );
  INV_X1 U9145 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n7909) );
  OR2_X1 U9146 ( .A1(n5839), .A2(n7909), .ZN(n7916) );
  INV_X1 U9147 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9836) );
  OAI21_X1 U9148 ( .B1(n7911), .B2(n9872), .A(n9836), .ZN(n7912) );
  NAND2_X1 U9149 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n7910) );
  NAND2_X1 U9150 ( .A1(n7912), .A2(n7938), .ZN(n9433) );
  OR2_X1 U9151 ( .A1(n8040), .A2(n9433), .ZN(n7915) );
  INV_X1 U9152 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7913) );
  OR2_X1 U9153 ( .A1(n8093), .A2(n7913), .ZN(n7914) );
  INV_X1 U9154 ( .A(n7918), .ZN(n9442) );
  AOI22_X1 U9155 ( .A1(n9447), .A2(n9189), .B1(n9188), .B2(n9442), .ZN(n7919)
         );
  NAND2_X1 U9156 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9255) );
  OAI211_X1 U9157 ( .C1(n9186), .C2(n9161), .A(n7919), .B(n9255), .ZN(n7920)
         );
  AOI21_X1 U9158 ( .B1(n10008), .B2(n9171), .A(n7920), .ZN(n7921) );
  OAI21_X1 U9159 ( .B1(n7922), .B2(n9195), .A(n7921), .ZN(P2_U3240) );
  OAI222_X1 U9160 ( .A1(P2_U3152), .A2(n7925), .B1(n10053), .B2(n7924), .C1(
        n7923), .C2(n9110), .ZN(P2_U3332) );
  NAND2_X1 U9161 ( .A1(n8132), .A2(n8693), .ZN(n7930) );
  AOI22_X1 U9162 ( .A1(n8685), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5819), .B2(
        n5856), .ZN(n7929) );
  XNOR2_X1 U9163 ( .A(n10005), .B(n8941), .ZN(n7934) );
  INV_X1 U9164 ( .A(n7934), .ZN(n7932) );
  NOR2_X1 U9165 ( .A1(n9186), .A2(n8940), .ZN(n7933) );
  INV_X1 U9166 ( .A(n7933), .ZN(n7931) );
  AND2_X1 U9167 ( .A1(n7934), .A2(n7933), .ZN(n8327) );
  NOR2_X1 U9168 ( .A1(n5139), .A2(n8327), .ZN(n7935) );
  XNOR2_X1 U9169 ( .A(n8328), .B(n7935), .ZN(n7948) );
  NAND2_X1 U9170 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9273) );
  OAI21_X1 U9171 ( .B1(n9467), .B2(n9159), .A(n9273), .ZN(n7946) );
  NAND2_X1 U9172 ( .A1(n8013), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7944) );
  INV_X1 U9173 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n7936) );
  OR2_X1 U9174 ( .A1(n5839), .A2(n7936), .ZN(n7943) );
  INV_X1 U9175 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U9176 ( .A1(n7938), .A2(n9650), .ZN(n7939) );
  NAND2_X1 U9177 ( .A1(n7988), .A2(n7939), .ZN(n9187) );
  OR2_X1 U9178 ( .A1(n8040), .A2(n9187), .ZN(n7942) );
  INV_X1 U9179 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7940) );
  OR2_X1 U9180 ( .A1(n8093), .A2(n7940), .ZN(n7941) );
  NAND4_X1 U9181 ( .A1(n7944), .A2(n7943), .A3(n7942), .A4(n7941), .ZN(n9394)
         );
  INV_X1 U9182 ( .A(n9394), .ZN(n9431) );
  OAI22_X1 U9183 ( .A1(n9431), .A2(n9161), .B1(n9206), .B2(n9433), .ZN(n7945)
         );
  AOI211_X1 U9184 ( .C1(n10005), .C2(n9171), .A(n7946), .B(n7945), .ZN(n7947)
         );
  OAI21_X1 U9185 ( .B1(n7948), .B2(n9195), .A(n7947), .ZN(P2_U3221) );
  AOI22_X1 U9186 ( .A1(n10679), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10682), .ZN(n7955) );
  AOI22_X1 U9187 ( .A1(n10674), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n7954) );
  INV_X1 U9188 ( .A(n5055), .ZN(n7949) );
  NAND3_X1 U9189 ( .A1(n7950), .A2(n7949), .A3(n6891), .ZN(n7951) );
  OAI211_X1 U9190 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10658), .A(n10670), .B(
        n7951), .ZN(n7952) );
  NAND2_X1 U9191 ( .A1(n7952), .A2(n10662), .ZN(n7953) );
  OAI211_X1 U9192 ( .C1(n7955), .C2(n10662), .A(n7954), .B(n7953), .ZN(
        P2_U3245) );
  OAI222_X1 U9193 ( .A1(n10528), .A2(n9679), .B1(n10532), .B2(n7956), .C1(
        n8619), .C2(P1_U3084), .ZN(P1_U3331) );
  INV_X1 U9194 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7976) );
  INV_X1 U9195 ( .A(n7964), .ZN(n7960) );
  AND2_X1 U9196 ( .A1(n7958), .A2(n7957), .ZN(n7959) );
  NOR2_X1 U9197 ( .A1(n7960), .A2(n7959), .ZN(n7967) );
  OR2_X1 U9198 ( .A1(n7961), .A2(n7967), .ZN(n7962) );
  AND2_X1 U9199 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  OR2_X1 U9200 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  MUX2_X1 U9201 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n8483), .Z(n7970) );
  INV_X1 U9202 ( .A(SI_28_), .ZN(n9564) );
  XNOR2_X1 U9203 ( .A(n7970), .B(n9564), .ZN(n8080) );
  INV_X1 U9204 ( .A(n7970), .ZN(n7971) );
  NAND2_X1 U9205 ( .A1(n7971), .A2(n9564), .ZN(n7972) );
  MUX2_X1 U9206 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n8483), .Z(n8469) );
  INV_X1 U9207 ( .A(SI_29_), .ZN(n7974) );
  XNOR2_X1 U9208 ( .A(n8469), .B(n7974), .ZN(n8467) );
  INV_X1 U9209 ( .A(n8684), .ZN(n9108) );
  OAI222_X1 U9210 ( .A1(n9110), .A2(n7976), .B1(n10053), .B2(n9108), .C1(n7975), .C2(P2_U3152), .ZN(P2_U3329) );
  NAND2_X1 U9211 ( .A1(n8231), .A2(n8693), .ZN(n7978) );
  NAND2_X1 U9212 ( .A1(n8685), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7977) );
  INV_X1 U9213 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9845) );
  INV_X1 U9214 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9620) );
  INV_X1 U9215 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9854) );
  INV_X1 U9216 ( .A(n8029), .ZN(n7980) );
  NAND2_X1 U9217 ( .A1(n7980), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8038) );
  INV_X1 U9218 ( .A(n8038), .ZN(n7981) );
  NAND2_X1 U9219 ( .A1(n7981), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8066) );
  XNOR2_X1 U9220 ( .A(n8066), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9124) );
  INV_X1 U9221 ( .A(n8040), .ZN(n8095) );
  INV_X1 U9222 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U9223 ( .A1(n6133), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7983) );
  NAND2_X1 U9224 ( .A1(n8013), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7982) );
  OAI211_X1 U9225 ( .C1(n7984), .C2(n8093), .A(n7983), .B(n7982), .ZN(n7985)
         );
  NAND2_X1 U9226 ( .A1(n9528), .A2(n9202), .ZN(n8835) );
  NAND2_X1 U9227 ( .A1(n8156), .A2(n8693), .ZN(n7987) );
  NAND2_X1 U9228 ( .A1(n8685), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U9229 ( .A1(n8013), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7994) );
  INV_X1 U9230 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9407) );
  OR2_X1 U9231 ( .A1(n5839), .A2(n9407), .ZN(n7993) );
  NAND2_X1 U9232 ( .A1(n7988), .A2(n9845), .ZN(n7989) );
  NAND2_X1 U9233 ( .A1(n8002), .A2(n7989), .ZN(n9406) );
  OR2_X1 U9234 ( .A1(n8040), .A2(n9406), .ZN(n7992) );
  INV_X1 U9235 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n7990) );
  OR2_X1 U9236 ( .A1(n8093), .A2(n7990), .ZN(n7991) );
  INV_X1 U9237 ( .A(n8346), .ZN(n9418) );
  INV_X1 U9238 ( .A(n10005), .ZN(n7996) );
  INV_X1 U9239 ( .A(n9465), .ZN(n9502) );
  NAND2_X1 U9240 ( .A1(n10023), .A2(n8969), .ZN(n9483) );
  NAND2_X1 U9241 ( .A1(n10020), .A2(n9465), .ZN(n8777) );
  NAND2_X1 U9242 ( .A1(n10015), .A2(n9447), .ZN(n8780) );
  NAND2_X1 U9243 ( .A1(n9453), .A2(n8781), .ZN(n9438) );
  XNOR2_X1 U9244 ( .A(n10008), .B(n9467), .ZN(n9445) );
  INV_X1 U9245 ( .A(n10008), .ZN(n9444) );
  NAND2_X1 U9246 ( .A1(n10005), .A2(n9186), .ZN(n8788) );
  NAND2_X1 U9247 ( .A1(n8789), .A2(n8788), .ZN(n9424) );
  NAND2_X1 U9248 ( .A1(n8145), .A2(n8693), .ZN(n7998) );
  NAND2_X1 U9249 ( .A1(n8685), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7997) );
  NOR2_X1 U9250 ( .A1(n9998), .A2(n9394), .ZN(n8798) );
  NAND2_X1 U9251 ( .A1(n9993), .A2(n8346), .ZN(n8807) );
  NAND2_X1 U9252 ( .A1(n8804), .A2(n8807), .ZN(n9398) );
  NAND2_X1 U9253 ( .A1(n8167), .A2(n8693), .ZN(n8000) );
  NAND2_X1 U9254 ( .A1(n8685), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U9255 ( .A1(n8013), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8008) );
  INV_X1 U9256 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8001) );
  OR2_X1 U9257 ( .A1(n5839), .A2(n8001), .ZN(n8007) );
  INV_X1 U9258 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U9259 ( .A1(n8002), .A2(n9867), .ZN(n8003) );
  NAND2_X1 U9260 ( .A1(n8011), .A2(n8003), .ZN(n8345) );
  OR2_X1 U9261 ( .A1(n8040), .A2(n8345), .ZN(n8006) );
  INV_X1 U9262 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8004) );
  OR2_X1 U9263 ( .A1(n8093), .A2(n8004), .ZN(n8005) );
  NAND2_X1 U9264 ( .A1(n9554), .A2(n9216), .ZN(n8808) );
  NAND2_X1 U9265 ( .A1(n8811), .A2(n8808), .ZN(n9386) );
  INV_X1 U9266 ( .A(n9554), .ZN(n9385) );
  NAND2_X1 U9267 ( .A1(n8178), .A2(n8693), .ZN(n8010) );
  NAND2_X1 U9268 ( .A1(n8685), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U9269 ( .A1(n8011), .A2(n9620), .ZN(n8012) );
  NAND2_X1 U9270 ( .A1(n8020), .A2(n8012), .ZN(n9372) );
  OR2_X1 U9271 ( .A1(n9372), .A2(n8040), .ZN(n8017) );
  NAND2_X1 U9272 ( .A1(n8013), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U9273 ( .A1(n6133), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U9274 ( .A1(n6134), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U9275 ( .A1(n9549), .A2(n9160), .ZN(n8815) );
  NAND2_X1 U9276 ( .A1(n8817), .A2(n8815), .ZN(n9369) );
  INV_X1 U9277 ( .A(n9549), .ZN(n9375) );
  NAND2_X1 U9278 ( .A1(n9371), .A2(n5696), .ZN(n9351) );
  NAND2_X1 U9279 ( .A1(n8191), .A2(n8693), .ZN(n8019) );
  NAND2_X1 U9280 ( .A1(n8685), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U9281 ( .A1(n8020), .A2(n9854), .ZN(n8021) );
  NAND2_X1 U9282 ( .A1(n8029), .A2(n8021), .ZN(n9158) );
  AOI22_X1 U9283 ( .A1(n8013), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n6133), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8023) );
  NAND2_X1 U9284 ( .A1(n6134), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8022) );
  OAI211_X1 U9285 ( .C1(n9158), .C2(n8040), .A(n8023), .B(n8022), .ZN(n9367)
         );
  NAND2_X1 U9286 ( .A1(n9543), .A2(n8024), .ZN(n8816) );
  NAND2_X1 U9287 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  NAND2_X1 U9288 ( .A1(n8203), .A2(n8693), .ZN(n8028) );
  NAND2_X1 U9289 ( .A1(n8685), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8027) );
  INV_X1 U9290 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U9291 ( .A1(n8029), .A2(n9634), .ZN(n8030) );
  AND2_X1 U9292 ( .A1(n8038), .A2(n8030), .ZN(n9343) );
  NAND2_X1 U9293 ( .A1(n9343), .A2(n8095), .ZN(n8033) );
  AOI22_X1 U9294 ( .A1(n6134), .A2(P2_REG1_REG_25__SCAN_IN), .B1(n6133), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U9295 ( .A1(n8013), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U9296 ( .A1(n9540), .A2(n9203), .ZN(n8825) );
  INV_X1 U9297 ( .A(n9203), .ZN(n9360) );
  NAND2_X1 U9298 ( .A1(n8218), .A2(n8693), .ZN(n8037) );
  NAND2_X1 U9299 ( .A1(n8685), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8036) );
  INV_X1 U9300 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U9301 ( .A1(n8038), .A2(n9877), .ZN(n8039) );
  NAND2_X1 U9302 ( .A1(n8066), .A2(n8039), .ZN(n9319) );
  OR2_X1 U9303 ( .A1(n9319), .A2(n8040), .ZN(n8046) );
  INV_X1 U9304 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U9305 ( .A1(n6133), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U9306 ( .A1(n8013), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8041) );
  OAI211_X1 U9307 ( .C1(n8093), .C2(n8043), .A(n8042), .B(n8041), .ZN(n8044)
         );
  INV_X1 U9308 ( .A(n8044), .ZN(n8045) );
  NAND2_X1 U9309 ( .A1(n8046), .A2(n8045), .ZN(n9215) );
  NAND2_X1 U9310 ( .A1(n9322), .A2(n9215), .ZN(n8829) );
  NAND2_X1 U9311 ( .A1(n9534), .A2(n9121), .ZN(n8060) );
  NAND2_X1 U9312 ( .A1(n8829), .A2(n8060), .ZN(n9324) );
  XOR2_X1 U9313 ( .A(n9292), .B(n9294), .Z(n9532) );
  INV_X1 U9314 ( .A(n9540), .ZN(n9346) );
  OR2_X1 U9315 ( .A1(n9491), .A2(n10023), .ZN(n9476) );
  OR2_X2 U9316 ( .A1(n9476), .A2(n10020), .ZN(n9474) );
  INV_X1 U9317 ( .A(n9993), .ZN(n9405) );
  NAND2_X1 U9318 ( .A1(n9401), .A2(n9405), .ZN(n9402) );
  NOR2_X1 U9319 ( .A1(n9549), .A2(n9381), .ZN(n9352) );
  NAND2_X1 U9320 ( .A1(n9346), .A2(n9353), .ZN(n9340) );
  INV_X1 U9321 ( .A(n9318), .ZN(n8047) );
  AOI21_X1 U9322 ( .B1(n9528), .B2(n8047), .A(n8085), .ZN(n9529) );
  AOI22_X1 U9323 ( .A1(n9124), .A2(n9492), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9426), .ZN(n8048) );
  OAI21_X1 U9324 ( .B1(n9127), .B2(n9495), .A(n8048), .ZN(n8077) );
  OR2_X1 U9325 ( .A1(n8973), .A2(n8366), .ZN(n8049) );
  INV_X1 U9326 ( .A(n8706), .ZN(n9482) );
  OAI211_X1 U9327 ( .C1(n9498), .C2(n9482), .A(n8777), .B(n9483), .ZN(n8051)
         );
  NAND2_X1 U9328 ( .A1(n8051), .A2(n8776), .ZN(n9463) );
  INV_X1 U9329 ( .A(n9454), .ZN(n9462) );
  INV_X1 U9330 ( .A(n9447), .ZN(n8052) );
  OR2_X1 U9331 ( .A1(n10015), .A2(n8052), .ZN(n8053) );
  INV_X1 U9332 ( .A(n9424), .ZN(n9428) );
  NAND2_X1 U9333 ( .A1(n9429), .A2(n9428), .ZN(n8054) );
  NAND2_X1 U9334 ( .A1(n9998), .A2(n9431), .ZN(n8055) );
  INV_X1 U9335 ( .A(n8807), .ZN(n8056) );
  INV_X1 U9336 ( .A(n9386), .ZN(n9379) );
  INV_X1 U9337 ( .A(n9357), .ZN(n8058) );
  NAND2_X1 U9338 ( .A1(n9335), .A2(n9333), .ZN(n8059) );
  AND2_X1 U9339 ( .A1(n8829), .A2(n9323), .ZN(n8827) );
  NAND2_X1 U9340 ( .A1(n9337), .A2(n8827), .ZN(n8062) );
  NAND2_X1 U9341 ( .A1(n8062), .A2(n8060), .ZN(n8064) );
  INV_X1 U9342 ( .A(n8060), .ZN(n8830) );
  NOR2_X1 U9343 ( .A1(n9292), .A2(n8830), .ZN(n8061) );
  NAND2_X1 U9344 ( .A1(n8062), .A2(n8061), .ZN(n8088) );
  INV_X1 U9345 ( .A(n8088), .ZN(n8063) );
  AOI211_X1 U9346 ( .C1(n9292), .C2(n8064), .A(n9486), .B(n8063), .ZN(n8075)
         );
  INV_X1 U9347 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9120) );
  INV_X1 U9348 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9837) );
  OAI21_X1 U9349 ( .B1(n8066), .B2(n9120), .A(n9837), .ZN(n8067) );
  NAND2_X1 U9350 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8065) );
  OR2_X1 U9351 ( .A1(n8066), .A2(n8065), .ZN(n8089) );
  NAND2_X1 U9352 ( .A1(n8907), .A2(n8095), .ZN(n8073) );
  INV_X1 U9353 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8070) );
  NAND2_X1 U9354 ( .A1(n6133), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U9355 ( .A1(n8013), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8068) );
  OAI211_X1 U9356 ( .C1(n8070), .C2(n8093), .A(n8069), .B(n8068), .ZN(n8071)
         );
  INV_X1 U9357 ( .A(n8071), .ZN(n8072) );
  OAI22_X1 U9358 ( .A1(n9308), .A2(n9468), .B1(n9121), .B2(n9466), .ZN(n8074)
         );
  NOR2_X1 U9359 ( .A1(n8075), .A2(n8074), .ZN(n9531) );
  NOR2_X1 U9360 ( .A1(n9531), .A2(n9504), .ZN(n8076) );
  AOI211_X1 U9361 ( .C1(n9507), .C2(n9529), .A(n8077), .B(n8076), .ZN(n8078)
         );
  OAI21_X1 U9362 ( .B1(n9532), .B2(n9509), .A(n8078), .ZN(P2_U3269) );
  NAND2_X1 U9363 ( .A1(n9127), .A2(n9202), .ZN(n9297) );
  NAND2_X1 U9364 ( .A1(n8079), .A2(n9297), .ZN(n8084) );
  NAND2_X1 U9365 ( .A1(n8392), .A2(n8693), .ZN(n8083) );
  NAND2_X1 U9366 ( .A1(n8685), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8082) );
  INV_X1 U9367 ( .A(n8085), .ZN(n8086) );
  INV_X1 U9368 ( .A(n9523), .ZN(n8839) );
  AOI21_X1 U9369 ( .B1(n9523), .B2(n8086), .A(n5078), .ZN(n9524) );
  AOI22_X1 U9370 ( .A1(n8907), .A2(n9492), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9426), .ZN(n8087) );
  OAI21_X1 U9371 ( .B1(n8839), .B2(n9495), .A(n8087), .ZN(n8098) );
  NAND2_X1 U9372 ( .A1(n8088), .A2(n8836), .ZN(n8683) );
  XNOR2_X1 U9373 ( .A(n8683), .B(n9290), .ZN(n8096) );
  INV_X1 U9374 ( .A(n8089), .ZN(n9310) );
  INV_X1 U9375 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U9376 ( .A1(n8013), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8091) );
  NAND2_X1 U9377 ( .A1(n6133), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8090) );
  OAI211_X1 U9378 ( .C1(n8093), .C2(n8092), .A(n8091), .B(n8090), .ZN(n8094)
         );
  AOI21_X1 U9379 ( .B1(n9310), .B2(n8095), .A(n8094), .ZN(n8909) );
  INV_X1 U9380 ( .A(n8909), .ZN(n9213) );
  INV_X1 U9381 ( .A(n9202), .ZN(n9214) );
  AOI211_X1 U9382 ( .C1(n9507), .C2(n9524), .A(n8098), .B(n8097), .ZN(n8099)
         );
  OAI21_X1 U9383 ( .B1(n9527), .B2(n9509), .A(n8099), .ZN(P2_U3268) );
  INV_X1 U9384 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U9385 ( .A1(n10224), .A2(n11039), .ZN(n8100) );
  NAND2_X1 U9386 ( .A1(n8102), .A2(n8487), .ZN(n8105) );
  AOI22_X1 U9387 ( .A1(n8472), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8133), .B2(
        n8103), .ZN(n8104) );
  NAND2_X1 U9388 ( .A1(n11061), .A2(n10214), .ZN(n8556) );
  NAND2_X1 U9389 ( .A1(n8555), .A2(n8556), .ZN(n11033) );
  NAND2_X1 U9390 ( .A1(n11061), .A2(n10424), .ZN(n8106) );
  NAND2_X1 U9391 ( .A1(n8107), .A2(n8487), .ZN(n8109) );
  AOI22_X1 U9392 ( .A1(n8472), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8133), .B2(
        n10246), .ZN(n8108) );
  NAND2_X1 U9393 ( .A1(n8162), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8117) );
  INV_X1 U9394 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10433) );
  OR2_X1 U9395 ( .A1(n6629), .A2(n10433), .ZN(n8116) );
  NAND2_X1 U9396 ( .A1(n8111), .A2(n8110), .ZN(n8112) );
  NAND2_X1 U9397 ( .A1(n8123), .A2(n8112), .ZN(n10432) );
  OR2_X1 U9398 ( .A1(n6203), .A2(n10432), .ZN(n8115) );
  INV_X1 U9399 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n8113) );
  OR2_X1 U9400 ( .A1(n8492), .A2(n8113), .ZN(n8114) );
  NAND4_X1 U9401 ( .A1(n8117), .A2(n8116), .A3(n8115), .A4(n8114), .ZN(n11038)
         );
  INV_X1 U9402 ( .A(n11038), .ZN(n10400) );
  NAND2_X1 U9403 ( .A1(n10500), .A2(n10400), .ZN(n8560) );
  NAND2_X1 U9404 ( .A1(n8559), .A2(n8560), .ZN(n10420) );
  OR2_X1 U9405 ( .A1(n10500), .A2(n11038), .ZN(n8118) );
  NAND2_X1 U9406 ( .A1(n10419), .A2(n8118), .ZN(n10403) );
  NAND2_X1 U9407 ( .A1(n8119), .A2(n8487), .ZN(n8121) );
  AOI22_X1 U9408 ( .A1(n8472), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8133), .B2(
        n10259), .ZN(n8120) );
  INV_X1 U9409 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U9410 ( .A1(n8123), .A2(n8122), .ZN(n8124) );
  NAND2_X1 U9411 ( .A1(n8149), .A2(n8124), .ZN(n10411) );
  OR2_X1 U9412 ( .A1(n10411), .A2(n8209), .ZN(n8129) );
  NAND2_X1 U9413 ( .A1(n8490), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8128) );
  INV_X1 U9414 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10237) );
  OR2_X1 U9415 ( .A1(n8496), .A2(n10237), .ZN(n8127) );
  INV_X1 U9416 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8125) );
  OR2_X1 U9417 ( .A1(n8492), .A2(n8125), .ZN(n8126) );
  NAND4_X1 U9418 ( .A1(n8129), .A2(n8128), .A3(n8127), .A4(n8126), .ZN(n10425)
         );
  INV_X1 U9419 ( .A(n10425), .ZN(n8130) );
  OR2_X1 U9420 ( .A1(n10494), .A2(n8130), .ZN(n8562) );
  NAND2_X1 U9421 ( .A1(n10494), .A2(n8130), .ZN(n8563) );
  NAND2_X1 U9422 ( .A1(n10494), .A2(n10425), .ZN(n8131) );
  NAND2_X1 U9423 ( .A1(n8132), .A2(n8487), .ZN(n8135) );
  AOI22_X1 U9424 ( .A1(n8472), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10789), 
        .B2(n8133), .ZN(n8134) );
  NAND2_X2 U9425 ( .A1(n8135), .A2(n8134), .ZN(n10489) );
  INV_X1 U9426 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U9427 ( .A1(n8238), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U9428 ( .A1(n8162), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8136) );
  OAI211_X1 U9429 ( .C1(n6629), .C2(n8138), .A(n8137), .B(n8136), .ZN(n8139)
         );
  INV_X1 U9430 ( .A(n8139), .ZN(n8141) );
  XNOR2_X1 U9431 ( .A(n8149), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n10386) );
  NAND2_X1 U9432 ( .A1(n10386), .A2(n8254), .ZN(n8140) );
  NAND2_X1 U9433 ( .A1(n8141), .A2(n8140), .ZN(n10376) );
  OR2_X1 U9434 ( .A1(n10489), .A2(n10376), .ZN(n8142) );
  NAND2_X1 U9435 ( .A1(n10489), .A2(n10376), .ZN(n8143) );
  NAND2_X1 U9436 ( .A1(n8144), .A2(n8143), .ZN(n10365) );
  NAND2_X1 U9437 ( .A1(n8145), .A2(n8487), .ZN(n8147) );
  NAND2_X1 U9438 ( .A1(n8472), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8146) );
  NAND2_X2 U9439 ( .A1(n8147), .A2(n8146), .ZN(n10484) );
  INV_X1 U9440 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8155) );
  INV_X1 U9441 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10091) );
  INV_X1 U9442 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8148) );
  OAI21_X1 U9443 ( .B1(n8149), .B2(n10091), .A(n8148), .ZN(n8150) );
  NAND2_X1 U9444 ( .A1(n8150), .A2(n8160), .ZN(n10368) );
  OR2_X1 U9445 ( .A1(n10368), .A2(n8209), .ZN(n8154) );
  NAND2_X1 U9446 ( .A1(n8490), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U9447 ( .A1(n8162), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8151) );
  AND2_X1 U9448 ( .A1(n8152), .A2(n8151), .ZN(n8153) );
  OAI211_X1 U9449 ( .C1(n8492), .C2(n8155), .A(n8154), .B(n8153), .ZN(n10394)
         );
  XNOR2_X1 U9450 ( .A(n10484), .B(n10394), .ZN(n10373) );
  NAND2_X1 U9451 ( .A1(n8156), .A2(n8487), .ZN(n8158) );
  NAND2_X1 U9452 ( .A1(n8472), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8157) );
  INV_X1 U9453 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8165) );
  INV_X1 U9454 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U9455 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  NAND2_X1 U9456 ( .A1(n8170), .A2(n8161), .ZN(n10361) );
  OR2_X1 U9457 ( .A1(n10361), .A2(n8209), .ZN(n8164) );
  AOI22_X1 U9458 ( .A1(n8162), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n8490), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n8163) );
  OAI211_X1 U9459 ( .C1(n8492), .C2(n8165), .A(n8164), .B(n8163), .ZN(n10375)
         );
  INV_X1 U9460 ( .A(n10375), .ZN(n8166) );
  NAND2_X1 U9461 ( .A1(n10479), .A2(n8166), .ZN(n8571) );
  NAND2_X1 U9462 ( .A1(n8167), .A2(n8487), .ZN(n8169) );
  NAND2_X1 U9463 ( .A1(n8472), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U9464 ( .A1(n8170), .A2(n10167), .ZN(n8171) );
  NAND2_X1 U9465 ( .A1(n8182), .A2(n8171), .ZN(n10339) );
  OR2_X1 U9466 ( .A1(n10339), .A2(n8209), .ZN(n8177) );
  INV_X1 U9467 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U9468 ( .A1(n8490), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8173) );
  NAND2_X1 U9469 ( .A1(n8238), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8172) );
  OAI211_X1 U9470 ( .C1(n8496), .C2(n8174), .A(n8173), .B(n8172), .ZN(n8175)
         );
  INV_X1 U9471 ( .A(n8175), .ZN(n8176) );
  NAND2_X1 U9472 ( .A1(n8177), .A2(n8176), .ZN(n10356) );
  NAND2_X1 U9473 ( .A1(n8178), .A2(n8487), .ZN(n8180) );
  NAND2_X1 U9474 ( .A1(n8472), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U9475 ( .A1(n8182), .A2(n8181), .ZN(n8183) );
  AND2_X1 U9476 ( .A1(n8195), .A2(n8183), .ZN(n10331) );
  NAND2_X1 U9477 ( .A1(n10331), .A2(n8254), .ZN(n8189) );
  INV_X1 U9478 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U9479 ( .A1(n8490), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U9480 ( .A1(n8238), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8184) );
  OAI211_X1 U9481 ( .C1(n8496), .C2(n8186), .A(n8185), .B(n8184), .ZN(n8187)
         );
  INV_X1 U9482 ( .A(n8187), .ZN(n8188) );
  NAND2_X1 U9483 ( .A1(n8189), .A2(n8188), .ZN(n10346) );
  NAND2_X1 U9484 ( .A1(n10469), .A2(n10346), .ZN(n8190) );
  NAND2_X1 U9485 ( .A1(n8472), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8192) );
  INV_X1 U9486 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U9487 ( .A1(n8195), .A2(n8194), .ZN(n8196) );
  NAND2_X1 U9488 ( .A1(n8207), .A2(n8196), .ZN(n10136) );
  OR2_X1 U9489 ( .A1(n10136), .A2(n6203), .ZN(n8202) );
  INV_X1 U9490 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U9491 ( .A1(n8490), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U9492 ( .A1(n8238), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8197) );
  OAI211_X1 U9493 ( .C1(n8496), .C2(n8199), .A(n8198), .B(n8197), .ZN(n8200)
         );
  INV_X1 U9494 ( .A(n8200), .ZN(n8201) );
  NAND2_X1 U9495 ( .A1(n8203), .A2(n8487), .ZN(n8205) );
  NAND2_X1 U9496 ( .A1(n8472), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8204) );
  INV_X1 U9497 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U9498 ( .A1(n8207), .A2(n8206), .ZN(n8208) );
  NAND2_X1 U9499 ( .A1(n8222), .A2(n8208), .ZN(n10311) );
  OR2_X1 U9500 ( .A1(n10311), .A2(n8209), .ZN(n8215) );
  INV_X1 U9501 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U9502 ( .A1(n8490), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U9503 ( .A1(n8238), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8210) );
  OAI211_X1 U9504 ( .C1(n8496), .C2(n8212), .A(n8211), .B(n8210), .ZN(n8213)
         );
  INV_X1 U9505 ( .A(n8213), .ZN(n8214) );
  INV_X1 U9506 ( .A(n10230), .ZN(n10294) );
  NAND2_X1 U9507 ( .A1(n10459), .A2(n10294), .ZN(n8590) );
  NAND2_X1 U9508 ( .A1(n8591), .A2(n8590), .ZN(n8585) );
  NAND2_X1 U9509 ( .A1(n10306), .A2(n8585), .ZN(n8217) );
  OR2_X1 U9510 ( .A1(n10230), .A2(n10459), .ZN(n8216) );
  NAND2_X1 U9511 ( .A1(n8472), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U9512 ( .A1(n8222), .A2(n8221), .ZN(n8223) );
  NAND2_X1 U9513 ( .A1(n10300), .A2(n8254), .ZN(n8229) );
  INV_X1 U9514 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U9515 ( .A1(n8490), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U9516 ( .A1(n8238), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8224) );
  OAI211_X1 U9517 ( .C1(n8496), .C2(n8226), .A(n8225), .B(n8224), .ZN(n8227)
         );
  INV_X1 U9518 ( .A(n8227), .ZN(n8228) );
  NOR2_X1 U9519 ( .A1(n10454), .A2(n10318), .ZN(n8230) );
  INV_X1 U9520 ( .A(n10454), .ZN(n10302) );
  NAND2_X1 U9521 ( .A1(n8472), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8232) );
  INV_X1 U9522 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8234) );
  NAND2_X1 U9523 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  NAND2_X1 U9524 ( .A1(n8248), .A2(n8236), .ZN(n10281) );
  INV_X1 U9525 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U9526 ( .A1(n8490), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U9527 ( .A1(n8238), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8239) );
  OAI211_X1 U9528 ( .C1(n8496), .C2(n8241), .A(n8240), .B(n8239), .ZN(n8242)
         );
  INV_X1 U9529 ( .A(n8242), .ZN(n8243) );
  NAND2_X1 U9530 ( .A1(n10449), .A2(n10295), .ZN(n8597) );
  NAND2_X1 U9531 ( .A1(n8392), .A2(n8487), .ZN(n8246) );
  NAND2_X1 U9532 ( .A1(n8472), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U9533 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  NAND2_X1 U9534 ( .A1(n8490), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U9535 ( .A1(n8238), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8251) );
  OAI211_X1 U9536 ( .C1(n8496), .C2(n8274), .A(n8252), .B(n8251), .ZN(n8253)
         );
  OR2_X1 U9537 ( .A1(n9099), .A2(n10058), .ZN(n8462) );
  NAND2_X1 U9538 ( .A1(n8255), .A2(n8662), .ZN(n8303) );
  NAND2_X1 U9539 ( .A1(n8303), .A2(n8256), .ZN(n8259) );
  NAND2_X1 U9540 ( .A1(n9099), .A2(n10908), .ZN(n8258) );
  INV_X1 U9541 ( .A(n10449), .ZN(n10284) );
  INV_X1 U9542 ( .A(n10459), .ZN(n10314) );
  INV_X1 U9543 ( .A(n10474), .ZN(n10342) );
  INV_X1 U9544 ( .A(n10494), .ZN(n10414) );
  INV_X1 U9545 ( .A(n10489), .ZN(n10388) );
  AOI21_X1 U9546 ( .B1(n10279), .B2(n9099), .A(n11043), .ZN(n8257) );
  NAND2_X1 U9547 ( .A1(n8257), .A2(n8309), .ZN(n8901) );
  OAI211_X1 U9548 ( .C1(n8259), .C2(n10911), .A(n8258), .B(n8901), .ZN(n8273)
         );
  NAND2_X1 U9549 ( .A1(n8260), .A2(n8656), .ZN(n8261) );
  INV_X1 U9550 ( .A(n11033), .ZN(n8655) );
  INV_X1 U9551 ( .A(n10420), .ZN(n10422) );
  INV_X1 U9552 ( .A(n10376), .ZN(n10401) );
  OR2_X1 U9553 ( .A1(n10489), .A2(n10401), .ZN(n8568) );
  NAND2_X1 U9554 ( .A1(n10489), .A2(n10401), .ZN(n8567) );
  NAND2_X1 U9555 ( .A1(n8562), .A2(n8559), .ZN(n8263) );
  AND2_X1 U9556 ( .A1(n8263), .A2(n8563), .ZN(n8447) );
  NOR2_X1 U9557 ( .A1(n10381), .A2(n8447), .ZN(n8264) );
  INV_X1 U9558 ( .A(n10394), .ZN(n10093) );
  NAND2_X1 U9559 ( .A1(n10354), .A2(n10355), .ZN(n10353) );
  NAND2_X1 U9560 ( .A1(n10353), .A2(n8571), .ZN(n10344) );
  INV_X1 U9561 ( .A(n10356), .ZN(n10082) );
  NAND2_X1 U9562 ( .A1(n10344), .A2(n10345), .ZN(n10343) );
  NAND2_X1 U9563 ( .A1(n10343), .A2(n8577), .ZN(n10325) );
  INV_X1 U9564 ( .A(n10346), .ZN(n10168) );
  OR2_X1 U9565 ( .A1(n10469), .A2(n10168), .ZN(n8453) );
  NAND2_X1 U9566 ( .A1(n10469), .A2(n10168), .ZN(n8419) );
  NAND2_X1 U9567 ( .A1(n10325), .A2(n10326), .ZN(n10324) );
  NAND2_X1 U9568 ( .A1(n10324), .A2(n8419), .ZN(n8281) );
  INV_X1 U9569 ( .A(n10327), .ZN(n8265) );
  NAND2_X1 U9570 ( .A1(n10464), .A2(n8265), .ZN(n8587) );
  NAND2_X1 U9571 ( .A1(n8281), .A2(n8660), .ZN(n8280) );
  NAND2_X1 U9572 ( .A1(n8280), .A2(n8587), .ZN(n10316) );
  NAND2_X1 U9573 ( .A1(n10316), .A2(n10317), .ZN(n10315) );
  NAND2_X1 U9574 ( .A1(n10315), .A2(n8590), .ZN(n10293) );
  NAND2_X1 U9575 ( .A1(n10293), .A2(n10296), .ZN(n10292) );
  NAND2_X1 U9576 ( .A1(n8629), .A2(n8597), .ZN(n10277) );
  INV_X1 U9577 ( .A(n10285), .ZN(n8266) );
  NOR2_X1 U9578 ( .A1(n10277), .A2(n8266), .ZN(n8267) );
  NAND2_X1 U9579 ( .A1(n10292), .A2(n8267), .ZN(n8268) );
  INV_X1 U9580 ( .A(n8662), .ZN(n8598) );
  OAI21_X1 U9581 ( .B1(n5092), .B2(n8598), .A(n8313), .ZN(n8270) );
  OAI22_X1 U9582 ( .A1(n9094), .A2(n10781), .B1(n10295), .B2(n10779), .ZN(
        n8269) );
  AOI21_X1 U9583 ( .B1(n8270), .B2(n11035), .A(n8269), .ZN(n8271) );
  NOR2_X1 U9584 ( .A1(n8273), .A2(n8900), .ZN(n10507) );
  MUX2_X1 U9585 ( .A(n8274), .B(n10507), .S(n11054), .Z(n8275) );
  INV_X1 U9586 ( .A(n8275), .ZN(P1_U3551) );
  XOR2_X1 U9587 ( .A(n8660), .B(n8276), .Z(n10467) );
  AOI211_X1 U9588 ( .C1(n10464), .C2(n10329), .A(n11043), .B(n10307), .ZN(
        n10463) );
  INV_X1 U9589 ( .A(n10464), .ZN(n8279) );
  INV_X1 U9590 ( .A(n10136), .ZN(n8277) );
  AOI22_X1 U9591 ( .A1(n8277), .A2(n11059), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n11070), .ZN(n8278) );
  OAI21_X1 U9592 ( .B1(n8279), .B2(n10430), .A(n8278), .ZN(n8284) );
  OAI21_X1 U9593 ( .B1(n8660), .B2(n8281), .A(n8280), .ZN(n8282) );
  AOI222_X1 U9594 ( .A1(n11035), .A2(n8282), .B1(n10230), .B2(n11037), .C1(
        n10346), .C2(n11040), .ZN(n10466) );
  NOR2_X1 U9595 ( .A1(n10466), .A2(n11070), .ZN(n8283) );
  AOI211_X1 U9596 ( .C1(n10463), .C2(n10291), .A(n8284), .B(n8283), .ZN(n8285)
         );
  OAI21_X1 U9597 ( .B1(n11064), .B2(n10467), .A(n8285), .ZN(P1_U3267) );
  NAND2_X1 U9598 ( .A1(n8286), .A2(n8287), .ZN(n8289) );
  XNOR2_X1 U9599 ( .A(n8289), .B(n8288), .ZN(n8292) );
  AOI22_X1 U9600 ( .A1(n10218), .A2(n6803), .B1(n8300), .B2(n10223), .ZN(n8291) );
  AOI22_X1 U9601 ( .A1(n10191), .A2(n8295), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n10179), .ZN(n8290) );
  OAI211_X1 U9602 ( .C1(n8292), .C2(n10226), .A(n8291), .B(n8290), .ZN(
        P1_U3220) );
  XNOR2_X1 U9603 ( .A(n8643), .B(n8293), .ZN(n10721) );
  XNOR2_X1 U9604 ( .A(n8643), .B(n8294), .ZN(n8296) );
  AOI222_X1 U9605 ( .A1(n11035), .A2(n8296), .B1(n8295), .B2(n11037), .C1(
        n6803), .C2(n11040), .ZN(n10719) );
  INV_X1 U9606 ( .A(n10719), .ZN(n8299) );
  OAI211_X1 U9607 ( .C1(n10720), .C2(n8297), .A(n10953), .B(n10726), .ZN(
        n10718) );
  INV_X1 U9608 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10633) );
  OAI22_X1 U9609 ( .A1(n10718), .A2(n10789), .B1(n10633), .B2(n10786), .ZN(
        n8298) );
  OAI21_X1 U9610 ( .B1(n8299), .B2(n8298), .A(n10795), .ZN(n8302) );
  AOI22_X1 U9611 ( .A1(n11060), .A2(n8300), .B1(n11070), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n8301) );
  OAI211_X1 U9612 ( .C1(n11064), .C2(n10721), .A(n8302), .B(n8301), .ZN(
        P1_U3290) );
  INV_X1 U9613 ( .A(n8303), .ZN(n8305) );
  NAND2_X1 U9614 ( .A1(n8684), .A2(n8487), .ZN(n8307) );
  NAND2_X1 U9615 ( .A1(n8472), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8306) );
  NOR2_X1 U9616 ( .A1(n10444), .A2(n9094), .ZN(n8603) );
  XNOR2_X1 U9617 ( .A(n8308), .B(n8665), .ZN(n10447) );
  AOI211_X1 U9618 ( .C1(n10444), .C2(n8309), .A(n11043), .B(n10273), .ZN(
        n10443) );
  INV_X1 U9619 ( .A(n10444), .ZN(n8312) );
  AOI22_X1 U9620 ( .A1(n8310), .A2(n11059), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n11070), .ZN(n8311) );
  OAI21_X1 U9621 ( .B1(n8312), .B2(n10430), .A(n8311), .ZN(n8324) );
  INV_X1 U9622 ( .A(n10058), .ZN(n10288) );
  INV_X1 U9623 ( .A(P1_B_REG_SCAN_IN), .ZN(n8315) );
  NOR2_X1 U9624 ( .A1(n6006), .A2(n8315), .ZN(n8316) );
  NOR2_X1 U9625 ( .A1(n10781), .A2(n8316), .ZN(n10268) );
  INV_X1 U9626 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U9627 ( .A1(n8490), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8319) );
  INV_X1 U9628 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8317) );
  OR2_X1 U9629 ( .A1(n8492), .A2(n8317), .ZN(n8318) );
  OAI211_X1 U9630 ( .C1(n8496), .C2(n8320), .A(n8319), .B(n8318), .ZN(n10228)
         );
  AOI22_X1 U9631 ( .A1(n10288), .A2(n11040), .B1(n10268), .B2(n10228), .ZN(
        n8322) );
  OAI222_X1 U9632 ( .A1(n9110), .A2(n8326), .B1(n10053), .B2(n8325), .C1(n5055), .C2(P2_U3152), .ZN(P2_U3331) );
  XNOR2_X1 U9633 ( .A(n9998), .B(n8941), .ZN(n8329) );
  AND2_X1 U9634 ( .A1(n9394), .A2(n8927), .ZN(n8330) );
  NAND2_X1 U9635 ( .A1(n8329), .A2(n8330), .ZN(n8333) );
  INV_X1 U9636 ( .A(n8329), .ZN(n9138) );
  INV_X1 U9637 ( .A(n8330), .ZN(n8331) );
  NAND2_X1 U9638 ( .A1(n9138), .A2(n8331), .ZN(n8332) );
  NAND2_X1 U9639 ( .A1(n8333), .A2(n8332), .ZN(n9184) );
  XNOR2_X1 U9640 ( .A(n9993), .B(n8941), .ZN(n8342) );
  NOR2_X1 U9641 ( .A1(n8346), .A2(n8940), .ZN(n8334) );
  NAND2_X1 U9642 ( .A1(n8342), .A2(n8334), .ZN(n8339) );
  INV_X1 U9643 ( .A(n8342), .ZN(n8336) );
  INV_X1 U9644 ( .A(n8334), .ZN(n8335) );
  NAND2_X1 U9645 ( .A1(n8336), .A2(n8335), .ZN(n8337) );
  AND2_X1 U9646 ( .A1(n8339), .A2(n8337), .ZN(n9137) );
  XNOR2_X1 U9647 ( .A(n9554), .B(n5877), .ZN(n8912) );
  NOR2_X1 U9648 ( .A1(n9216), .A2(n8940), .ZN(n8910) );
  XNOR2_X1 U9649 ( .A(n8912), .B(n8910), .ZN(n8344) );
  AND2_X1 U9650 ( .A1(n8344), .A2(n8339), .ZN(n8340) );
  NAND3_X1 U9651 ( .A1(n8342), .A2(n9128), .A3(n9418), .ZN(n8343) );
  OAI21_X1 U9652 ( .B1(n8341), .B2(n9195), .A(n8343), .ZN(n8351) );
  INV_X1 U9653 ( .A(n8344), .ZN(n8350) );
  INV_X1 U9654 ( .A(n8345), .ZN(n9383) );
  AOI22_X1 U9655 ( .A1(n9188), .A2(n9383), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8348) );
  OAI22_X1 U9656 ( .A1(n9160), .A2(n9468), .B1(n8346), .B2(n9466), .ZN(n9388)
         );
  NAND2_X1 U9657 ( .A1(n9388), .A2(n9208), .ZN(n8347) );
  OAI211_X1 U9658 ( .C1(n9385), .C2(n9211), .A(n8348), .B(n8347), .ZN(n8349)
         );
  AOI21_X1 U9659 ( .B1(n8351), .B2(n8350), .A(n8349), .ZN(n8352) );
  OAI21_X1 U9660 ( .B1(n8913), .B2(n9195), .A(n8352), .ZN(P2_U3237) );
  INV_X1 U9661 ( .A(n9221), .ZN(n8356) );
  AOI22_X1 U9662 ( .A1(n9223), .A2(n9189), .B1(n9188), .B2(n8353), .ZN(n8355)
         );
  OAI211_X1 U9663 ( .C1(n8356), .C2(n9161), .A(n8355), .B(n8354), .ZN(n8362)
         );
  INV_X1 U9664 ( .A(n8967), .ZN(n8360) );
  AOI22_X1 U9665 ( .A1(n8357), .A2(n9167), .B1(n9223), .B2(n9128), .ZN(n8359)
         );
  NOR3_X1 U9666 ( .A1(n8360), .A2(n8359), .A3(n8358), .ZN(n8361) );
  AOI211_X1 U9667 ( .C1(n9171), .C2(n8363), .A(n8362), .B(n8361), .ZN(n8364)
         );
  OAI21_X1 U9668 ( .B1(n8365), .B2(n9195), .A(n8364), .ZN(P2_U3241) );
  NAND2_X1 U9669 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10668) );
  OAI21_X1 U9670 ( .B1(n8366), .B2(n9161), .A(n10668), .ZN(n8369) );
  OAI22_X1 U9671 ( .A1(n8372), .A2(n9159), .B1(n9206), .B2(n8367), .ZN(n8368)
         );
  AOI211_X1 U9672 ( .C1(n8370), .C2(n9171), .A(n8369), .B(n8368), .ZN(n8377)
         );
  INV_X1 U9673 ( .A(n8371), .ZN(n8375) );
  OAI22_X1 U9674 ( .A1(n8373), .A2(n9195), .B1(n8372), .B2(n9198), .ZN(n8374)
         );
  NAND3_X1 U9675 ( .A1(n8391), .A2(n8375), .A3(n8374), .ZN(n8376) );
  OAI211_X1 U9676 ( .C1(n8979), .C2(n9195), .A(n8377), .B(n8376), .ZN(P2_U3236) );
  NAND3_X1 U9677 ( .A1(n8378), .A2(n9128), .A3(n9219), .ZN(n8379) );
  OAI21_X1 U9678 ( .B1(n8380), .B2(n9195), .A(n8379), .ZN(n8383) );
  INV_X1 U9679 ( .A(n8381), .ZN(n8382) );
  NAND2_X1 U9680 ( .A1(n8383), .A2(n8382), .ZN(n8390) );
  OAI21_X1 U9681 ( .B1(n8975), .B2(n9161), .A(n8384), .ZN(n8388) );
  OAI22_X1 U9682 ( .A1(n8386), .A2(n9159), .B1(n9206), .B2(n8385), .ZN(n8387)
         );
  AOI211_X1 U9683 ( .C1(n10976), .C2(n9171), .A(n8388), .B(n8387), .ZN(n8389)
         );
  OAI211_X1 U9684 ( .C1(n9195), .C2(n8391), .A(n8390), .B(n8389), .ZN(P2_U3226) );
  INV_X1 U9685 ( .A(n8392), .ZN(n9105) );
  INV_X1 U9686 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8393) );
  OAI222_X1 U9687 ( .A1(n10532), .A2(n9105), .B1(n6007), .B2(P1_U3084), .C1(
        n8393), .C2(n10528), .ZN(P1_U3325) );
  OAI222_X1 U9688 ( .A1(n10528), .A2(n9683), .B1(n10532), .B2(n8394), .C1(
        n10359), .C2(P1_U3084), .ZN(P1_U3334) );
  NAND2_X1 U9689 ( .A1(n8601), .A2(n8597), .ZN(n8628) );
  AOI21_X1 U9690 ( .B1(n10732), .B2(n10720), .A(n8667), .ZN(n8399) );
  INV_X1 U9691 ( .A(n8395), .ZN(n8398) );
  INV_X1 U9692 ( .A(n8396), .ZN(n8397) );
  AOI211_X1 U9693 ( .C1(n8399), .C2(n8398), .A(n8397), .B(n10730), .ZN(n8403)
         );
  INV_X1 U9694 ( .A(n8400), .ZN(n8402) );
  OAI21_X1 U9695 ( .B1(n8403), .B2(n8402), .A(n8401), .ZN(n8405) );
  OAI211_X1 U9696 ( .C1(n8407), .C2(n8406), .A(n8405), .B(n8404), .ZN(n8410)
         );
  NAND3_X1 U9697 ( .A1(n8410), .A2(n8409), .A3(n8408), .ZN(n8413) );
  INV_X1 U9698 ( .A(n8505), .ZN(n8411) );
  AOI21_X1 U9699 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8418) );
  AND2_X1 U9700 ( .A1(n8506), .A2(n8414), .ZN(n8504) );
  INV_X1 U9701 ( .A(n8504), .ZN(n8417) );
  NAND2_X1 U9702 ( .A1(n8446), .A2(n5066), .ZN(n8415) );
  AND2_X1 U9703 ( .A1(n8415), .A2(n8571), .ZN(n8573) );
  NAND3_X1 U9704 ( .A1(n8573), .A2(n8577), .A3(n8567), .ZN(n8622) );
  INV_X1 U9705 ( .A(n8622), .ZN(n8416) );
  OAI21_X1 U9706 ( .B1(n8418), .B2(n8417), .A(n8416), .ZN(n8458) );
  AND2_X1 U9707 ( .A1(n8587), .A2(n8419), .ZN(n8582) );
  AND2_X1 U9708 ( .A1(n8590), .A2(n8582), .ZN(n8452) );
  INV_X1 U9709 ( .A(n8452), .ZN(n8431) );
  AND2_X1 U9710 ( .A1(n8560), .A2(n8556), .ZN(n8420) );
  AND2_X1 U9711 ( .A1(n8563), .A2(n8420), .ZN(n8444) );
  INV_X1 U9712 ( .A(n8444), .ZN(n8430) );
  NAND2_X1 U9713 ( .A1(n8525), .A2(n8421), .ZN(n8422) );
  NAND2_X1 U9714 ( .A1(n8422), .A2(n8526), .ZN(n8423) );
  NOR2_X1 U9715 ( .A1(n8424), .A2(n8423), .ZN(n8425) );
  AND2_X1 U9716 ( .A1(n8535), .A2(n8425), .ZN(n8426) );
  NAND2_X1 U9717 ( .A1(n8436), .A2(n8426), .ZN(n8433) );
  INV_X1 U9718 ( .A(n8433), .ZN(n8427) );
  NAND4_X1 U9719 ( .A1(n8552), .A2(n8428), .A3(n8427), .A4(n8546), .ZN(n8429)
         );
  OR3_X1 U9720 ( .A1(n8431), .A2(n8430), .A3(n8429), .ZN(n8624) );
  INV_X1 U9721 ( .A(n8432), .ZN(n8513) );
  NOR2_X1 U9722 ( .A1(n8521), .A2(n8513), .ZN(n8434) );
  AOI21_X1 U9723 ( .B1(n8434), .B2(n8525), .A(n8433), .ZN(n8441) );
  INV_X1 U9724 ( .A(n8435), .ZN(n8437) );
  OAI211_X1 U9725 ( .C1(n8438), .C2(n8437), .A(n8436), .B(n8535), .ZN(n8439)
         );
  NAND3_X1 U9726 ( .A1(n8544), .A2(n8537), .A3(n8439), .ZN(n8440) );
  OAI211_X1 U9727 ( .C1(n8441), .C2(n8440), .A(n8552), .B(n8546), .ZN(n8442)
         );
  NAND3_X1 U9728 ( .A1(n8555), .A2(n8551), .A3(n8442), .ZN(n8443) );
  NAND2_X1 U9729 ( .A1(n8444), .A2(n8443), .ZN(n8450) );
  OR2_X1 U9730 ( .A1(n10484), .A2(n10093), .ZN(n8445) );
  NAND2_X1 U9731 ( .A1(n8446), .A2(n8445), .ZN(n8572) );
  INV_X1 U9732 ( .A(n8447), .ZN(n10389) );
  OAI21_X1 U9733 ( .B1(n10389), .B2(n5490), .A(n8568), .ZN(n8448) );
  OAI211_X1 U9734 ( .C1(n8572), .C2(n8448), .A(n8573), .B(n8577), .ZN(n8449)
         );
  OAI211_X1 U9735 ( .C1(n8622), .C2(n8450), .A(n8580), .B(n8449), .ZN(n8451)
         );
  NAND2_X1 U9736 ( .A1(n8452), .A2(n8451), .ZN(n8456) );
  AND2_X1 U9737 ( .A1(n8586), .A2(n8453), .ZN(n8578) );
  INV_X1 U9738 ( .A(n8578), .ZN(n8454) );
  NAND3_X1 U9739 ( .A1(n8590), .A2(n8587), .A3(n8454), .ZN(n8455) );
  NAND4_X1 U9740 ( .A1(n8456), .A2(n8594), .A3(n8591), .A4(n8455), .ZN(n8625)
         );
  INV_X1 U9741 ( .A(n8625), .ZN(n8457) );
  OAI211_X1 U9742 ( .C1(n8458), .C2(n8624), .A(n8457), .B(n10286), .ZN(n8461)
         );
  INV_X1 U9743 ( .A(n8629), .ZN(n8459) );
  NOR2_X1 U9744 ( .A1(n8459), .A2(n10285), .ZN(n8627) );
  INV_X1 U9745 ( .A(n8627), .ZN(n8460) );
  NAND2_X1 U9746 ( .A1(n8461), .A2(n8460), .ZN(n8465) );
  INV_X1 U9747 ( .A(n8462), .ZN(n8463) );
  OR2_X1 U9748 ( .A1(n8603), .A2(n8463), .ZN(n8633) );
  INV_X1 U9749 ( .A(n8633), .ZN(n8464) );
  OAI21_X1 U9750 ( .B1(n8628), .B2(n8465), .A(n8464), .ZN(n8476) );
  INV_X1 U9751 ( .A(n8466), .ZN(n8632) );
  OR2_X1 U9752 ( .A1(n8469), .A2(SI_29_), .ZN(n8470) );
  MUX2_X1 U9753 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8483), .Z(n8479) );
  INV_X1 U9754 ( .A(SI_30_), .ZN(n9559) );
  XNOR2_X1 U9755 ( .A(n8479), .B(n9559), .ZN(n8477) );
  NAND2_X1 U9756 ( .A1(n9109), .A2(n8487), .ZN(n8474) );
  NAND2_X1 U9757 ( .A1(n8472), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8473) );
  INV_X1 U9758 ( .A(n10228), .ZN(n8475) );
  OR2_X1 U9759 ( .A1(n8609), .A2(n8475), .ZN(n8663) );
  AOI21_X1 U9760 ( .B1(n8476), .B2(n8632), .A(n5439), .ZN(n8499) );
  NAND2_X1 U9761 ( .A1(n8478), .A2(n8477), .ZN(n8482) );
  INV_X1 U9762 ( .A(n8479), .ZN(n8480) );
  NAND2_X1 U9763 ( .A1(n8480), .A2(n9559), .ZN(n8481) );
  NAND2_X1 U9764 ( .A1(n8482), .A2(n8481), .ZN(n8486) );
  MUX2_X1 U9765 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8483), .Z(n8484) );
  INV_X1 U9766 ( .A(SI_31_), .ZN(n9767) );
  XNOR2_X1 U9767 ( .A(n8484), .B(n9767), .ZN(n8485) );
  NAND2_X1 U9768 ( .A1(n10045), .A2(n8487), .ZN(n8489) );
  NAND2_X1 U9769 ( .A1(n8472), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8488) );
  INV_X1 U9770 ( .A(n10439), .ZN(n8498) );
  INV_X1 U9771 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U9772 ( .A1(n8490), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8494) );
  INV_X1 U9773 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8491) );
  OR2_X1 U9774 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  OAI211_X1 U9775 ( .C1(n8496), .C2(n8495), .A(n8494), .B(n8493), .ZN(n10269)
         );
  INV_X1 U9776 ( .A(n10269), .ZN(n8611) );
  NOR2_X1 U9777 ( .A1(n8498), .A2(n8611), .ZN(n8635) );
  INV_X1 U9778 ( .A(n8635), .ZN(n8497) );
  OAI21_X1 U9779 ( .B1(n10442), .B2(n10228), .A(n8497), .ZN(n8669) );
  NAND2_X1 U9780 ( .A1(n8498), .A2(n8611), .ZN(n8666) );
  OAI21_X1 U9781 ( .B1(n8499), .B2(n8669), .A(n8666), .ZN(n8500) );
  XNOR2_X1 U9782 ( .A(n8500), .B(n10359), .ZN(n8677) );
  INV_X1 U9783 ( .A(n8501), .ZN(n8616) );
  INV_X1 U9784 ( .A(n8613), .ZN(n8610) );
  XNOR2_X1 U9785 ( .A(n10802), .B(n8613), .ZN(n8502) );
  NAND2_X1 U9786 ( .A1(n8502), .A2(n10801), .ZN(n8509) );
  INV_X1 U9787 ( .A(n10844), .ZN(n8503) );
  AOI21_X1 U9788 ( .B1(n8509), .B2(n8504), .A(n8503), .ZN(n8511) );
  AND2_X1 U9789 ( .A1(n10844), .A2(n8505), .ZN(n8508) );
  INV_X1 U9790 ( .A(n8506), .ZN(n8507) );
  AOI21_X1 U9791 ( .B1(n8509), .B2(n8508), .A(n8507), .ZN(n8510) );
  AOI21_X1 U9792 ( .B1(n8512), .B2(n10846), .A(n8646), .ZN(n8517) );
  NOR2_X1 U9793 ( .A1(n8514), .A2(n8613), .ZN(n8516) );
  NAND3_X1 U9794 ( .A1(n8514), .A2(n8513), .A3(n8610), .ZN(n8515) );
  OAI21_X1 U9795 ( .B1(n8517), .B2(n8516), .A(n8515), .ZN(n8519) );
  NAND2_X1 U9796 ( .A1(n8521), .A2(n8613), .ZN(n8518) );
  NAND2_X1 U9797 ( .A1(n8519), .A2(n8518), .ZN(n8524) );
  OR3_X1 U9798 ( .A1(n8521), .A2(n8610), .A3(n8520), .ZN(n8523) );
  AOI21_X1 U9799 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n8534) );
  MUX2_X1 U9800 ( .A(n10958), .B(n10907), .S(n8610), .Z(n8530) );
  MUX2_X1 U9801 ( .A(n8526), .B(n8525), .S(n8610), .Z(n8527) );
  OAI21_X1 U9802 ( .B1(n8530), .B2(n8528), .A(n8527), .ZN(n8533) );
  INV_X1 U9803 ( .A(n10956), .ZN(n8532) );
  NAND2_X1 U9804 ( .A1(n8530), .A2(n8529), .ZN(n8531) );
  MUX2_X1 U9805 ( .A(n8536), .B(n8535), .S(n8613), .Z(n8539) );
  INV_X1 U9806 ( .A(n8537), .ZN(n8545) );
  MUX2_X1 U9807 ( .A(n8543), .B(n8545), .S(n8613), .Z(n8538) );
  AOI21_X1 U9808 ( .B1(n8540), .B2(n8539), .A(n8538), .ZN(n8542) );
  MUX2_X1 U9809 ( .A(n8546), .B(n8544), .S(n8613), .Z(n8541) );
  OAI21_X1 U9810 ( .B1(n8542), .B2(n8653), .A(n8541), .ZN(n8550) );
  NAND2_X1 U9811 ( .A1(n8544), .A2(n8543), .ZN(n8548) );
  NAND2_X1 U9812 ( .A1(n8546), .A2(n8545), .ZN(n8547) );
  MUX2_X1 U9813 ( .A(n8548), .B(n8547), .S(n8610), .Z(n8549) );
  NAND3_X1 U9814 ( .A1(n8550), .A2(n8656), .A3(n8549), .ZN(n8554) );
  MUX2_X1 U9815 ( .A(n8552), .B(n8551), .S(n8613), .Z(n8553) );
  NAND3_X1 U9816 ( .A1(n8554), .A2(n8655), .A3(n8553), .ZN(n8558) );
  MUX2_X1 U9817 ( .A(n8556), .B(n8555), .S(n8610), .Z(n8557) );
  AOI21_X1 U9818 ( .B1(n8558), .B2(n8557), .A(n10420), .ZN(n8566) );
  MUX2_X1 U9819 ( .A(n8560), .B(n8559), .S(n8610), .Z(n8561) );
  NAND2_X1 U9820 ( .A1(n10402), .A2(n8561), .ZN(n8565) );
  INV_X1 U9821 ( .A(n10381), .ZN(n10392) );
  MUX2_X1 U9822 ( .A(n8563), .B(n8562), .S(n8613), .Z(n8564) );
  OAI211_X1 U9823 ( .C1(n8566), .C2(n8565), .A(n10392), .B(n8564), .ZN(n8570)
         );
  MUX2_X1 U9824 ( .A(n8568), .B(n8567), .S(n8613), .Z(n8569) );
  NAND2_X1 U9825 ( .A1(n8572), .A2(n8571), .ZN(n8574) );
  NAND3_X1 U9826 ( .A1(n8576), .A2(n10345), .A3(n8575), .ZN(n8581) );
  NAND3_X1 U9827 ( .A1(n8581), .A2(n10326), .A3(n8577), .ZN(n8579) );
  NAND2_X1 U9828 ( .A1(n8579), .A2(n8578), .ZN(n8584) );
  NAND3_X1 U9829 ( .A1(n8581), .A2(n10326), .A3(n8580), .ZN(n8583) );
  MUX2_X1 U9830 ( .A(n8587), .B(n8586), .S(n8613), .Z(n8588) );
  NAND3_X1 U9831 ( .A1(n8589), .A2(n10317), .A3(n8588), .ZN(n8593) );
  MUX2_X1 U9832 ( .A(n8591), .B(n8590), .S(n8613), .Z(n8592) );
  NAND3_X1 U9833 ( .A1(n8593), .A2(n10296), .A3(n8592), .ZN(n8596) );
  NAND3_X1 U9834 ( .A1(n8596), .A2(n10286), .A3(n8595), .ZN(n8600) );
  MUX2_X1 U9835 ( .A(n8629), .B(n8597), .S(n8613), .Z(n8599) );
  NAND3_X1 U9836 ( .A1(n8602), .A2(n8632), .A3(n8601), .ZN(n8605) );
  INV_X1 U9837 ( .A(n8603), .ZN(n8604) );
  OAI21_X1 U9838 ( .B1(n8606), .B2(n8633), .A(n8632), .ZN(n8607) );
  NAND2_X1 U9839 ( .A1(n10269), .A2(n10228), .ZN(n8608) );
  NAND2_X1 U9840 ( .A1(n8609), .A2(n8608), .ZN(n8631) );
  INV_X1 U9841 ( .A(n8666), .ZN(n8614) );
  OR2_X1 U9842 ( .A1(n8663), .A2(n8611), .ZN(n8612) );
  AND2_X1 U9843 ( .A1(n8666), .A2(n8612), .ZN(n8636) );
  NAND2_X1 U9844 ( .A1(n8619), .A2(n8618), .ZN(n8620) );
  INV_X1 U9845 ( .A(n10845), .ZN(n8623) );
  NOR3_X1 U9846 ( .A1(n8624), .A2(n8623), .A3(n8622), .ZN(n8626) );
  NOR2_X1 U9847 ( .A1(n8626), .A2(n8625), .ZN(n8630) );
  AOI211_X1 U9848 ( .C1(n8630), .C2(n8629), .A(n8628), .B(n8627), .ZN(n8634)
         );
  OAI211_X1 U9849 ( .C1(n8634), .C2(n8633), .A(n8632), .B(n8631), .ZN(n8637)
         );
  AOI211_X1 U9850 ( .C1(n8637), .C2(n8636), .A(n8667), .B(n8635), .ZN(n8638)
         );
  NOR2_X1 U9851 ( .A1(n8638), .A2(n10789), .ZN(n8671) );
  INV_X1 U9852 ( .A(n10355), .ZN(n10352) );
  AND4_X1 U9853 ( .A1(n8642), .A2(n8641), .A3(n8640), .A4(n8639), .ZN(n8644)
         );
  NAND4_X1 U9854 ( .A1(n8644), .A2(n10801), .A3(n10774), .A4(n8643), .ZN(n8647) );
  INV_X1 U9855 ( .A(n10846), .ZN(n10839) );
  NOR4_X1 U9856 ( .A1(n8647), .A2(n8646), .A3(n10839), .A4(n8645), .ZN(n8650)
         );
  NAND3_X1 U9857 ( .A1(n8650), .A2(n8649), .A3(n8648), .ZN(n8651) );
  NOR4_X1 U9858 ( .A1(n8653), .A2(n8652), .A3(n10956), .A4(n8651), .ZN(n8654)
         );
  NAND4_X1 U9859 ( .A1(n10422), .A2(n8656), .A3(n8655), .A4(n8654), .ZN(n8657)
         );
  NOR4_X1 U9860 ( .A1(n10352), .A2(n5273), .A3(n10381), .A4(n8657), .ZN(n8658)
         );
  AND4_X1 U9861 ( .A1(n10326), .A2(n10345), .A3(n8658), .A4(n10373), .ZN(n8659) );
  NAND4_X1 U9862 ( .A1(n10296), .A2(n10317), .A3(n8660), .A4(n8659), .ZN(n8661) );
  NOR3_X1 U9863 ( .A1(n8662), .A2(n10277), .A3(n8661), .ZN(n8664) );
  NAND4_X1 U9864 ( .A1(n8666), .A2(n8665), .A3(n8664), .A4(n8663), .ZN(n8668)
         );
  OAI21_X1 U9865 ( .B1(n8669), .B2(n8668), .A(n8667), .ZN(n8670) );
  MUX2_X1 U9866 ( .A(n10789), .B(n8671), .S(n8670), .Z(n8672) );
  MUX2_X1 U9867 ( .A(n8677), .B(n8676), .S(n8675), .Z(n8682) );
  NOR4_X1 U9868 ( .A1(n8678), .A2(n10521), .A3(n6007), .A4(n6006), .ZN(n8680)
         );
  OAI21_X1 U9869 ( .B1(n6465), .B2(n8681), .A(P1_B_REG_SCAN_IN), .ZN(n8679) );
  OAI22_X1 U9870 ( .A1(n8682), .A2(n8681), .B1(n8680), .B2(n8679), .ZN(
        P1_U3240) );
  NAND2_X1 U9871 ( .A1(n8684), .A2(n8693), .ZN(n8687) );
  NAND2_X1 U9872 ( .A1(n8685), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8686) );
  NAND2_X1 U9873 ( .A1(n9521), .A2(n8909), .ZN(n8845) );
  NAND2_X1 U9874 ( .A1(n9109), .A2(n8693), .ZN(n8689) );
  INV_X1 U9875 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9111) );
  OR2_X1 U9876 ( .A1(n5858), .A2(n9111), .ZN(n8688) );
  NOR2_X1 U9877 ( .A1(n9514), .A2(n9306), .ZN(n8702) );
  INV_X1 U9878 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8692) );
  INV_X1 U9879 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9282) );
  OR2_X1 U9880 ( .A1(n5839), .A2(n9282), .ZN(n8691) );
  NAND2_X1 U9881 ( .A1(n6134), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8690) );
  OAI211_X1 U9882 ( .C1(n5506), .C2(n8692), .A(n8691), .B(n8690), .ZN(n9212)
         );
  NAND2_X1 U9883 ( .A1(n10045), .A2(n8693), .ZN(n8695) );
  INV_X1 U9884 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10048) );
  OR2_X1 U9885 ( .A1(n5858), .A2(n10048), .ZN(n8694) );
  INV_X1 U9886 ( .A(n9212), .ZN(n9281) );
  OR2_X1 U9887 ( .A1(n9510), .A2(n9281), .ZN(n8696) );
  NAND2_X1 U9888 ( .A1(n9514), .A2(n9306), .ZN(n8848) );
  AND2_X1 U9889 ( .A1(n9510), .A2(n9281), .ZN(n8701) );
  XNOR2_X1 U9890 ( .A(n8698), .B(n5819), .ZN(n8699) );
  AOI21_X1 U9891 ( .B1(n8700), .B2(n8927), .A(n8699), .ZN(n8892) );
  INV_X1 U9892 ( .A(n8701), .ZN(n8703) );
  INV_X1 U9893 ( .A(n8702), .ZN(n8849) );
  AND2_X1 U9894 ( .A1(n8703), .A2(n8849), .ZN(n8882) );
  AND2_X1 U9895 ( .A1(n5819), .A2(n8887), .ZN(n8705) );
  NAND2_X1 U9896 ( .A1(n8705), .A2(n8704), .ZN(n8850) );
  MUX2_X1 U9897 ( .A(n8883), .B(n8882), .S(n8850), .Z(n8853) );
  MUX2_X1 U9898 ( .A(n8706), .B(n9483), .S(n8840), .Z(n8775) );
  INV_X1 U9899 ( .A(n8710), .ZN(n8711) );
  MUX2_X1 U9900 ( .A(n8713), .B(n8712), .S(n8840), .Z(n8714) );
  NAND2_X1 U9901 ( .A1(n8714), .A2(n8860), .ZN(n8715) );
  AOI21_X1 U9902 ( .B1(n8716), .B2(n5529), .A(n8715), .ZN(n8726) );
  MUX2_X1 U9903 ( .A(n8718), .B(n8717), .S(n8850), .Z(n8720) );
  NAND2_X1 U9904 ( .A1(n8720), .A2(n8719), .ZN(n8725) );
  AND2_X1 U9905 ( .A1(n9224), .A2(n8840), .ZN(n8722) );
  NOR2_X1 U9906 ( .A1(n9224), .A2(n8840), .ZN(n8721) );
  MUX2_X1 U9907 ( .A(n8722), .B(n8721), .S(n9170), .Z(n8723) );
  INV_X1 U9908 ( .A(n8723), .ZN(n8724) );
  OAI21_X1 U9909 ( .B1(n8726), .B2(n8725), .A(n8724), .ZN(n8728) );
  INV_X1 U9910 ( .A(n8861), .ZN(n8727) );
  NAND2_X1 U9911 ( .A1(n8728), .A2(n8727), .ZN(n8732) );
  MUX2_X1 U9912 ( .A(n8730), .B(n8729), .S(n8840), .Z(n8731) );
  NAND3_X1 U9913 ( .A1(n8732), .A2(n8865), .A3(n8731), .ZN(n8741) );
  MUX2_X1 U9914 ( .A(n8734), .B(n8733), .S(n8850), .Z(n8736) );
  NOR2_X1 U9915 ( .A1(n8736), .A2(n8735), .ZN(n8740) );
  AOI21_X1 U9916 ( .B1(n8744), .B2(n8737), .A(n8840), .ZN(n8745) );
  AOI21_X1 U9917 ( .B1(n8742), .B2(n8738), .A(n8850), .ZN(n8739) );
  AOI211_X1 U9918 ( .C1(n8741), .C2(n8740), .A(n8745), .B(n8739), .ZN(n8751)
         );
  MUX2_X1 U9919 ( .A(n8742), .B(n8746), .S(n8840), .Z(n8743) );
  OAI211_X1 U9920 ( .C1(n8745), .C2(n8744), .A(n8748), .B(n8743), .ZN(n8750)
         );
  AND2_X1 U9921 ( .A1(n8752), .A2(n8746), .ZN(n8747) );
  MUX2_X1 U9922 ( .A(n8748), .B(n8747), .S(n8850), .Z(n8749) );
  OAI211_X1 U9923 ( .C1(n8751), .C2(n8750), .A(n8753), .B(n8749), .ZN(n8757)
         );
  AND2_X1 U9924 ( .A1(n8758), .A2(n8752), .ZN(n8755) );
  AND2_X1 U9925 ( .A1(n8760), .A2(n8753), .ZN(n8754) );
  MUX2_X1 U9926 ( .A(n8755), .B(n8754), .S(n8850), .Z(n8756) );
  NAND3_X1 U9927 ( .A1(n8757), .A2(n8872), .A3(n8756), .ZN(n8767) );
  NAND2_X1 U9928 ( .A1(n8762), .A2(n8758), .ZN(n8759) );
  NAND2_X1 U9929 ( .A1(n8759), .A2(n8761), .ZN(n8765) );
  NAND2_X1 U9930 ( .A1(n8761), .A2(n8760), .ZN(n8763) );
  NAND2_X1 U9931 ( .A1(n8763), .A2(n8762), .ZN(n8764) );
  MUX2_X1 U9932 ( .A(n8765), .B(n8764), .S(n8840), .Z(n8766) );
  NAND3_X1 U9933 ( .A1(n8767), .A2(n8873), .A3(n8766), .ZN(n8771) );
  MUX2_X1 U9934 ( .A(n8769), .B(n8768), .S(n8850), .Z(n8770) );
  NAND2_X1 U9935 ( .A1(n9500), .A2(n8840), .ZN(n8773) );
  OR2_X1 U9936 ( .A1(n9500), .A2(n8840), .ZN(n8772) );
  MUX2_X1 U9937 ( .A(n8773), .B(n8772), .S(n8973), .Z(n8774) );
  MUX2_X1 U9938 ( .A(n8777), .B(n8776), .S(n8840), .Z(n8778) );
  MUX2_X1 U9939 ( .A(n9447), .B(n10015), .S(n8850), .Z(n8779) );
  INV_X1 U9940 ( .A(n8781), .ZN(n8782) );
  NAND2_X1 U9941 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  NAND2_X1 U9942 ( .A1(n8785), .A2(n8784), .ZN(n8795) );
  MUX2_X1 U9943 ( .A(n9467), .B(n9444), .S(n8840), .Z(n8796) );
  OR2_X1 U9944 ( .A1(n8795), .A2(n8796), .ZN(n8792) );
  AND2_X1 U9945 ( .A1(n8789), .A2(n10008), .ZN(n8787) );
  INV_X1 U9946 ( .A(n8788), .ZN(n8786) );
  AOI21_X1 U9947 ( .B1(n8792), .B2(n8787), .A(n8786), .ZN(n8794) );
  INV_X1 U9948 ( .A(n9467), .ZN(n9217) );
  AND2_X1 U9949 ( .A1(n8788), .A2(n9217), .ZN(n8791) );
  INV_X1 U9950 ( .A(n8789), .ZN(n8790) );
  AOI21_X1 U9951 ( .B1(n8792), .B2(n8791), .A(n8790), .ZN(n8793) );
  NAND3_X1 U9952 ( .A1(n9428), .A2(n8796), .A3(n8795), .ZN(n8797) );
  MUX2_X1 U9953 ( .A(n9394), .B(n9998), .S(n8840), .Z(n8799) );
  INV_X1 U9954 ( .A(n8799), .ZN(n8800) );
  NAND2_X1 U9955 ( .A1(n8802), .A2(n8801), .ZN(n8803) );
  AOI21_X1 U9956 ( .B1(n8811), .B2(n8804), .A(n8850), .ZN(n8805) );
  OAI21_X1 U9957 ( .B1(n8806), .B2(n8805), .A(n8808), .ZN(n8810) );
  NAND2_X1 U9958 ( .A1(n8808), .A2(n8807), .ZN(n8809) );
  AOI21_X1 U9959 ( .B1(n8817), .B2(n8811), .A(n8840), .ZN(n8813) );
  INV_X1 U9960 ( .A(n8815), .ZN(n8812) );
  NOR2_X1 U9961 ( .A1(n8813), .A2(n8812), .ZN(n8814) );
  AND2_X1 U9962 ( .A1(n8816), .A2(n8815), .ZN(n8819) );
  AND2_X1 U9963 ( .A1(n9333), .A2(n8817), .ZN(n8818) );
  MUX2_X1 U9964 ( .A(n8819), .B(n8818), .S(n8840), .Z(n8820) );
  INV_X1 U9965 ( .A(n9323), .ZN(n8821) );
  OAI211_X1 U9966 ( .C1(n9367), .C2(n8850), .A(n8822), .B(n9333), .ZN(n8823)
         );
  OAI211_X1 U9967 ( .C1(n8824), .C2(n8850), .A(n8825), .B(n8823), .ZN(n8834)
         );
  INV_X1 U9968 ( .A(n8825), .ZN(n8826) );
  NOR2_X1 U9969 ( .A1(n8830), .A2(n8826), .ZN(n8828) );
  MUX2_X1 U9970 ( .A(n8828), .B(n8827), .S(n8850), .Z(n8833) );
  INV_X1 U9971 ( .A(n8829), .ZN(n8831) );
  MUX2_X1 U9972 ( .A(n8831), .B(n8830), .S(n8850), .Z(n8832) );
  AOI21_X1 U9973 ( .B1(n8834), .B2(n8833), .A(n8832), .ZN(n8838) );
  MUX2_X1 U9974 ( .A(n8836), .B(n8835), .S(n8850), .Z(n8837) );
  OAI211_X1 U9975 ( .C1(n8838), .C2(n9292), .A(n8880), .B(n8837), .ZN(n8844)
         );
  INV_X1 U9976 ( .A(n9303), .ZN(n8843) );
  INV_X1 U9977 ( .A(n9308), .ZN(n9289) );
  NAND3_X1 U9978 ( .A1(n8839), .A2(n9289), .A3(n8850), .ZN(n8842) );
  NAND3_X1 U9979 ( .A1(n9523), .A2(n9308), .A3(n8840), .ZN(n8841) );
  MUX2_X1 U9980 ( .A(n8846), .B(n8845), .S(n8850), .Z(n8847) );
  NAND2_X1 U9981 ( .A1(n9510), .A2(n9212), .ZN(n8852) );
  MUX2_X1 U9982 ( .A(n9510), .B(n9212), .S(n8850), .Z(n8851) );
  NOR3_X1 U9983 ( .A1(n8855), .A2(n8859), .A3(n5462), .ZN(n8891) );
  INV_X1 U9984 ( .A(n8856), .ZN(n8888) );
  NAND4_X1 U9985 ( .A1(n8860), .A2(n5529), .A3(n8859), .A4(n8858), .ZN(n8864)
         );
  NOR4_X1 U9986 ( .A1(n8864), .A2(n8863), .A3(n8862), .A4(n8861), .ZN(n8867)
         );
  NAND4_X1 U9987 ( .A1(n8867), .A2(n8866), .A3(n5521), .A4(n8865), .ZN(n8870)
         );
  NOR4_X1 U9988 ( .A1(n8870), .A2(n10920), .A3(n8869), .A4(n7417), .ZN(n8871)
         );
  NAND4_X1 U9989 ( .A1(n8874), .A2(n8873), .A3(n8872), .A4(n8871), .ZN(n8875)
         );
  NOR4_X1 U9990 ( .A1(n9454), .A2(n5176), .A3(n9497), .A4(n8875), .ZN(n8876)
         );
  NAND3_X1 U9991 ( .A1(n9428), .A2(n8876), .A3(n5641), .ZN(n8877) );
  NOR4_X1 U9992 ( .A1(n9386), .A2(n9416), .A3(n9398), .A4(n8877), .ZN(n8878)
         );
  NAND4_X1 U9993 ( .A1(n9332), .A2(n9357), .A3(n8057), .A4(n8878), .ZN(n8879)
         );
  NOR4_X1 U9994 ( .A1(n9303), .A2(n9292), .A3(n9324), .A4(n8879), .ZN(n8881)
         );
  NAND4_X1 U9995 ( .A1(n8883), .A2(n8882), .A3(n8881), .A4(n8880), .ZN(n8885)
         );
  XNOR2_X1 U9996 ( .A(n8885), .B(n8884), .ZN(n8886) );
  AOI211_X1 U9997 ( .C1(n8889), .C2(n8888), .A(n8887), .B(n8886), .ZN(n8890)
         );
  NOR4_X1 U9998 ( .A1(n8894), .A2(n9466), .A3(n8893), .A4(n5055), .ZN(n8897)
         );
  OAI21_X1 U9999 ( .B1(n8898), .B2(n8895), .A(P2_B_REG_SCAN_IN), .ZN(n8896) );
  OAI22_X1 U10000 ( .A1(n8899), .A2(n8898), .B1(n8897), .B2(n8896), .ZN(
        P2_U3244) );
  NAND2_X1 U10001 ( .A1(n8900), .A2(n10795), .ZN(n8906) );
  INV_X1 U10002 ( .A(n8901), .ZN(n8904) );
  AOI22_X1 U10003 ( .A1(n9091), .A2(n11059), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n11070), .ZN(n8902) );
  OAI21_X1 U10004 ( .B1(n5378), .B2(n10430), .A(n8902), .ZN(n8903) );
  AOI21_X1 U10005 ( .B1(n8904), .B2(n10291), .A(n8903), .ZN(n8905) );
  OAI211_X1 U10006 ( .C1(n10415), .C2(n8259), .A(n8906), .B(n8905), .ZN(
        P1_U3263) );
  AOI22_X1 U10007 ( .A1(n8907), .A2(n9188), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8908) );
  OAI21_X1 U10008 ( .B1(n8909), .B2(n9161), .A(n8908), .ZN(n8945) );
  INV_X1 U10009 ( .A(n8910), .ZN(n8911) );
  XNOR2_X1 U10010 ( .A(n9549), .B(n5877), .ZN(n8916) );
  XNOR2_X1 U10011 ( .A(n9543), .B(n5877), .ZN(n9154) );
  NAND2_X1 U10012 ( .A1(n9367), .A2(n8927), .ZN(n9156) );
  AND2_X1 U10013 ( .A1(n9154), .A2(n9156), .ZN(n8914) );
  OAI22_X1 U10014 ( .A1(n5693), .A2(n8914), .B1(n9154), .B2(n9156), .ZN(n8915)
         );
  INV_X1 U10015 ( .A(n8915), .ZN(n8921) );
  INV_X1 U10016 ( .A(n8916), .ZN(n8917) );
  XNOR2_X1 U10017 ( .A(n8918), .B(n8917), .ZN(n9131) );
  INV_X1 U10018 ( .A(n9160), .ZN(n9359) );
  NAND2_X1 U10019 ( .A1(n9359), .A2(n8927), .ZN(n9129) );
  AOI21_X1 U10020 ( .B1(n9154), .B2(n8024), .A(n9129), .ZN(n8919) );
  NAND2_X1 U10021 ( .A1(n9131), .A2(n8919), .ZN(n8920) );
  XNOR2_X1 U10022 ( .A(n9540), .B(n8941), .ZN(n8922) );
  NOR2_X1 U10023 ( .A1(n9203), .A2(n8940), .ZN(n8923) );
  NAND2_X1 U10024 ( .A1(n8922), .A2(n8923), .ZN(n8926) );
  INV_X1 U10025 ( .A(n8922), .ZN(n9199) );
  INV_X1 U10026 ( .A(n8923), .ZN(n8924) );
  NAND2_X1 U10027 ( .A1(n9199), .A2(n8924), .ZN(n8925) );
  AND2_X1 U10028 ( .A1(n8926), .A2(n8925), .ZN(n9146) );
  XNOR2_X1 U10029 ( .A(n9322), .B(n5877), .ZN(n8928) );
  AND2_X1 U10030 ( .A1(n9215), .A2(n8927), .ZN(n8929) );
  NAND2_X1 U10031 ( .A1(n8928), .A2(n8929), .ZN(n8932) );
  INV_X1 U10032 ( .A(n8928), .ZN(n9116) );
  INV_X1 U10033 ( .A(n8929), .ZN(n8930) );
  NAND2_X1 U10034 ( .A1(n9116), .A2(n8930), .ZN(n8931) );
  AND2_X1 U10035 ( .A1(n8932), .A2(n8931), .ZN(n9194) );
  NAND2_X1 U10036 ( .A1(n9113), .A2(n8932), .ZN(n8938) );
  XNOR2_X1 U10037 ( .A(n9528), .B(n8941), .ZN(n8933) );
  NOR2_X1 U10038 ( .A1(n9202), .A2(n8940), .ZN(n8934) );
  NAND2_X1 U10039 ( .A1(n8933), .A2(n8934), .ZN(n8939) );
  INV_X1 U10040 ( .A(n8933), .ZN(n8936) );
  INV_X1 U10041 ( .A(n8934), .ZN(n8935) );
  NAND2_X1 U10042 ( .A1(n8936), .A2(n8935), .ZN(n8937) );
  AND2_X1 U10043 ( .A1(n8939), .A2(n8937), .ZN(n9114) );
  NOR2_X1 U10044 ( .A1(n9308), .A2(n8940), .ZN(n8942) );
  MUX2_X1 U10045 ( .A(n8942), .B(n9308), .S(n8941), .Z(n8943) );
  INV_X1 U10046 ( .A(n8946), .ZN(n9493) );
  AOI22_X1 U10047 ( .A1(n9500), .A2(n9189), .B1(n9188), .B2(n9493), .ZN(n8948)
         );
  OAI211_X1 U10048 ( .C1(n9465), .C2(n9161), .A(n8948), .B(n8947), .ZN(n8954)
         );
  INV_X1 U10049 ( .A(n8982), .ZN(n8952) );
  AOI22_X1 U10050 ( .A1(n8949), .A2(n9167), .B1(n9128), .B2(n9500), .ZN(n8951)
         );
  NOR3_X1 U10051 ( .A1(n8952), .A2(n8951), .A3(n8950), .ZN(n8953) );
  AOI211_X1 U10052 ( .C1(n9171), .C2(n10023), .A(n8954), .B(n8953), .ZN(n8955)
         );
  OAI21_X1 U10053 ( .B1(n8956), .B2(n9195), .A(n8955), .ZN(P2_U3243) );
  NAND2_X1 U10054 ( .A1(n8957), .A2(n9208), .ZN(n8959) );
  OAI211_X1 U10055 ( .C1(n9206), .C2(n8960), .A(n8959), .B(n8958), .ZN(n8964)
         );
  INV_X1 U10056 ( .A(n9166), .ZN(n8963) );
  AOI22_X1 U10057 ( .A1(n9167), .A2(n8961), .B1(n9224), .B2(n9128), .ZN(n8962)
         );
  AOI211_X1 U10058 ( .C1(n9171), .C2(n8965), .A(n8964), .B(n5133), .ZN(n8966)
         );
  OAI21_X1 U10059 ( .B1(n8967), .B2(n9195), .A(n8966), .ZN(P2_U3229) );
  OAI21_X1 U10060 ( .B1(n8969), .B2(n9161), .A(n8968), .ZN(n8972) );
  OAI22_X1 U10061 ( .A1(n8975), .A2(n9159), .B1(n9206), .B2(n8970), .ZN(n8971)
         );
  AOI211_X1 U10062 ( .C1(n8973), .C2(n9171), .A(n8972), .B(n8971), .ZN(n8981)
         );
  INV_X1 U10063 ( .A(n8974), .ZN(n8978) );
  OAI22_X1 U10064 ( .A1(n8976), .A2(n9195), .B1(n8975), .B2(n9198), .ZN(n8977)
         );
  NAND3_X1 U10065 ( .A1(n8979), .A2(n8978), .A3(n8977), .ZN(n8980) );
  OAI211_X1 U10066 ( .C1(n8982), .C2(n9195), .A(n8981), .B(n8980), .ZN(
        P2_U3217) );
  AOI22_X1 U10067 ( .A1(n10474), .A2(n9086), .B1(n9085), .B2(n10356), .ZN(
        n9056) );
  NAND2_X1 U10068 ( .A1(n10474), .A2(n7122), .ZN(n8984) );
  NAND2_X1 U10069 ( .A1(n10356), .A2(n9080), .ZN(n8983) );
  NAND2_X1 U10070 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  XNOR2_X1 U10071 ( .A(n8985), .B(n9076), .ZN(n9054) );
  INV_X1 U10072 ( .A(n9054), .ZN(n9055) );
  AOI22_X1 U10073 ( .A1(n10479), .A2(n9086), .B1(n9085), .B2(n10375), .ZN(
        n9053) );
  NAND2_X1 U10074 ( .A1(n10479), .A2(n7122), .ZN(n8987) );
  NAND2_X1 U10075 ( .A1(n10375), .A2(n9086), .ZN(n8986) );
  NAND2_X1 U10076 ( .A1(n8987), .A2(n8986), .ZN(n8988) );
  XNOR2_X1 U10077 ( .A(n8988), .B(n9076), .ZN(n9051) );
  INV_X1 U10078 ( .A(n9051), .ZN(n9052) );
  NAND2_X1 U10079 ( .A1(n10489), .A2(n7122), .ZN(n8990) );
  NAND2_X1 U10080 ( .A1(n10376), .A2(n9080), .ZN(n8989) );
  NAND2_X1 U10081 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  XNOR2_X1 U10082 ( .A(n8991), .B(n9076), .ZN(n9043) );
  AND2_X1 U10083 ( .A1(n10376), .A2(n9085), .ZN(n8992) );
  AOI21_X1 U10084 ( .B1(n10489), .B2(n9080), .A(n8992), .ZN(n9041) );
  INV_X1 U10085 ( .A(n9041), .ZN(n9042) );
  OAI21_X1 U10086 ( .B1(n8995), .B2(n8994), .A(n8993), .ZN(n8997) );
  NAND2_X1 U10087 ( .A1(n8995), .A2(n8994), .ZN(n8996) );
  NAND2_X1 U10088 ( .A1(n10984), .A2(n7122), .ZN(n8999) );
  NAND2_X1 U10089 ( .A1(n10959), .A2(n9080), .ZN(n8998) );
  NAND2_X1 U10090 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  XNOR2_X1 U10091 ( .A(n9000), .B(n9076), .ZN(n9003) );
  NAND2_X1 U10092 ( .A1(n10984), .A2(n9080), .ZN(n9002) );
  NAND2_X1 U10093 ( .A1(n10959), .A2(n9085), .ZN(n9001) );
  NAND2_X1 U10094 ( .A1(n9002), .A2(n9001), .ZN(n9004) );
  INV_X1 U10095 ( .A(n9003), .ZN(n9006) );
  INV_X1 U10096 ( .A(n9004), .ZN(n9005) );
  NAND2_X1 U10097 ( .A1(n9006), .A2(n9005), .ZN(n10153) );
  NAND2_X1 U10098 ( .A1(n10074), .A2(n7122), .ZN(n9008) );
  NAND2_X1 U10099 ( .A1(n10231), .A2(n9080), .ZN(n9007) );
  NAND2_X1 U10100 ( .A1(n9008), .A2(n9007), .ZN(n9009) );
  AND2_X1 U10101 ( .A1(n10153), .A2(n5061), .ZN(n9010) );
  OR2_X1 U10102 ( .A1(n10150), .A2(n5061), .ZN(n9011) );
  OR2_X1 U10103 ( .A1(n5061), .A2(n10153), .ZN(n10063) );
  NAND2_X1 U10104 ( .A1(n10074), .A2(n9080), .ZN(n9013) );
  NAND2_X1 U10105 ( .A1(n10231), .A2(n9085), .ZN(n9012) );
  NAND2_X1 U10106 ( .A1(n9013), .A2(n9012), .ZN(n10067) );
  AND2_X1 U10107 ( .A1(n10063), .A2(n10067), .ZN(n9014) );
  NAND2_X1 U10108 ( .A1(n10224), .A2(n7122), .ZN(n9016) );
  NAND2_X1 U10109 ( .A1(n11039), .A2(n9086), .ZN(n9015) );
  NAND2_X1 U10110 ( .A1(n9016), .A2(n9015), .ZN(n9017) );
  NAND2_X1 U10111 ( .A1(n10224), .A2(n9080), .ZN(n9019) );
  NAND2_X1 U10112 ( .A1(n11039), .A2(n9085), .ZN(n9018) );
  NAND2_X1 U10113 ( .A1(n9019), .A2(n9018), .ZN(n10212) );
  NAND2_X1 U10114 ( .A1(n11061), .A2(n7122), .ZN(n9021) );
  NAND2_X1 U10115 ( .A1(n10424), .A2(n9080), .ZN(n9020) );
  NAND2_X1 U10116 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  XNOR2_X1 U10117 ( .A(n9022), .B(n9076), .ZN(n9024) );
  AND2_X1 U10118 ( .A1(n10424), .A2(n9085), .ZN(n9023) );
  AOI21_X1 U10119 ( .B1(n11061), .B2(n9086), .A(n9023), .ZN(n9025) );
  XNOR2_X1 U10120 ( .A(n9024), .B(n9025), .ZN(n10114) );
  INV_X1 U10121 ( .A(n9024), .ZN(n9026) );
  NAND2_X1 U10122 ( .A1(n9026), .A2(n9025), .ZN(n9027) );
  NAND2_X1 U10123 ( .A1(n10500), .A2(n7122), .ZN(n9029) );
  NAND2_X1 U10124 ( .A1(n11038), .A2(n9086), .ZN(n9028) );
  NAND2_X1 U10125 ( .A1(n9029), .A2(n9028), .ZN(n9030) );
  XNOR2_X1 U10126 ( .A(n9030), .B(n9083), .ZN(n10123) );
  AND2_X1 U10127 ( .A1(n11038), .A2(n9085), .ZN(n9031) );
  AOI21_X1 U10128 ( .B1(n10500), .B2(n9086), .A(n9031), .ZN(n9032) );
  INV_X1 U10129 ( .A(n10123), .ZN(n9033) );
  INV_X1 U10130 ( .A(n9032), .ZN(n10122) );
  NAND2_X1 U10131 ( .A1(n9033), .A2(n10122), .ZN(n9034) );
  NAND2_X1 U10132 ( .A1(n10494), .A2(n7122), .ZN(n9037) );
  NAND2_X1 U10133 ( .A1(n10425), .A2(n9080), .ZN(n9036) );
  NAND2_X1 U10134 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  XNOR2_X1 U10135 ( .A(n9038), .B(n9076), .ZN(n10183) );
  NAND2_X1 U10136 ( .A1(n10494), .A2(n9080), .ZN(n9040) );
  NAND2_X1 U10137 ( .A1(n10425), .A2(n9085), .ZN(n9039) );
  NAND2_X1 U10138 ( .A1(n9040), .A2(n9039), .ZN(n10188) );
  XNOR2_X1 U10139 ( .A(n9043), .B(n9041), .ZN(n10088) );
  NAND2_X1 U10140 ( .A1(n10484), .A2(n7122), .ZN(n9045) );
  NAND2_X1 U10141 ( .A1(n10394), .A2(n9086), .ZN(n9044) );
  NAND2_X1 U10142 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  XNOR2_X1 U10143 ( .A(n9046), .B(n9076), .ZN(n9050) );
  NAND2_X1 U10144 ( .A1(n10484), .A2(n9086), .ZN(n9048) );
  NAND2_X1 U10145 ( .A1(n10394), .A2(n9085), .ZN(n9047) );
  NAND2_X1 U10146 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  NOR2_X1 U10147 ( .A1(n9050), .A2(n9049), .ZN(n10140) );
  NAND2_X1 U10148 ( .A1(n9050), .A2(n9049), .ZN(n10141) );
  XOR2_X1 U10149 ( .A(n9053), .B(n9051), .Z(n10098) );
  XOR2_X1 U10150 ( .A(n9056), .B(n9054), .Z(n10165) );
  AOI22_X1 U10151 ( .A1(n10469), .A2(n7122), .B1(n9080), .B2(n10346), .ZN(
        n9057) );
  AOI22_X1 U10152 ( .A1(n10469), .A2(n9080), .B1(n9085), .B2(n10346), .ZN(
        n10077) );
  AOI22_X1 U10153 ( .A1(n10464), .A2(n9086), .B1(n9085), .B2(n10327), .ZN(
        n9061) );
  NAND2_X1 U10154 ( .A1(n10464), .A2(n7122), .ZN(n9059) );
  NAND2_X1 U10155 ( .A1(n10327), .A2(n9080), .ZN(n9058) );
  NAND2_X1 U10156 ( .A1(n9059), .A2(n9058), .ZN(n9060) );
  XNOR2_X1 U10157 ( .A(n9060), .B(n9076), .ZN(n9063) );
  XOR2_X1 U10158 ( .A(n9061), .B(n9063), .Z(n10133) );
  INV_X1 U10159 ( .A(n9061), .ZN(n9062) );
  NAND2_X1 U10160 ( .A1(n10459), .A2(n7122), .ZN(n9065) );
  NAND2_X1 U10161 ( .A1(n10230), .A2(n9086), .ZN(n9064) );
  NAND2_X1 U10162 ( .A1(n9065), .A2(n9064), .ZN(n9066) );
  XNOR2_X1 U10163 ( .A(n9066), .B(n9076), .ZN(n9067) );
  AOI22_X1 U10164 ( .A1(n10459), .A2(n9080), .B1(n9085), .B2(n10230), .ZN(
        n9068) );
  XNOR2_X1 U10165 ( .A(n9067), .B(n9068), .ZN(n10105) );
  INV_X1 U10166 ( .A(n9067), .ZN(n9069) );
  AOI22_X1 U10167 ( .A1(n10454), .A2(n9086), .B1(n9085), .B2(n10318), .ZN(
        n9072) );
  AOI22_X1 U10168 ( .A1(n10454), .A2(n7122), .B1(n9080), .B2(n10318), .ZN(
        n9070) );
  XNOR2_X1 U10169 ( .A(n9070), .B(n9076), .ZN(n9071) );
  XOR2_X1 U10170 ( .A(n9072), .B(n9071), .Z(n10199) );
  INV_X1 U10171 ( .A(n9071), .ZN(n9074) );
  INV_X1 U10172 ( .A(n9072), .ZN(n9073) );
  NAND2_X1 U10173 ( .A1(n9074), .A2(n9073), .ZN(n9075) );
  AOI22_X1 U10174 ( .A1(n10449), .A2(n7122), .B1(n9080), .B2(n10229), .ZN(
        n9077) );
  XNOR2_X1 U10175 ( .A(n9077), .B(n9076), .ZN(n10055) );
  AND2_X1 U10176 ( .A1(n10229), .A2(n9085), .ZN(n9078) );
  AOI21_X1 U10177 ( .B1(n10449), .B2(n9080), .A(n9078), .ZN(n10056) );
  NAND2_X1 U10178 ( .A1(n10055), .A2(n10056), .ZN(n9079) );
  NAND2_X1 U10179 ( .A1(n10057), .A2(n9079), .ZN(n9103) );
  NAND2_X1 U10180 ( .A1(n9099), .A2(n7122), .ZN(n9082) );
  OR2_X1 U10181 ( .A1(n10058), .A2(n6027), .ZN(n9081) );
  NAND2_X1 U10182 ( .A1(n9082), .A2(n9081), .ZN(n9084) );
  XNOR2_X1 U10183 ( .A(n9084), .B(n9083), .ZN(n9089) );
  NAND2_X1 U10184 ( .A1(n9099), .A2(n9086), .ZN(n9087) );
  OAI21_X1 U10185 ( .B1(n10058), .B2(n5360), .A(n9087), .ZN(n9088) );
  XNOR2_X1 U10186 ( .A(n9089), .B(n9088), .ZN(n9096) );
  INV_X1 U10187 ( .A(n9096), .ZN(n9090) );
  NAND2_X1 U10188 ( .A1(n9090), .A2(n10197), .ZN(n9102) );
  OR2_X1 U10189 ( .A1(n10055), .A2(n10056), .ZN(n9095) );
  NAND2_X1 U10190 ( .A1(n9103), .A2(n5694), .ZN(n9101) );
  AOI22_X1 U10191 ( .A1(n10218), .A2(n10229), .B1(n9091), .B2(n10203), .ZN(
        n9093) );
  NAND2_X1 U10192 ( .A1(P1_U3084), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9092) );
  OAI211_X1 U10193 ( .C1(n9094), .C2(n10215), .A(n9093), .B(n9092), .ZN(n9098)
         );
  NOR3_X1 U10194 ( .A1(n9096), .A2(n10226), .A3(n9095), .ZN(n9097) );
  AOI211_X1 U10195 ( .C1(n9099), .C2(n10223), .A(n9098), .B(n9097), .ZN(n9100)
         );
  OAI211_X1 U10196 ( .C1(n9103), .C2(n9102), .A(n9101), .B(n9100), .ZN(
        P1_U3218) );
  INV_X1 U10197 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9106) );
  OAI222_X1 U10198 ( .A1(n9110), .A2(n9106), .B1(n6076), .B2(n9105), .C1(n9104), .C2(P2_U3152), .ZN(P2_U3330) );
  INV_X1 U10199 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9107) );
  OAI222_X1 U10200 ( .A1(n10532), .A2(n9108), .B1(n6013), .B2(P1_U3084), .C1(
        n9107), .C2(n10528), .ZN(P1_U3324) );
  INV_X1 U10201 ( .A(n9109), .ZN(n10531) );
  INV_X1 U10202 ( .A(n9114), .ZN(n9115) );
  AOI21_X1 U10203 ( .B1(n9113), .B2(n9115), .A(n9195), .ZN(n9119) );
  NOR3_X1 U10204 ( .A1(n9116), .A2(n9121), .A3(n9198), .ZN(n9118) );
  OAI21_X1 U10205 ( .B1(n9119), .B2(n9118), .A(n9117), .ZN(n9126) );
  OAI22_X1 U10206 ( .A1(n9121), .A2(n9159), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9120), .ZN(n9123) );
  NOR2_X1 U10207 ( .A1(n9308), .A2(n9161), .ZN(n9122) );
  AOI211_X1 U10208 ( .C1(n9188), .C2(n9124), .A(n9123), .B(n9122), .ZN(n9125)
         );
  OAI211_X1 U10209 ( .C1(n9127), .C2(n9211), .A(n9126), .B(n9125), .ZN(
        P2_U3216) );
  AOI22_X1 U10210 ( .A1(n9131), .A2(n9167), .B1(n9128), .B2(n9359), .ZN(n9136)
         );
  INV_X1 U10211 ( .A(n9129), .ZN(n9130) );
  NAND2_X1 U10212 ( .A1(n9131), .A2(n9130), .ZN(n9152) );
  INV_X1 U10213 ( .A(n9152), .ZN(n9135) );
  OAI22_X1 U10214 ( .A1(n8024), .A2(n9161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9620), .ZN(n9133) );
  OAI22_X1 U10215 ( .A1(n9216), .A2(n9159), .B1(n9206), .B2(n9372), .ZN(n9132)
         );
  AOI211_X1 U10216 ( .C1(n9549), .C2(n9171), .A(n9133), .B(n9132), .ZN(n9134)
         );
  OAI21_X1 U10217 ( .B1(n9136), .B2(n9135), .A(n9134), .ZN(P2_U3218) );
  AOI21_X1 U10218 ( .B1(n9181), .B2(n5421), .A(n9195), .ZN(n9140) );
  NOR3_X1 U10219 ( .A1(n9138), .A2(n9431), .A3(n9198), .ZN(n9139) );
  OAI21_X1 U10220 ( .B1(n9140), .B2(n9139), .A(n8341), .ZN(n9144) );
  OAI22_X1 U10221 ( .A1(n9216), .A2(n9161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9845), .ZN(n9142) );
  OAI22_X1 U10222 ( .A1(n9431), .A2(n9159), .B1(n9206), .B2(n9406), .ZN(n9141)
         );
  AOI211_X1 U10223 ( .C1(n9993), .C2(n9171), .A(n9142), .B(n9141), .ZN(n9143)
         );
  NAND2_X1 U10224 ( .A1(n9144), .A2(n9143), .ZN(P2_U3225) );
  OAI211_X1 U10225 ( .C1(n9146), .C2(n9145), .A(n9197), .B(n9167), .ZN(n9151)
         );
  AOI22_X1 U10226 ( .A1(n9215), .A2(n9501), .B1(n9499), .B2(n9367), .ZN(n9338)
         );
  AOI22_X1 U10227 ( .A1(n9343), .A2(n9188), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n9147) );
  OAI21_X1 U10228 ( .B1(n9338), .B2(n9148), .A(n9147), .ZN(n9149) );
  INV_X1 U10229 ( .A(n9149), .ZN(n9150) );
  OAI211_X1 U10230 ( .C1(n9346), .C2(n9211), .A(n9151), .B(n9150), .ZN(
        P2_U3227) );
  NAND2_X1 U10231 ( .A1(n9152), .A2(n5693), .ZN(n9153) );
  XOR2_X1 U10232 ( .A(n9154), .B(n9153), .Z(n9157) );
  OAI22_X1 U10233 ( .A1(n9157), .A2(n9195), .B1(n8024), .B2(n9198), .ZN(n9155)
         );
  OAI21_X1 U10234 ( .B1(n9157), .B2(n9156), .A(n9155), .ZN(n9165) );
  INV_X1 U10235 ( .A(n9158), .ZN(n9355) );
  OAI22_X1 U10236 ( .A1(n9160), .A2(n9159), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9854), .ZN(n9163) );
  NOR2_X1 U10237 ( .A1(n9203), .A2(n9161), .ZN(n9162) );
  AOI211_X1 U10238 ( .C1(n9188), .C2(n9355), .A(n9163), .B(n9162), .ZN(n9164)
         );
  OAI211_X1 U10239 ( .C1(n8025), .C2(n9211), .A(n9165), .B(n9164), .ZN(
        P2_U3231) );
  OAI21_X1 U10240 ( .B1(n5401), .B2(n9174), .A(n9166), .ZN(n9168) );
  NAND2_X1 U10241 ( .A1(n9168), .A2(n9167), .ZN(n9180) );
  AOI22_X1 U10242 ( .A1(n9223), .A2(n9185), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n9179) );
  INV_X1 U10243 ( .A(n9169), .ZN(n9172) );
  AOI22_X1 U10244 ( .A1(n9188), .A2(n9172), .B1(n9171), .B2(n9170), .ZN(n9178)
         );
  NOR3_X1 U10245 ( .A1(n9174), .A2(n9173), .A3(n9198), .ZN(n9176) );
  OAI21_X1 U10246 ( .B1(n9176), .B2(n9189), .A(n9175), .ZN(n9177) );
  NAND4_X1 U10247 ( .A1(n9180), .A2(n9179), .A3(n9178), .A4(n9177), .ZN(
        P2_U3232) );
  INV_X1 U10248 ( .A(n9181), .ZN(n9182) );
  AOI211_X1 U10249 ( .C1(n9184), .C2(n9183), .A(n9195), .B(n9182), .ZN(n9193)
         );
  INV_X1 U10250 ( .A(n9998), .ZN(n9415) );
  AOI22_X1 U10251 ( .A1(n9418), .A2(n9185), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n9191) );
  INV_X1 U10252 ( .A(n9186), .ZN(n9448) );
  INV_X1 U10253 ( .A(n9187), .ZN(n9413) );
  AOI22_X1 U10254 ( .A1(n9448), .A2(n9189), .B1(n9413), .B2(n9188), .ZN(n9190)
         );
  OAI211_X1 U10255 ( .C1(n9415), .C2(n9211), .A(n9191), .B(n9190), .ZN(n9192)
         );
  OR2_X1 U10256 ( .A1(n9193), .A2(n9192), .ZN(P2_U3235) );
  INV_X1 U10257 ( .A(n9194), .ZN(n9196) );
  AOI21_X1 U10258 ( .B1(n9197), .B2(n9196), .A(n9195), .ZN(n9201) );
  NOR3_X1 U10259 ( .A1(n9199), .A2(n9203), .A3(n9198), .ZN(n9200) );
  OAI21_X1 U10260 ( .B1(n9201), .B2(n9200), .A(n9113), .ZN(n9210) );
  OR2_X1 U10261 ( .A1(n9202), .A2(n9468), .ZN(n9205) );
  OR2_X1 U10262 ( .A1(n9203), .A2(n9466), .ZN(n9204) );
  NAND2_X1 U10263 ( .A1(n9205), .A2(n9204), .ZN(n9326) );
  OAI22_X1 U10264 ( .A1(n9319), .A2(n9206), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9877), .ZN(n9207) );
  AOI21_X1 U10265 ( .B1(n9326), .B2(n9208), .A(n9207), .ZN(n9209) );
  OAI211_X1 U10266 ( .C1(n9322), .C2(n9211), .A(n9210), .B(n9209), .ZN(
        P2_U3242) );
  MUX2_X1 U10267 ( .A(n9212), .B(P2_DATAO_REG_31__SCAN_IN), .S(n9226), .Z(
        P2_U3583) );
  MUX2_X1 U10268 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9213), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10269 ( .A(n9289), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9226), .Z(
        P2_U3580) );
  MUX2_X1 U10270 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9214), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10271 ( .A(n9215), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9226), .Z(
        P2_U3578) );
  MUX2_X1 U10272 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9360), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10273 ( .A(n9367), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9226), .Z(
        P2_U3576) );
  MUX2_X1 U10274 ( .A(n9359), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9226), .Z(
        P2_U3575) );
  INV_X1 U10275 ( .A(n9216), .ZN(n9395) );
  MUX2_X1 U10276 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9395), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10277 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9418), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10278 ( .A(n9394), .B(P2_DATAO_REG_20__SCAN_IN), .S(n9226), .Z(
        P2_U3572) );
  MUX2_X1 U10279 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9448), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10280 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9217), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10281 ( .A(n9447), .B(P2_DATAO_REG_17__SCAN_IN), .S(n9226), .Z(
        P2_U3569) );
  MUX2_X1 U10282 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9502), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10283 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9218), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10284 ( .A(n9500), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9226), .Z(
        P2_U3566) );
  MUX2_X1 U10285 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9219), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10286 ( .A(n9220), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9226), .Z(
        P2_U3560) );
  MUX2_X1 U10287 ( .A(n9221), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9226), .Z(
        P2_U3559) );
  MUX2_X1 U10288 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n9222), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10289 ( .A(n9223), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9226), .Z(
        P2_U3557) );
  MUX2_X1 U10290 ( .A(n9224), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9226), .Z(
        P2_U3556) );
  MUX2_X1 U10291 ( .A(n9225), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9226), .Z(
        P2_U3554) );
  MUX2_X1 U10292 ( .A(n6531), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9226), .Z(
        P2_U3553) );
  MUX2_X1 U10293 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9227), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI211_X1 U10294 ( .C1(n9230), .C2(n9229), .A(n10679), .B(n9228), .ZN(n9240)
         );
  AOI21_X1 U10295 ( .B1(n10674), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9231), .ZN(
        n9239) );
  NAND2_X1 U10296 ( .A1(n10660), .A2(n9232), .ZN(n9238) );
  OAI21_X1 U10297 ( .B1(n9235), .B2(n9234), .A(n9233), .ZN(n9236) );
  OR2_X1 U10298 ( .A1(n10658), .A2(n9236), .ZN(n9237) );
  NAND4_X1 U10299 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(
        P2_U3255) );
  OR2_X1 U10300 ( .A1(n9262), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U10301 ( .A1(n9262), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9241) );
  NAND2_X1 U10302 ( .A1(n9242), .A2(n9241), .ZN(n9247) );
  AOI21_X1 U10303 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9244), .A(n9243), .ZN(
        n9245) );
  INV_X1 U10304 ( .A(n9245), .ZN(n9246) );
  NOR2_X1 U10305 ( .A1(n9247), .A2(n9246), .ZN(n9264) );
  AOI21_X1 U10306 ( .B1(n9247), .B2(n9246), .A(n9264), .ZN(n9261) );
  OAI21_X1 U10307 ( .B1(n9250), .B2(n9249), .A(n9248), .ZN(n9253) );
  OR2_X1 U10308 ( .A1(n9262), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U10309 ( .A1(n9262), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U10310 ( .A1(n9267), .A2(n9251), .ZN(n9252) );
  NOR2_X1 U10311 ( .A1(n9252), .A2(n9253), .ZN(n9269) );
  AOI21_X1 U10312 ( .B1(n9253), .B2(n9252), .A(n9269), .ZN(n9254) );
  NOR2_X1 U10313 ( .A1(n10658), .A2(n9254), .ZN(n9259) );
  INV_X1 U10314 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9256) );
  OAI21_X1 U10315 ( .B1(n9257), .B2(n9256), .A(n9255), .ZN(n9258) );
  AOI211_X1 U10316 ( .C1(n10660), .C2(n9262), .A(n9259), .B(n9258), .ZN(n9260)
         );
  OAI21_X1 U10317 ( .B1(n9261), .B2(n9278), .A(n9260), .ZN(P2_U3263) );
  MUX2_X1 U10318 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n7909), .S(n5819), .Z(n9266) );
  NOR2_X1 U10319 ( .A1(n9262), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9263) );
  NOR2_X1 U10320 ( .A1(n9264), .A2(n9263), .ZN(n9265) );
  XNOR2_X1 U10321 ( .A(n9266), .B(n9265), .ZN(n9277) );
  INV_X1 U10322 ( .A(n9267), .ZN(n9268) );
  OR2_X1 U10323 ( .A1(n9269), .A2(n9268), .ZN(n9271) );
  XNOR2_X1 U10324 ( .A(n5819), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9270) );
  XNOR2_X1 U10325 ( .A(n9271), .B(n9270), .ZN(n9274) );
  NAND2_X1 U10326 ( .A1(n10674), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9272) );
  OAI211_X1 U10327 ( .C1(n10658), .C2(n9274), .A(n9273), .B(n9272), .ZN(n9275)
         );
  AOI21_X1 U10328 ( .B1(n5819), .B2(n10660), .A(n9275), .ZN(n9276) );
  OAI21_X1 U10329 ( .B1(n9278), .B2(n9277), .A(n9276), .ZN(P2_U3264) );
  NOR2_X1 U10330 ( .A1(n9514), .A2(n5054), .ZN(n9279) );
  XOR2_X1 U10331 ( .A(n9279), .B(n9510), .Z(n9512) );
  OAI21_X1 U10332 ( .B1(n5055), .B2(n9280), .A(n9501), .ZN(n9307) );
  NOR2_X1 U10333 ( .A1(n9281), .A2(n9307), .ZN(n9513) );
  NAND2_X1 U10334 ( .A1(n9513), .A2(n10946), .ZN(n9285) );
  OAI21_X1 U10335 ( .B1(n10946), .B2(n9282), .A(n9285), .ZN(n9283) );
  AOI21_X1 U10336 ( .B1(n9510), .B2(n9427), .A(n9283), .ZN(n9284) );
  OAI21_X1 U10337 ( .B1(n9512), .B2(n9309), .A(n9284), .ZN(P2_U3265) );
  XNOR2_X1 U10338 ( .A(n5054), .B(n9514), .ZN(n9516) );
  INV_X1 U10339 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9286) );
  OAI21_X1 U10340 ( .B1(n10946), .B2(n9286), .A(n9285), .ZN(n9287) );
  AOI21_X1 U10341 ( .B1(n9514), .B2(n9427), .A(n9287), .ZN(n9288) );
  OAI21_X1 U10342 ( .B1(n9516), .B2(n9309), .A(n9288), .ZN(P2_U3266) );
  OR2_X1 U10343 ( .A1(n9523), .A2(n9289), .ZN(n9296) );
  INV_X1 U10344 ( .A(n9296), .ZN(n9291) );
  OR2_X1 U10345 ( .A1(n9291), .A2(n9290), .ZN(n9295) );
  AND2_X1 U10346 ( .A1(n9292), .A2(n9295), .ZN(n9293) );
  NAND2_X1 U10347 ( .A1(n9294), .A2(n9293), .ZN(n9301) );
  INV_X1 U10348 ( .A(n9295), .ZN(n9299) );
  AND2_X1 U10349 ( .A1(n9297), .A2(n9296), .ZN(n9298) );
  NAND2_X1 U10350 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  XNOR2_X1 U10351 ( .A(n9302), .B(n9303), .ZN(n9517) );
  INV_X1 U10352 ( .A(n9517), .ZN(n9316) );
  XNOR2_X1 U10353 ( .A(n9304), .B(n9303), .ZN(n9305) );
  INV_X1 U10354 ( .A(n9521), .ZN(n9312) );
  OAI21_X1 U10355 ( .B1(n9312), .B2(n5078), .A(n5054), .ZN(n9518) );
  NOR2_X1 U10356 ( .A1(n9518), .A2(n9309), .ZN(n9314) );
  AOI22_X1 U10357 ( .A1(n9310), .A2(n9492), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9426), .ZN(n9311) );
  OAI21_X1 U10358 ( .B1(n9312), .B2(n9495), .A(n9311), .ZN(n9313) );
  AOI211_X1 U10359 ( .C1(n9519), .C2(n10946), .A(n9314), .B(n9313), .ZN(n9315)
         );
  OAI21_X1 U10360 ( .B1(n9316), .B2(n9509), .A(n9315), .ZN(P2_U3267) );
  XOR2_X1 U10361 ( .A(n9324), .B(n9317), .Z(n9537) );
  AOI211_X1 U10362 ( .C1(n9534), .C2(n9340), .A(n11011), .B(n9318), .ZN(n9533)
         );
  INV_X1 U10363 ( .A(n9319), .ZN(n9320) );
  AOI22_X1 U10364 ( .A1(n9320), .A2(n9492), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n9426), .ZN(n9321) );
  OAI21_X1 U10365 ( .B1(n9322), .B2(n9495), .A(n9321), .ZN(n9329) );
  NAND2_X1 U10366 ( .A1(n9337), .A2(n9323), .ZN(n9325) );
  XNOR2_X1 U10367 ( .A(n9325), .B(n9324), .ZN(n9327) );
  AOI21_X1 U10368 ( .B1(n9327), .B2(n10923), .A(n9326), .ZN(n9536) );
  NOR2_X1 U10369 ( .A1(n9536), .A2(n9504), .ZN(n9328) );
  AOI211_X1 U10370 ( .C1(n9533), .C2(n9481), .A(n9329), .B(n9328), .ZN(n9330)
         );
  OAI21_X1 U10371 ( .B1(n9537), .B2(n9509), .A(n9330), .ZN(P2_U3270) );
  XNOR2_X1 U10372 ( .A(n9331), .B(n9332), .ZN(n9542) );
  NAND3_X1 U10373 ( .A1(n9335), .A2(n9334), .A3(n9333), .ZN(n9336) );
  NAND3_X1 U10374 ( .A1(n9337), .A2(n10923), .A3(n9336), .ZN(n9339) );
  NAND2_X1 U10375 ( .A1(n9339), .A2(n9338), .ZN(n9538) );
  INV_X1 U10376 ( .A(n9353), .ZN(n9342) );
  INV_X1 U10377 ( .A(n9340), .ZN(n9341) );
  AOI211_X1 U10378 ( .C1(n9540), .C2(n9342), .A(n11011), .B(n9341), .ZN(n9539)
         );
  NAND2_X1 U10379 ( .A1(n9539), .A2(n9481), .ZN(n9345) );
  AOI22_X1 U10380 ( .A1(n9343), .A2(n9492), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9426), .ZN(n9344) );
  OAI211_X1 U10381 ( .C1(n9346), .C2(n9495), .A(n9345), .B(n9344), .ZN(n9347)
         );
  AOI21_X1 U10382 ( .B1(n9538), .B2(n10946), .A(n9347), .ZN(n9348) );
  OAI21_X1 U10383 ( .B1(n9542), .B2(n9509), .A(n9348), .ZN(P2_U3271) );
  INV_X1 U10384 ( .A(n9349), .ZN(n9350) );
  AOI21_X1 U10385 ( .B1(n9357), .B2(n9351), .A(n9350), .ZN(n9547) );
  INV_X1 U10386 ( .A(n9352), .ZN(n9354) );
  AOI21_X1 U10387 ( .B1(n9543), .B2(n9354), .A(n9353), .ZN(n9544) );
  AOI22_X1 U10388 ( .A1(n9355), .A2(n9492), .B1(n9426), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n9356) );
  OAI21_X1 U10389 ( .B1(n8025), .B2(n9495), .A(n9356), .ZN(n9363) );
  XNOR2_X1 U10390 ( .A(n9358), .B(n9357), .ZN(n9361) );
  AOI222_X1 U10391 ( .A1(n10923), .A2(n9361), .B1(n9360), .B2(n9501), .C1(
        n9359), .C2(n9499), .ZN(n9546) );
  NOR2_X1 U10392 ( .A1(n9546), .A2(n9504), .ZN(n9362) );
  AOI211_X1 U10393 ( .C1(n9544), .C2(n9507), .A(n9363), .B(n9362), .ZN(n9364)
         );
  OAI21_X1 U10394 ( .B1(n9547), .B2(n9509), .A(n9364), .ZN(P2_U3272) );
  OAI21_X1 U10395 ( .B1(n9366), .B2(n8057), .A(n9365), .ZN(n9368) );
  AOI222_X1 U10396 ( .A1(n10923), .A2(n9368), .B1(n9367), .B2(n9501), .C1(
        n9395), .C2(n9499), .ZN(n9552) );
  OR2_X1 U10397 ( .A1(n9370), .A2(n9369), .ZN(n9548) );
  NAND3_X1 U10398 ( .A1(n9548), .A2(n9371), .A3(n9400), .ZN(n9378) );
  XNOR2_X1 U10399 ( .A(n9375), .B(n9381), .ZN(n9550) );
  INV_X1 U10400 ( .A(n9372), .ZN(n9373) );
  AOI22_X1 U10401 ( .A1(n9426), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9373), .B2(
        n9492), .ZN(n9374) );
  OAI21_X1 U10402 ( .B1(n9375), .B2(n9495), .A(n9374), .ZN(n9376) );
  AOI21_X1 U10403 ( .B1(n9550), .B2(n9507), .A(n9376), .ZN(n9377) );
  OAI211_X1 U10404 ( .C1(n9504), .C2(n9552), .A(n9378), .B(n9377), .ZN(
        P2_U3273) );
  XNOR2_X1 U10405 ( .A(n9380), .B(n9379), .ZN(n9558) );
  INV_X1 U10406 ( .A(n9381), .ZN(n9382) );
  AOI21_X1 U10407 ( .B1(n9554), .B2(n9402), .A(n9382), .ZN(n9555) );
  AOI22_X1 U10408 ( .A1(n9426), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9383), .B2(
        n9492), .ZN(n9384) );
  OAI21_X1 U10409 ( .B1(n9385), .B2(n9495), .A(n9384), .ZN(n9391) );
  XNOR2_X1 U10410 ( .A(n9387), .B(n9386), .ZN(n9389) );
  AOI21_X1 U10411 ( .B1(n9389), .B2(n10923), .A(n9388), .ZN(n9557) );
  NOR2_X1 U10412 ( .A1(n9557), .A2(n9504), .ZN(n9390) );
  AOI211_X1 U10413 ( .C1(n9555), .C2(n9507), .A(n9391), .B(n9390), .ZN(n9392)
         );
  OAI21_X1 U10414 ( .B1(n9558), .B2(n9509), .A(n9392), .ZN(P2_U3274) );
  XOR2_X1 U10415 ( .A(n9398), .B(n9393), .Z(n9396) );
  AOI222_X1 U10416 ( .A1(n10923), .A2(n9396), .B1(n9395), .B2(n9501), .C1(
        n9394), .C2(n9499), .ZN(n9996) );
  OAI21_X1 U10417 ( .B1(n9399), .B2(n9398), .A(n9397), .ZN(n9992) );
  NAND2_X1 U10418 ( .A1(n9992), .A2(n9400), .ZN(n9411) );
  INV_X1 U10419 ( .A(n9401), .ZN(n9404) );
  INV_X1 U10420 ( .A(n9402), .ZN(n9403) );
  AOI21_X1 U10421 ( .B1(n9993), .B2(n9404), .A(n9403), .ZN(n9994) );
  NOR2_X1 U10422 ( .A1(n9405), .A2(n9495), .ZN(n9409) );
  OAI22_X1 U10423 ( .A1(n10946), .A2(n9407), .B1(n9406), .B2(n10935), .ZN(
        n9408) );
  AOI211_X1 U10424 ( .C1(n9994), .C2(n9507), .A(n9409), .B(n9408), .ZN(n9410)
         );
  OAI211_X1 U10425 ( .C1(n9504), .C2(n9996), .A(n9411), .B(n9410), .ZN(
        P2_U3275) );
  OAI21_X1 U10426 ( .B1(n9416), .B2(n9412), .A(n5124), .ZN(n10002) );
  XOR2_X1 U10427 ( .A(n9998), .B(n9432), .Z(n9999) );
  AOI22_X1 U10428 ( .A1(n9426), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9413), .B2(
        n9492), .ZN(n9414) );
  OAI21_X1 U10429 ( .B1(n9415), .B2(n9495), .A(n9414), .ZN(n9421) );
  XNOR2_X1 U10430 ( .A(n9417), .B(n9416), .ZN(n9419) );
  AOI222_X1 U10431 ( .A1(n10923), .A2(n9419), .B1(n9418), .B2(n9501), .C1(
        n9448), .C2(n9499), .ZN(n10001) );
  NOR2_X1 U10432 ( .A1(n10001), .A2(n9504), .ZN(n9420) );
  AOI211_X1 U10433 ( .C1(n9999), .C2(n9507), .A(n9421), .B(n9420), .ZN(n9422)
         );
  OAI21_X1 U10434 ( .B1(n10002), .B2(n9509), .A(n9422), .ZN(P2_U3276) );
  OAI21_X1 U10435 ( .B1(n9425), .B2(n9424), .A(n9423), .ZN(n10007) );
  AOI22_X1 U10436 ( .A1(n10005), .A2(n9427), .B1(P2_REG2_REG_19__SCAN_IN), 
        .B2(n9426), .ZN(n9437) );
  XNOR2_X1 U10437 ( .A(n9429), .B(n9428), .ZN(n9430) );
  OAI222_X1 U10438 ( .A1(n9468), .A2(n9431), .B1(n9466), .B2(n9467), .C1(n9486), .C2(n9430), .ZN(n10003) );
  AOI211_X1 U10439 ( .C1(n10005), .C2(n9439), .A(n11011), .B(n5468), .ZN(
        n10004) );
  INV_X1 U10440 ( .A(n10004), .ZN(n9434) );
  OAI22_X1 U10441 ( .A1(n9434), .A2(n5819), .B1(n10935), .B2(n9433), .ZN(n9435) );
  OAI21_X1 U10442 ( .B1(n10003), .B2(n9435), .A(n10946), .ZN(n9436) );
  OAI211_X1 U10443 ( .C1(n10007), .C2(n9509), .A(n9437), .B(n9436), .ZN(
        P2_U3277) );
  XNOR2_X1 U10444 ( .A(n9438), .B(n5641), .ZN(n10012) );
  INV_X1 U10445 ( .A(n9457), .ZN(n9441) );
  INV_X1 U10446 ( .A(n9439), .ZN(n9440) );
  AOI21_X1 U10447 ( .B1(n10008), .B2(n9441), .A(n9440), .ZN(n10009) );
  AOI22_X1 U10448 ( .A1(n9426), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9442), .B2(
        n9492), .ZN(n9443) );
  OAI21_X1 U10449 ( .B1(n9444), .B2(n9495), .A(n9443), .ZN(n9451) );
  XNOR2_X1 U10450 ( .A(n9446), .B(n9445), .ZN(n9449) );
  AOI222_X1 U10451 ( .A1(n10923), .A2(n9449), .B1(n9448), .B2(n9501), .C1(
        n9447), .C2(n9499), .ZN(n10011) );
  NOR2_X1 U10452 ( .A1(n10011), .A2(n9504), .ZN(n9450) );
  AOI211_X1 U10453 ( .C1(n10009), .C2(n9507), .A(n9451), .B(n9450), .ZN(n9452)
         );
  OAI21_X1 U10454 ( .B1(n10012), .B2(n9509), .A(n9452), .ZN(P2_U3278) );
  OAI21_X1 U10455 ( .B1(n9455), .B2(n9454), .A(n9453), .ZN(n9456) );
  INV_X1 U10456 ( .A(n9456), .ZN(n10017) );
  AOI211_X1 U10457 ( .C1(n10015), .C2(n9474), .A(n11011), .B(n9457), .ZN(
        n10014) );
  INV_X1 U10458 ( .A(n10015), .ZN(n9458) );
  NOR2_X1 U10459 ( .A1(n9458), .A2(n9495), .ZN(n9461) );
  OAI22_X1 U10460 ( .A1(n10946), .A2(n7588), .B1(n9459), .B2(n10935), .ZN(
        n9460) );
  AOI211_X1 U10461 ( .C1(n10014), .C2(n9481), .A(n9461), .B(n9460), .ZN(n9470)
         );
  XNOR2_X1 U10462 ( .A(n9463), .B(n9462), .ZN(n9464) );
  OAI222_X1 U10463 ( .A1(n9468), .A2(n9467), .B1(n9466), .B2(n9465), .C1(n9464), .C2(n9486), .ZN(n10013) );
  NAND2_X1 U10464 ( .A1(n10013), .A2(n10946), .ZN(n9469) );
  OAI211_X1 U10465 ( .C1(n10017), .C2(n9509), .A(n9470), .B(n9469), .ZN(
        P2_U3279) );
  AOI21_X1 U10466 ( .B1(n9472), .B2(n9471), .A(n5126), .ZN(n9473) );
  INV_X1 U10467 ( .A(n9473), .ZN(n10022) );
  INV_X1 U10468 ( .A(n9474), .ZN(n9475) );
  AOI211_X1 U10469 ( .C1(n10020), .C2(n9476), .A(n11011), .B(n9475), .ZN(
        n10019) );
  INV_X1 U10470 ( .A(n10020), .ZN(n9477) );
  NOR2_X1 U10471 ( .A1(n9477), .A2(n9495), .ZN(n9480) );
  OAI22_X1 U10472 ( .A1(n10946), .A2(n7255), .B1(n9478), .B2(n10935), .ZN(
        n9479) );
  AOI211_X1 U10473 ( .C1(n10019), .C2(n9481), .A(n9480), .B(n9479), .ZN(n9489)
         );
  AOI21_X1 U10474 ( .B1(n9498), .B2(n9483), .A(n9482), .ZN(n9484) );
  XNOR2_X1 U10475 ( .A(n9484), .B(n5176), .ZN(n9487) );
  OAI21_X1 U10476 ( .B1(n9487), .B2(n9486), .A(n9485), .ZN(n10018) );
  NAND2_X1 U10477 ( .A1(n10018), .A2(n10946), .ZN(n9488) );
  OAI211_X1 U10478 ( .C1(n10022), .C2(n9509), .A(n9489), .B(n9488), .ZN(
        P2_U3280) );
  XNOR2_X1 U10479 ( .A(n9490), .B(n9497), .ZN(n10027) );
  XOR2_X1 U10480 ( .A(n10023), .B(n9491), .Z(n10024) );
  INV_X1 U10481 ( .A(n10023), .ZN(n9496) );
  AOI22_X1 U10482 ( .A1(n9426), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9493), .B2(
        n9492), .ZN(n9494) );
  OAI21_X1 U10483 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9506) );
  XNOR2_X1 U10484 ( .A(n9498), .B(n9497), .ZN(n9503) );
  AOI222_X1 U10485 ( .A1(n10923), .A2(n9503), .B1(n9502), .B2(n9501), .C1(
        n9500), .C2(n9499), .ZN(n10026) );
  NOR2_X1 U10486 ( .A1(n10026), .A2(n9504), .ZN(n9505) );
  AOI211_X1 U10487 ( .C1(n10024), .C2(n9507), .A(n9506), .B(n9505), .ZN(n9508)
         );
  OAI21_X1 U10488 ( .B1(n10027), .B2(n9509), .A(n9508), .ZN(P2_U3281) );
  AOI21_X1 U10489 ( .B1(n9510), .B2(n10925), .A(n9513), .ZN(n9511) );
  OAI21_X1 U10490 ( .B1(n9512), .B2(n11011), .A(n9511), .ZN(n10028) );
  MUX2_X1 U10491 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n10028), .S(n11018), .Z(
        P2_U3551) );
  AOI21_X1 U10492 ( .B1(n9514), .B2(n10925), .A(n9513), .ZN(n9515) );
  OAI21_X1 U10493 ( .B1(n9516), .B2(n11011), .A(n9515), .ZN(n10029) );
  MUX2_X1 U10494 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n10029), .S(n11018), .Z(
        P2_U3550) );
  NAND2_X1 U10495 ( .A1(n9517), .A2(n11015), .ZN(n9522) );
  NOR2_X1 U10496 ( .A1(n9518), .A2(n11011), .ZN(n9520) );
  AOI22_X1 U10497 ( .A1(n9524), .A2(n10927), .B1(n9523), .B2(n10925), .ZN(
        n9525) );
  OAI211_X1 U10498 ( .C1(n9527), .C2(n10992), .A(n9526), .B(n9525), .ZN(n10031) );
  MUX2_X1 U10499 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n10031), .S(n11018), .Z(
        P2_U3548) );
  AOI22_X1 U10500 ( .A1(n9529), .A2(n10927), .B1(n9528), .B2(n10925), .ZN(
        n9530) );
  OAI211_X1 U10501 ( .C1(n9532), .C2(n10992), .A(n9531), .B(n9530), .ZN(n10032) );
  MUX2_X1 U10502 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n10032), .S(n11018), .Z(
        P2_U3547) );
  AOI21_X1 U10503 ( .B1(n9534), .B2(n10925), .A(n9533), .ZN(n9535) );
  OAI211_X1 U10504 ( .C1(n9537), .C2(n10992), .A(n9536), .B(n9535), .ZN(n10033) );
  MUX2_X1 U10505 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n10033), .S(n11018), .Z(
        P2_U3546) );
  AOI211_X1 U10506 ( .C1(n9540), .C2(n10925), .A(n9539), .B(n9538), .ZN(n9541)
         );
  OAI21_X1 U10507 ( .B1(n9542), .B2(n10992), .A(n9541), .ZN(n10034) );
  MUX2_X1 U10508 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n10034), .S(n11018), .Z(
        P2_U3545) );
  AOI22_X1 U10509 ( .A1(n9544), .A2(n10927), .B1(n9543), .B2(n10925), .ZN(
        n9545) );
  OAI211_X1 U10510 ( .C1(n9547), .C2(n10992), .A(n9546), .B(n9545), .ZN(n10035) );
  MUX2_X1 U10511 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n10035), .S(n11018), .Z(
        P2_U3544) );
  NAND3_X1 U10512 ( .A1(n9548), .A2(n9371), .A3(n11015), .ZN(n9553) );
  AOI22_X1 U10513 ( .A1(n9550), .A2(n10927), .B1(n9549), .B2(n10925), .ZN(
        n9551) );
  NAND3_X1 U10514 ( .A1(n9553), .A2(n9552), .A3(n9551), .ZN(n10036) );
  MUX2_X1 U10515 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n10036), .S(n11018), .Z(
        P2_U3543) );
  AOI22_X1 U10516 ( .A1(n9555), .A2(n10927), .B1(n9554), .B2(n10925), .ZN(
        n9556) );
  OAI211_X1 U10517 ( .C1(n9558), .C2(n10992), .A(n9557), .B(n9556), .ZN(n10037) );
  MUX2_X1 U10518 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n10037), .S(n11018), .Z(
        n9991) );
  XOR2_X1 U10519 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n9563) );
  XNOR2_X1 U10520 ( .A(n9559), .B(keyinput_130), .ZN(n9562) );
  XNOR2_X1 U10521 ( .A(n9767), .B(keyinput_129), .ZN(n9561) );
  XNOR2_X1 U10522 ( .A(SI_29_), .B(keyinput_131), .ZN(n9560) );
  NAND4_X1 U10523 ( .A1(n9563), .A2(n9562), .A3(n9561), .A4(n9560), .ZN(n9567)
         );
  XNOR2_X1 U10524 ( .A(n9564), .B(keyinput_132), .ZN(n9566) );
  XNOR2_X1 U10525 ( .A(n9772), .B(keyinput_133), .ZN(n9565) );
  NAND3_X1 U10526 ( .A1(n9567), .A2(n9566), .A3(n9565), .ZN(n9575) );
  XNOR2_X1 U10527 ( .A(n9776), .B(keyinput_134), .ZN(n9574) );
  XNOR2_X1 U10528 ( .A(n9568), .B(keyinput_136), .ZN(n9572) );
  XNOR2_X1 U10529 ( .A(n9777), .B(keyinput_135), .ZN(n9571) );
  XNOR2_X1 U10530 ( .A(n9569), .B(keyinput_137), .ZN(n9570) );
  NAND3_X1 U10531 ( .A1(n9572), .A2(n9571), .A3(n9570), .ZN(n9573) );
  AOI21_X1 U10532 ( .B1(n9575), .B2(n9574), .A(n9573), .ZN(n9578) );
  XNOR2_X1 U10533 ( .A(SI_22_), .B(keyinput_138), .ZN(n9577) );
  XNOR2_X1 U10534 ( .A(SI_21_), .B(keyinput_139), .ZN(n9576) );
  NOR3_X1 U10535 ( .A1(n9578), .A2(n9577), .A3(n9576), .ZN(n9587) );
  XNOR2_X1 U10536 ( .A(n9579), .B(keyinput_143), .ZN(n9586) );
  XNOR2_X1 U10537 ( .A(SI_18_), .B(keyinput_142), .ZN(n9585) );
  XNOR2_X1 U10538 ( .A(SI_20_), .B(keyinput_140), .ZN(n9583) );
  XNOR2_X1 U10539 ( .A(SI_16_), .B(keyinput_144), .ZN(n9582) );
  XNOR2_X1 U10540 ( .A(SI_19_), .B(keyinput_141), .ZN(n9581) );
  XNOR2_X1 U10541 ( .A(SI_15_), .B(keyinput_145), .ZN(n9580) );
  NAND4_X1 U10542 ( .A1(n9583), .A2(n9582), .A3(n9581), .A4(n9580), .ZN(n9584)
         );
  NOR4_X1 U10543 ( .A1(n9587), .A2(n9586), .A3(n9585), .A4(n9584), .ZN(n9592)
         );
  XNOR2_X1 U10544 ( .A(n9588), .B(keyinput_146), .ZN(n9591) );
  XNOR2_X1 U10545 ( .A(n9589), .B(keyinput_147), .ZN(n9590) );
  OAI21_X1 U10546 ( .B1(n9592), .B2(n9591), .A(n9590), .ZN(n9595) );
  XNOR2_X1 U10547 ( .A(SI_12_), .B(keyinput_148), .ZN(n9594) );
  XNOR2_X1 U10548 ( .A(n9800), .B(keyinput_149), .ZN(n9593) );
  AOI21_X1 U10549 ( .B1(n9595), .B2(n9594), .A(n9593), .ZN(n9598) );
  XNOR2_X1 U10550 ( .A(SI_10_), .B(keyinput_150), .ZN(n9597) );
  XNOR2_X1 U10551 ( .A(SI_9_), .B(keyinput_151), .ZN(n9596) );
  NOR3_X1 U10552 ( .A1(n9598), .A2(n9597), .A3(n9596), .ZN(n9601) );
  XNOR2_X1 U10553 ( .A(n9808), .B(keyinput_152), .ZN(n9600) );
  XNOR2_X1 U10554 ( .A(SI_7_), .B(keyinput_153), .ZN(n9599) );
  NOR3_X1 U10555 ( .A1(n9601), .A2(n9600), .A3(n9599), .ZN(n9610) );
  XOR2_X1 U10556 ( .A(SI_6_), .B(keyinput_154), .Z(n9606) );
  XNOR2_X1 U10557 ( .A(n9602), .B(keyinput_157), .ZN(n9605) );
  XNOR2_X1 U10558 ( .A(SI_4_), .B(keyinput_156), .ZN(n9604) );
  XNOR2_X1 U10559 ( .A(SI_5_), .B(keyinput_155), .ZN(n9603) );
  NAND4_X1 U10560 ( .A1(n9606), .A2(n9605), .A3(n9604), .A4(n9603), .ZN(n9609)
         );
  XNOR2_X1 U10561 ( .A(n9817), .B(keyinput_159), .ZN(n9608) );
  XNOR2_X1 U10562 ( .A(SI_2_), .B(keyinput_158), .ZN(n9607) );
  OAI211_X1 U10563 ( .C1(n9610), .C2(n9609), .A(n9608), .B(n9607), .ZN(n9618)
         );
  XNOR2_X1 U10564 ( .A(n9611), .B(keyinput_161), .ZN(n9615) );
  XNOR2_X1 U10565 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n9614)
         );
  XNOR2_X1 U10566 ( .A(SI_0_), .B(keyinput_160), .ZN(n9613) );
  XNOR2_X1 U10567 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_162), .ZN(n9612) );
  NOR4_X1 U10568 ( .A1(n9615), .A2(n9614), .A3(n9613), .A4(n9612), .ZN(n9617)
         );
  XNOR2_X1 U10569 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n9616)
         );
  AOI21_X1 U10570 ( .B1(n9618), .B2(n9617), .A(n9616), .ZN(n9623) );
  XNOR2_X1 U10571 ( .A(n9619), .B(keyinput_165), .ZN(n9622) );
  XNOR2_X1 U10572 ( .A(n9620), .B(keyinput_166), .ZN(n9621) );
  OAI21_X1 U10573 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9627) );
  XNOR2_X1 U10574 ( .A(n9624), .B(keyinput_167), .ZN(n9626) );
  XOR2_X1 U10575 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .Z(n9625) );
  AOI21_X1 U10576 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(n9630) );
  XNOR2_X1 U10577 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n9629)
         );
  XNOR2_X1 U10578 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n9628)
         );
  OAI21_X1 U10579 ( .B1(n9630), .B2(n9629), .A(n9628), .ZN(n9633) );
  XNOR2_X1 U10580 ( .A(n9841), .B(keyinput_171), .ZN(n9632) );
  XNOR2_X1 U10581 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n9631)
         );
  NAND3_X1 U10582 ( .A1(n9633), .A2(n9632), .A3(n9631), .ZN(n9640) );
  XNOR2_X1 U10583 ( .A(n9845), .B(keyinput_173), .ZN(n9639) );
  XNOR2_X1 U10584 ( .A(n9846), .B(keyinput_176), .ZN(n9637) );
  XNOR2_X1 U10585 ( .A(n9634), .B(keyinput_175), .ZN(n9636) );
  XNOR2_X1 U10586 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n9635)
         );
  NAND3_X1 U10587 ( .A1(n9637), .A2(n9636), .A3(n9635), .ZN(n9638) );
  AOI21_X1 U10588 ( .B1(n9640), .B2(n9639), .A(n9638), .ZN(n9649) );
  XOR2_X1 U10589 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .Z(n9644) );
  XNOR2_X1 U10590 ( .A(n9853), .B(keyinput_177), .ZN(n9643) );
  XNOR2_X1 U10591 ( .A(n9854), .B(keyinput_179), .ZN(n9642) );
  XNOR2_X1 U10592 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n9641)
         );
  NAND4_X1 U10593 ( .A1(n9644), .A2(n9643), .A3(n9642), .A4(n9641), .ZN(n9648)
         );
  XNOR2_X1 U10594 ( .A(n9645), .B(keyinput_181), .ZN(n9647) );
  XNOR2_X1 U10595 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n9646)
         );
  OAI211_X1 U10596 ( .C1(n9649), .C2(n9648), .A(n9647), .B(n9646), .ZN(n9653)
         );
  XNOR2_X1 U10597 ( .A(n9650), .B(keyinput_183), .ZN(n9652) );
  XNOR2_X1 U10598 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n9651)
         );
  AOI21_X1 U10599 ( .B1(n9653), .B2(n9652), .A(n9651), .ZN(n9656) );
  XNOR2_X1 U10600 ( .A(n9867), .B(keyinput_185), .ZN(n9655) );
  XNOR2_X1 U10601 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n9654)
         );
  OAI21_X1 U10602 ( .B1(n9656), .B2(n9655), .A(n9654), .ZN(n9660) );
  XOR2_X1 U10603 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n9659) );
  XNOR2_X1 U10604 ( .A(n9871), .B(keyinput_189), .ZN(n9658) );
  XNOR2_X1 U10605 ( .A(n9872), .B(keyinput_188), .ZN(n9657) );
  NAND4_X1 U10606 ( .A1(n9660), .A2(n9659), .A3(n9658), .A4(n9657), .ZN(n9663)
         );
  XNOR2_X1 U10607 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_190), .ZN(n9662)
         );
  XNOR2_X1 U10608 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n9661)
         );
  AOI21_X1 U10609 ( .B1(n9663), .B2(n9662), .A(n9661), .ZN(n9674) );
  XOR2_X1 U10610 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .Z(n9667) );
  XOR2_X1 U10611 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .Z(n9666)
         );
  XNOR2_X1 U10612 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n9665)
         );
  XNOR2_X1 U10613 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n9664)
         );
  NAND4_X1 U10614 ( .A1(n9667), .A2(n9666), .A3(n9665), .A4(n9664), .ZN(n9673)
         );
  XNOR2_X1 U10615 ( .A(n9887), .B(keyinput_197), .ZN(n9672) );
  OAI22_X1 U10616 ( .A1(n9670), .A2(keyinput_198), .B1(keyinput_196), .B2(
        P2_DATAO_REG_28__SCAN_IN), .ZN(n9669) );
  AND2_X1 U10617 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_196), .ZN(n9668) );
  AOI211_X1 U10618 ( .C1(keyinput_198), .C2(n9670), .A(n9669), .B(n9668), .ZN(
        n9671) );
  OAI211_X1 U10619 ( .C1(n9674), .C2(n9673), .A(n9672), .B(n9671), .ZN(n9678)
         );
  XNOR2_X1 U10620 ( .A(n9892), .B(keyinput_199), .ZN(n9677) );
  XOR2_X1 U10621 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .Z(n9676)
         );
  XNOR2_X1 U10622 ( .A(n9893), .B(keyinput_201), .ZN(n9675) );
  AOI211_X1 U10623 ( .C1(n9678), .C2(n9677), .A(n9676), .B(n9675), .ZN(n9682)
         );
  XNOR2_X1 U10624 ( .A(n9679), .B(keyinput_202), .ZN(n9681) );
  XOR2_X1 U10625 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n9680)
         );
  OAI21_X1 U10626 ( .B1(n9682), .B2(n9681), .A(n9680), .ZN(n9688) );
  XNOR2_X1 U10627 ( .A(n9683), .B(keyinput_205), .ZN(n9687) );
  XNOR2_X1 U10628 ( .A(n9684), .B(keyinput_204), .ZN(n9686) );
  XOR2_X1 U10629 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .Z(n9685)
         );
  NAND4_X1 U10630 ( .A1(n9688), .A2(n9687), .A3(n9686), .A4(n9685), .ZN(n9691)
         );
  XNOR2_X1 U10631 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n9690)
         );
  XNOR2_X1 U10632 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .ZN(n9689)
         );
  NAND3_X1 U10633 ( .A1(n9691), .A2(n9690), .A3(n9689), .ZN(n9694) );
  XNOR2_X1 U10634 ( .A(n9908), .B(keyinput_209), .ZN(n9693) );
  XNOR2_X1 U10635 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .ZN(n9692)
         );
  AOI21_X1 U10636 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9698) );
  XNOR2_X1 U10637 ( .A(n9912), .B(keyinput_211), .ZN(n9697) );
  XNOR2_X1 U10638 ( .A(n9695), .B(keyinput_212), .ZN(n9696) );
  OAI21_X1 U10639 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9701) );
  XOR2_X1 U10640 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .Z(n9700)
         );
  XNOR2_X1 U10641 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n9699)
         );
  NAND3_X1 U10642 ( .A1(n9701), .A2(n9700), .A3(n9699), .ZN(n9704) );
  XNOR2_X1 U10643 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .ZN(n9703)
         );
  XNOR2_X1 U10644 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .ZN(n9702)
         );
  NAND3_X1 U10645 ( .A1(n9704), .A2(n9703), .A3(n9702), .ZN(n9707) );
  XNOR2_X1 U10646 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .ZN(n9706)
         );
  XNOR2_X1 U10647 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_218), .ZN(n9705)
         );
  AOI21_X1 U10648 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9710) );
  XNOR2_X1 U10649 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_220), .ZN(n9709) );
  XNOR2_X1 U10650 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_219), .ZN(n9708) );
  NOR3_X1 U10651 ( .A1(n9710), .A2(n9709), .A3(n9708), .ZN(n9717) );
  XNOR2_X1 U10652 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_222), .ZN(n9714) );
  XNOR2_X1 U10653 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_221), .ZN(n9713) );
  XNOR2_X1 U10654 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_223), .ZN(n9712) );
  XNOR2_X1 U10655 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_224), .ZN(n9711) );
  NAND4_X1 U10656 ( .A1(n9714), .A2(n9713), .A3(n9712), .A4(n9711), .ZN(n9716)
         );
  XNOR2_X1 U10657 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_225), .ZN(n9715) );
  OAI21_X1 U10658 ( .B1(n9717), .B2(n9716), .A(n9715), .ZN(n9724) );
  XNOR2_X1 U10659 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_227), .ZN(n9719) );
  XNOR2_X1 U10660 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_226), .ZN(n9718) );
  NOR2_X1 U10661 ( .A1(n9719), .A2(n9718), .ZN(n9723) );
  XNOR2_X1 U10662 ( .A(n9720), .B(keyinput_229), .ZN(n9722) );
  XOR2_X1 U10663 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_228), .Z(n9721) );
  AOI211_X1 U10664 ( .C1(n9724), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9728)
         );
  XNOR2_X1 U10665 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_230), .ZN(n9727) );
  XNOR2_X1 U10666 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_231), .ZN(n9726) );
  XNOR2_X1 U10667 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_232), .ZN(n9725) );
  NOR4_X1 U10668 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n9732)
         );
  XNOR2_X1 U10669 ( .A(n9729), .B(keyinput_233), .ZN(n9731) );
  XNOR2_X1 U10670 ( .A(n5746), .B(keyinput_234), .ZN(n9730) );
  OAI21_X1 U10671 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9737) );
  XNOR2_X1 U10672 ( .A(n9733), .B(keyinput_235), .ZN(n9736) );
  XNOR2_X1 U10673 ( .A(n9734), .B(keyinput_236), .ZN(n9735) );
  AOI21_X1 U10674 ( .B1(n9737), .B2(n9736), .A(n9735), .ZN(n9742) );
  XNOR2_X1 U10675 ( .A(n9738), .B(keyinput_238), .ZN(n9741) );
  XNOR2_X1 U10676 ( .A(n9954), .B(keyinput_239), .ZN(n9740) );
  XNOR2_X1 U10677 ( .A(n9956), .B(keyinput_237), .ZN(n9739) );
  NOR4_X1 U10678 ( .A1(n9742), .A2(n9741), .A3(n9740), .A4(n9739), .ZN(n9751)
         );
  XNOR2_X1 U10679 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_243), .ZN(n9750) );
  XNOR2_X1 U10680 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_240), .ZN(n9749) );
  XNOR2_X1 U10681 ( .A(n9743), .B(keyinput_244), .ZN(n9747) );
  XNOR2_X1 U10682 ( .A(n9744), .B(keyinput_241), .ZN(n9746) );
  XNOR2_X1 U10683 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_242), .ZN(n9745) );
  NAND3_X1 U10684 ( .A1(n9747), .A2(n9746), .A3(n9745), .ZN(n9748) );
  NOR4_X1 U10685 ( .A1(n9751), .A2(n9750), .A3(n9749), .A4(n9748), .ZN(n9754)
         );
  XNOR2_X1 U10686 ( .A(n9967), .B(keyinput_246), .ZN(n9753) );
  XNOR2_X1 U10687 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_245), .ZN(n9752) );
  NOR3_X1 U10688 ( .A1(n9754), .A2(n9753), .A3(n9752), .ZN(n9758) );
  XNOR2_X1 U10689 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_247), .ZN(n9757) );
  XOR2_X1 U10690 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_249), .Z(n9756) );
  XNOR2_X1 U10691 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_248), .ZN(n9755) );
  OAI211_X1 U10692 ( .C1(n9758), .C2(n9757), .A(n9756), .B(n9755), .ZN(n9760)
         );
  XNOR2_X1 U10693 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_250), .ZN(n9759) );
  NAND2_X1 U10694 ( .A1(n9760), .A2(n9759), .ZN(n9766) );
  INV_X1 U10695 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10535) );
  OAI22_X1 U10696 ( .A1(n10535), .A2(keyinput_253), .B1(keyinput_252), .B2(
        P1_D_REG_1__SCAN_IN), .ZN(n9761) );
  AOI221_X1 U10697 ( .B1(n10535), .B2(keyinput_253), .C1(P1_D_REG_1__SCAN_IN), 
        .C2(keyinput_252), .A(n9761), .ZN(n9765) );
  XOR2_X1 U10698 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_255), .Z(n9764) );
  INV_X1 U10699 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10536) );
  OAI22_X1 U10700 ( .A1(n10536), .A2(keyinput_254), .B1(P1_D_REG_0__SCAN_IN), 
        .B2(keyinput_251), .ZN(n9762) );
  AOI221_X1 U10701 ( .B1(n10536), .B2(keyinput_254), .C1(keyinput_251), .C2(
        P1_D_REG_0__SCAN_IN), .A(n9762), .ZN(n9763) );
  NAND4_X1 U10702 ( .A1(n9766), .A2(n9765), .A3(n9764), .A4(n9763), .ZN(n9989)
         );
  XOR2_X1 U10703 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n9771) );
  XNOR2_X1 U10704 ( .A(n9767), .B(keyinput_1), .ZN(n9770) );
  XNOR2_X1 U10705 ( .A(SI_30_), .B(keyinput_2), .ZN(n9769) );
  XNOR2_X1 U10706 ( .A(SI_29_), .B(keyinput_3), .ZN(n9768) );
  NAND4_X1 U10707 ( .A1(n9771), .A2(n9770), .A3(n9769), .A4(n9768), .ZN(n9775)
         );
  XNOR2_X1 U10708 ( .A(n9772), .B(keyinput_5), .ZN(n9774) );
  XNOR2_X1 U10709 ( .A(SI_28_), .B(keyinput_4), .ZN(n9773) );
  NAND3_X1 U10710 ( .A1(n9775), .A2(n9774), .A3(n9773), .ZN(n9783) );
  XNOR2_X1 U10711 ( .A(n9776), .B(keyinput_6), .ZN(n9782) );
  XNOR2_X1 U10712 ( .A(n9777), .B(keyinput_7), .ZN(n9780) );
  XNOR2_X1 U10713 ( .A(SI_23_), .B(keyinput_9), .ZN(n9779) );
  XNOR2_X1 U10714 ( .A(SI_24_), .B(keyinput_8), .ZN(n9778) );
  NAND3_X1 U10715 ( .A1(n9780), .A2(n9779), .A3(n9778), .ZN(n9781) );
  AOI21_X1 U10716 ( .B1(n9783), .B2(n9782), .A(n9781), .ZN(n9787) );
  XNOR2_X1 U10717 ( .A(n9784), .B(keyinput_10), .ZN(n9786) );
  XNOR2_X1 U10718 ( .A(SI_21_), .B(keyinput_11), .ZN(n9785) );
  NOR3_X1 U10719 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(n9795) );
  XNOR2_X1 U10720 ( .A(SI_15_), .B(keyinput_17), .ZN(n9794) );
  XNOR2_X1 U10721 ( .A(SI_20_), .B(keyinput_12), .ZN(n9793) );
  XNOR2_X1 U10722 ( .A(SI_17_), .B(keyinput_15), .ZN(n9791) );
  XNOR2_X1 U10723 ( .A(SI_18_), .B(keyinput_14), .ZN(n9790) );
  XNOR2_X1 U10724 ( .A(SI_19_), .B(keyinput_13), .ZN(n9789) );
  XNOR2_X1 U10725 ( .A(SI_16_), .B(keyinput_16), .ZN(n9788) );
  NAND4_X1 U10726 ( .A1(n9791), .A2(n9790), .A3(n9789), .A4(n9788), .ZN(n9792)
         );
  NOR4_X1 U10727 ( .A1(n9795), .A2(n9794), .A3(n9793), .A4(n9792), .ZN(n9798)
         );
  XNOR2_X1 U10728 ( .A(SI_14_), .B(keyinput_18), .ZN(n9797) );
  XNOR2_X1 U10729 ( .A(SI_13_), .B(keyinput_19), .ZN(n9796) );
  OAI21_X1 U10730 ( .B1(n9798), .B2(n9797), .A(n9796), .ZN(n9803) );
  XNOR2_X1 U10731 ( .A(n9799), .B(keyinput_20), .ZN(n9802) );
  XNOR2_X1 U10732 ( .A(n9800), .B(keyinput_21), .ZN(n9801) );
  AOI21_X1 U10733 ( .B1(n9803), .B2(n9802), .A(n9801), .ZN(n9807) );
  XNOR2_X1 U10734 ( .A(n9804), .B(keyinput_23), .ZN(n9806) );
  XNOR2_X1 U10735 ( .A(SI_10_), .B(keyinput_22), .ZN(n9805) );
  NOR3_X1 U10736 ( .A1(n9807), .A2(n9806), .A3(n9805), .ZN(n9811) );
  XNOR2_X1 U10737 ( .A(n9808), .B(keyinput_24), .ZN(n9810) );
  XOR2_X1 U10738 ( .A(SI_7_), .B(keyinput_25), .Z(n9809) );
  NOR3_X1 U10739 ( .A1(n9811), .A2(n9810), .A3(n9809), .ZN(n9822) );
  XNOR2_X1 U10740 ( .A(n9812), .B(keyinput_28), .ZN(n9816) );
  XNOR2_X1 U10741 ( .A(SI_6_), .B(keyinput_26), .ZN(n9815) );
  XNOR2_X1 U10742 ( .A(SI_3_), .B(keyinput_29), .ZN(n9814) );
  XNOR2_X1 U10743 ( .A(SI_5_), .B(keyinput_27), .ZN(n9813) );
  NAND4_X1 U10744 ( .A1(n9816), .A2(n9815), .A3(n9814), .A4(n9813), .ZN(n9821)
         );
  XNOR2_X1 U10745 ( .A(n9817), .B(keyinput_31), .ZN(n9820) );
  XNOR2_X1 U10746 ( .A(n9818), .B(keyinput_30), .ZN(n9819) );
  OAI211_X1 U10747 ( .C1(n9822), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9829)
         );
  XOR2_X1 U10748 ( .A(SI_0_), .B(keyinput_32), .Z(n9826) );
  XNOR2_X1 U10749 ( .A(P2_U3152), .B(keyinput_34), .ZN(n9825) );
  XNOR2_X1 U10750 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n9824) );
  XNOR2_X1 U10751 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n9823) );
  NOR4_X1 U10752 ( .A1(n9826), .A2(n9825), .A3(n9824), .A4(n9823), .ZN(n9828)
         );
  XOR2_X1 U10753 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .Z(n9827) );
  AOI21_X1 U10754 ( .B1(n9829), .B2(n9828), .A(n9827), .ZN(n9832) );
  XNOR2_X1 U10755 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n9831)
         );
  XNOR2_X1 U10756 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n9830)
         );
  OAI21_X1 U10757 ( .B1(n9832), .B2(n9831), .A(n9830), .ZN(n9835) );
  XNOR2_X1 U10758 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n9834)
         );
  XNOR2_X1 U10759 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n9833) );
  AOI21_X1 U10760 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9840) );
  XNOR2_X1 U10761 ( .A(n9836), .B(keyinput_41), .ZN(n9839) );
  XNOR2_X1 U10762 ( .A(n9837), .B(keyinput_42), .ZN(n9838) );
  OAI21_X1 U10763 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9844) );
  XOR2_X1 U10764 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n9843) );
  XNOR2_X1 U10765 ( .A(n9841), .B(keyinput_43), .ZN(n9842) );
  NAND3_X1 U10766 ( .A1(n9844), .A2(n9843), .A3(n9842), .ZN(n9852) );
  XNOR2_X1 U10767 ( .A(n9845), .B(keyinput_45), .ZN(n9851) );
  XNOR2_X1 U10768 ( .A(n9846), .B(keyinput_48), .ZN(n9849) );
  XNOR2_X1 U10769 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n9848)
         );
  XNOR2_X1 U10770 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n9847)
         );
  NAND3_X1 U10771 ( .A1(n9849), .A2(n9848), .A3(n9847), .ZN(n9850) );
  AOI21_X1 U10772 ( .B1(n9852), .B2(n9851), .A(n9850), .ZN(n9863) );
  XNOR2_X1 U10773 ( .A(n9853), .B(keyinput_49), .ZN(n9859) );
  XNOR2_X1 U10774 ( .A(n9854), .B(keyinput_51), .ZN(n9858) );
  XNOR2_X1 U10775 ( .A(n9855), .B(keyinput_50), .ZN(n9857) );
  XNOR2_X1 U10776 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n9856) );
  NAND4_X1 U10777 ( .A1(n9859), .A2(n9858), .A3(n9857), .A4(n9856), .ZN(n9862)
         );
  XNOR2_X1 U10778 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n9861) );
  XNOR2_X1 U10779 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n9860) );
  OAI211_X1 U10780 ( .C1(n9863), .C2(n9862), .A(n9861), .B(n9860), .ZN(n9866)
         );
  XNOR2_X1 U10781 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n9865)
         );
  XNOR2_X1 U10782 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .ZN(n9864)
         );
  AOI21_X1 U10783 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(n9870) );
  XNOR2_X1 U10784 ( .A(n9867), .B(keyinput_57), .ZN(n9869) );
  XNOR2_X1 U10785 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n9868)
         );
  OAI21_X1 U10786 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9876) );
  XNOR2_X1 U10787 ( .A(n9871), .B(keyinput_61), .ZN(n9875) );
  XOR2_X1 U10788 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .Z(n9874) );
  XNOR2_X1 U10789 ( .A(n9872), .B(keyinput_60), .ZN(n9873) );
  NAND4_X1 U10790 ( .A1(n9876), .A2(n9875), .A3(n9874), .A4(n9873), .ZN(n9880)
         );
  XNOR2_X1 U10791 ( .A(n9877), .B(keyinput_62), .ZN(n9879) );
  XNOR2_X1 U10792 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_63), .ZN(n9878)
         );
  AOI21_X1 U10793 ( .B1(n9880), .B2(n9879), .A(n9878), .ZN(n9891) );
  XOR2_X1 U10794 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n9884) );
  XOR2_X1 U10795 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .Z(n9883) );
  XNOR2_X1 U10796 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .ZN(n9882)
         );
  XNOR2_X1 U10797 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .ZN(n9881) );
  NAND4_X1 U10798 ( .A1(n9884), .A2(n9883), .A3(n9882), .A4(n9881), .ZN(n9890)
         );
  OAI22_X1 U10799 ( .A1(n9887), .A2(keyinput_69), .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_70), .ZN(n9886) );
  AND2_X1 U10800 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_70), .ZN(n9885)
         );
  AOI211_X1 U10801 ( .C1(keyinput_69), .C2(n9887), .A(n9886), .B(n9885), .ZN(
        n9889) );
  XNOR2_X1 U10802 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .ZN(n9888)
         );
  OAI211_X1 U10803 ( .C1(n9891), .C2(n9890), .A(n9889), .B(n9888), .ZN(n9897)
         );
  XNOR2_X1 U10804 ( .A(n9892), .B(keyinput_71), .ZN(n9896) );
  XOR2_X1 U10805 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n9895) );
  XNOR2_X1 U10806 ( .A(n9893), .B(keyinput_73), .ZN(n9894) );
  AOI211_X1 U10807 ( .C1(n9897), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9900)
         );
  XNOR2_X1 U10808 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n9899)
         );
  XNOR2_X1 U10809 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .ZN(n9898)
         );
  OAI21_X1 U10810 ( .B1(n9900), .B2(n9899), .A(n9898), .ZN(n9904) );
  XNOR2_X1 U10811 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n9903)
         );
  XNOR2_X1 U10812 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n9902)
         );
  XNOR2_X1 U10813 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n9901)
         );
  NAND4_X1 U10814 ( .A1(n9904), .A2(n9903), .A3(n9902), .A4(n9901), .ZN(n9907)
         );
  XOR2_X1 U10815 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .Z(n9906) );
  XNOR2_X1 U10816 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n9905)
         );
  NAND3_X1 U10817 ( .A1(n9907), .A2(n9906), .A3(n9905), .ZN(n9911) );
  XNOR2_X1 U10818 ( .A(n9908), .B(keyinput_81), .ZN(n9910) );
  XNOR2_X1 U10819 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n9909)
         );
  AOI21_X1 U10820 ( .B1(n9911), .B2(n9910), .A(n9909), .ZN(n9915) );
  XNOR2_X1 U10821 ( .A(n9912), .B(keyinput_83), .ZN(n9914) );
  XNOR2_X1 U10822 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n9913)
         );
  OAI21_X1 U10823 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9919) );
  XNOR2_X1 U10824 ( .A(n9916), .B(keyinput_86), .ZN(n9918) );
  XNOR2_X1 U10825 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n9917)
         );
  NAND3_X1 U10826 ( .A1(n9919), .A2(n9918), .A3(n9917), .ZN(n9922) );
  XNOR2_X1 U10827 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .ZN(n9921)
         );
  XNOR2_X1 U10828 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n9920)
         );
  NAND3_X1 U10829 ( .A1(n9922), .A2(n9921), .A3(n9920), .ZN(n9925) );
  XNOR2_X1 U10830 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n9924)
         );
  XOR2_X1 U10831 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .Z(n9923) );
  AOI21_X1 U10832 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9928) );
  XNOR2_X1 U10833 ( .A(n10584), .B(keyinput_91), .ZN(n9927) );
  XNOR2_X1 U10834 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_92), .ZN(n9926) );
  NOR3_X1 U10835 ( .A1(n9928), .A2(n9927), .A3(n9926), .ZN(n9935) );
  XNOR2_X1 U10836 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_95), .ZN(n9932) );
  XNOR2_X1 U10837 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_94), .ZN(n9931) );
  XNOR2_X1 U10838 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_93), .ZN(n9930) );
  XNOR2_X1 U10839 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .ZN(n9929) );
  NAND4_X1 U10840 ( .A1(n9932), .A2(n9931), .A3(n9930), .A4(n9929), .ZN(n9934)
         );
  XNOR2_X1 U10841 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_97), .ZN(n9933) );
  OAI21_X1 U10842 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9939) );
  XNOR2_X1 U10843 ( .A(n9936), .B(keyinput_98), .ZN(n9938) );
  XNOR2_X1 U10844 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_99), .ZN(n9937) );
  NAND3_X1 U10845 ( .A1(n9939), .A2(n9938), .A3(n9937), .ZN(n9942) );
  XOR2_X1 U10846 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_100), .Z(n9941) );
  XNOR2_X1 U10847 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_101), .ZN(n9940) );
  NAND3_X1 U10848 ( .A1(n9942), .A2(n9941), .A3(n9940), .ZN(n9947) );
  XNOR2_X1 U10849 ( .A(n9943), .B(keyinput_103), .ZN(n9946) );
  XNOR2_X1 U10850 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_102), .ZN(n9945) );
  XNOR2_X1 U10851 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_104), .ZN(n9944) );
  NAND4_X1 U10852 ( .A1(n9947), .A2(n9946), .A3(n9945), .A4(n9944), .ZN(n9950)
         );
  XNOR2_X1 U10853 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_105), .ZN(n9949) );
  XNOR2_X1 U10854 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_106), .ZN(n9948) );
  AOI21_X1 U10855 ( .B1(n9950), .B2(n9949), .A(n9948), .ZN(n9953) );
  XNOR2_X1 U10856 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_107), .ZN(n9952) );
  XNOR2_X1 U10857 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_108), .ZN(n9951) );
  OAI21_X1 U10858 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9960) );
  XNOR2_X1 U10859 ( .A(n9954), .B(keyinput_111), .ZN(n9959) );
  OAI22_X1 U10860 ( .A1(n9956), .A2(keyinput_109), .B1(keyinput_110), .B2(
        P1_IR_REG_19__SCAN_IN), .ZN(n9955) );
  AOI21_X1 U10861 ( .B1(n9956), .B2(keyinput_109), .A(n9955), .ZN(n9958) );
  NAND2_X1 U10862 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_110), .ZN(n9957)
         );
  NAND4_X1 U10863 ( .A1(n9960), .A2(n9959), .A3(n9958), .A4(n9957), .ZN(n9971)
         );
  XNOR2_X1 U10864 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_112), .ZN(n9966) );
  XNOR2_X1 U10865 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_116), .ZN(n9962) );
  XNOR2_X1 U10866 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_114), .ZN(n9961) );
  NAND2_X1 U10867 ( .A1(n9962), .A2(n9961), .ZN(n9965) );
  XNOR2_X1 U10868 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_113), .ZN(n9964) );
  XNOR2_X1 U10869 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_115), .ZN(n9963) );
  NOR4_X1 U10870 ( .A1(n9966), .A2(n9965), .A3(n9964), .A4(n9963), .ZN(n9970)
         );
  XNOR2_X1 U10871 ( .A(n9967), .B(keyinput_118), .ZN(n9969) );
  XNOR2_X1 U10872 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_117), .ZN(n9968) );
  AOI211_X1 U10873 ( .C1(n9971), .C2(n9970), .A(n9969), .B(n9968), .ZN(n9977)
         );
  XNOR2_X1 U10874 ( .A(n9972), .B(keyinput_119), .ZN(n9976) );
  XNOR2_X1 U10875 ( .A(n9973), .B(keyinput_120), .ZN(n9975) );
  XNOR2_X1 U10876 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_121), .ZN(n9974) );
  OAI211_X1 U10877 ( .C1(n9977), .C2(n9976), .A(n9975), .B(n9974), .ZN(n9987)
         );
  XNOR2_X1 U10878 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .ZN(n9986) );
  INV_X1 U10879 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U10880 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_123), .B1(n10537), 
        .B2(keyinput_127), .ZN(n9978) );
  OAI221_X1 U10881 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_123), .C1(n10537), 
        .C2(keyinput_127), .A(n9978), .ZN(n9985) );
  INV_X1 U10882 ( .A(keyinput_124), .ZN(n9983) );
  OAI22_X1 U10883 ( .A1(n10535), .A2(keyinput_125), .B1(n9979), .B2(
        keyinput_124), .ZN(n9980) );
  AOI21_X1 U10884 ( .B1(n10535), .B2(keyinput_125), .A(n9980), .ZN(n9982) );
  XNOR2_X1 U10885 ( .A(keyinput_126), .B(P1_D_REG_3__SCAN_IN), .ZN(n9981) );
  OAI211_X1 U10886 ( .C1(P1_D_REG_1__SCAN_IN), .C2(n9983), .A(n9982), .B(n9981), .ZN(n9984) );
  AOI211_X1 U10887 ( .C1(n9987), .C2(n9986), .A(n9985), .B(n9984), .ZN(n9988)
         );
  NAND2_X1 U10888 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  XNOR2_X1 U10889 ( .A(n9991), .B(n9990), .ZN(P2_U3542) );
  INV_X1 U10890 ( .A(n9992), .ZN(n9997) );
  AOI22_X1 U10891 ( .A1(n9994), .A2(n10927), .B1(n9993), .B2(n10925), .ZN(
        n9995) );
  OAI211_X1 U10892 ( .C1(n9997), .C2(n10992), .A(n9996), .B(n9995), .ZN(n10038) );
  MUX2_X1 U10893 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n10038), .S(n11018), .Z(
        P2_U3541) );
  AOI22_X1 U10894 ( .A1(n9999), .A2(n10927), .B1(n9998), .B2(n10925), .ZN(
        n10000) );
  OAI211_X1 U10895 ( .C1(n10002), .C2(n10992), .A(n10001), .B(n10000), .ZN(
        n10039) );
  MUX2_X1 U10896 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n10039), .S(n11018), .Z(
        P2_U3540) );
  AOI211_X1 U10897 ( .C1(n10005), .C2(n10925), .A(n10004), .B(n10003), .ZN(
        n10006) );
  OAI21_X1 U10898 ( .B1(n10007), .B2(n10992), .A(n10006), .ZN(n10040) );
  MUX2_X1 U10899 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n10040), .S(n11018), .Z(
        P2_U3539) );
  AOI22_X1 U10900 ( .A1(n10009), .A2(n10927), .B1(n10008), .B2(n10925), .ZN(
        n10010) );
  OAI211_X1 U10901 ( .C1(n10012), .C2(n10992), .A(n10011), .B(n10010), .ZN(
        n10041) );
  MUX2_X1 U10902 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n10041), .S(n11018), .Z(
        P2_U3538) );
  AOI211_X1 U10903 ( .C1(n10015), .C2(n10925), .A(n10014), .B(n10013), .ZN(
        n10016) );
  OAI21_X1 U10904 ( .B1(n10017), .B2(n10992), .A(n10016), .ZN(n10042) );
  MUX2_X1 U10905 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n10042), .S(n11018), .Z(
        P2_U3537) );
  AOI211_X1 U10906 ( .C1(n10020), .C2(n10925), .A(n10019), .B(n10018), .ZN(
        n10021) );
  OAI21_X1 U10907 ( .B1(n10022), .B2(n10992), .A(n10021), .ZN(n10043) );
  MUX2_X1 U10908 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n10043), .S(n11018), .Z(
        P2_U3536) );
  AOI22_X1 U10909 ( .A1(n10024), .A2(n10927), .B1(n10023), .B2(n10925), .ZN(
        n10025) );
  OAI211_X1 U10910 ( .C1(n10027), .C2(n10992), .A(n10026), .B(n10025), .ZN(
        n10044) );
  MUX2_X1 U10911 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n10044), .S(n11018), .Z(
        P2_U3535) );
  MUX2_X1 U10912 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n10028), .S(n11001), .Z(
        P2_U3519) );
  MUX2_X1 U10913 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n10029), .S(n11001), .Z(
        P2_U3518) );
  MUX2_X1 U10914 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n10031), .S(n11001), .Z(
        P2_U3516) );
  MUX2_X1 U10915 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n10032), .S(n11001), .Z(
        P2_U3515) );
  MUX2_X1 U10916 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n10033), .S(n11001), .Z(
        P2_U3514) );
  MUX2_X1 U10917 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n10034), .S(n11001), .Z(
        P2_U3513) );
  MUX2_X1 U10918 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n10035), .S(n11001), .Z(
        P2_U3512) );
  MUX2_X1 U10919 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n10036), .S(n11001), .Z(
        P2_U3511) );
  MUX2_X1 U10920 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n10037), .S(n11001), .Z(
        P2_U3510) );
  MUX2_X1 U10921 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n10038), .S(n11001), .Z(
        P2_U3509) );
  MUX2_X1 U10922 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n10039), .S(n11001), .Z(
        P2_U3508) );
  MUX2_X1 U10923 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n10040), .S(n11001), .Z(
        P2_U3507) );
  MUX2_X1 U10924 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n10041), .S(n11001), .Z(
        P2_U3505) );
  MUX2_X1 U10925 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n10042), .S(n11001), .Z(
        P2_U3502) );
  MUX2_X1 U10926 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n10043), .S(n11001), .Z(
        P2_U3499) );
  MUX2_X1 U10927 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n10044), .S(n11001), .Z(
        P2_U3496) );
  INV_X1 U10928 ( .A(n10045), .ZN(n10527) );
  NAND3_X1 U10929 ( .A1(n10046), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n10049) );
  OAI22_X1 U10930 ( .A1(n10050), .A2(n10049), .B1(n10048), .B2(n10047), .ZN(
        n10051) );
  INV_X1 U10931 ( .A(n10051), .ZN(n10052) );
  OAI21_X1 U10932 ( .B1(n10527), .B2(n10053), .A(n10052), .ZN(P2_U3327) );
  MUX2_X1 U10933 ( .A(n10054), .B(n10662), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3358) );
  NOR2_X1 U10934 ( .A1(n10058), .A2(n10215), .ZN(n10061) );
  AOI22_X1 U10935 ( .A1(n10318), .A2(n10218), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10059) );
  OAI21_X1 U10936 ( .B1(n10221), .B2(n10281), .A(n10059), .ZN(n10060) );
  AOI211_X1 U10937 ( .C1(n10449), .C2(n10223), .A(n10061), .B(n10060), .ZN(
        n10062) );
  AND2_X1 U10938 ( .A1(n5702), .A2(n10063), .ZN(n10064) );
  NAND2_X1 U10939 ( .A1(n10065), .A2(n10064), .ZN(n10066) );
  XOR2_X1 U10940 ( .A(n10067), .B(n10066), .Z(n10076) );
  NOR2_X1 U10941 ( .A1(n10215), .A2(n10068), .ZN(n10069) );
  AOI211_X1 U10942 ( .C1(n10218), .C2(n10959), .A(n10070), .B(n10069), .ZN(
        n10071) );
  OAI21_X1 U10943 ( .B1(n10221), .B2(n10072), .A(n10071), .ZN(n10073) );
  AOI21_X1 U10944 ( .B1(n10074), .B2(n10223), .A(n10073), .ZN(n10075) );
  OAI21_X1 U10945 ( .B1(n10076), .B2(n10226), .A(n10075), .ZN(P1_U3213) );
  XNOR2_X1 U10946 ( .A(n10078), .B(n10077), .ZN(n10079) );
  XNOR2_X1 U10947 ( .A(n5089), .B(n10079), .ZN(n10085) );
  AOI22_X1 U10948 ( .A1(n10327), .A2(n10191), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10081) );
  NAND2_X1 U10949 ( .A1(n10203), .A2(n10331), .ZN(n10080) );
  OAI211_X1 U10950 ( .C1(n10082), .C2(n10126), .A(n10081), .B(n10080), .ZN(
        n10083) );
  AOI21_X1 U10951 ( .B1(n10469), .B2(n10223), .A(n10083), .ZN(n10084) );
  OAI21_X1 U10952 ( .B1(n10085), .B2(n10226), .A(n10084), .ZN(P1_U3214) );
  INV_X1 U10953 ( .A(n10086), .ZN(n10090) );
  AOI21_X1 U10954 ( .B1(n10087), .B2(n10187), .A(n10088), .ZN(n10089) );
  OAI21_X1 U10955 ( .B1(n10090), .B2(n10089), .A(n10197), .ZN(n10096) );
  NOR2_X1 U10956 ( .A1(n10091), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10264) );
  AOI21_X1 U10957 ( .B1(n10218), .B2(n10425), .A(n10264), .ZN(n10092) );
  OAI21_X1 U10958 ( .B1(n10093), .B2(n10215), .A(n10092), .ZN(n10094) );
  AOI21_X1 U10959 ( .B1(n10386), .B2(n10203), .A(n10094), .ZN(n10095) );
  OAI211_X1 U10960 ( .C1(n10388), .C2(n10206), .A(n10096), .B(n10095), .ZN(
        P1_U3217) );
  AOI21_X1 U10961 ( .B1(n10098), .B2(n10097), .A(n5102), .ZN(n10103) );
  AOI22_X1 U10962 ( .A1(n10356), .A2(n10191), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10100) );
  NAND2_X1 U10963 ( .A1(n10218), .A2(n10394), .ZN(n10099) );
  OAI211_X1 U10964 ( .C1(n10221), .C2(n10361), .A(n10100), .B(n10099), .ZN(
        n10101) );
  AOI21_X1 U10965 ( .B1(n10479), .B2(n10223), .A(n10101), .ZN(n10102) );
  OAI21_X1 U10966 ( .B1(n10103), .B2(n10226), .A(n10102), .ZN(P1_U3221) );
  XOR2_X1 U10967 ( .A(n10105), .B(n10104), .Z(n10111) );
  NOR2_X1 U10968 ( .A1(n10311), .A2(n10221), .ZN(n10109) );
  AOI22_X1 U10969 ( .A1(n10327), .A2(n10218), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10106) );
  OAI21_X1 U10970 ( .B1(n10107), .B2(n10215), .A(n10106), .ZN(n10108) );
  AOI211_X1 U10971 ( .C1(n10459), .C2(n10223), .A(n10109), .B(n10108), .ZN(
        n10110) );
  OAI21_X1 U10972 ( .B1(n10111), .B2(n10226), .A(n10110), .ZN(P1_U3223) );
  INV_X1 U10973 ( .A(n11061), .ZN(n11048) );
  OAI21_X1 U10974 ( .B1(n10114), .B2(n10112), .A(n10113), .ZN(n10115) );
  NAND2_X1 U10975 ( .A1(n10115), .A2(n10197), .ZN(n10120) );
  INV_X1 U10976 ( .A(n10116), .ZN(n11058) );
  AOI22_X1 U10977 ( .A1(n10218), .A2(n11039), .B1(P1_REG3_REG_16__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10117) );
  OAI21_X1 U10978 ( .B1(n10400), .B2(n10215), .A(n10117), .ZN(n10118) );
  AOI21_X1 U10979 ( .B1(n11058), .B2(n10203), .A(n10118), .ZN(n10119) );
  OAI211_X1 U10980 ( .C1(n11048), .C2(n10206), .A(n10120), .B(n10119), .ZN(
        P1_U3224) );
  XNOR2_X1 U10981 ( .A(n10123), .B(n10122), .ZN(n10124) );
  XNOR2_X1 U10982 ( .A(n10121), .B(n10124), .ZN(n10131) );
  OAI21_X1 U10983 ( .B1(n10126), .B2(n10214), .A(n10125), .ZN(n10127) );
  AOI21_X1 U10984 ( .B1(n10191), .B2(n10425), .A(n10127), .ZN(n10128) );
  OAI21_X1 U10985 ( .B1(n10221), .B2(n10432), .A(n10128), .ZN(n10129) );
  AOI21_X1 U10986 ( .B1(n10500), .B2(n10223), .A(n10129), .ZN(n10130) );
  OAI21_X1 U10987 ( .B1(n10131), .B2(n10226), .A(n10130), .ZN(P1_U3226) );
  XOR2_X1 U10988 ( .A(n10133), .B(n10132), .Z(n10139) );
  AOI22_X1 U10989 ( .A1(n10230), .A2(n10191), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10135) );
  NAND2_X1 U10990 ( .A1(n10346), .A2(n10218), .ZN(n10134) );
  OAI211_X1 U10991 ( .C1(n10221), .C2(n10136), .A(n10135), .B(n10134), .ZN(
        n10137) );
  AOI21_X1 U10992 ( .B1(n10464), .B2(n10223), .A(n10137), .ZN(n10138) );
  OAI21_X1 U10993 ( .B1(n10139), .B2(n10226), .A(n10138), .ZN(P1_U3227) );
  NAND2_X1 U10994 ( .A1(n5679), .A2(n10141), .ZN(n10142) );
  XNOR2_X1 U10995 ( .A(n10143), .B(n10142), .ZN(n10148) );
  AOI22_X1 U10996 ( .A1(n10218), .A2(n10376), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10145) );
  NAND2_X1 U10997 ( .A1(n10191), .A2(n10375), .ZN(n10144) );
  OAI211_X1 U10998 ( .C1(n10221), .C2(n10368), .A(n10145), .B(n10144), .ZN(
        n10146) );
  AOI21_X1 U10999 ( .B1(n10484), .B2(n10223), .A(n10146), .ZN(n10147) );
  OAI21_X1 U11000 ( .B1(n10148), .B2(n10226), .A(n10147), .ZN(P1_U3231) );
  INV_X1 U11001 ( .A(n10149), .ZN(n10154) );
  NAND2_X1 U11002 ( .A1(n5368), .A2(n10153), .ZN(n10151) );
  AOI22_X1 U11003 ( .A1(n10154), .A2(n10153), .B1(n10152), .B2(n10151), .ZN(
        n10163) );
  INV_X1 U11004 ( .A(n10155), .ZN(n10158) );
  NOR2_X1 U11005 ( .A1(n10215), .A2(n10156), .ZN(n10157) );
  AOI211_X1 U11006 ( .C1(n10218), .C2(n10232), .A(n10158), .B(n10157), .ZN(
        n10159) );
  OAI21_X1 U11007 ( .B1(n10221), .B2(n10160), .A(n10159), .ZN(n10161) );
  AOI21_X1 U11008 ( .B1(n10984), .B2(n10223), .A(n10161), .ZN(n10162) );
  OAI21_X1 U11009 ( .B1(n10163), .B2(n10226), .A(n10162), .ZN(P1_U3232) );
  AOI21_X1 U11010 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(n10173) );
  OAI22_X1 U11011 ( .A1(n10168), .A2(n10215), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10167), .ZN(n10169) );
  AOI21_X1 U11012 ( .B1(n10218), .B2(n10375), .A(n10169), .ZN(n10170) );
  OAI21_X1 U11013 ( .B1(n10221), .B2(n10339), .A(n10170), .ZN(n10171) );
  AOI21_X1 U11014 ( .B1(n10474), .B2(n10223), .A(n10171), .ZN(n10172) );
  OAI21_X1 U11015 ( .B1(n10173), .B2(n10226), .A(n10172), .ZN(P1_U3233) );
  OAI21_X1 U11016 ( .B1(n10176), .B2(n10175), .A(n10174), .ZN(n10177) );
  NAND2_X1 U11017 ( .A1(n10177), .A2(n10197), .ZN(n10182) );
  AOI22_X1 U11018 ( .A1(n10218), .A2(n10732), .B1(n10740), .B2(n10223), .ZN(
        n10181) );
  AOI22_X1 U11019 ( .A1(n10191), .A2(n10731), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10179), .ZN(n10180) );
  NAND3_X1 U11020 ( .A1(n10182), .A2(n10181), .A3(n10180), .ZN(P1_U3235) );
  XNOR2_X1 U11021 ( .A(n10184), .B(n10183), .ZN(n10186) );
  INV_X1 U11022 ( .A(n10188), .ZN(n10185) );
  NAND2_X1 U11023 ( .A1(n10186), .A2(n10185), .ZN(n10190) );
  INV_X1 U11024 ( .A(n10187), .ZN(n10189) );
  AOI22_X1 U11025 ( .A1(n10190), .A2(n10087), .B1(n10189), .B2(n10188), .ZN(
        n10196) );
  AOI22_X1 U11026 ( .A1(n10191), .A2(n10376), .B1(P1_REG3_REG_18__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10193) );
  NAND2_X1 U11027 ( .A1(n10218), .A2(n11038), .ZN(n10192) );
  OAI211_X1 U11028 ( .C1(n10221), .C2(n10411), .A(n10193), .B(n10192), .ZN(
        n10194) );
  AOI21_X1 U11029 ( .B1(n10494), .B2(n10223), .A(n10194), .ZN(n10195) );
  OAI21_X1 U11030 ( .B1(n10196), .B2(n10226), .A(n10195), .ZN(P1_U3236) );
  OAI211_X1 U11031 ( .C1(n10200), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        n10205) );
  AOI22_X1 U11032 ( .A1(n10230), .A2(n10218), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10201) );
  OAI21_X1 U11033 ( .B1(n10295), .B2(n10215), .A(n10201), .ZN(n10202) );
  AOI21_X1 U11034 ( .B1(n10300), .B2(n10203), .A(n10202), .ZN(n10204) );
  OAI211_X1 U11035 ( .C1(n10302), .C2(n10206), .A(n10205), .B(n10204), .ZN(
        P1_U3238) );
  INV_X1 U11036 ( .A(n10207), .ZN(n10209) );
  NAND2_X1 U11037 ( .A1(n10209), .A2(n10208), .ZN(n10211) );
  AOI22_X1 U11038 ( .A1(n10212), .A2(n10211), .B1(n10112), .B2(n10210), .ZN(
        n10227) );
  INV_X1 U11039 ( .A(n10213), .ZN(n10217) );
  NOR2_X1 U11040 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  AOI211_X1 U11041 ( .C1(n10218), .C2(n10231), .A(n10217), .B(n10216), .ZN(
        n10219) );
  OAI21_X1 U11042 ( .B1(n10221), .B2(n10220), .A(n10219), .ZN(n10222) );
  AOI21_X1 U11043 ( .B1(n10224), .B2(n10223), .A(n10222), .ZN(n10225) );
  OAI21_X1 U11044 ( .B1(n10227), .B2(n10226), .A(n10225), .ZN(P1_U3239) );
  MUX2_X1 U11045 ( .A(n10269), .B(P1_DATAO_REG_31__SCAN_IN), .S(n10236), .Z(
        P1_U3586) );
  MUX2_X1 U11046 ( .A(n10228), .B(P1_DATAO_REG_30__SCAN_IN), .S(n10236), .Z(
        P1_U3585) );
  MUX2_X1 U11047 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10288), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U11048 ( .A(n10229), .B(P1_DATAO_REG_27__SCAN_IN), .S(n10236), .Z(
        P1_U3582) );
  MUX2_X1 U11049 ( .A(n10318), .B(P1_DATAO_REG_26__SCAN_IN), .S(n10236), .Z(
        P1_U3581) );
  MUX2_X1 U11050 ( .A(n10230), .B(P1_DATAO_REG_25__SCAN_IN), .S(n10236), .Z(
        P1_U3580) );
  MUX2_X1 U11051 ( .A(n10327), .B(P1_DATAO_REG_24__SCAN_IN), .S(n10236), .Z(
        P1_U3579) );
  MUX2_X1 U11052 ( .A(n10346), .B(P1_DATAO_REG_23__SCAN_IN), .S(n10236), .Z(
        P1_U3578) );
  MUX2_X1 U11053 ( .A(n10356), .B(P1_DATAO_REG_22__SCAN_IN), .S(n10236), .Z(
        P1_U3577) );
  MUX2_X1 U11054 ( .A(n10375), .B(P1_DATAO_REG_21__SCAN_IN), .S(n10236), .Z(
        P1_U3576) );
  MUX2_X1 U11055 ( .A(n10394), .B(P1_DATAO_REG_20__SCAN_IN), .S(n10236), .Z(
        P1_U3575) );
  MUX2_X1 U11056 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10376), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U11057 ( .A(n10425), .B(P1_DATAO_REG_18__SCAN_IN), .S(n10236), .Z(
        P1_U3573) );
  MUX2_X1 U11058 ( .A(n11038), .B(P1_DATAO_REG_17__SCAN_IN), .S(n10236), .Z(
        P1_U3572) );
  MUX2_X1 U11059 ( .A(n10424), .B(P1_DATAO_REG_16__SCAN_IN), .S(n10236), .Z(
        P1_U3571) );
  MUX2_X1 U11060 ( .A(n11039), .B(P1_DATAO_REG_15__SCAN_IN), .S(n10236), .Z(
        P1_U3570) );
  MUX2_X1 U11061 ( .A(n10231), .B(P1_DATAO_REG_14__SCAN_IN), .S(n10236), .Z(
        P1_U3569) );
  MUX2_X1 U11062 ( .A(n10959), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10236), .Z(
        P1_U3568) );
  MUX2_X1 U11063 ( .A(n10232), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10236), .Z(
        P1_U3567) );
  MUX2_X1 U11064 ( .A(n10958), .B(P1_DATAO_REG_11__SCAN_IN), .S(n10236), .Z(
        P1_U3566) );
  MUX2_X1 U11065 ( .A(n10233), .B(P1_DATAO_REG_10__SCAN_IN), .S(n10236), .Z(
        P1_U3565) );
  MUX2_X1 U11066 ( .A(n10849), .B(P1_DATAO_REG_9__SCAN_IN), .S(n10236), .Z(
        P1_U3564) );
  MUX2_X1 U11067 ( .A(n10848), .B(P1_DATAO_REG_7__SCAN_IN), .S(n10236), .Z(
        P1_U3562) );
  MUX2_X1 U11068 ( .A(n10234), .B(P1_DATAO_REG_6__SCAN_IN), .S(n10236), .Z(
        P1_U3561) );
  MUX2_X1 U11069 ( .A(n10803), .B(P1_DATAO_REG_5__SCAN_IN), .S(n10236), .Z(
        P1_U3560) );
  MUX2_X1 U11070 ( .A(n10235), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10236), .Z(
        P1_U3559) );
  MUX2_X1 U11071 ( .A(n10731), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10236), .Z(
        P1_U3558) );
  MUX2_X1 U11072 ( .A(n10732), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10236), .Z(
        P1_U3556) );
  MUX2_X1 U11073 ( .A(n6803), .B(P1_DATAO_REG_0__SCAN_IN), .S(n10236), .Z(
        P1_U3555) );
  XNOR2_X1 U11074 ( .A(n10259), .B(n10237), .ZN(n10240) );
  AOI21_X1 U11075 ( .B1(n10246), .B2(P1_REG1_REG_17__SCAN_IN), .A(n10238), 
        .ZN(n10239) );
  NAND2_X1 U11076 ( .A1(n10239), .A2(n10240), .ZN(n10255) );
  OAI21_X1 U11077 ( .B1(n10240), .B2(n10239), .A(n10255), .ZN(n10253) );
  INV_X1 U11078 ( .A(n10259), .ZN(n10244) );
  NAND2_X1 U11079 ( .A1(n10696), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n10243) );
  NAND2_X1 U11080 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3084), .ZN(n10242)
         );
  OAI211_X1 U11081 ( .C1(n10692), .C2(n10244), .A(n10243), .B(n10242), .ZN(
        n10252) );
  AOI21_X1 U11082 ( .B1(n10246), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10245), 
        .ZN(n10250) );
  INV_X1 U11083 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10248) );
  NOR2_X1 U11084 ( .A1(n10259), .A2(n10248), .ZN(n10247) );
  AOI21_X1 U11085 ( .B1(n10259), .B2(n10248), .A(n10247), .ZN(n10249) );
  NOR2_X1 U11086 ( .A1(n10250), .A2(n10249), .ZN(n10258) );
  AOI211_X1 U11087 ( .C1(n10250), .C2(n10249), .A(n10258), .B(n10701), .ZN(
        n10251) );
  AOI211_X1 U11088 ( .C1(n10636), .C2(n10253), .A(n10252), .B(n10251), .ZN(
        n10254) );
  INV_X1 U11089 ( .A(n10254), .ZN(P1_U3259) );
  XNOR2_X1 U11090 ( .A(n10359), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10257) );
  OAI21_X1 U11091 ( .B1(n10259), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10255), 
        .ZN(n10256) );
  XNOR2_X1 U11092 ( .A(n10257), .B(n10256), .ZN(n10263) );
  MUX2_X1 U11093 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8138), .S(n10789), .Z(
        n10261) );
  AOI21_X1 U11094 ( .B1(n10259), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10258), 
        .ZN(n10260) );
  XNOR2_X1 U11095 ( .A(n10261), .B(n10260), .ZN(n10262) );
  AOI22_X1 U11096 ( .A1(n10636), .A2(n10263), .B1(n10640), .B2(n10262), .ZN(
        n10266) );
  AOI21_X1 U11097 ( .B1(n10605), .B2(n10789), .A(n10264), .ZN(n10265) );
  NAND2_X1 U11098 ( .A1(n10442), .A2(n10273), .ZN(n10272) );
  XNOR2_X1 U11099 ( .A(n10439), .B(n10272), .ZN(n10267) );
  NAND2_X1 U11100 ( .A1(n10267), .A2(n10953), .ZN(n10438) );
  NAND2_X1 U11101 ( .A1(n10269), .A2(n10268), .ZN(n10440) );
  NOR2_X1 U11102 ( .A1(n11070), .A2(n10440), .ZN(n10275) );
  NOR2_X1 U11103 ( .A1(n10439), .A2(n10430), .ZN(n10270) );
  AOI211_X1 U11104 ( .C1(n11070), .C2(P1_REG2_REG_31__SCAN_IN), .A(n10275), 
        .B(n10270), .ZN(n10271) );
  OAI21_X1 U11105 ( .B1(n11063), .B2(n10438), .A(n10271), .ZN(P1_U3261) );
  OAI211_X1 U11106 ( .C1(n10442), .C2(n10273), .A(n10953), .B(n10272), .ZN(
        n10441) );
  NOR2_X1 U11107 ( .A1(n10442), .A2(n10430), .ZN(n10274) );
  AOI211_X1 U11108 ( .C1(n11070), .C2(P1_REG2_REG_30__SCAN_IN), .A(n10275), 
        .B(n10274), .ZN(n10276) );
  OAI21_X1 U11109 ( .B1(n11063), .B2(n10441), .A(n10276), .ZN(P1_U3262) );
  XNOR2_X1 U11110 ( .A(n10278), .B(n10277), .ZN(n10452) );
  INV_X1 U11111 ( .A(n10279), .ZN(n10280) );
  AOI211_X1 U11112 ( .C1(n10449), .C2(n5382), .A(n11043), .B(n10280), .ZN(
        n10448) );
  INV_X1 U11113 ( .A(n10281), .ZN(n10282) );
  AOI22_X1 U11114 ( .A1(n10282), .A2(n11059), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n11070), .ZN(n10283) );
  OAI21_X1 U11115 ( .B1(n10284), .B2(n10430), .A(n10283), .ZN(n10290) );
  NAND2_X1 U11116 ( .A1(n10292), .A2(n10285), .ZN(n10287) );
  XNOR2_X1 U11117 ( .A(n10287), .B(n10286), .ZN(n10289) );
  OAI21_X1 U11118 ( .B1(n10296), .B2(n10293), .A(n10292), .ZN(n10298) );
  OAI22_X1 U11119 ( .A1(n10295), .A2(n10781), .B1(n10294), .B2(n10779), .ZN(
        n10297) );
  AOI211_X1 U11120 ( .C1(n10454), .C2(n10308), .A(n11043), .B(n10299), .ZN(
        n10453) );
  AOI22_X1 U11121 ( .A1(n10300), .A2(n11059), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n11070), .ZN(n10301) );
  OAI21_X1 U11122 ( .B1(n10302), .B2(n10430), .A(n10301), .ZN(n10304) );
  NOR2_X1 U11123 ( .A1(n10457), .A2(n10415), .ZN(n10303) );
  AOI211_X1 U11124 ( .C1(n10453), .C2(n10291), .A(n10304), .B(n10303), .ZN(
        n10305) );
  OAI21_X1 U11125 ( .B1(n10456), .B2(n11070), .A(n10305), .ZN(P1_U3265) );
  XNOR2_X1 U11126 ( .A(n10306), .B(n10317), .ZN(n10462) );
  INV_X1 U11127 ( .A(n10307), .ZN(n10310) );
  INV_X1 U11128 ( .A(n10308), .ZN(n10309) );
  AOI211_X1 U11129 ( .C1(n10459), .C2(n10310), .A(n11043), .B(n10309), .ZN(
        n10458) );
  INV_X1 U11130 ( .A(n10311), .ZN(n10312) );
  AOI22_X1 U11131 ( .A1(n10312), .A2(n11059), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n11070), .ZN(n10313) );
  OAI21_X1 U11132 ( .B1(n10314), .B2(n10430), .A(n10313), .ZN(n10321) );
  OAI21_X1 U11133 ( .B1(n10317), .B2(n10316), .A(n10315), .ZN(n10319) );
  AOI222_X1 U11134 ( .A1(n11035), .A2(n10319), .B1(n10318), .B2(n11037), .C1(
        n10327), .C2(n11040), .ZN(n10461) );
  NOR2_X1 U11135 ( .A1(n10461), .A2(n11070), .ZN(n10320) );
  AOI211_X1 U11136 ( .C1(n10458), .C2(n10291), .A(n10321), .B(n10320), .ZN(
        n10322) );
  OAI21_X1 U11137 ( .B1(n10462), .B2(n11064), .A(n10322), .ZN(P1_U3266) );
  XNOR2_X1 U11138 ( .A(n10323), .B(n10326), .ZN(n10472) );
  OAI21_X1 U11139 ( .B1(n10326), .B2(n10325), .A(n10324), .ZN(n10328) );
  AOI222_X1 U11140 ( .A1(n11035), .A2(n10328), .B1(n10327), .B2(n11037), .C1(
        n10356), .C2(n11040), .ZN(n10471) );
  INV_X1 U11141 ( .A(n10329), .ZN(n10330) );
  AOI211_X1 U11142 ( .C1(n10469), .C2(n10337), .A(n11043), .B(n10330), .ZN(
        n10468) );
  AOI22_X1 U11143 ( .A1(n10468), .A2(n10359), .B1(n11059), .B2(n10331), .ZN(
        n10332) );
  AOI21_X1 U11144 ( .B1(n10471), .B2(n10332), .A(n11070), .ZN(n10333) );
  INV_X1 U11145 ( .A(n10333), .ZN(n10335) );
  AOI22_X1 U11146 ( .A1(n10469), .A2(n11060), .B1(n11070), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n10334) );
  OAI211_X1 U11147 ( .C1(n10472), .C2(n11064), .A(n10335), .B(n10334), .ZN(
        P1_U3268) );
  XOR2_X1 U11148 ( .A(n10345), .B(n10336), .Z(n10477) );
  INV_X1 U11149 ( .A(n10337), .ZN(n10338) );
  AOI211_X1 U11150 ( .C1(n10474), .C2(n5388), .A(n11043), .B(n10338), .ZN(
        n10473) );
  INV_X1 U11151 ( .A(n10339), .ZN(n10340) );
  AOI22_X1 U11152 ( .A1(n11070), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10340), 
        .B2(n11059), .ZN(n10341) );
  OAI21_X1 U11153 ( .B1(n10342), .B2(n10430), .A(n10341), .ZN(n10349) );
  OAI21_X1 U11154 ( .B1(n10345), .B2(n10344), .A(n10343), .ZN(n10347) );
  AOI222_X1 U11155 ( .A1(n11035), .A2(n10347), .B1(n10346), .B2(n11037), .C1(
        n10375), .C2(n11040), .ZN(n10476) );
  NOR2_X1 U11156 ( .A1(n10476), .A2(n11070), .ZN(n10348) );
  AOI211_X1 U11157 ( .C1(n10473), .C2(n10291), .A(n10349), .B(n10348), .ZN(
        n10350) );
  OAI21_X1 U11158 ( .B1(n11064), .B2(n10477), .A(n10350), .ZN(P1_U3269) );
  OAI21_X1 U11159 ( .B1(n5097), .B2(n10352), .A(n10351), .ZN(n10482) );
  AOI22_X1 U11160 ( .A1(n10479), .A2(n11060), .B1(n11070), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n10364) );
  OAI21_X1 U11161 ( .B1(n10355), .B2(n10354), .A(n10353), .ZN(n10357) );
  AOI222_X1 U11162 ( .A1(n11035), .A2(n10357), .B1(n10356), .B2(n11037), .C1(
        n10394), .C2(n11040), .ZN(n10481) );
  AOI211_X1 U11163 ( .C1(n10479), .C2(n10366), .A(n11043), .B(n10358), .ZN(
        n10478) );
  NAND2_X1 U11164 ( .A1(n10478), .A2(n10359), .ZN(n10360) );
  OAI211_X1 U11165 ( .C1(n10786), .C2(n10361), .A(n10481), .B(n10360), .ZN(
        n10362) );
  NAND2_X1 U11166 ( .A1(n10362), .A2(n10795), .ZN(n10363) );
  OAI211_X1 U11167 ( .C1(n10482), .C2(n11064), .A(n10364), .B(n10363), .ZN(
        P1_U3270) );
  XOR2_X1 U11168 ( .A(n10365), .B(n10373), .Z(n10487) );
  INV_X1 U11169 ( .A(n10366), .ZN(n10367) );
  AOI211_X1 U11170 ( .C1(n10484), .C2(n10383), .A(n11043), .B(n10367), .ZN(
        n10483) );
  INV_X1 U11171 ( .A(n10484), .ZN(n10371) );
  INV_X1 U11172 ( .A(n10368), .ZN(n10369) );
  AOI22_X1 U11173 ( .A1(n11070), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10369), 
        .B2(n11059), .ZN(n10370) );
  OAI21_X1 U11174 ( .B1(n10371), .B2(n10430), .A(n10370), .ZN(n10379) );
  OAI21_X1 U11175 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(n10377) );
  AOI222_X1 U11176 ( .A1(n11035), .A2(n10377), .B1(n10376), .B2(n11040), .C1(
        n10375), .C2(n11037), .ZN(n10486) );
  NOR2_X1 U11177 ( .A1(n10486), .A2(n11070), .ZN(n10378) );
  AOI211_X1 U11178 ( .C1(n10483), .C2(n10291), .A(n10379), .B(n10378), .ZN(
        n10380) );
  OAI21_X1 U11179 ( .B1(n10487), .B2(n11064), .A(n10380), .ZN(P1_U3271) );
  XNOR2_X1 U11180 ( .A(n10382), .B(n10381), .ZN(n10492) );
  INV_X1 U11181 ( .A(n10409), .ZN(n10385) );
  INV_X1 U11182 ( .A(n10383), .ZN(n10384) );
  AOI211_X1 U11183 ( .C1(n10489), .C2(n10385), .A(n11043), .B(n10384), .ZN(
        n10488) );
  AOI22_X1 U11184 ( .A1(n11070), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10386), 
        .B2(n11059), .ZN(n10387) );
  OAI21_X1 U11185 ( .B1(n10388), .B2(n10430), .A(n10387), .ZN(n10397) );
  AND2_X1 U11186 ( .A1(n10390), .A2(n10389), .ZN(n10393) );
  OAI21_X1 U11187 ( .B1(n10393), .B2(n10392), .A(n10391), .ZN(n10395) );
  AOI222_X1 U11188 ( .A1(n11035), .A2(n10395), .B1(n10425), .B2(n11040), .C1(
        n10394), .C2(n11037), .ZN(n10491) );
  NOR2_X1 U11189 ( .A1(n10491), .A2(n11070), .ZN(n10396) );
  AOI211_X1 U11190 ( .C1(n10488), .C2(n10291), .A(n10397), .B(n10396), .ZN(
        n10398) );
  OAI21_X1 U11191 ( .B1(n11064), .B2(n10492), .A(n10398), .ZN(P1_U3272) );
  XNOR2_X1 U11192 ( .A(n10399), .B(n5273), .ZN(n10408) );
  OAI22_X1 U11193 ( .A1(n10401), .A2(n10781), .B1(n10400), .B2(n10779), .ZN(
        n10407) );
  NAND2_X1 U11194 ( .A1(n10403), .A2(n10402), .ZN(n10404) );
  NAND2_X1 U11195 ( .A1(n10405), .A2(n10404), .ZN(n10497) );
  NOR2_X1 U11196 ( .A1(n10497), .A2(n10851), .ZN(n10406) );
  AOI211_X1 U11197 ( .C1(n11035), .C2(n10408), .A(n10407), .B(n10406), .ZN(
        n10496) );
  INV_X1 U11198 ( .A(n10429), .ZN(n10410) );
  AOI211_X1 U11199 ( .C1(n10494), .C2(n10410), .A(n11043), .B(n10409), .ZN(
        n10493) );
  INV_X1 U11200 ( .A(n10411), .ZN(n10412) );
  AOI22_X1 U11201 ( .A1(n11070), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10412), 
        .B2(n11059), .ZN(n10413) );
  OAI21_X1 U11202 ( .B1(n10414), .B2(n10430), .A(n10413), .ZN(n10417) );
  NOR2_X1 U11203 ( .A1(n10497), .A2(n10415), .ZN(n10416) );
  AOI211_X1 U11204 ( .C1(n10493), .C2(n10291), .A(n10417), .B(n10416), .ZN(
        n10418) );
  OAI21_X1 U11205 ( .B1(n10496), .B2(n11070), .A(n10418), .ZN(P1_U3273) );
  OAI21_X1 U11206 ( .B1(n10421), .B2(n10420), .A(n10419), .ZN(n10498) );
  XNOR2_X1 U11207 ( .A(n10423), .B(n10422), .ZN(n10427) );
  AOI22_X1 U11208 ( .A1(n11037), .A2(n10425), .B1(n10424), .B2(n11040), .ZN(
        n10426) );
  OAI21_X1 U11209 ( .B1(n10427), .B2(n10777), .A(n10426), .ZN(n10428) );
  AOI21_X1 U11210 ( .B1(n10498), .B2(n10913), .A(n10428), .ZN(n10502) );
  AOI211_X1 U11211 ( .C1(n10500), .C2(n11045), .A(n11043), .B(n10429), .ZN(
        n10499) );
  INV_X1 U11212 ( .A(n10500), .ZN(n10431) );
  NOR2_X1 U11213 ( .A1(n10431), .A2(n10430), .ZN(n10435) );
  OAI22_X1 U11214 ( .A1(n10795), .A2(n10433), .B1(n10432), .B2(n10786), .ZN(
        n10434) );
  AOI211_X1 U11215 ( .C1(n10499), .C2(n10291), .A(n10435), .B(n10434), .ZN(
        n10437) );
  NAND2_X1 U11216 ( .A1(n10498), .A2(n10863), .ZN(n10436) );
  OAI211_X1 U11217 ( .C1(n10502), .C2(n11070), .A(n10437), .B(n10436), .ZN(
        P1_U3274) );
  OAI211_X1 U11218 ( .C1(n10439), .C2(n11047), .A(n10438), .B(n10440), .ZN(
        n10504) );
  MUX2_X1 U11219 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10504), .S(n11054), .Z(
        P1_U3554) );
  OAI211_X1 U11220 ( .C1(n10442), .C2(n11047), .A(n10441), .B(n10440), .ZN(
        n10505) );
  MUX2_X1 U11221 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10505), .S(n11054), .Z(
        P1_U3553) );
  AOI21_X1 U11222 ( .B1(n10908), .B2(n10444), .A(n10443), .ZN(n10445) );
  OAI211_X1 U11223 ( .C1(n10447), .C2(n10769), .A(n10446), .B(n10445), .ZN(
        n10506) );
  MUX2_X1 U11224 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10506), .S(n11054), .Z(
        P1_U3552) );
  AOI21_X1 U11225 ( .B1(n10908), .B2(n10449), .A(n10448), .ZN(n10450) );
  OAI211_X1 U11226 ( .C1(n10452), .C2(n10769), .A(n10451), .B(n10450), .ZN(
        n10510) );
  MUX2_X1 U11227 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10510), .S(n11054), .Z(
        P1_U3550) );
  AOI21_X1 U11228 ( .B1(n10908), .B2(n10454), .A(n10453), .ZN(n10455) );
  OAI211_X1 U11229 ( .C1(n10457), .C2(n10911), .A(n10456), .B(n10455), .ZN(
        n10511) );
  MUX2_X1 U11230 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10511), .S(n11054), .Z(
        P1_U3549) );
  AOI21_X1 U11231 ( .B1(n10908), .B2(n10459), .A(n10458), .ZN(n10460) );
  OAI211_X1 U11232 ( .C1(n10462), .C2(n10769), .A(n10461), .B(n10460), .ZN(
        n10512) );
  MUX2_X1 U11233 ( .A(n10512), .B(P1_REG1_REG_25__SCAN_IN), .S(n11052), .Z(
        P1_U3548) );
  AOI21_X1 U11234 ( .B1(n10908), .B2(n10464), .A(n10463), .ZN(n10465) );
  OAI211_X1 U11235 ( .C1(n10467), .C2(n10769), .A(n10466), .B(n10465), .ZN(
        n10513) );
  MUX2_X1 U11236 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10513), .S(n11054), .Z(
        P1_U3547) );
  AOI21_X1 U11237 ( .B1(n10908), .B2(n10469), .A(n10468), .ZN(n10470) );
  OAI211_X1 U11238 ( .C1(n10472), .C2(n10769), .A(n10471), .B(n10470), .ZN(
        n10514) );
  MUX2_X1 U11239 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10514), .S(n11054), .Z(
        P1_U3546) );
  AOI21_X1 U11240 ( .B1(n10908), .B2(n10474), .A(n10473), .ZN(n10475) );
  OAI211_X1 U11241 ( .C1(n10477), .C2(n10769), .A(n10476), .B(n10475), .ZN(
        n10515) );
  MUX2_X1 U11242 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10515), .S(n11054), .Z(
        P1_U3545) );
  AOI21_X1 U11243 ( .B1(n10908), .B2(n10479), .A(n10478), .ZN(n10480) );
  OAI211_X1 U11244 ( .C1(n10482), .C2(n10769), .A(n10481), .B(n10480), .ZN(
        n10516) );
  MUX2_X1 U11245 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10516), .S(n11054), .Z(
        P1_U3544) );
  AOI21_X1 U11246 ( .B1(n10908), .B2(n10484), .A(n10483), .ZN(n10485) );
  OAI211_X1 U11247 ( .C1(n10487), .C2(n10769), .A(n10486), .B(n10485), .ZN(
        n10517) );
  MUX2_X1 U11248 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10517), .S(n11054), .Z(
        P1_U3543) );
  AOI21_X1 U11249 ( .B1(n10908), .B2(n10489), .A(n10488), .ZN(n10490) );
  OAI211_X1 U11250 ( .C1(n10492), .C2(n10769), .A(n10491), .B(n10490), .ZN(
        n10518) );
  MUX2_X1 U11251 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10518), .S(n11054), .Z(
        P1_U3542) );
  AOI21_X1 U11252 ( .B1(n10908), .B2(n10494), .A(n10493), .ZN(n10495) );
  OAI211_X1 U11253 ( .C1(n10911), .C2(n10497), .A(n10496), .B(n10495), .ZN(
        n10519) );
  MUX2_X1 U11254 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10519), .S(n11054), .Z(
        P1_U3541) );
  INV_X1 U11255 ( .A(n10498), .ZN(n10503) );
  AOI21_X1 U11256 ( .B1(n10908), .B2(n10500), .A(n10499), .ZN(n10501) );
  OAI211_X1 U11257 ( .C1(n10503), .C2(n10911), .A(n10502), .B(n10501), .ZN(
        n10520) );
  MUX2_X1 U11258 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10520), .S(n11054), .Z(
        P1_U3540) );
  MUX2_X1 U11259 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10504), .S(n11057), .Z(
        P1_U3522) );
  MUX2_X1 U11260 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10505), .S(n11057), .Z(
        P1_U3521) );
  MUX2_X1 U11261 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10506), .S(n11057), .Z(
        P1_U3520) );
  INV_X1 U11262 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10508) );
  MUX2_X1 U11263 ( .A(n10508), .B(n10507), .S(n11057), .Z(n10509) );
  INV_X1 U11264 ( .A(n10509), .ZN(P1_U3519) );
  MUX2_X1 U11265 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10510), .S(n11057), .Z(
        P1_U3518) );
  MUX2_X1 U11266 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10511), .S(n11057), .Z(
        P1_U3517) );
  MUX2_X1 U11267 ( .A(n10512), .B(P1_REG0_REG_25__SCAN_IN), .S(n11055), .Z(
        P1_U3516) );
  MUX2_X1 U11268 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10513), .S(n11057), .Z(
        P1_U3515) );
  MUX2_X1 U11269 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10514), .S(n11057), .Z(
        P1_U3514) );
  MUX2_X1 U11270 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10515), .S(n11057), .Z(
        P1_U3513) );
  MUX2_X1 U11271 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10516), .S(n11057), .Z(
        P1_U3512) );
  MUX2_X1 U11272 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10517), .S(n11057), .Z(
        P1_U3511) );
  MUX2_X1 U11273 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10518), .S(n11057), .Z(
        P1_U3510) );
  MUX2_X1 U11274 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10519), .S(n11057), .Z(
        P1_U3508) );
  MUX2_X1 U11275 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10520), .S(n11057), .Z(
        P1_U3505) );
  MUX2_X1 U11276 ( .A(n10522), .B(P1_D_REG_1__SCAN_IN), .S(n10521), .Z(
        P1_U3441) );
  NOR4_X1 U11277 ( .A1(n10523), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n6374), .ZN(n10524) );
  AOI21_X1 U11278 ( .B1(n10525), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10524), 
        .ZN(n10526) );
  OAI21_X1 U11279 ( .B1(n10527), .B2(n10532), .A(n10526), .ZN(P1_U3322) );
  INV_X1 U11280 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10529) );
  OAI222_X1 U11281 ( .A1(n10532), .A2(n10531), .B1(n10530), .B2(P1_U3084), 
        .C1(n10529), .C2(n10528), .ZN(P1_U3323) );
  INV_X1 U11282 ( .A(n10533), .ZN(n10534) );
  MUX2_X1 U11283 ( .A(n10534), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11284 ( .A1(n10538), .A2(n10535), .ZN(P1_U3321) );
  NOR2_X1 U11285 ( .A1(n10538), .A2(n10536), .ZN(P1_U3320) );
  NOR2_X1 U11286 ( .A1(n10538), .A2(n10537), .ZN(P1_U3319) );
  AND2_X1 U11287 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10539), .ZN(P1_U3318) );
  AND2_X1 U11288 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10539), .ZN(P1_U3317) );
  AND2_X1 U11289 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10539), .ZN(P1_U3316) );
  AND2_X1 U11290 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10539), .ZN(P1_U3315) );
  AND2_X1 U11291 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10539), .ZN(P1_U3314) );
  AND2_X1 U11292 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10539), .ZN(P1_U3313) );
  AND2_X1 U11293 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10539), .ZN(P1_U3312) );
  AND2_X1 U11294 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10539), .ZN(P1_U3311) );
  AND2_X1 U11295 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10539), .ZN(P1_U3310) );
  AND2_X1 U11296 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10539), .ZN(P1_U3309) );
  AND2_X1 U11297 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10539), .ZN(P1_U3308) );
  AND2_X1 U11298 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10539), .ZN(P1_U3307) );
  AND2_X1 U11299 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10539), .ZN(P1_U3306) );
  AND2_X1 U11300 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10539), .ZN(P1_U3305) );
  AND2_X1 U11301 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10539), .ZN(P1_U3304) );
  AND2_X1 U11302 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10539), .ZN(P1_U3303) );
  AND2_X1 U11303 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10539), .ZN(P1_U3302) );
  AND2_X1 U11304 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10539), .ZN(P1_U3301) );
  AND2_X1 U11305 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10539), .ZN(P1_U3300) );
  AND2_X1 U11306 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10539), .ZN(P1_U3299) );
  AND2_X1 U11307 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10539), .ZN(P1_U3298) );
  AND2_X1 U11308 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10539), .ZN(P1_U3297) );
  AND2_X1 U11309 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10539), .ZN(P1_U3296) );
  AND2_X1 U11310 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10539), .ZN(P1_U3295) );
  AND2_X1 U11311 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10539), .ZN(P1_U3294) );
  AND2_X1 U11312 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10539), .ZN(P1_U3293) );
  AND2_X1 U11313 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10539), .ZN(P1_U3292) );
  NOR2_X1 U11314 ( .A1(n10541), .A2(n10540), .ZN(n10545) );
  INV_X1 U11315 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10544) );
  AOI22_X1 U11316 ( .A1(n10649), .A2(n10545), .B1(n10544), .B2(n10646), .ZN(
        P2_U3438) );
  AND2_X1 U11317 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10646), .ZN(P2_U3326) );
  AND2_X1 U11318 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10646), .ZN(P2_U3325) );
  AND2_X1 U11319 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10646), .ZN(P2_U3324) );
  AND2_X1 U11320 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10646), .ZN(P2_U3323) );
  AND2_X1 U11321 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10646), .ZN(P2_U3322) );
  AND2_X1 U11322 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10646), .ZN(P2_U3321) );
  AND2_X1 U11323 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10646), .ZN(P2_U3320) );
  AND2_X1 U11324 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10646), .ZN(P2_U3319) );
  AND2_X1 U11325 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10646), .ZN(P2_U3318) );
  AND2_X1 U11326 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10646), .ZN(P2_U3317) );
  AND2_X1 U11327 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10646), .ZN(P2_U3316) );
  AND2_X1 U11328 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10646), .ZN(P2_U3315) );
  AND2_X1 U11329 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10646), .ZN(P2_U3314) );
  AND2_X1 U11330 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10646), .ZN(P2_U3313) );
  AND2_X1 U11331 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10646), .ZN(P2_U3312) );
  AND2_X1 U11332 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10646), .ZN(P2_U3311) );
  AND2_X1 U11333 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10646), .ZN(P2_U3310) );
  AND2_X1 U11334 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10646), .ZN(P2_U3309) );
  AND2_X1 U11335 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10646), .ZN(P2_U3308) );
  AND2_X1 U11336 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10646), .ZN(P2_U3307) );
  AND2_X1 U11337 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10646), .ZN(P2_U3306) );
  AND2_X1 U11338 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10646), .ZN(P2_U3305) );
  AND2_X1 U11339 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10646), .ZN(P2_U3304) );
  AND2_X1 U11340 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10646), .ZN(P2_U3303) );
  AND2_X1 U11341 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10646), .ZN(P2_U3302) );
  AND2_X1 U11342 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10646), .ZN(P2_U3301) );
  AND2_X1 U11343 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10646), .ZN(P2_U3300) );
  AND2_X1 U11344 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10646), .ZN(P2_U3299) );
  AND2_X1 U11345 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10646), .ZN(P2_U3298) );
  AND2_X1 U11346 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10646), .ZN(P2_U3297) );
  XOR2_X1 U11347 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11348 ( .A(n10546), .ZN(n10547) );
  NAND2_X1 U11349 ( .A1(n10548), .A2(n10547), .ZN(n10549) );
  XNOR2_X1 U11350 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10549), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11351 ( .A(n10551), .B(n10550), .Z(ADD_1071_U54) );
  XOR2_X1 U11352 ( .A(n10553), .B(n10552), .Z(ADD_1071_U53) );
  XNOR2_X1 U11353 ( .A(n10555), .B(n10554), .ZN(ADD_1071_U52) );
  NOR2_X1 U11354 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  XOR2_X1 U11355 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10558), .Z(ADD_1071_U51) );
  XOR2_X1 U11356 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10559), .Z(ADD_1071_U50) );
  XOR2_X1 U11357 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10560), .Z(ADD_1071_U49) );
  XOR2_X1 U11358 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10561), .Z(ADD_1071_U48) );
  XOR2_X1 U11359 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10562), .Z(ADD_1071_U47) );
  XOR2_X1 U11360 ( .A(n10564), .B(n10563), .Z(ADD_1071_U63) );
  XOR2_X1 U11361 ( .A(n10566), .B(n10565), .Z(ADD_1071_U62) );
  XNOR2_X1 U11362 ( .A(n10568), .B(n10567), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11363 ( .A(n10570), .B(n10569), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11364 ( .A(n10572), .B(n10571), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11365 ( .A(n10574), .B(n10573), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11366 ( .A(n10576), .B(n10575), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11367 ( .A(n10578), .B(n10577), .ZN(ADD_1071_U56) );
  NOR2_X1 U11368 ( .A1(n10580), .A2(n10579), .ZN(n10581) );
  XOR2_X1 U11369 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10581), .Z(ADD_1071_U55)
         );
  OAI21_X1 U11370 ( .B1(n10583), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10582), .ZN(
        n10585) );
  XNOR2_X1 U11371 ( .A(n10585), .B(n10584), .ZN(n10588) );
  AOI22_X1 U11372 ( .A1(n10696), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10586) );
  OAI21_X1 U11373 ( .B1(n10588), .B2(n10587), .A(n10586), .ZN(P1_U3241) );
  INV_X1 U11374 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10589) );
  OR2_X1 U11375 ( .A1(n10618), .A2(n10589), .ZN(n10592) );
  INV_X1 U11376 ( .A(n10590), .ZN(n10591) );
  OAI211_X1 U11377 ( .C1(n10692), .C2(n10593), .A(n10592), .B(n10591), .ZN(
        n10594) );
  INV_X1 U11378 ( .A(n10594), .ZN(n10603) );
  OAI211_X1 U11379 ( .C1(n10597), .C2(n10596), .A(n10640), .B(n10595), .ZN(
        n10602) );
  OAI211_X1 U11380 ( .C1(n10600), .C2(n10599), .A(n10636), .B(n10598), .ZN(
        n10601) );
  NAND3_X1 U11381 ( .A1(n10603), .A2(n10602), .A3(n10601), .ZN(P1_U3247) );
  AOI22_X1 U11382 ( .A1(n10696), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n10605), 
        .B2(n10604), .ZN(n10616) );
  AOI21_X1 U11383 ( .B1(n10608), .B2(n10607), .A(n10606), .ZN(n10609) );
  OR2_X1 U11384 ( .A1(n10609), .A2(n10693), .ZN(n10614) );
  OAI211_X1 U11385 ( .C1(n10612), .C2(n10611), .A(n10640), .B(n10610), .ZN(
        n10613) );
  NAND4_X1 U11386 ( .A1(n10616), .A2(n10615), .A3(n10614), .A4(n10613), .ZN(
        P1_U3250) );
  INV_X1 U11387 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10617) );
  OR2_X1 U11388 ( .A1(n10618), .A2(n10617), .ZN(n10621) );
  INV_X1 U11389 ( .A(n10619), .ZN(n10620) );
  OAI211_X1 U11390 ( .C1(n10692), .C2(n10622), .A(n10621), .B(n10620), .ZN(
        n10623) );
  INV_X1 U11391 ( .A(n10623), .ZN(n10632) );
  OAI211_X1 U11392 ( .C1(n10626), .C2(n10625), .A(n10640), .B(n10624), .ZN(
        n10631) );
  OAI211_X1 U11393 ( .C1(n10629), .C2(n10628), .A(n10636), .B(n10627), .ZN(
        n10630) );
  NAND3_X1 U11394 ( .A1(n10632), .A2(n10631), .A3(n10630), .ZN(P1_U3244) );
  OAI22_X1 U11395 ( .A1(n10692), .A2(n5491), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10633), .ZN(n10634) );
  AOI21_X1 U11396 ( .B1(n10696), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n10634), .ZN(
        n10645) );
  OAI211_X1 U11397 ( .C1(n10638), .C2(n10637), .A(n10636), .B(n10635), .ZN(
        n10644) );
  OAI211_X1 U11398 ( .C1(n10642), .C2(n10641), .A(n10640), .B(n10639), .ZN(
        n10643) );
  NAND3_X1 U11399 ( .A1(n10645), .A2(n10644), .A3(n10643), .ZN(P1_U3242) );
  INV_X1 U11400 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U11401 ( .A1(n10649), .A2(n10648), .B1(n10647), .B2(n10646), .ZN(
        P2_U3437) );
  NAND2_X1 U11402 ( .A1(n10651), .A2(n10650), .ZN(n10654) );
  INV_X1 U11403 ( .A(n10652), .ZN(n10653) );
  NAND2_X1 U11404 ( .A1(n10654), .A2(n10653), .ZN(n10657) );
  NAND2_X1 U11405 ( .A1(P2_U3152), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n10656) );
  NAND2_X1 U11406 ( .A1(n10674), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10655) );
  OAI211_X1 U11407 ( .C1(n10658), .C2(n10657), .A(n10656), .B(n10655), .ZN(
        n10659) );
  AOI21_X1 U11408 ( .B1(n10661), .B2(n10660), .A(n10659), .ZN(n10667) );
  NOR2_X1 U11409 ( .A1(n5253), .A2(n6891), .ZN(n10665) );
  OAI211_X1 U11410 ( .C1(n10665), .C2(n10664), .A(n10679), .B(n10663), .ZN(
        n10666) );
  NAND2_X1 U11411 ( .A1(n10667), .A2(n10666), .ZN(P2_U3246) );
  INV_X1 U11412 ( .A(n10668), .ZN(n10673) );
  NAND3_X1 U11413 ( .A1(n10669), .A2(n10679), .A3(P2_REG2_REG_13__SCAN_IN), 
        .ZN(n10671) );
  AOI21_X1 U11414 ( .B1(n10671), .B2(n10670), .A(n10676), .ZN(n10672) );
  AOI211_X1 U11415 ( .C1(n10674), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n10673), 
        .B(n10672), .ZN(n10687) );
  NAND3_X1 U11416 ( .A1(n10677), .A2(n10676), .A3(n10675), .ZN(n10678) );
  NAND3_X1 U11417 ( .A1(n10680), .A2(n10679), .A3(n10678), .ZN(n10686) );
  OAI211_X1 U11418 ( .C1(n10684), .C2(n10683), .A(n10682), .B(n10681), .ZN(
        n10685) );
  NAND3_X1 U11419 ( .A1(n10687), .A2(n10686), .A3(n10685), .ZN(P2_U3258) );
  XNOR2_X1 U11420 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11421 ( .B1(n10690), .B2(n10689), .A(n10688), .ZN(n10694) );
  OAI22_X1 U11422 ( .A1(n10694), .A2(n10693), .B1(n10692), .B2(n10691), .ZN(
        n10695) );
  AOI21_X1 U11423 ( .B1(n10696), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n10695), .ZN(
        n10705) );
  AOI21_X1 U11424 ( .B1(n10699), .B2(n10698), .A(n10697), .ZN(n10700) );
  OR2_X1 U11425 ( .A1(n10701), .A2(n10700), .ZN(n10702) );
  NAND4_X1 U11426 ( .A1(n10705), .A2(n10704), .A3(n10703), .A4(n10702), .ZN(
        P1_U3245) );
  INV_X1 U11427 ( .A(n10706), .ZN(n10710) );
  AOI21_X1 U11428 ( .B1(n10789), .B2(n10708), .A(n10707), .ZN(n10709) );
  NOR2_X1 U11429 ( .A1(n10710), .A2(n10709), .ZN(n10712) );
  AOI22_X1 U11430 ( .A1(n11059), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n11070), .ZN(n10711) );
  OAI21_X1 U11431 ( .B1(n11070), .B2(n10712), .A(n10711), .ZN(P1_U3291) );
  AOI211_X1 U11432 ( .C1(n11015), .C2(n10715), .A(n5147), .B(n10714), .ZN(
        n10717) );
  INV_X1 U11433 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U11434 ( .A1(n11018), .A2(n10717), .B1(n10716), .B2(n11017), .ZN(
        P2_U3520) );
  AOI22_X1 U11435 ( .A1(n11001), .A2(n10717), .B1(n5825), .B2(n11019), .ZN(
        P2_U3451) );
  OAI211_X1 U11436 ( .C1(n10720), .C2(n11047), .A(n10719), .B(n10718), .ZN(
        n10723) );
  AOI21_X1 U11437 ( .B1(n10851), .B2(n10911), .A(n10721), .ZN(n10722) );
  NOR2_X1 U11438 ( .A1(n10723), .A2(n10722), .ZN(n10724) );
  AOI22_X1 U11439 ( .A1(n11054), .A2(n10724), .B1(n6467), .B2(n11052), .ZN(
        P1_U3524) );
  AOI22_X1 U11440 ( .A1(n11057), .A2(n10724), .B1(n6468), .B2(n11055), .ZN(
        P1_U3457) );
  INV_X1 U11441 ( .A(n10911), .ZN(n11028) );
  XNOR2_X1 U11442 ( .A(n10725), .B(n10729), .ZN(n10743) );
  OAI211_X1 U11443 ( .C1(n5373), .C2(n10728), .A(n10953), .B(n10727), .ZN(
        n10741) );
  OAI21_X1 U11444 ( .B1(n10728), .B2(n11047), .A(n10741), .ZN(n10737) );
  XNOR2_X1 U11445 ( .A(n10730), .B(n10729), .ZN(n10734) );
  AOI22_X1 U11446 ( .A1(n11040), .A2(n10732), .B1(n10731), .B2(n11037), .ZN(
        n10733) );
  OAI21_X1 U11447 ( .B1(n10734), .B2(n10777), .A(n10733), .ZN(n10735) );
  AOI21_X1 U11448 ( .B1(n10913), .B2(n10743), .A(n10735), .ZN(n10746) );
  INV_X1 U11449 ( .A(n10746), .ZN(n10736) );
  AOI211_X1 U11450 ( .C1(n11028), .C2(n10743), .A(n10737), .B(n10736), .ZN(
        n10739) );
  AOI22_X1 U11451 ( .A1(n11054), .A2(n10739), .B1(n10738), .B2(n11052), .ZN(
        P1_U3525) );
  AOI22_X1 U11452 ( .A1(n11057), .A2(n10739), .B1(n6204), .B2(n11055), .ZN(
        P1_U3460) );
  AOI222_X1 U11453 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n11070), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n11059), .C1(n10740), .C2(n11060), .ZN(
        n10745) );
  INV_X1 U11454 ( .A(n10741), .ZN(n10742) );
  AOI22_X1 U11455 ( .A1(n10743), .A2(n10863), .B1(n10291), .B2(n10742), .ZN(
        n10744) );
  OAI211_X1 U11456 ( .C1(n11070), .C2(n10746), .A(n10745), .B(n10744), .ZN(
        P1_U3289) );
  OAI211_X1 U11457 ( .C1(n10749), .C2(n11047), .A(n10748), .B(n10747), .ZN(
        n10752) );
  AOI21_X1 U11458 ( .B1(n10851), .B2(n10911), .A(n10750), .ZN(n10751) );
  NOR2_X1 U11459 ( .A1(n10752), .A2(n10751), .ZN(n10753) );
  AOI22_X1 U11460 ( .A1(n11054), .A2(n10753), .B1(n6231), .B2(n11052), .ZN(
        P1_U3526) );
  AOI22_X1 U11461 ( .A1(n11057), .A2(n10753), .B1(n6570), .B2(n11055), .ZN(
        P1_U3463) );
  OAI22_X1 U11462 ( .A1(n10755), .A2(n11011), .B1(n10754), .B2(n11010), .ZN(
        n10757) );
  AOI211_X1 U11463 ( .C1(n10884), .C2(n10758), .A(n10757), .B(n10756), .ZN(
        n10759) );
  AOI22_X1 U11464 ( .A1(n11018), .A2(n10759), .B1(n6297), .B2(n11017), .ZN(
        P2_U3523) );
  AOI22_X1 U11465 ( .A1(n11001), .A2(n10759), .B1(n5866), .B2(n11019), .ZN(
        P2_U3460) );
  OAI211_X1 U11466 ( .C1(n10762), .C2(n11047), .A(n10761), .B(n10760), .ZN(
        n10765) );
  AOI21_X1 U11467 ( .B1(n10851), .B2(n10911), .A(n10763), .ZN(n10764) );
  NOR2_X1 U11468 ( .A1(n10765), .A2(n10764), .ZN(n10768) );
  AOI22_X1 U11469 ( .A1(n11054), .A2(n10768), .B1(n10766), .B2(n11052), .ZN(
        P1_U3527) );
  INV_X1 U11470 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U11471 ( .A1(n11057), .A2(n10768), .B1(n10767), .B2(n11055), .ZN(
        P1_U3466) );
  XOR2_X1 U11472 ( .A(n10774), .B(n10770), .Z(n10793) );
  INV_X1 U11473 ( .A(n10771), .ZN(n10772) );
  OAI211_X1 U11474 ( .C1(n10772), .C2(n10773), .A(n10953), .B(n10808), .ZN(
        n10790) );
  OAI21_X1 U11475 ( .B1(n10773), .B2(n11047), .A(n10790), .ZN(n10782) );
  XNOR2_X1 U11476 ( .A(n10775), .B(n10774), .ZN(n10776) );
  OAI222_X1 U11477 ( .A1(n10781), .A2(n10780), .B1(n10779), .B2(n10778), .C1(
        n10777), .C2(n10776), .ZN(n10791) );
  AOI211_X1 U11478 ( .C1(n11050), .C2(n10793), .A(n10782), .B(n10791), .ZN(
        n10783) );
  AOI22_X1 U11479 ( .A1(n11054), .A2(n10783), .B1(n6689), .B2(n11052), .ZN(
        P1_U3528) );
  AOI22_X1 U11480 ( .A1(n11057), .A2(n10783), .B1(n6688), .B2(n11055), .ZN(
        P1_U3469) );
  NAND2_X1 U11481 ( .A1(n6460), .A2(n10784), .ZN(n10788) );
  OR2_X1 U11482 ( .A1(n10786), .A2(n10785), .ZN(n10787) );
  OAI211_X1 U11483 ( .C1(n10790), .C2(n10789), .A(n10788), .B(n10787), .ZN(
        n10792) );
  AOI211_X1 U11484 ( .C1(n10794), .C2(n10793), .A(n10792), .B(n10791), .ZN(
        n10796) );
  AOI22_X1 U11485 ( .A1(n11070), .A2(n10797), .B1(n10796), .B2(n10795), .ZN(
        P1_U3286) );
  INV_X1 U11486 ( .A(n10798), .ZN(n10799) );
  AOI21_X1 U11487 ( .B1(n10801), .B2(n10800), .A(n10799), .ZN(n10815) );
  XNOR2_X1 U11488 ( .A(n10802), .B(n10801), .ZN(n10806) );
  AOI22_X1 U11489 ( .A1(n11040), .A2(n10803), .B1(n10848), .B2(n11037), .ZN(
        n10804) );
  OAI21_X1 U11490 ( .B1(n10815), .B2(n10851), .A(n10804), .ZN(n10805) );
  AOI21_X1 U11491 ( .B1(n10806), .B2(n11035), .A(n10805), .ZN(n10820) );
  AOI211_X1 U11492 ( .C1(n10814), .C2(n10808), .A(n11043), .B(n10807), .ZN(
        n10816) );
  AOI21_X1 U11493 ( .B1(n10908), .B2(n10814), .A(n10816), .ZN(n10809) );
  OAI211_X1 U11494 ( .C1(n10815), .C2(n10911), .A(n10820), .B(n10809), .ZN(
        n10810) );
  INV_X1 U11495 ( .A(n10810), .ZN(n10811) );
  AOI22_X1 U11496 ( .A1(n11054), .A2(n10811), .B1(n6924), .B2(n11052), .ZN(
        P1_U3529) );
  AOI22_X1 U11497 ( .A1(n11057), .A2(n10811), .B1(n6927), .B2(n11055), .ZN(
        P1_U3472) );
  INV_X1 U11498 ( .A(n10812), .ZN(n10813) );
  AOI222_X1 U11499 ( .A1(n10814), .A2(n11060), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n11070), .C1(n11059), .C2(n10813), .ZN(n10819) );
  INV_X1 U11500 ( .A(n10815), .ZN(n10817) );
  AOI22_X1 U11501 ( .A1(n10817), .A2(n10863), .B1(n10291), .B2(n10816), .ZN(
        n10818) );
  OAI211_X1 U11502 ( .C1(n11070), .C2(n10820), .A(n10819), .B(n10818), .ZN(
        P1_U3285) );
  OAI211_X1 U11503 ( .C1(n10823), .C2(n11047), .A(n10822), .B(n10821), .ZN(
        n10826) );
  AOI21_X1 U11504 ( .B1(n10851), .B2(n10911), .A(n10824), .ZN(n10825) );
  NOR2_X1 U11505 ( .A1(n10826), .A2(n10825), .ZN(n10829) );
  AOI22_X1 U11506 ( .A1(n11054), .A2(n10829), .B1(n10827), .B2(n11052), .ZN(
        P1_U3530) );
  INV_X1 U11507 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U11508 ( .A1(n11057), .A2(n10829), .B1(n10828), .B2(n11055), .ZN(
        P1_U3475) );
  AOI22_X1 U11509 ( .A1(n10831), .A2(n10927), .B1(n10830), .B2(n10925), .ZN(
        n10832) );
  OAI211_X1 U11510 ( .C1(n10992), .C2(n10834), .A(n10833), .B(n10832), .ZN(
        n10835) );
  INV_X1 U11511 ( .A(n10835), .ZN(n10837) );
  AOI22_X1 U11512 ( .A1(n11018), .A2(n10837), .B1(n6310), .B2(n11017), .ZN(
        P2_U3527) );
  INV_X1 U11513 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U11514 ( .A1(n11001), .A2(n10837), .B1(n10836), .B2(n11019), .ZN(
        P2_U3472) );
  OAI21_X1 U11515 ( .B1(n10840), .B2(n10839), .A(n10838), .ZN(n10852) );
  INV_X1 U11516 ( .A(n10852), .ZN(n10864) );
  OAI211_X1 U11517 ( .C1(n10842), .C2(n10843), .A(n10953), .B(n10841), .ZN(
        n10861) );
  OAI21_X1 U11518 ( .B1(n10843), .B2(n11047), .A(n10861), .ZN(n10856) );
  NAND2_X1 U11519 ( .A1(n10845), .A2(n10844), .ZN(n10847) );
  XNOR2_X1 U11520 ( .A(n10847), .B(n10846), .ZN(n10854) );
  AOI22_X1 U11521 ( .A1(n11037), .A2(n10849), .B1(n10848), .B2(n11040), .ZN(
        n10850) );
  OAI21_X1 U11522 ( .B1(n10852), .B2(n10851), .A(n10850), .ZN(n10853) );
  AOI21_X1 U11523 ( .B1(n10854), .B2(n11035), .A(n10853), .ZN(n10867) );
  INV_X1 U11524 ( .A(n10867), .ZN(n10855) );
  AOI211_X1 U11525 ( .C1(n11028), .C2(n10864), .A(n10856), .B(n10855), .ZN(
        n10857) );
  AOI22_X1 U11526 ( .A1(n11054), .A2(n10857), .B1(n6179), .B2(n11052), .ZN(
        P1_U3531) );
  AOI22_X1 U11527 ( .A1(n11057), .A2(n10857), .B1(n6184), .B2(n11055), .ZN(
        P1_U3478) );
  INV_X1 U11528 ( .A(n10858), .ZN(n10859) );
  AOI222_X1 U11529 ( .A1(n10860), .A2(n11060), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n11070), .C1(n11059), .C2(n10859), .ZN(n10866) );
  INV_X1 U11530 ( .A(n10861), .ZN(n10862) );
  AOI22_X1 U11531 ( .A1(n10864), .A2(n10863), .B1(n10291), .B2(n10862), .ZN(
        n10865) );
  OAI211_X1 U11532 ( .C1(n11070), .C2(n10867), .A(n10866), .B(n10865), .ZN(
        P1_U3283) );
  NAND3_X1 U11533 ( .A1(n10869), .A2(n10868), .A3(n11015), .ZN(n10871) );
  OAI211_X1 U11534 ( .C1(n10872), .C2(n11010), .A(n10871), .B(n10870), .ZN(
        n10873) );
  NOR2_X1 U11535 ( .A1(n10874), .A2(n10873), .ZN(n10876) );
  AOI22_X1 U11536 ( .A1(n11018), .A2(n10876), .B1(n6307), .B2(n11017), .ZN(
        P2_U3528) );
  INV_X1 U11537 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U11538 ( .A1(n11001), .A2(n10876), .B1(n10875), .B2(n11019), .ZN(
        P2_U3475) );
  INV_X1 U11539 ( .A(n10877), .ZN(n10883) );
  INV_X1 U11540 ( .A(n10878), .ZN(n10879) );
  OAI22_X1 U11541 ( .A1(n10880), .A2(n11011), .B1(n10879), .B2(n11010), .ZN(
        n10882) );
  AOI211_X1 U11542 ( .C1(n10884), .C2(n10883), .A(n10882), .B(n10881), .ZN(
        n10886) );
  AOI22_X1 U11543 ( .A1(n11018), .A2(n10886), .B1(n6157), .B2(n11017), .ZN(
        P2_U3529) );
  INV_X1 U11544 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U11545 ( .A1(n11001), .A2(n10886), .B1(n10885), .B2(n11019), .ZN(
        P2_U3478) );
  NAND2_X1 U11546 ( .A1(n10887), .A2(n10908), .ZN(n10888) );
  NAND2_X1 U11547 ( .A1(n10889), .A2(n10888), .ZN(n10890) );
  AOI21_X1 U11548 ( .B1(n10891), .B2(n11028), .A(n10890), .ZN(n10892) );
  AOI22_X1 U11549 ( .A1(n11054), .A2(n10896), .B1(n10894), .B2(n11052), .ZN(
        P1_U3533) );
  INV_X1 U11550 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U11551 ( .A1(n11057), .A2(n10896), .B1(n10895), .B2(n11055), .ZN(
        P1_U3484) );
  NOR2_X1 U11552 ( .A1(n10897), .A2(n10992), .ZN(n10902) );
  OAI22_X1 U11553 ( .A1(n10899), .A2(n11011), .B1(n10898), .B2(n11010), .ZN(
        n10901) );
  AOI211_X1 U11554 ( .C1(n10902), .C2(n7680), .A(n10901), .B(n10900), .ZN(
        n10904) );
  AOI22_X1 U11555 ( .A1(n11018), .A2(n10904), .B1(n6547), .B2(n11017), .ZN(
        P2_U3530) );
  INV_X1 U11556 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U11557 ( .A1(n11001), .A2(n10904), .B1(n10903), .B2(n11019), .ZN(
        P2_U3481) );
  INV_X1 U11558 ( .A(n10910), .ZN(n10914) );
  AOI211_X1 U11559 ( .C1(n10908), .C2(n10907), .A(n10906), .B(n10905), .ZN(
        n10909) );
  OAI21_X1 U11560 ( .B1(n10911), .B2(n10910), .A(n10909), .ZN(n10912) );
  AOI21_X1 U11561 ( .B1(n10914), .B2(n10913), .A(n10912), .ZN(n10916) );
  AOI22_X1 U11562 ( .A1(n11054), .A2(n10916), .B1(n10915), .B2(n11052), .ZN(
        P1_U3534) );
  AOI22_X1 U11563 ( .A1(n11057), .A2(n10916), .B1(n7358), .B2(n11055), .ZN(
        P1_U3487) );
  OAI21_X1 U11564 ( .B1(n10918), .B2(n10920), .A(n10917), .ZN(n10919) );
  INV_X1 U11565 ( .A(n10919), .ZN(n10945) );
  INV_X1 U11566 ( .A(n10920), .ZN(n10921) );
  XNOR2_X1 U11567 ( .A(n10922), .B(n10921), .ZN(n10924) );
  NAND2_X1 U11568 ( .A1(n10924), .A2(n10923), .ZN(n10941) );
  AOI21_X1 U11569 ( .B1(n10939), .B2(n10925), .A(n10936), .ZN(n10930) );
  OAI211_X1 U11570 ( .C1(n10929), .C2(n10928), .A(n10927), .B(n10926), .ZN(
        n10942) );
  NAND3_X1 U11571 ( .A1(n10941), .A2(n10930), .A3(n10942), .ZN(n10931) );
  AOI21_X1 U11572 ( .B1(n10945), .B2(n11015), .A(n10931), .ZN(n10933) );
  AOI22_X1 U11573 ( .A1(n11018), .A2(n10933), .B1(n7163), .B2(n11017), .ZN(
        P2_U3531) );
  INV_X1 U11574 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U11575 ( .A1(n11001), .A2(n10933), .B1(n10932), .B2(n11019), .ZN(
        P2_U3484) );
  NOR2_X1 U11576 ( .A1(n10935), .A2(n10934), .ZN(n10937) );
  AOI211_X1 U11577 ( .C1(n10939), .C2(n10938), .A(n10937), .B(n10936), .ZN(
        n10940) );
  OAI211_X1 U11578 ( .C1(n5819), .C2(n10942), .A(n10941), .B(n10940), .ZN(
        n10943) );
  AOI21_X1 U11579 ( .B1(n10945), .B2(n10944), .A(n10943), .ZN(n10947) );
  AOI22_X1 U11580 ( .A1(n9426), .A2(n10948), .B1(n10947), .B2(n10946), .ZN(
        P2_U3285) );
  OR2_X1 U11581 ( .A1(n10949), .A2(n10956), .ZN(n10950) );
  AND2_X1 U11582 ( .A1(n10951), .A2(n10950), .ZN(n10972) );
  OAI211_X1 U11583 ( .C1(n10954), .C2(n10955), .A(n10953), .B(n10952), .ZN(
        n10969) );
  OAI21_X1 U11584 ( .B1(n10955), .B2(n11047), .A(n10969), .ZN(n10962) );
  XNOR2_X1 U11585 ( .A(n10957), .B(n10956), .ZN(n10960) );
  AOI222_X1 U11586 ( .A1(n11035), .A2(n10960), .B1(n10959), .B2(n11037), .C1(
        n10958), .C2(n11040), .ZN(n10975) );
  INV_X1 U11587 ( .A(n10975), .ZN(n10961) );
  AOI211_X1 U11588 ( .C1(n10972), .C2(n11050), .A(n10962), .B(n10961), .ZN(
        n10965) );
  AOI22_X1 U11589 ( .A1(n11054), .A2(n10965), .B1(n10963), .B2(n11052), .ZN(
        P1_U3535) );
  INV_X1 U11590 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U11591 ( .A1(n11057), .A2(n10965), .B1(n10964), .B2(n11055), .ZN(
        P1_U3490) );
  INV_X1 U11592 ( .A(n10966), .ZN(n10967) );
  AOI222_X1 U11593 ( .A1(n10968), .A2(n11060), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n11070), .C1(n11059), .C2(n10967), .ZN(n10974) );
  NOR2_X1 U11594 ( .A1(n10969), .A2(n11063), .ZN(n10970) );
  AOI21_X1 U11595 ( .B1(n10972), .B2(n10971), .A(n10970), .ZN(n10973) );
  OAI211_X1 U11596 ( .C1(n11070), .C2(n10975), .A(n10974), .B(n10973), .ZN(
        P1_U3279) );
  INV_X1 U11597 ( .A(n10976), .ZN(n10977) );
  OAI22_X1 U11598 ( .A1(n10978), .A2(n11011), .B1(n10977), .B2(n11010), .ZN(
        n10980) );
  AOI211_X1 U11599 ( .C1(n11015), .C2(n10981), .A(n10980), .B(n10979), .ZN(
        n10983) );
  AOI22_X1 U11600 ( .A1(n11018), .A2(n10983), .B1(n6164), .B2(n11017), .ZN(
        P2_U3532) );
  INV_X1 U11601 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U11602 ( .A1(n11001), .A2(n10983), .B1(n10982), .B2(n11019), .ZN(
        P2_U3487) );
  INV_X1 U11603 ( .A(n10984), .ZN(n10987) );
  OAI211_X1 U11604 ( .C1(n10987), .C2(n11047), .A(n10986), .B(n10985), .ZN(
        n10988) );
  AOI21_X1 U11605 ( .B1(n11050), .B2(n10989), .A(n10988), .ZN(n10991) );
  AOI22_X1 U11606 ( .A1(n11054), .A2(n10991), .B1(n10990), .B2(n11052), .ZN(
        P1_U3536) );
  AOI22_X1 U11607 ( .A1(n11057), .A2(n10991), .B1(n7715), .B2(n11055), .ZN(
        P1_U3493) );
  NOR2_X1 U11608 ( .A1(n10993), .A2(n10992), .ZN(n10998) );
  OAI22_X1 U11609 ( .A1(n10995), .A2(n11011), .B1(n10994), .B2(n11010), .ZN(
        n10997) );
  AOI211_X1 U11610 ( .C1(n10998), .C2(n7777), .A(n10997), .B(n10996), .ZN(
        n11000) );
  AOI22_X1 U11611 ( .A1(n11018), .A2(n11000), .B1(n6997), .B2(n11017), .ZN(
        P2_U3533) );
  INV_X1 U11612 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U11613 ( .A1(n11001), .A2(n11000), .B1(n10999), .B2(n11019), .ZN(
        P2_U3490) );
  OAI211_X1 U11614 ( .C1(n5390), .C2(n11047), .A(n11003), .B(n11002), .ZN(
        n11004) );
  AOI21_X1 U11615 ( .B1(n11050), .B2(n11005), .A(n11004), .ZN(n11008) );
  AOI22_X1 U11616 ( .A1(n11054), .A2(n11008), .B1(n11006), .B2(n11052), .ZN(
        P1_U3537) );
  INV_X1 U11617 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11007) );
  AOI22_X1 U11618 ( .A1(n11057), .A2(n11008), .B1(n11007), .B2(n11055), .ZN(
        P1_U3496) );
  INV_X1 U11619 ( .A(n11009), .ZN(n11016) );
  OAI22_X1 U11620 ( .A1(n11012), .A2(n11011), .B1(n5472), .B2(n11010), .ZN(
        n11013) );
  AOI211_X1 U11621 ( .C1(n11016), .C2(n11015), .A(n11014), .B(n11013), .ZN(
        n11021) );
  AOI22_X1 U11622 ( .A1(n11018), .A2(n11021), .B1(n7619), .B2(n11017), .ZN(
        P2_U3534) );
  INV_X1 U11623 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U11624 ( .A1(n11001), .A2(n11021), .B1(n11020), .B2(n11019), .ZN(
        P2_U3493) );
  INV_X1 U11625 ( .A(n11022), .ZN(n11027) );
  OAI21_X1 U11626 ( .B1(n11024), .B2(n11047), .A(n11023), .ZN(n11026) );
  AOI211_X1 U11627 ( .C1(n11028), .C2(n11027), .A(n11026), .B(n11025), .ZN(
        n11030) );
  AOI22_X1 U11628 ( .A1(n11054), .A2(n11030), .B1(n11029), .B2(n11052), .ZN(
        P1_U3538) );
  AOI22_X1 U11629 ( .A1(n11057), .A2(n11030), .B1(n7806), .B2(n11055), .ZN(
        P1_U3499) );
  OAI21_X1 U11630 ( .B1(n11032), .B2(n11033), .A(n11031), .ZN(n11065) );
  INV_X1 U11631 ( .A(n11065), .ZN(n11051) );
  XNOR2_X1 U11632 ( .A(n11034), .B(n11033), .ZN(n11036) );
  NAND2_X1 U11633 ( .A1(n11036), .A2(n11035), .ZN(n11042) );
  AOI22_X1 U11634 ( .A1(n11040), .A2(n11039), .B1(n11038), .B2(n11037), .ZN(
        n11041) );
  AOI21_X1 U11635 ( .B1(n11044), .B2(n11061), .A(n11043), .ZN(n11046) );
  NAND2_X1 U11636 ( .A1(n11046), .A2(n11045), .ZN(n11062) );
  OAI211_X1 U11637 ( .C1(n11048), .C2(n11047), .A(n11069), .B(n11062), .ZN(
        n11049) );
  AOI21_X1 U11638 ( .B1(n11051), .B2(n11050), .A(n11049), .ZN(n11056) );
  AOI22_X1 U11639 ( .A1(n11054), .A2(n11056), .B1(n11053), .B2(n11052), .ZN(
        P1_U3539) );
  AOI22_X1 U11640 ( .A1(n11057), .A2(n11056), .B1(n7856), .B2(n11055), .ZN(
        P1_U3502) );
  AOI222_X1 U11641 ( .A1(n11061), .A2(n11060), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n11070), .C1(n11059), .C2(n11058), .ZN(n11068) );
  OAI22_X1 U11642 ( .A1(n11065), .A2(n11064), .B1(n11063), .B2(n11062), .ZN(
        n11066) );
  INV_X1 U11643 ( .A(n11066), .ZN(n11067) );
  OAI211_X1 U11644 ( .C1(n11070), .C2(n11069), .A(n11068), .B(n11067), .ZN(
        P1_U3275) );
  XNOR2_X1 U11645 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X2 U5136 ( .A(n6600), .Z(n9086) );
  CLKBUF_X1 U5180 ( .A(n6571), .Z(n8490) );
  INV_X1 U5193 ( .A(n6609), .ZN(n7011) );
  CLKBUF_X1 U5194 ( .A(n5882), .Z(n8040) );
  OR2_X1 U5258 ( .A1(n10713), .A2(n8859), .ZN(n11011) );
  OAI211_X1 U5370 ( .C1(n7005), .C2(n6581), .A(n6580), .B(n6579), .ZN(n8406)
         );
endmodule

