

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3104, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068;

  INV_X1 U3536 ( .A(n3130), .ZN(n3093) );
  XNOR2_X1 U3537 ( .A(n4359), .B(n4358), .ZN(n5333) );
  CLKBUF_X2 U3538 ( .A(n6324), .Z(n3130) );
  INV_X2 U3539 ( .A(n6329), .ZN(n6360) );
  OR2_X1 U3540 ( .A1(n4267), .A2(n4253), .ZN(n4976) );
  OAI21_X1 U3541 ( .B1(n3711), .B2(n3822), .A(n3710), .ZN(n4666) );
  NAND2_X1 U3542 ( .A1(n3417), .A2(n3394), .ZN(n4589) );
  OR2_X1 U3544 ( .A1(n3355), .A2(n3354), .ZN(n3356) );
  NAND2_X1 U3545 ( .A1(n3309), .A2(n3308), .ZN(n3355) );
  OR2_X1 U3546 ( .A1(n3285), .A2(n3317), .ZN(n4340) );
  INV_X1 U3547 ( .A(n4657), .ZN(n5023) );
  CLKBUF_X2 U3548 ( .A(n4288), .Z(n4313) );
  CLKBUF_X2 U3549 ( .A(n3365), .Z(n4070) );
  CLKBUF_X2 U3550 ( .A(n3338), .Z(n3360) );
  CLKBUF_X2 U3551 ( .A(n3396), .Z(n3096) );
  CLKBUF_X2 U3552 ( .A(n3329), .Z(n4291) );
  BUF_X1 U3553 ( .A(n3283), .Z(n4239) );
  INV_X1 U3554 ( .A(n4724), .ZN(n4256) );
  INV_X1 U3555 ( .A(n3283), .ZN(n3290) );
  AND2_X2 U3557 ( .A1(n4552), .A2(n4442), .ZN(n3429) );
  AND2_X2 U3558 ( .A1(n4630), .A2(n3154), .ZN(n3329) );
  AND2_X2 U3559 ( .A1(n4552), .A2(n4553), .ZN(n3396) );
  AND2_X2 U3560 ( .A1(n4442), .A2(n4601), .ZN(n3365) );
  CLKBUF_X2 U3561 ( .A(n3359), .Z(n3097) );
  AND2_X2 U3562 ( .A1(n4553), .A2(n4601), .ZN(n3339) );
  NOR2_X1 U3563 ( .A1(n3124), .A2(n5169), .ZN(n4228) );
  XNOR2_X1 U3564 ( .A(n3572), .B(n3483), .ZN(n3724) );
  BUF_X1 U3565 ( .A(n5169), .Z(n3131) );
  NAND2_X1 U3566 ( .A1(n3553), .A2(n3476), .ZN(n3572) );
  AND2_X1 U3567 ( .A1(n3537), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6467)
         );
  OAI21_X1 U3568 ( .B1(n3679), .B2(STATE2_REG_0__SCAN_IN), .A(n3375), .ZN(
        n3376) );
  OR2_X1 U3570 ( .A1(n6470), .A2(n6467), .ZN(n3538) );
  INV_X1 U3571 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6782) );
  NOR2_X1 U3572 ( .A1(n4308), .A2(n5012), .ZN(n4393) );
  INV_X1 U3573 ( .A(n6478), .ZN(n5632) );
  NAND2_X2 U3574 ( .A1(n3112), .A2(n3356), .ZN(n3679) );
  OR2_X1 U3575 ( .A1(n4267), .A2(n4136), .ZN(n6515) );
  OR2_X1 U3576 ( .A1(n4267), .A2(n4571), .ZN(n6521) );
  AND2_X1 U3577 ( .A1(n3294), .A2(n4724), .ZN(n3088) );
  AND4_X1 U3578 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n3089)
         );
  AND2_X1 U3579 ( .A1(n3111), .A2(n3108), .ZN(n3090) );
  AND2_X1 U3581 ( .A1(n4552), .A2(n4553), .ZN(n3091) );
  XNOR2_X1 U3582 ( .A(n3515), .B(n3514), .ZN(n3517) );
  AOI21_X2 U3583 ( .B1(n5002), .B2(n6779), .A(n5001), .ZN(n5003) );
  XNOR2_X2 U3584 ( .A(n3550), .B(n4255), .ZN(n4737) );
  NAND2_X2 U3585 ( .A1(n3549), .A2(n3548), .ZN(n3550) );
  AOI21_X2 U3586 ( .B1(n3314), .B2(n4251), .A(n3313), .ZN(n4250) );
  INV_X1 U3587 ( .A(n4119), .ZN(n3092) );
  AOI211_X2 U3588 ( .C1(n5502), .C2(n5476), .A(n5475), .B(n5474), .ZN(n5699)
         );
  AND2_X1 U3589 ( .A1(n5139), .A2(n5138), .ZN(n5141) );
  OR2_X1 U3590 ( .A1(n5074), .A2(n4374), .ZN(n5051) );
  AND2_X1 U3591 ( .A1(n3115), .A2(n3116), .ZN(n5126) );
  NOR2_X1 U3592 ( .A1(n5184), .A2(n5188), .ZN(n5167) );
  NAND2_X1 U3593 ( .A1(n3690), .A2(n4517), .ZN(n4530) );
  NAND2_X1 U3594 ( .A1(n4980), .A2(n4187), .ZN(n4981) );
  NOR2_X2 U3595 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  MUX2_X1 U3596 ( .A(n4228), .B(n3131), .S(EBX_REG_3__SCAN_IN), .Z(n4153) );
  OAI21_X1 U3597 ( .B1(n5169), .B2(EBX_REG_0__SCAN_IN), .A(n4138), .ZN(n4499)
         );
  OR2_X1 U3598 ( .A1(n4239), .A2(n4647), .ZN(n3423) );
  CLKBUF_X2 U3599 ( .A(n4147), .Z(n4349) );
  INV_X1 U3600 ( .A(n4127), .ZN(n3094) );
  OR2_X1 U3601 ( .A1(n4137), .A2(n3128), .ZN(n4210) );
  INV_X2 U3602 ( .A(n4147), .ZN(n5169) );
  CLKBUF_X2 U3603 ( .A(n3358), .Z(n4311) );
  BUF_X2 U3604 ( .A(n3429), .Z(n3095) );
  CLKBUF_X2 U3605 ( .A(n3367), .Z(n4296) );
  MUX2_X1 U3606 ( .A(n4383), .B(n5002), .S(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .Z(n4104) );
  OAI21_X1 U3607 ( .B1(n4393), .B2(n4395), .A(n4394), .ZN(n5019) );
  XNOR2_X1 U3608 ( .A(n4394), .B(n4339), .ZN(n5042) );
  OAI21_X1 U3609 ( .B1(n5141), .B2(n5124), .A(n5123), .ZN(n5487) );
  INV_X1 U3610 ( .A(n3111), .ZN(n5066) );
  NAND2_X1 U3611 ( .A1(n3592), .A2(n3591), .ZN(n4962) );
  INV_X1 U3612 ( .A(n4355), .ZN(n4359) );
  NOR3_X1 U3613 ( .A1(n5005), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6843), 
        .ZN(n4263) );
  AOI211_X1 U3614 ( .C1(EBX_REG_5__SCAN_IN), .C2(n6358), .A(n6354), .B(n6353), 
        .ZN(n6355) );
  NOR4_X1 U3615 ( .A1(n5051), .A2(REIP_REG_31__SCAN_IN), .A3(n6797), .A4(n6703), .ZN(n4380) );
  NAND2_X1 U3616 ( .A1(n3730), .A2(n3729), .ZN(n4835) );
  NOR2_X1 U3617 ( .A1(n5184), .A2(n5188), .ZN(n3115) );
  CLKBUF_X1 U3618 ( .A(n3567), .Z(n3098) );
  NAND2_X1 U3619 ( .A1(n5532), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5533) );
  XNOR2_X1 U3620 ( .A(n3539), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4948)
         );
  NAND2_X1 U3621 ( .A1(n3694), .A2(n3693), .ZN(n4618) );
  CLKBUF_X1 U3622 ( .A(n3695), .Z(n5855) );
  CLKBUF_X1 U3623 ( .A(n5387), .Z(n6388) );
  AND2_X2 U3624 ( .A1(n5299), .A2(n4364), .ZN(n6329) );
  AND2_X1 U3625 ( .A1(n5293), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5299) );
  AND2_X1 U3626 ( .A1(n4132), .A2(n4131), .ZN(n4267) );
  INV_X2 U3627 ( .A(n5436), .ZN(n6387) );
  AND2_X2 U3628 ( .A1(n5368), .A2(n5264), .ZN(n4980) );
  XNOR2_X1 U3629 ( .A(n4589), .B(n4590), .ZN(n4550) );
  OR2_X2 U3630 ( .A1(n5278), .A2(n5280), .ZN(n5367) );
  CLKBUF_X1 U3631 ( .A(n4641), .Z(n5906) );
  INV_X1 U3632 ( .A(n3413), .ZN(n3528) );
  OR3_X2 U3633 ( .A1(n4525), .A2(n4130), .A3(n4256), .ZN(n4131) );
  XNOR2_X1 U3634 ( .A(n3517), .B(n3376), .ZN(n4641) );
  NAND2_X1 U3635 ( .A1(n4838), .A2(n5379), .ZN(n5278) );
  CLKBUF_X1 U3636 ( .A(n4567), .Z(n5848) );
  AOI21_X1 U3637 ( .B1(n4567), .B2(n4647), .A(n3412), .ZN(n3413) );
  OR2_X2 U3638 ( .A1(n4420), .A2(n6646), .ZN(n4525) );
  AND2_X1 U3639 ( .A1(n4793), .A2(n4839), .ZN(n4838) );
  AOI21_X1 U3640 ( .B1(n3645), .B2(n3644), .A(n3643), .ZN(n3652) );
  NAND2_X1 U3641 ( .A1(n4520), .A2(n4519), .ZN(n4518) );
  OAI211_X1 U3642 ( .C1(n3353), .C2(n3424), .A(n3352), .B(n3492), .ZN(n3514)
         );
  AND2_X2 U3643 ( .A1(n3337), .A2(n4239), .ZN(n3638) );
  AND2_X1 U3644 ( .A1(n4150), .A2(n4149), .ZN(n4533) );
  NAND2_X1 U3645 ( .A1(n3094), .A2(n3088), .ZN(n3286) );
  INV_X1 U3646 ( .A(n4210), .ZN(n4220) );
  CLKBUF_X1 U3647 ( .A(n3677), .Z(n4717) );
  CLKBUF_X1 U3648 ( .A(n3290), .Z(n4685) );
  AND2_X1 U3649 ( .A1(n4349), .A2(n4210), .ZN(n4498) );
  CLKBUF_X1 U3650 ( .A(n3294), .Z(n4698) );
  OR2_X1 U3651 ( .A1(n3350), .A2(n3349), .ZN(n3575) );
  AND4_X2 U3652 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n4724)
         );
  NAND3_X1 U3653 ( .A1(n3178), .A2(n3177), .A3(n3139), .ZN(n3284) );
  AND3_X1 U3654 ( .A1(n3238), .A2(n3237), .A3(n3236), .ZN(n3254) );
  AND4_X1 U3655 ( .A1(n3196), .A2(n3195), .A3(n3194), .A4(n3193), .ZN(n3197)
         );
  AND4_X1 U3656 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3199)
         );
  AND4_X1 U3657 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3252)
         );
  AND4_X1 U3658 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), .ZN(n3251)
         );
  AND4_X1 U3659 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3233)
         );
  AND4_X1 U3660 ( .A1(n3242), .A2(n3241), .A3(n3240), .A4(n3239), .ZN(n3253)
         );
  AND4_X1 U3661 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3169)
         );
  AND4_X1 U3662 ( .A1(n3225), .A2(n3224), .A3(n3223), .A4(n3222), .ZN(n3231)
         );
  AND4_X1 U3663 ( .A1(n3167), .A2(n3166), .A3(n3165), .A4(n3164), .ZN(n3168)
         );
  CLKBUF_X2 U3664 ( .A(n3339), .Z(n4321) );
  INV_X2 U3665 ( .A(n6746), .ZN(n6734) );
  AND2_X2 U3666 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4601) );
  NOR2_X1 U3669 ( .A1(n5452), .A2(n3101), .ZN(n5002) );
  OR2_X1 U3670 ( .A1(n3141), .A2(n5653), .ZN(n3101) );
  NAND2_X1 U3671 ( .A1(n3572), .A2(n3477), .ZN(n3707) );
  OR2_X1 U3672 ( .A1(n3292), .A2(n3127), .ZN(n3123) );
  AOI211_X2 U3673 ( .C1(n5632), .C2(n5526), .A(n5525), .B(n5524), .ZN(n5527)
         );
  NOR2_X2 U3675 ( .A1(n5687), .A2(n5678), .ZN(n5666) );
  AND2_X2 U3676 ( .A1(n3291), .A2(n3201), .ZN(n3674) );
  OAI21_X1 U3677 ( .B1(n3679), .B2(STATE2_REG_0__SCAN_IN), .A(n3496), .ZN(
        n3502) );
  INV_X2 U3678 ( .A(n4254), .ZN(n3292) );
  AND2_X1 U3681 ( .A1(n3305), .A2(n3384), .ZN(n3104) );
  CLKBUF_X1 U3683 ( .A(n5637), .Z(n3106) );
  NAND2_X1 U3684 ( .A1(n5535), .A2(n5534), .ZN(n3107) );
  AND2_X2 U3685 ( .A1(n3107), .A2(n5533), .ZN(n5544) );
  NAND2_X1 U3686 ( .A1(n3491), .A2(n3490), .ZN(n3539) );
  OAI22_X2 U3687 ( .A1(n5565), .A2(n5566), .B1(n3597), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5535) );
  AOI21_X2 U3688 ( .B1(n5554), .B2(n5536), .A(n5544), .ZN(n5537) );
  NAND2_X1 U3689 ( .A1(n3538), .A2(n6468), .ZN(n4949) );
  OR2_X1 U3690 ( .A1(n5002), .A2(n4383), .ZN(n4384) );
  OAI21_X1 U3691 ( .B1(n3707), .B2(n3822), .A(n3706), .ZN(n4788) );
  AND2_X1 U3692 ( .A1(n4091), .A2(n3108), .ZN(n3109) );
  INV_X1 U3693 ( .A(n5067), .ZN(n3108) );
  AND2_X1 U3694 ( .A1(n3109), .A2(n4051), .ZN(n3110) );
  AND2_X1 U3695 ( .A1(n5093), .A2(n4051), .ZN(n3111) );
  NAND2_X1 U3696 ( .A1(n3355), .A2(n3354), .ZN(n3112) );
  INV_X1 U3697 ( .A(n3692), .ZN(n3113) );
  NAND2_X1 U3698 ( .A1(n3355), .A2(n3354), .ZN(n3383) );
  AOI21_X1 U3699 ( .B1(n5042), .B2(n6472), .A(n5040), .ZN(n5041) );
  NOR2_X2 U3700 ( .A1(n3969), .A2(n6955), .ZN(n3963) );
  NOR2_X2 U3701 ( .A1(n3785), .A2(n5282), .ZN(n3745) );
  NOR2_X2 U3702 ( .A1(n3791), .A2(n5266), .ZN(n3805) );
  NAND2_X1 U3703 ( .A1(n3607), .A2(n3606), .ZN(n5462) );
  XNOR2_X1 U3704 ( .A(n3415), .B(n3394), .ZN(n4567) );
  NAND2_X1 U3705 ( .A1(n5042), .A2(n3093), .ZN(n3114) );
  NAND2_X1 U3706 ( .A1(n3114), .A2(n4382), .ZN(U2796) );
  AND2_X1 U3707 ( .A1(n3117), .A2(n4206), .ZN(n3116) );
  INV_X1 U3708 ( .A(n5154), .ZN(n3117) );
  AND2_X1 U3709 ( .A1(n4196), .A2(n4195), .ZN(n3118) );
  AND2_X1 U3710 ( .A1(n4674), .A2(n3120), .ZN(n3121) );
  INV_X1 U3711 ( .A(n4532), .ZN(n3119) );
  INV_X1 U3712 ( .A(n4621), .ZN(n3120) );
  AND2_X1 U3713 ( .A1(n3119), .A2(n3120), .ZN(n4620) );
  OR2_X1 U3714 ( .A1(n4137), .A2(n3128), .ZN(n3122) );
  AND2_X2 U3715 ( .A1(n4554), .A2(n4442), .ZN(n3357) );
  NAND2_X1 U3716 ( .A1(n4196), .A2(n4195), .ZN(n5215) );
  OR2_X1 U3717 ( .A1(n3292), .A2(n3127), .ZN(n3124) );
  NAND2_X1 U3719 ( .A1(n4152), .A2(n4151), .ZN(n4532) );
  AND2_X2 U3720 ( .A1(n5099), .A2(n4223), .ZN(n5081) );
  AND2_X2 U3721 ( .A1(n3310), .A2(n3088), .ZN(n4126) );
  AND2_X2 U3722 ( .A1(n3714), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3703)
         );
  NOR2_X2 U3723 ( .A1(n3713), .A2(n6835), .ZN(n3714) );
  AND2_X1 U3724 ( .A1(n5385), .A2(n4254), .ZN(n4119) );
  NAND2_X1 U3725 ( .A1(n4137), .A2(n4254), .ZN(n4147) );
  AOI211_X2 U3726 ( .C1(n5089), .C2(REIP_REG_27__SCAN_IN), .A(n5076), .B(n5075), .ZN(n5077) );
  AOI211_X2 U3727 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5174), .A(n5161), .B(n5160), .ZN(n5162) );
  AND4_X1 U3728 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3127)
         );
  AND4_X1 U3729 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3128)
         );
  AOI211_X2 U3730 ( .C1(REIP_REG_25__SCAN_IN), .C2(n5134), .A(n5108), .B(n5107), .ZN(n5109) );
  INV_X2 U3731 ( .A(n5027), .ZN(n3129) );
  NAND2_X4 U3732 ( .A1(n5039), .A2(n3146), .ZN(n5027) );
  NAND2_X1 U3733 ( .A1(n5293), .A2(n4348), .ZN(n6324) );
  NOR2_X2 U3734 ( .A1(n4670), .A2(n4792), .ZN(n4793) );
  XNOR2_X2 U3735 ( .A(n4238), .B(n4354), .ZN(n4960) );
  CLKBUF_X1 U3736 ( .A(n3323), .Z(n4312) );
  INV_X1 U3738 ( .A(n3620), .ZN(n3337) );
  CLKBUF_X1 U3739 ( .A(n3357), .Z(n4314) );
  OR2_X1 U3740 ( .A1(n5532), .A2(n5788), .ZN(n5531) );
  OR2_X1 U3741 ( .A1(n3373), .A2(n3372), .ZN(n3519) );
  NAND2_X2 U3742 ( .A1(n3673), .A2(n3672), .ZN(n4420) );
  NAND2_X1 U3743 ( .A1(n3670), .A2(n3669), .ZN(n3673) );
  NOR2_X1 U3744 ( .A1(n5907), .A2(n5906), .ZN(n5957) );
  AOI22_X1 U3745 ( .A1(n3429), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3155) );
  CLKBUF_X1 U3746 ( .A(n3323), .Z(n4290) );
  NOR2_X1 U3747 ( .A1(n3184), .A2(n3144), .ZN(n3200) );
  NAND2_X1 U3748 ( .A1(n3638), .A2(n4119), .ZN(n3660) );
  INV_X1 U3749 ( .A(n3638), .ZN(n3657) );
  OR2_X1 U3750 ( .A1(n3435), .A2(n3434), .ZN(n3489) );
  OR2_X1 U3751 ( .A1(n4049), .A2(n5152), .ZN(n5110) );
  AND2_X1 U3752 ( .A1(n5228), .A2(n5230), .ZN(n5212) );
  NOR2_X1 U3753 ( .A1(n5247), .A2(n5248), .ZN(n5228) );
  NAND2_X1 U3754 ( .A1(n3840), .A2(n3839), .ZN(n5247) );
  INV_X1 U3755 ( .A(n5355), .ZN(n3839) );
  INV_X1 U3756 ( .A(n5354), .ZN(n3840) );
  NAND3_X1 U3757 ( .A1(n4624), .A2(n4788), .A3(n3723), .ZN(n4789) );
  AND2_X1 U3758 ( .A1(n4666), .A2(n4623), .ZN(n3723) );
  INV_X1 U3759 ( .A(n4342), .ZN(n4334) );
  INV_X1 U3760 ( .A(n3687), .ZN(n4083) );
  INV_X1 U3761 ( .A(n5216), .ZN(n4200) );
  AND2_X1 U3762 ( .A1(n3500), .A2(n3499), .ZN(n3504) );
  INV_X1 U3763 ( .A(n3495), .ZN(n3496) );
  NAND3_X1 U3764 ( .A1(n3276), .A2(n3094), .A3(n4256), .ZN(n3285) );
  NAND2_X1 U3765 ( .A1(n3422), .A2(n3421), .ZN(n4590) );
  OR2_X2 U3766 ( .A1(n3211), .A2(n3210), .ZN(n4137) );
  INV_X1 U3767 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4756) );
  CLKBUF_X1 U3768 ( .A(n3284), .Z(n4512) );
  AOI21_X1 U3770 ( .B1(n3678), .B2(n4717), .A(n6782), .ZN(n4511) );
  NOR2_X1 U3771 ( .A1(n4333), .A2(n5014), .ZN(n4345) );
  NAND2_X1 U3772 ( .A1(n4393), .A2(n4395), .ZN(n4394) );
  NAND2_X1 U3773 ( .A1(n4087), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4333)
         );
  INV_X1 U3774 ( .A(n4498), .ZN(n4356) );
  AND2_X1 U3775 ( .A1(n3596), .A2(n3595), .ZN(n3600) );
  CLKBUF_X1 U3776 ( .A(n4550), .Z(n4551) );
  INV_X1 U3777 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U3778 ( .A1(n4648), .A2(n4647), .ZN(n5840) );
  INV_X1 U3779 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6864) );
  INV_X1 U3780 ( .A(n6120), .ZN(n5956) );
  AND2_X1 U3781 ( .A1(n5436), .A2(n4526), .ZN(n6385) );
  AND2_X1 U3782 ( .A1(n5436), .A2(n4527), .ZN(n5434) );
  OR2_X1 U3783 ( .A1(n5395), .A2(n6178), .ZN(n4099) );
  NAND2_X1 U3784 ( .A1(n5625), .A2(n4093), .ZN(n5630) );
  INV_X1 U3785 ( .A(n6498), .ZN(n6465) );
  INV_X1 U3786 ( .A(n5630), .ZN(n6466) );
  OR2_X1 U3787 ( .A1(n5006), .A2(n5037), .ZN(n5007) );
  INV_X1 U3788 ( .A(n6515), .ZN(n6502) );
  OR2_X1 U3789 ( .A1(n4267), .A2(n4242), .ZN(n6500) );
  OR2_X1 U3790 ( .A1(n4973), .A2(n4972), .ZN(n5765) );
  CLKBUF_X1 U3791 ( .A(n3678), .Z(n6120) );
  INV_X1 U3792 ( .A(n5998), .ZN(n6186) );
  INV_X1 U3793 ( .A(n4551), .ZN(n6070) );
  BUF_X1 U3794 ( .A(n4639), .Z(n5852) );
  NAND2_X1 U3795 ( .A1(n5023), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3620) );
  INV_X1 U3797 ( .A(n3409), .ZN(n3532) );
  AOI22_X1 U3798 ( .A1(n3357), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3429), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U3799 ( .A1(n3442), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U3800 ( .A1(n3357), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U3801 ( .A1(n3358), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U3802 ( .A1(n3323), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3151) );
  CLKBUF_X1 U3803 ( .A(n3357), .Z(n3344) );
  OR2_X1 U3804 ( .A1(n3473), .A2(n3472), .ZN(n3484) );
  OR2_X1 U3805 ( .A1(n3448), .A2(n3447), .ZN(n3545) );
  INV_X1 U3806 ( .A(n4502), .ZN(n3180) );
  OR2_X1 U3807 ( .A1(n3335), .A2(n3334), .ZN(n3518) );
  AND2_X1 U3808 ( .A1(n3657), .A2(n4111), .ZN(n3651) );
  NAND2_X1 U3809 ( .A1(n4502), .A2(n3284), .ZN(n4127) );
  INV_X1 U3810 ( .A(n3423), .ZN(n4504) );
  NAND2_X1 U3811 ( .A1(n3293), .A2(n3292), .ZN(n3508) );
  INV_X1 U3812 ( .A(n4657), .ZN(n3293) );
  NAND2_X1 U3813 ( .A1(n5093), .A2(n3110), .ZN(n4308) );
  OR2_X1 U3814 ( .A1(n4050), .A2(n5110), .ZN(n5094) );
  OR2_X1 U3815 ( .A1(n5163), .A2(n5164), .ZN(n5152) );
  NOR2_X1 U3816 ( .A1(n4834), .A2(n3790), .ZN(n5260) );
  NAND2_X1 U3817 ( .A1(n3731), .A2(n4835), .ZN(n4834) );
  INV_X1 U3818 ( .A(n4789), .ZN(n3731) );
  OR2_X1 U3819 ( .A1(n3553), .A2(n3476), .ZN(n3477) );
  INV_X1 U3820 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6835) );
  AND2_X1 U3821 ( .A1(n5627), .A2(n5626), .ZN(n3566) );
  NAND4_X1 U3822 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .ZN(n3283)
         );
  AND4_X1 U3823 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n3198)
         );
  INV_X1 U3824 ( .A(n3660), .ZN(n3668) );
  AND2_X1 U3825 ( .A1(n3667), .A2(n3666), .ZN(n4113) );
  INV_X1 U3826 ( .A(n3436), .ZN(n3437) );
  NOR2_X1 U3827 ( .A1(n5852), .A2(n5906), .ZN(n4842) );
  OR2_X1 U3828 ( .A1(n5852), .A2(n4759), .ZN(n4683) );
  INV_X1 U3829 ( .A(n5906), .ZN(n4759) );
  AND2_X1 U3830 ( .A1(n5852), .A2(n4755), .ZN(n5861) );
  INV_X1 U3831 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7026) );
  OR2_X1 U3832 ( .A1(n6722), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4092) );
  AND2_X1 U3833 ( .A1(n5183), .A2(n4367), .ZN(n5133) );
  OR3_X1 U3834 ( .A1(n6738), .A2(n6465), .A3(n4344), .ZN(n5293) );
  CLKBUF_X1 U3835 ( .A(n4127), .Z(n5043) );
  OR2_X1 U3836 ( .A1(n4525), .A2(n4426), .ZN(n4465) );
  OR2_X1 U3837 ( .A1(n3952), .A2(n5457), .ZN(n3944) );
  OR2_X1 U3838 ( .A1(n3954), .A2(n5116), .ZN(n3952) );
  NAND2_X1 U3839 ( .A1(n3963), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3954)
         );
  AND2_X1 U3840 ( .A1(n4000), .A2(n3999), .ZN(n5153) );
  NOR2_X1 U3841 ( .A1(n5213), .A2(n5152), .ZN(n5166) );
  INV_X1 U3842 ( .A(n4017), .ZN(n3942) );
  OR2_X1 U3843 ( .A1(n4032), .A2(n7007), .ZN(n4034) );
  OR2_X1 U3844 ( .A1(n5213), .A2(n5199), .ZN(n5197) );
  NAND2_X1 U3845 ( .A1(n3874), .A2(n3873), .ZN(n4015) );
  NAND2_X1 U3846 ( .A1(n3868), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3872)
         );
  CLKBUF_X1 U3847 ( .A(n5212), .Z(n5232) );
  AND3_X1 U3848 ( .A1(n3855), .A2(n3854), .A3(n3853), .ZN(n5248) );
  CLKBUF_X1 U3849 ( .A(n5228), .Z(n5229) );
  NAND2_X1 U3850 ( .A1(n3825), .A2(n3824), .ZN(n5354) );
  INV_X1 U3851 ( .A(n4990), .ZN(n3825) );
  AND3_X1 U3852 ( .A1(n3838), .A2(n3837), .A3(n3836), .ZN(n5355) );
  NAND2_X1 U3853 ( .A1(n3805), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3806)
         );
  NOR2_X2 U3854 ( .A1(n6959), .A2(n3806), .ZN(n3852) );
  CLKBUF_X1 U3855 ( .A(n4990), .Z(n5362) );
  NAND2_X1 U3856 ( .A1(n3745), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3791)
         );
  CLKBUF_X1 U3857 ( .A(n5260), .Z(n5261) );
  NAND2_X1 U3858 ( .A1(n3771), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3785)
         );
  AND2_X1 U3859 ( .A1(n3726), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3771)
         );
  AND2_X1 U3861 ( .A1(n3703), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3726)
         );
  INV_X1 U3862 ( .A(n3696), .ZN(n3697) );
  NAND2_X1 U3863 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3697), .ZN(n3713)
         );
  NAND2_X1 U3864 ( .A1(n3702), .A2(n3701), .ZN(n4617) );
  NAND2_X1 U3865 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3696) );
  NAND2_X1 U3866 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5653) );
  BUF_X1 U3867 ( .A(n5068), .Z(n5084) );
  OAI21_X1 U3868 ( .B1(n5519), .B2(n3603), .A(n5532), .ZN(n3607) );
  NAND2_X1 U3869 ( .A1(n5462), .A2(n5461), .ZN(n5460) );
  BUF_X1 U3870 ( .A(n5099), .Z(n5129) );
  AND2_X1 U3871 ( .A1(n5532), .A2(n5743), .ZN(n5466) );
  OR3_X1 U3872 ( .A1(n5532), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5536) );
  CLKBUF_X1 U3873 ( .A(n5184), .Z(n5218) );
  INV_X1 U3874 ( .A(n5238), .ZN(n4196) );
  AND2_X1 U3875 ( .A1(n5532), .A2(n5788), .ZN(n5530) );
  AND2_X1 U3876 ( .A1(n4982), .A2(n5359), .ZN(n4187) );
  AND2_X1 U3877 ( .A1(n5597), .A2(n3588), .ZN(n3589) );
  NAND2_X1 U3878 ( .A1(n6495), .A2(n4984), .ZN(n5795) );
  OR2_X1 U3879 ( .A1(n5532), .A2(n5807), .ZN(n5597) );
  CLKBUF_X1 U3880 ( .A(n5600), .Z(n5619) );
  AND2_X1 U3881 ( .A1(n4167), .A2(n4166), .ZN(n4792) );
  OR2_X1 U3882 ( .A1(n4453), .A2(n4259), .ZN(n4556) );
  INV_X1 U3883 ( .A(n4672), .ZN(n4162) );
  INV_X1 U3884 ( .A(n4534), .ZN(n4152) );
  INV_X1 U3885 ( .A(n3286), .ZN(n3278) );
  INV_X1 U3886 ( .A(n3504), .ZN(n3501) );
  CLKBUF_X1 U3887 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4568) );
  INV_X1 U3888 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4566) );
  OR2_X1 U3889 ( .A1(n5848), .A2(n4799), .ZN(n5992) );
  INV_X1 U3890 ( .A(n4683), .ZN(n4696) );
  OR2_X1 U3891 ( .A1(n5846), .A2(n5998), .ZN(n4695) );
  AND4_X1 U3892 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3230)
         );
  AND4_X1 U3893 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n3232)
         );
  OR2_X1 U3894 ( .A1(n5840), .A2(n6864), .ZN(n4725) );
  AND2_X1 U3895 ( .A1(n5861), .A2(n5906), .ZN(n6179) );
  AND2_X1 U3896 ( .A1(n4599), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4503) );
  INV_X1 U3897 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5282) );
  INV_X1 U3898 ( .A(n6363), .ZN(n6348) );
  AND2_X1 U3899 ( .A1(n5293), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6363) );
  INV_X1 U3900 ( .A(n6346), .ZN(n6362) );
  INV_X1 U3901 ( .A(n6366), .ZN(n6335) );
  INV_X1 U3902 ( .A(n5236), .ZN(n5326) );
  NAND2_X1 U3903 ( .A1(n4237), .A2(n4236), .ZN(n4238) );
  NAND2_X1 U3904 ( .A1(n5058), .A2(n4350), .ZN(n4236) );
  OR2_X1 U3905 ( .A1(n5058), .A2(n3131), .ZN(n4237) );
  OAI211_X2 U3906 ( .C1(n4525), .C2(n4555), .A(n4524), .B(n7065), .ZN(n5436)
         );
  INV_X2 U3907 ( .A(n6385), .ZN(n5438) );
  NAND2_X1 U3908 ( .A1(n4345), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4347)
         );
  INV_X2 U3909 ( .A(n6178), .ZN(n6472) );
  CLKBUF_X1 U3910 ( .A(n5519), .Z(n5520) );
  INV_X1 U3911 ( .A(n5796), .ZN(n6496) );
  CLKBUF_X1 U3912 ( .A(n4435), .Z(n4436) );
  OR2_X1 U3913 ( .A1(n4420), .A2(n6864), .ZN(n6712) );
  INV_X1 U3914 ( .A(n5899), .ZN(n4829) );
  AND2_X1 U3915 ( .A1(n4905), .A2(n4904), .ZN(n4930) );
  NOR2_X1 U3916 ( .A1(n5912), .A2(n5956), .ZN(n5958) );
  OR3_X1 U3917 ( .A1(n6538), .A2(n6537), .A3(n6536), .ZN(n6572) );
  OR2_X1 U3918 ( .A1(n5907), .A2(n4650), .ZN(n6596) );
  INV_X1 U3919 ( .A(n6602), .ZN(n6534) );
  INV_X1 U3920 ( .A(n5994), .ZN(n6026) );
  OAI211_X1 U3921 ( .C1(n6040), .C2(n6039), .A(n6123), .B(n6038), .ZN(n6062)
         );
  INV_X1 U3922 ( .A(n6092), .ZN(n6606) );
  INV_X1 U3923 ( .A(n6108), .ZN(n6627) );
  OAI211_X1 U3924 ( .C1(n6186), .C2(n6073), .A(n4758), .B(n6182), .ZN(n4782)
         );
  INV_X1 U3925 ( .A(n6088), .ZN(n6578) );
  NAND2_X1 U3926 ( .A1(n6179), .A2(n5956), .ZN(n6223) );
  OAI21_X1 U3927 ( .B1(n5019), .B2(n6178), .A(n4398), .ZN(n4399) );
  NAND2_X1 U3928 ( .A1(n5651), .A2(n6474), .ZN(n4101) );
  AOI21_X1 U3929 ( .B1(n5333), .B2(n6518), .A(n5007), .ZN(n5011) );
  AND2_X1 U3930 ( .A1(n4283), .A2(n3138), .ZN(n4284) );
  AND2_X1 U3931 ( .A1(n4389), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4390)
         );
  AOI21_X1 U3932 ( .B1(n3388), .B2(n4568), .A(n3393), .ZN(n3416) );
  NAND2_X2 U3933 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  OR2_X2 U3934 ( .A1(n5722), .A2(n5469), .ZN(n3132) );
  AND2_X1 U3935 ( .A1(n3675), .A2(n4137), .ZN(n3133) );
  AND2_X1 U3936 ( .A1(n3462), .A2(n3461), .ZN(n3134) );
  AND2_X2 U3937 ( .A1(n3674), .A2(n3213), .ZN(n3310) );
  AND2_X1 U3938 ( .A1(n4508), .A2(n4507), .ZN(n5373) );
  AND2_X1 U3939 ( .A1(n5128), .A2(n5143), .ZN(n3135) );
  INV_X1 U3940 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3635) );
  INV_X1 U3941 ( .A(n4991), .ZN(n3824) );
  OAI21_X1 U3942 ( .B1(n4467), .B2(n6868), .A(n4466), .ZN(n6462) );
  INV_X1 U3943 ( .A(n3573), .ZN(n3597) );
  AND4_X1 U3944 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n3136)
         );
  NOR2_X1 U3945 ( .A1(n4391), .A2(n4390), .ZN(n3137) );
  OR2_X1 U3946 ( .A1(n5008), .A2(n4103), .ZN(n3138) );
  AND3_X1 U3947 ( .A1(n3176), .A2(n3175), .A3(n3174), .ZN(n3139) );
  NOR2_X1 U3948 ( .A1(n5848), .A2(n4436), .ZN(n3140) );
  OR2_X1 U3949 ( .A1(n3597), .A2(n4224), .ZN(n3141) );
  NAND2_X1 U3950 ( .A1(n5531), .A2(n3599), .ZN(n3142) );
  AND2_X1 U3952 ( .A1(n5587), .A2(n5579), .ZN(n3143) );
  NOR2_X1 U3953 ( .A1(n4512), .A2(n6782), .ZN(n4337) );
  AND2_X1 U3954 ( .A1(n3329), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3144) );
  XOR2_X1 U3955 ( .A(n5003), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .Z(n3145) );
  AND2_X1 U3956 ( .A1(n5293), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3146) );
  INV_X1 U3957 ( .A(n4110), .ZN(n3627) );
  NAND2_X1 U3958 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  NAND2_X1 U3959 ( .A1(n3630), .A2(n3629), .ZN(n3634) );
  NAND2_X1 U3960 ( .A1(n3634), .A2(n3633), .ZN(n3645) );
  AOI22_X1 U3961 ( .A1(n3442), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3175) );
  AND2_X1 U3962 ( .A1(n3574), .A2(n5604), .ZN(n3580) );
  OR2_X1 U3963 ( .A1(n3407), .A2(n3406), .ZN(n3409) );
  NAND2_X1 U3964 ( .A1(n4504), .A2(n5169), .ZN(n3299) );
  OAI21_X1 U3965 ( .B1(n3494), .B2(n4647), .A(n3503), .ZN(n3495) );
  AND2_X1 U3966 ( .A1(n6072), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3618)
         );
  AOI22_X1 U3967 ( .A1(n3429), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U3968 ( .A1(n3396), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3160) );
  OR2_X1 U3969 ( .A1(n3498), .A2(n4647), .ZN(n3570) );
  AND4_X1 U3970 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3178)
         );
  AND2_X2 U3971 ( .A1(n3180), .A2(n3312), .ZN(n3315) );
  INV_X1 U3972 ( .A(n4034), .ZN(n3943) );
  BUF_X1 U3973 ( .A(n4289), .Z(n4319) );
  OR2_X1 U3974 ( .A1(n3665), .A2(n3664), .ZN(n3667) );
  INV_X1 U3975 ( .A(n5473), .ZN(n3601) );
  OR2_X1 U3976 ( .A1(n3584), .A2(n3583), .ZN(n3585) );
  BUF_X1 U3977 ( .A(n3384), .Z(n3385) );
  OR2_X1 U3978 ( .A1(n4147), .A2(EBX_REG_1__SCAN_IN), .ZN(n4140) );
  AND2_X1 U3979 ( .A1(n3235), .A2(n3234), .ZN(n3236) );
  NAND2_X1 U3980 ( .A1(n3329), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U3981 ( .A1(n3943), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3969)
         );
  INV_X1 U3982 ( .A(n3872), .ZN(n3874) );
  INV_X1 U3983 ( .A(n4337), .ZN(n3687) );
  OR2_X1 U3984 ( .A1(n3460), .A2(n3459), .ZN(n3559) );
  OR2_X1 U3985 ( .A1(n3318), .A2(n4147), .ZN(n4437) );
  NAND2_X1 U3986 ( .A1(n3502), .A2(n3501), .ZN(n3506) );
  AND2_X1 U3987 ( .A1(n5133), .A2(n5098), .ZN(n5087) );
  AND2_X1 U3988 ( .A1(n6329), .A2(n4365), .ZN(n5237) );
  INV_X1 U3989 ( .A(n5240), .ZN(n4195) );
  AND2_X1 U3990 ( .A1(n5079), .A2(n5078), .ZN(n4051) );
  INV_X1 U3991 ( .A(n3963), .ZN(n3971) );
  INV_X1 U3992 ( .A(n3822), .ZN(n3849) );
  NOR2_X1 U3993 ( .A1(n5460), .A2(n5000), .ZN(n5001) );
  INV_X1 U3994 ( .A(n3679), .ZN(n5952) );
  XNOR2_X1 U3995 ( .A(n3488), .B(n4755), .ZN(n3695) );
  INV_X1 U3996 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6072) );
  CLKBUF_X1 U3997 ( .A(n3508), .Z(n6740) );
  INV_X1 U3998 ( .A(n6358), .ZN(n6310) );
  INV_X2 U3999 ( .A(n3508), .ZN(n4467) );
  OR2_X1 U4000 ( .A1(n5213), .A2(n5094), .ZN(n5114) );
  NAND2_X1 U4001 ( .A1(n3725), .A2(n3849), .ZN(n3730) );
  INV_X1 U4002 ( .A(n4357), .ZN(n4358) );
  INV_X1 U4003 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4103) );
  OAI21_X1 U4004 ( .B1(n5513), .B2(n5483), .A(n5482), .ZN(n5504) );
  OR2_X1 U4005 ( .A1(n4267), .A2(n4556), .ZN(n5796) );
  INV_X1 U4006 ( .A(n4092), .ZN(n4094) );
  OR2_X1 U4007 ( .A1(n4802), .A2(n5956), .ZN(n5899) );
  INV_X1 U4008 ( .A(n5958), .ZN(n5985) );
  OR2_X1 U4009 ( .A1(n5854), .A2(n5998), .ZN(n4654) );
  NAND2_X1 U4010 ( .A1(n6712), .A2(n4646), .ZN(n4648) );
  OR2_X1 U4012 ( .A1(n4725), .A2(n5386), .ZN(n6632) );
  OR2_X1 U4013 ( .A1(n4551), .A2(n5998), .ZN(n6529) );
  AOI21_X1 U4014 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6072), .A(n5840), .ZN(
        n6182) );
  NAND2_X1 U4015 ( .A1(n4465), .A2(n6230), .ZN(n6738) );
  OR2_X1 U4016 ( .A1(n4380), .A2(n4379), .ZN(n4381) );
  NOR2_X1 U4017 ( .A1(n5204), .A2(n6685), .ZN(n5183) );
  NOR2_X1 U4018 ( .A1(n5039), .A2(n4599), .ZN(n4348) );
  NAND2_X1 U4019 ( .A1(n5026), .A2(n5025), .ZN(n6358) );
  AND2_X1 U4020 ( .A1(n5381), .A2(n4512), .ZN(n6379) );
  AND2_X1 U4021 ( .A1(n6418), .A2(n6735), .ZN(n6413) );
  INV_X1 U4022 ( .A(n6420), .ZN(n7062) );
  AND2_X1 U4023 ( .A1(n5114), .A2(n5113), .ZN(n5480) );
  NOR2_X1 U4024 ( .A1(n5377), .A2(n5378), .ZN(n5376) );
  INV_X1 U4025 ( .A(n5625), .ZN(n6474) );
  OR2_X1 U4026 ( .A1(n5710), .A2(n4280), .ZN(n5697) );
  INV_X1 U4027 ( .A(n6500), .ZN(n6518) );
  INV_X1 U4028 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4599) );
  INV_X1 U4029 ( .A(n6223), .ZN(n5901) );
  OAI211_X1 U4030 ( .C1(n6186), .C2(n5865), .A(n4806), .B(n6182), .ZN(n4830)
         );
  OAI211_X1 U4031 ( .C1(n4902), .C2(n4906), .A(n6123), .B(n6080), .ZN(n4928)
         );
  AND2_X1 U4032 ( .A1(n4684), .A2(n4696), .ZN(n4932) );
  OAI211_X1 U4033 ( .C1(n6186), .C2(n5963), .A(n5962), .B(n6182), .ZN(n5987)
         );
  AND2_X1 U4034 ( .A1(n5957), .A2(n5956), .ZN(n6570) );
  INV_X1 U4035 ( .A(n6596), .ZN(n4879) );
  OAI211_X1 U4036 ( .C1(n6002), .C2(n6001), .A(n6182), .B(n6000), .ZN(n6027)
         );
  NOR2_X1 U4037 ( .A1(n5995), .A2(n6120), .ZN(n6065) );
  AND2_X1 U4038 ( .A1(n3140), .A2(n4551), .ZN(n6039) );
  INV_X1 U4039 ( .A(n6104), .ZN(n6591) );
  OAI21_X1 U4040 ( .B1(n6078), .B2(n6077), .A(n6076), .ZN(n6112) );
  INV_X1 U4041 ( .A(n6069), .ZN(n6117) );
  AND2_X1 U4042 ( .A1(n6179), .A2(n6120), .ZN(n6225) );
  AOI211_X1 U4043 ( .C1(n5134), .C2(REIP_REG_24__SCAN_IN), .A(n5121), .B(n5120), .ZN(n5122) );
  AND2_X1 U4044 ( .A1(n5292), .A2(n6324), .ZN(n6370) );
  INV_X1 U4045 ( .A(n5480), .ZN(n5405) );
  OR2_X1 U4046 ( .A1(n4667), .A2(n4625), .ZN(n6371) );
  INV_X1 U4047 ( .A(n5434), .ZN(n5437) );
  INV_X1 U4048 ( .A(n6394), .ZN(n4496) );
  OR3_X1 U4049 ( .A1(n4525), .A2(n4463), .A3(n4462), .ZN(n6418) );
  INV_X1 U4050 ( .A(n6413), .ZN(n6419) );
  INV_X1 U4051 ( .A(n6462), .ZN(n6420) );
  OR3_X2 U4052 ( .A1(n4525), .A2(n4468), .A3(READY_N), .ZN(n7065) );
  AND2_X1 U4053 ( .A1(n4099), .A2(n4098), .ZN(n4100) );
  OR2_X1 U4054 ( .A1(n4525), .A2(n4597), .ZN(n5625) );
  NAND2_X1 U4055 ( .A1(n5630), .A2(n5647), .ZN(n6478) );
  XNOR2_X1 U4056 ( .A(n4384), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5018)
         );
  INV_X1 U4057 ( .A(n4899), .ZN(n4935) );
  INV_X1 U4058 ( .A(n5905), .ZN(n5947) );
  NAND3_X1 U4059 ( .A1(n4649), .A2(n5906), .A3(n6120), .ZN(n6602) );
  OR2_X1 U4060 ( .A1(n5995), .A2(n5956), .ZN(n5994) );
  AOI21_X1 U4061 ( .B1(n6035), .B2(n6039), .A(n6034), .ZN(n6068) );
  NAND2_X1 U4062 ( .A1(n4697), .A2(n4696), .ZN(n6641) );
  NAND2_X1 U4063 ( .A1(n4689), .A2(n5855), .ZN(n6634) );
  INV_X1 U4064 ( .A(n6121), .ZN(n6171) );
  AOI21_X1 U4065 ( .B1(n6185), .B2(n6184), .A(n6183), .ZN(n6228) );
  OAI21_X1 U4066 ( .B1(n5018), .B2(n6515), .A(n3137), .ZN(U2989) );
  NAND2_X1 U4067 ( .A1(n6864), .A2(n4599), .ZN(n6722) );
  XNOR2_X1 U4068 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6033) );
  OAI22_X1 U4069 ( .A1(n4092), .A2(n6033), .B1(n4503), .B2(n4756), .ZN(n3301)
         );
  INV_X2 U4070 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4577) );
  AND2_X4 U4071 ( .A1(n4577), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4441)
         );
  INV_X1 U4072 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3147) );
  AND2_X4 U4073 ( .A1(n3147), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4554)
         );
  AND2_X4 U4074 ( .A1(n4441), .A2(n4554), .ZN(n4288) );
  INV_X1 U4075 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3148) );
  AND2_X4 U4076 ( .A1(n3148), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4552)
         );
  AND2_X4 U4077 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4553) );
  AOI22_X1 U4078 ( .A1(n4288), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3152) );
  NOR2_X4 U4079 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4630) );
  AND2_X2 U4080 ( .A1(n4552), .A2(n4630), .ZN(n3323) );
  AND2_X2 U4081 ( .A1(n4554), .A2(n4630), .ZN(n3324) );
  AND2_X4 U4082 ( .A1(n4441), .A2(n4552), .ZN(n3358) );
  AND2_X4 U4083 ( .A1(n4441), .A2(n4601), .ZN(n3255) );
  NOR2_X4 U4084 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4085 ( .A1(n3329), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3149) );
  AND2_X4 U4086 ( .A1(n4441), .A2(n3154), .ZN(n3442) );
  INV_X1 U4087 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3153) );
  AND2_X4 U4090 ( .A1(n4630), .A2(n4601), .ZN(n3359) );
  AOI22_X1 U4091 ( .A1(n3338), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3359), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3157) );
  AND2_X4 U4092 ( .A1(n3154), .A2(n4553), .ZN(n3367) );
  AND2_X4 U4093 ( .A1(n4554), .A2(n4553), .ZN(n3401) );
  NAND2_X2 U4094 ( .A1(n3159), .A2(n3089), .ZN(n4502) );
  INV_X1 U4095 ( .A(n4502), .ZN(n3677) );
  AOI22_X1 U4096 ( .A1(n4288), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4097 ( .A1(n3255), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4098 ( .A1(n3358), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4099 ( .A1(n3338), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3359), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4100 ( .A1(n3401), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4101 ( .A1(n3442), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3164) );
  NAND2_X2 U4102 ( .A1(n3169), .A2(n3168), .ZN(n3312) );
  AOI22_X1 U4103 ( .A1(n3255), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4104 ( .A1(n3323), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4105 ( .A1(n3365), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4106 ( .A1(n3358), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4107 ( .A1(n3338), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3359), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4108 ( .A1(n3357), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3174) );
  OAI21_X1 U4109 ( .B1(n3677), .B2(n3312), .A(n3284), .ZN(n3179) );
  INV_X1 U4110 ( .A(n3179), .ZN(n3291) );
  NAND2_X1 U4111 ( .A1(n3323), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U4112 ( .A1(n3324), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U4113 ( .A1(n3358), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3181) );
  NAND3_X1 U4114 ( .A1(n3183), .A2(n3182), .A3(n3181), .ZN(n3184) );
  NAND2_X1 U4115 ( .A1(n3442), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3188) );
  NAND2_X1 U4116 ( .A1(n3255), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3187)
         );
  NAND2_X1 U4117 ( .A1(n3396), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U4118 ( .A1(n3365), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3185)
         );
  NAND2_X1 U4119 ( .A1(n3357), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U4120 ( .A1(n3429), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U4121 ( .A1(n3338), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U4122 ( .A1(n3359), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3189)
         );
  NAND2_X1 U4123 ( .A1(n4288), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U4124 ( .A1(n3401), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3195)
         );
  NAND2_X1 U4125 ( .A1(n3339), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3194)
         );
  NAND2_X1 U4126 ( .A1(n3367), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U4127 ( .A1(n3315), .A2(n3290), .ZN(n3201) );
  AOI22_X1 U4128 ( .A1(n3255), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4129 ( .A1(n3442), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4130 ( .A1(n3429), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3203) );
  AOI22_X1 U4131 ( .A1(n3365), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3202) );
  NAND4_X1 U4132 ( .A1(n3205), .A2(n3204), .A3(n3203), .A4(n3202), .ZN(n3211)
         );
  AOI22_X1 U4133 ( .A1(n3358), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4134 ( .A1(n4288), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3208) );
  AOI22_X1 U4135 ( .A1(n3396), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3359), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U4136 ( .A1(n3357), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3206) );
  NAND4_X1 U4137 ( .A1(n3209), .A2(n3208), .A3(n3207), .A4(n3206), .ZN(n3210)
         );
  OAI21_X1 U4138 ( .B1(n3315), .B2(n3290), .A(n4137), .ZN(n3212) );
  INV_X1 U4139 ( .A(n3212), .ZN(n3213) );
  INV_X1 U4140 ( .A(n3312), .ZN(n3294) );
  NAND2_X1 U4141 ( .A1(n3358), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4142 ( .A1(n3255), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3216)
         );
  NAND2_X1 U4143 ( .A1(n3323), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4144 ( .A1(n3324), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4145 ( .A1(n4288), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3221)
         );
  NAND2_X1 U4146 ( .A1(n3396), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U4147 ( .A1(n3339), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3219)
         );
  NAND2_X1 U4148 ( .A1(n3329), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4149 ( .A1(n3429), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4150 ( .A1(n3357), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4151 ( .A1(n3401), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3223)
         );
  NAND2_X1 U4152 ( .A1(n3367), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4153 ( .A1(n3442), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4154 ( .A1(n3365), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3228)
         );
  NAND2_X1 U4155 ( .A1(n3338), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4156 ( .A1(n3359), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3226)
         );
  NAND2_X1 U4157 ( .A1(n4288), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3237)
         );
  NAND2_X1 U4158 ( .A1(n3091), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4159 ( .A1(n3339), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3234)
         );
  NAND2_X1 U4160 ( .A1(n3358), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U4161 ( .A1(n3255), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3241)
         );
  NAND2_X1 U4162 ( .A1(n3323), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4163 ( .A1(n3324), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4164 ( .A1(n3429), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4165 ( .A1(n3357), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3245) );
  NAND2_X1 U4166 ( .A1(n3401), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3244)
         );
  NAND2_X1 U4167 ( .A1(n3367), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3243) );
  NAND2_X1 U4168 ( .A1(n3442), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U4169 ( .A1(n3365), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3249)
         );
  NAND2_X1 U4170 ( .A1(n3338), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3248) );
  NAND2_X1 U4171 ( .A1(n3359), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3247)
         );
  AND4_X4 U4172 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n4657)
         );
  NAND2_X1 U4173 ( .A1(n3358), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3259) );
  NAND2_X1 U4174 ( .A1(n3255), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3258)
         );
  NAND2_X1 U4175 ( .A1(n4288), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3257)
         );
  NAND2_X1 U4176 ( .A1(n3323), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3256) );
  NAND2_X1 U4178 ( .A1(n3429), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3263) );
  NAND2_X1 U4179 ( .A1(n3338), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3262) );
  NAND2_X1 U4180 ( .A1(n3357), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4181 ( .A1(n3401), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3260)
         );
  NAND2_X1 U4183 ( .A1(n3442), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3267) );
  NAND2_X1 U4184 ( .A1(n3365), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3266)
         );
  NAND2_X1 U4185 ( .A1(n3367), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3265) );
  NAND2_X1 U4186 ( .A1(n3359), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3264)
         );
  NAND2_X1 U4188 ( .A1(n3396), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4189 ( .A1(n3324), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U4190 ( .A1(n3329), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4191 ( .A1(n3339), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3268)
         );
  XNOR2_X1 U4194 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4105) );
  NAND2_X1 U4195 ( .A1(n3292), .A2(n4105), .ZN(n3295) );
  AND2_X1 U4196 ( .A1(n3337), .A2(n3295), .ZN(n3281) );
  NAND2_X1 U4197 ( .A1(n3290), .A2(n3312), .ZN(n3318) );
  INV_X1 U4198 ( .A(n3318), .ZN(n3276) );
  INV_X1 U4199 ( .A(n4137), .ZN(n4661) );
  NAND2_X1 U4200 ( .A1(n4661), .A2(n4657), .ZN(n3317) );
  NAND2_X1 U4201 ( .A1(n3292), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3279) );
  NOR2_X1 U4202 ( .A1(n4421), .A2(n4137), .ZN(n3277) );
  NAND2_X1 U4203 ( .A1(n3278), .A2(n3277), .ZN(n4240) );
  INV_X2 U4204 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n4647) );
  AOI21_X2 U4206 ( .B1(n4126), .B2(n3281), .A(n3280), .ZN(n3304) );
  INV_X1 U4207 ( .A(n3304), .ZN(n3282) );
  OAI21_X1 U4208 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3301), .A(n3282), 
        .ZN(n3305) );
  NAND4_X1 U4209 ( .A1(n4239), .A2(n4724), .A3(n3677), .A4(n3284), .ZN(n3856)
         );
  NAND4_X1 U4210 ( .A1(n3286), .A2(n3285), .A3(n4657), .A4(n3856), .ZN(n3289)
         );
  NAND2_X1 U4211 ( .A1(n4657), .A2(n4137), .ZN(n3509) );
  NAND2_X1 U4212 ( .A1(n4657), .A2(n4254), .ZN(n5297) );
  OAI21_X1 U4213 ( .B1(n3315), .B2(n3509), .A(n5297), .ZN(n3287) );
  INV_X1 U4214 ( .A(n3287), .ZN(n3288) );
  NAND2_X1 U4215 ( .A1(n3291), .A2(n4685), .ZN(n4118) );
  NAND2_X1 U4216 ( .A1(n4118), .A2(n4467), .ZN(n3297) );
  AOI21_X1 U4217 ( .B1(n4698), .B2(n3295), .A(n4256), .ZN(n3296) );
  NAND4_X1 U4218 ( .A1(n3311), .A2(n3310), .A3(n3297), .A4(n3296), .ZN(n3298)
         );
  NAND2_X1 U4219 ( .A1(n3298), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3300) );
  NAND2_X1 U4220 ( .A1(n3300), .A2(n3299), .ZN(n3387) );
  NAND2_X1 U4221 ( .A1(n3387), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3303) );
  INV_X1 U4222 ( .A(n3301), .ZN(n3302) );
  NAND3_X1 U4223 ( .A1(n3304), .A2(n3303), .A3(n3302), .ZN(n3384) );
  NAND2_X1 U4224 ( .A1(n3305), .A2(n3384), .ZN(n3382) );
  NAND2_X1 U4225 ( .A1(n3387), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3309) );
  INV_X1 U4226 ( .A(n4503), .ZN(n3306) );
  MUX2_X1 U4227 ( .A(n3306), .B(n4094), .S(n6072), .Z(n3307) );
  INV_X1 U4228 ( .A(n3307), .ZN(n3308) );
  INV_X1 U4229 ( .A(n3311), .ZN(n3314) );
  NAND2_X1 U4230 ( .A1(n4119), .A2(n4685), .ZN(n4251) );
  NOR2_X1 U4231 ( .A1(n4657), .A2(n4724), .ZN(n3313) );
  INV_X1 U4232 ( .A(n4118), .ZN(n3316) );
  INV_X1 U4233 ( .A(n4115), .ZN(n3675) );
  NAND2_X1 U4234 ( .A1(n3316), .A2(n3133), .ZN(n3321) );
  OR2_X1 U4235 ( .A1(n3856), .A2(n3317), .ZN(n4569) );
  OR2_X1 U4236 ( .A1(n6722), .A2(n4647), .ZN(n6647) );
  INV_X1 U4237 ( .A(n6647), .ZN(n3319) );
  NAND3_X1 U4238 ( .A1(n4569), .A2(n3319), .A3(n4437), .ZN(n3320) );
  AOI21_X1 U4239 ( .B1(n3321), .B2(n4467), .A(n3320), .ZN(n3322) );
  OAI211_X1 U4240 ( .C1(n3292), .C2(n3310), .A(n4250), .B(n3322), .ZN(n3354)
         );
  XNOR2_X2 U4241 ( .A(n3382), .B(n3383), .ZN(n4435) );
  AOI22_X1 U4243 ( .A1(n4312), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4244 ( .A1(n4313), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4245 ( .A1(n3095), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4246 ( .A1(n4314), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3325) );
  NAND4_X1 U4247 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3335)
         );
  BUF_X1 U4248 ( .A(n3255), .Z(n3395) );
  AOI22_X1 U4249 ( .A1(n4311), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4250 ( .A1(n3467), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4251 ( .A1(n4291), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4252 ( .A1(n4296), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3330) );
  NAND4_X1 U4253 ( .A1(n3333), .A2(n3332), .A3(n3331), .A4(n3330), .ZN(n3334)
         );
  NAND2_X1 U4254 ( .A1(n4504), .A2(n3518), .ZN(n3336) );
  OAI21_X4 U4255 ( .B1(n4435), .B2(STATE2_REG_0__SCAN_IN), .A(n3336), .ZN(
        n3515) );
  INV_X1 U4256 ( .A(n3518), .ZN(n3353) );
  NAND2_X1 U4257 ( .A1(n4657), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3424) );
  NAND2_X1 U4258 ( .A1(n3638), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4259 ( .A1(n3358), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3323), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4260 ( .A1(n4313), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4261 ( .A1(n4069), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4262 ( .A1(n4291), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3340) );
  NAND4_X1 U4263 ( .A1(n3343), .A2(n3342), .A3(n3341), .A4(n3340), .ZN(n3350)
         );
  AOI22_X1 U4264 ( .A1(n3395), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4289), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4265 ( .A1(n3096), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4266 ( .A1(n3095), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4267 ( .A1(n3344), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3345) );
  NAND4_X1 U4268 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n3345), .ZN(n3349)
         );
  INV_X1 U4269 ( .A(n3575), .ZN(n3351) );
  NAND2_X1 U4270 ( .A1(n4504), .A2(n3351), .ZN(n3492) );
  NAND2_X1 U4271 ( .A1(n3515), .A2(n3514), .ZN(n3377) );
  AOI22_X1 U4272 ( .A1(n3467), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4273 ( .A1(n3344), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4274 ( .A1(n3358), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4289), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4275 ( .A1(n3360), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3361) );
  NAND4_X1 U4276 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3373)
         );
  AOI22_X1 U4277 ( .A1(n3395), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4312), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4278 ( .A1(n4313), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4279 ( .A1(n4291), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4280 ( .A1(n4069), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3368) );
  NAND4_X1 U4281 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  NAND2_X1 U4282 ( .A1(n4657), .A2(n3519), .ZN(n3497) );
  NAND2_X1 U4283 ( .A1(n4685), .A2(n3575), .ZN(n3498) );
  OAI21_X1 U4284 ( .B1(n3423), .B2(n3497), .A(n3570), .ZN(n3374) );
  INV_X1 U4285 ( .A(n3374), .ZN(n3375) );
  INV_X1 U4286 ( .A(n3376), .ZN(n3516) );
  NAND2_X1 U4287 ( .A1(n3377), .A2(n3516), .ZN(n3381) );
  INV_X1 U4288 ( .A(n3515), .ZN(n3379) );
  INV_X1 U4289 ( .A(n3514), .ZN(n3378) );
  NAND2_X1 U4290 ( .A1(n3379), .A2(n3378), .ZN(n3380) );
  NAND2_X1 U4291 ( .A1(n3381), .A2(n3380), .ZN(n3527) );
  INV_X1 U4292 ( .A(n3527), .ZN(n3414) );
  NAND2_X1 U4293 ( .A1(n3104), .A2(n3112), .ZN(n3386) );
  NAND2_X1 U4294 ( .A1(n3386), .A2(n3385), .ZN(n3415) );
  AND2_X1 U4296 ( .A1(n7026), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6784)
         );
  NAND2_X1 U4297 ( .A1(n6784), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4298 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3389) );
  NAND2_X1 U4299 ( .A1(n3389), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4300 ( .A1(n3391), .A2(n3390), .ZN(n4850) );
  NAND2_X1 U4301 ( .A1(n4094), .A2(n4850), .ZN(n3392) );
  OAI21_X1 U4302 ( .B1(n4503), .B2(n7026), .A(n3392), .ZN(n3393) );
  INV_X1 U4303 ( .A(n3416), .ZN(n3394) );
  AOI22_X1 U4304 ( .A1(n4311), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4305 ( .A1(n4313), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4306 ( .A1(n4290), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3398) );
  INV_X1 U4307 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6850) );
  AOI22_X1 U4308 ( .A1(n4291), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3397) );
  NAND4_X1 U4309 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3407)
         );
  AOI22_X1 U4310 ( .A1(n3467), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3405) );
  BUF_X1 U4311 ( .A(n3401), .Z(n4069) );
  AOI22_X1 U4312 ( .A1(n3095), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4313 ( .A1(n3360), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4314 ( .A1(n4314), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3402) );
  NAND4_X1 U4315 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3406)
         );
  NAND2_X1 U4316 ( .A1(n3638), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3408) );
  OAI21_X1 U4317 ( .B1(n3532), .B2(n3424), .A(n3408), .ZN(n3411) );
  NAND2_X1 U4318 ( .A1(n4504), .A2(n3409), .ZN(n3410) );
  XNOR2_X1 U4319 ( .A(n3411), .B(n3410), .ZN(n3412) );
  NAND2_X1 U4320 ( .A1(n3414), .A2(n3528), .ZN(n3488) );
  INV_X1 U4321 ( .A(n3415), .ZN(n3417) );
  NAND2_X1 U4322 ( .A1(n3388), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3422) );
  NAND3_X1 U4323 ( .A1(n6535), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6530) );
  INV_X1 U4324 ( .A(n6530), .ZN(n3418) );
  NAND2_X1 U4325 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3418), .ZN(n6595) );
  NAND2_X1 U4326 ( .A1(n6535), .A2(n6595), .ZN(n3419) );
  NAND3_X1 U4327 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6125) );
  INV_X1 U4328 ( .A(n6125), .ZN(n6188) );
  NAND2_X1 U4329 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6188), .ZN(n6191) );
  NAND2_X1 U4330 ( .A1(n3419), .A2(n6191), .ZN(n6079) );
  OAI22_X1 U4331 ( .A1(n4092), .A2(n6079), .B1(n4503), .B2(n6535), .ZN(n3420)
         );
  INV_X1 U4332 ( .A(n3420), .ZN(n3421) );
  NAND2_X2 U4333 ( .A1(n3424), .A2(n3423), .ZN(n3671) );
  AOI22_X1 U4334 ( .A1(n4311), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4335 ( .A1(n3467), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4336 ( .A1(n3401), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4337 ( .A1(n4291), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3425) );
  NAND4_X1 U4338 ( .A1(n3428), .A2(n3427), .A3(n3426), .A4(n3425), .ZN(n3435)
         );
  AOI22_X1 U4339 ( .A1(n3395), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4312), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4340 ( .A1(n4313), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4341 ( .A1(n3095), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4342 ( .A1(n4314), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3430) );
  NAND4_X1 U4343 ( .A1(n3433), .A2(n3432), .A3(n3431), .A4(n3430), .ZN(n3434)
         );
  AOI22_X1 U4344 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n3638), .B1(n3671), 
        .B2(n3489), .ZN(n3436) );
  AOI21_X2 U4345 ( .B1(n4550), .B2(n4647), .A(n3437), .ZN(n4640) );
  NOR2_X2 U4346 ( .A1(n3488), .A2(n4640), .ZN(n3541) );
  NAND2_X1 U4347 ( .A1(n3638), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4348 ( .A1(n4311), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4349 ( .A1(n4313), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4350 ( .A1(n4290), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3439) );
  INV_X1 U4351 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n7014) );
  AOI22_X1 U4352 ( .A1(n4291), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3438) );
  NAND4_X1 U4353 ( .A1(n3441), .A2(n3440), .A3(n3439), .A4(n3438), .ZN(n3448)
         );
  AOI22_X1 U4355 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3442), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4356 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3095), .B1(n3401), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4357 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3360), .B1(n3097), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4358 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4314), .B1(n4296), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3443) );
  NAND4_X1 U4359 ( .A1(n3446), .A2(n3445), .A3(n3444), .A4(n3443), .ZN(n3447)
         );
  NAND2_X1 U4360 ( .A1(n3671), .A2(n3545), .ZN(n3449) );
  NAND2_X1 U4361 ( .A1(n3450), .A2(n3449), .ZN(n3543) );
  NAND2_X1 U4362 ( .A1(n3541), .A2(n3543), .ZN(n3554) );
  NAND2_X1 U4363 ( .A1(n3638), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4364 ( .A1(n4311), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4312), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4365 ( .A1(n4313), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4366 ( .A1(n3467), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4367 ( .A1(n4291), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3451) );
  NAND4_X1 U4368 ( .A1(n3454), .A2(n3453), .A3(n3452), .A4(n3451), .ZN(n3460)
         );
  AOI22_X1 U4369 ( .A1(n3395), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4370 ( .A1(n3095), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4371 ( .A1(n4070), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4372 ( .A1(n4314), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3455) );
  NAND4_X1 U4373 ( .A1(n3458), .A2(n3457), .A3(n3456), .A4(n3455), .ZN(n3459)
         );
  NAND2_X1 U4374 ( .A1(n3671), .A2(n3559), .ZN(n3461) );
  NOR2_X2 U4375 ( .A1(n3554), .A2(n3134), .ZN(n3553) );
  NAND2_X1 U4376 ( .A1(n3638), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4377 ( .A1(n4311), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4378 ( .A1(n4313), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3465) );
  INV_X1 U4379 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6799) );
  AOI22_X1 U4380 ( .A1(n4290), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4381 ( .A1(n4291), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4382 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3473)
         );
  AOI22_X1 U4383 ( .A1(n3467), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4384 ( .A1(n3095), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4385 ( .A1(n3360), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4386 ( .A1(n4314), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3468) );
  NAND4_X1 U4387 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3472)
         );
  NAND2_X1 U4388 ( .A1(n3671), .A2(n3484), .ZN(n3474) );
  NAND2_X1 U4389 ( .A1(n3475), .A2(n3474), .ZN(n3476) );
  NAND2_X1 U4390 ( .A1(n3518), .A2(n3519), .ZN(n3531) );
  NAND2_X1 U4391 ( .A1(n3531), .A2(n3532), .ZN(n3530) );
  NAND2_X1 U4392 ( .A1(n3530), .A2(n3489), .ZN(n3546) );
  INV_X1 U4393 ( .A(n3545), .ZN(n3478) );
  NOR2_X1 U4394 ( .A1(n3546), .A2(n3478), .ZN(n3560) );
  NAND2_X1 U4395 ( .A1(n3560), .A2(n3559), .ZN(n3558) );
  XNOR2_X1 U4396 ( .A(n3558), .B(n3484), .ZN(n3479) );
  NAND2_X1 U4397 ( .A1(n3479), .A2(n4467), .ZN(n3480) );
  OAI21_X2 U4398 ( .B1(n3707), .B2(n3092), .A(n3480), .ZN(n3481) );
  INV_X1 U4399 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4164) );
  XNOR2_X1 U4400 ( .A(n3481), .B(n4164), .ZN(n5635) );
  INV_X1 U4401 ( .A(n5635), .ZN(n3482) );
  NAND2_X1 U4402 ( .A1(n3481), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3564)
         );
  NAND2_X1 U4403 ( .A1(n3482), .A2(n3564), .ZN(n5627) );
  AOI22_X1 U4404 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n3638), .B1(n3671), 
        .B2(n3575), .ZN(n3483) );
  INV_X1 U4405 ( .A(n3558), .ZN(n3485) );
  NAND2_X1 U4406 ( .A1(n3485), .A2(n3484), .ZN(n3577) );
  XNOR2_X1 U4407 ( .A(n3577), .B(n3575), .ZN(n3486) );
  NAND2_X1 U4408 ( .A1(n3486), .A2(n4467), .ZN(n3487) );
  OAI21_X2 U4409 ( .B1(n3724), .B2(n3092), .A(n3487), .ZN(n3567) );
  INV_X1 U4410 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5822) );
  XNOR2_X1 U4411 ( .A(n3567), .B(n5822), .ZN(n5626) );
  INV_X1 U4412 ( .A(n4640), .ZN(n4755) );
  NAND2_X1 U4413 ( .A1(n4119), .A2(n3695), .ZN(n3491) );
  OAI211_X1 U4414 ( .C1(n3489), .C2(n3530), .A(n3546), .B(n4467), .ZN(n3490)
         );
  OR2_X1 U4415 ( .A1(n3498), .A2(n3519), .ZN(n3494) );
  INV_X1 U4416 ( .A(n3492), .ZN(n3493) );
  NAND2_X1 U4417 ( .A1(n3493), .A2(n3519), .ZN(n3503) );
  NAND2_X1 U4418 ( .A1(n3638), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3500) );
  AND3_X1 U4419 ( .A1(n3498), .A2(n3497), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3499) );
  NAND2_X1 U4420 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  NAND2_X1 U4421 ( .A1(n3506), .A2(n3505), .ZN(n3678) );
  INV_X1 U4422 ( .A(n3678), .ZN(n3507) );
  NAND2_X1 U4423 ( .A1(n3507), .A2(n4119), .ZN(n3513) );
  CLKBUF_X1 U4424 ( .A(n3509), .Z(n3510) );
  OAI21_X1 U4425 ( .B1(n6740), .B2(n3519), .A(n3510), .ZN(n3511) );
  INV_X1 U4426 ( .A(n3511), .ZN(n3512) );
  NAND2_X1 U4427 ( .A1(n3513), .A2(n3512), .ZN(n5646) );
  NAND2_X1 U4428 ( .A1(n5646), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3525)
         );
  XNOR2_X1 U4429 ( .A(n3525), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4541)
         );
  NAND2_X1 U4430 ( .A1(n4641), .A2(n7068), .ZN(n3524) );
  OAI21_X1 U4431 ( .B1(n3519), .B2(n3518), .A(n3531), .ZN(n3521) );
  NAND2_X1 U4432 ( .A1(n4724), .A2(n4137), .ZN(n4245) );
  INV_X1 U4433 ( .A(n4245), .ZN(n3520) );
  OAI211_X1 U4434 ( .C1(n3521), .C2(n6740), .A(n3520), .B(n5385), .ZN(n3522)
         );
  INV_X1 U4435 ( .A(n3522), .ZN(n3523) );
  NAND2_X1 U4436 ( .A1(n3524), .A2(n3523), .ZN(n4540) );
  NAND2_X1 U4437 ( .A1(n4541), .A2(n4540), .ZN(n4539) );
  INV_X1 U4438 ( .A(n3525), .ZN(n6513) );
  NAND2_X1 U4439 ( .A1(n6513), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3526)
         );
  NAND2_X1 U4440 ( .A1(n4539), .A2(n3526), .ZN(n6470) );
  BUF_X1 U4441 ( .A(n3527), .Z(n3529) );
  XNOR2_X2 U4442 ( .A(n3529), .B(n3528), .ZN(n4639) );
  NAND2_X1 U4443 ( .A1(n4639), .A2(n4119), .ZN(n3536) );
  OAI21_X1 U4444 ( .B1(n3532), .B2(n3531), .A(n3530), .ZN(n3534) );
  INV_X1 U4445 ( .A(n3510), .ZN(n3533) );
  AOI21_X1 U4446 ( .B1(n3534), .B2(n4467), .A(n3533), .ZN(n3535) );
  NAND2_X1 U4447 ( .A1(n3536), .A2(n3535), .ZN(n3537) );
  OR2_X1 U4448 ( .A1(n3537), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6468)
         );
  INV_X1 U4449 ( .A(n3539), .ZN(n3540) );
  INV_X1 U4450 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6837) );
  OAI22_X1 U4451 ( .A1(n4948), .A2(n4949), .B1(n3540), .B2(n6837), .ZN(n4735)
         );
  BUF_X1 U4452 ( .A(n3541), .Z(n3542) );
  INV_X1 U4453 ( .A(n3542), .ZN(n3544) );
  XNOR2_X1 U4454 ( .A(n3544), .B(n3543), .ZN(n3712) );
  NAND2_X1 U4455 ( .A1(n3712), .A2(n4119), .ZN(n3549) );
  XNOR2_X1 U4456 ( .A(n3546), .B(n3545), .ZN(n3547) );
  NAND2_X1 U4457 ( .A1(n3547), .A2(n4467), .ZN(n3548) );
  INV_X1 U4458 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U4459 ( .A1(n4735), .A2(n4737), .ZN(n3552) );
  NAND2_X1 U4460 ( .A1(n3550), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3551)
         );
  NAND2_X1 U4461 ( .A1(n3552), .A2(n3551), .ZN(n4882) );
  INV_X1 U4462 ( .A(n3553), .ZN(n3556) );
  NAND2_X1 U4463 ( .A1(n3554), .A2(n3134), .ZN(n3555) );
  NAND2_X1 U4464 ( .A1(n3556), .A2(n3555), .ZN(n3711) );
  INV_X1 U4465 ( .A(n3711), .ZN(n3557) );
  NAND2_X1 U4466 ( .A1(n3557), .A2(n4119), .ZN(n3562) );
  OAI211_X1 U4467 ( .C1(n3560), .C2(n3559), .A(n3558), .B(n4467), .ZN(n3561)
         );
  NAND2_X1 U4468 ( .A1(n3562), .A2(n3561), .ZN(n3563) );
  INV_X1 U4469 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4893) );
  XNOR2_X1 U4470 ( .A(n3563), .B(n4893), .ZN(n4883) );
  NAND2_X1 U4471 ( .A1(n4882), .A2(n4883), .ZN(n5637) );
  NAND2_X1 U4472 ( .A1(n3563), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5638)
         );
  AND2_X1 U4473 ( .A1(n5638), .A2(n3564), .ZN(n3565) );
  NAND2_X1 U4474 ( .A1(n5637), .A2(n3565), .ZN(n5628) );
  NAND2_X1 U4475 ( .A1(n3566), .A2(n5628), .ZN(n3569) );
  NAND2_X1 U4476 ( .A1(n3098), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3568)
         );
  NAND2_X1 U4477 ( .A1(n3569), .A2(n3568), .ZN(n5600) );
  NOR2_X1 U4478 ( .A1(n3570), .A2(n3092), .ZN(n3571) );
  INV_X1 U4479 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5807) );
  AND2_X1 U4480 ( .A1(n3573), .A2(n5807), .ZN(n5598) );
  INV_X1 U4481 ( .A(n5598), .ZN(n3574) );
  INV_X1 U4482 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U4483 ( .A1(n3573), .A2(n5808), .ZN(n5604) );
  NAND2_X1 U4484 ( .A1(n4467), .A2(n3575), .ZN(n3576) );
  OR2_X1 U4485 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  NAND2_X1 U4486 ( .A1(n3573), .A2(n3578), .ZN(n3581) );
  INV_X1 U4487 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5815) );
  XNOR2_X1 U4488 ( .A(n3581), .B(n5815), .ZN(n5620) );
  AND2_X1 U4489 ( .A1(n3580), .A2(n5620), .ZN(n3579) );
  NAND2_X1 U4490 ( .A1(n5600), .A2(n3579), .ZN(n3586) );
  INV_X1 U4491 ( .A(n3580), .ZN(n3584) );
  NAND2_X1 U4492 ( .A1(n3581), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5601)
         );
  INV_X1 U4493 ( .A(n5601), .ZN(n3582) );
  NOR2_X1 U4494 ( .A1(n3573), .A2(n5808), .ZN(n5603) );
  NOR2_X1 U4495 ( .A1(n3582), .A2(n5603), .ZN(n3583) );
  NAND2_X1 U4496 ( .A1(n3586), .A2(n3585), .ZN(n5577) );
  INV_X1 U4497 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U4498 ( .A1(n5532), .A2(n6486), .ZN(n5587) );
  CLKBUF_X3 U4499 ( .A(n3573), .Z(n5532) );
  INV_X1 U4500 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U4501 ( .A1(n5532), .A2(n5580), .ZN(n5579) );
  NAND2_X1 U4502 ( .A1(n5577), .A2(n3143), .ZN(n3590) );
  NOR2_X1 U4503 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3587) );
  OR2_X1 U4504 ( .A1(n5532), .A2(n3587), .ZN(n3588) );
  NAND2_X1 U4505 ( .A1(n3590), .A2(n3589), .ZN(n4961) );
  INV_X1 U4506 ( .A(n4961), .ZN(n3592) );
  INV_X1 U4507 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6948) );
  XNOR2_X1 U4508 ( .A(n5532), .B(n6948), .ZN(n4964) );
  INV_X1 U4509 ( .A(n4964), .ZN(n3591) );
  NAND2_X1 U4510 ( .A1(n5532), .A2(n6948), .ZN(n5528) );
  NAND3_X1 U4511 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(INSTADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n3593) );
  NAND2_X1 U4512 ( .A1(n5532), .A2(n3593), .ZN(n3594) );
  AND2_X1 U4513 ( .A1(n5528), .A2(n3594), .ZN(n3596) );
  NAND2_X1 U4514 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4274) );
  NAND2_X1 U4515 ( .A1(n5532), .A2(n4274), .ZN(n3595) );
  INV_X1 U4516 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5788) );
  INV_X1 U4517 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5768) );
  INV_X1 U4518 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6942) );
  INV_X1 U4519 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6928) );
  INV_X1 U4520 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5728) );
  NAND4_X1 U4521 ( .A1(n5768), .A2(n6942), .A3(n6928), .A4(n5728), .ZN(n3598)
         );
  NAND2_X1 U4522 ( .A1(n3597), .A2(n3598), .ZN(n3599) );
  AOI21_X2 U4523 ( .B1(n4962), .B2(n3600), .A(n3142), .ZN(n5519) );
  AND2_X1 U4524 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5723) );
  AND2_X1 U4525 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U4526 ( .A1(n5723), .A2(n5467), .ZN(n5485) );
  INV_X1 U4527 ( .A(n5485), .ZN(n3602) );
  NAND2_X1 U4528 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U4529 ( .A1(n3602), .A2(n3601), .ZN(n3603) );
  INV_X1 U4530 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6999) );
  INV_X1 U4531 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6925) );
  INV_X1 U4532 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5708) );
  INV_X1 U4533 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5692) );
  NAND4_X1 U4534 ( .A1(n6999), .A2(n6925), .A3(n5708), .A4(n5692), .ZN(n3604)
         );
  INV_X1 U4535 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5743) );
  INV_X1 U4536 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U4537 ( .A1(n5743), .A2(n5733), .ZN(n3608) );
  NOR2_X1 U4538 ( .A1(n3604), .A2(n3608), .ZN(n3605) );
  NAND2_X1 U4539 ( .A1(n5519), .A2(n3605), .ZN(n3606) );
  NOR2_X1 U4540 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5676) );
  NAND3_X1 U4541 ( .A1(n5462), .A2(n3597), .A3(n5676), .ZN(n5441) );
  INV_X1 U4542 ( .A(n3608), .ZN(n5724) );
  NOR2_X1 U4543 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3610) );
  NOR2_X1 U4544 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3609) );
  NAND4_X1 U4545 ( .A1(n5724), .A2(n3610), .A3(n3609), .A4(n5708), .ZN(n3611)
         );
  NAND2_X1 U4546 ( .A1(n3597), .A2(n3611), .ZN(n3612) );
  NAND2_X1 U4547 ( .A1(n5519), .A2(n3612), .ZN(n3615) );
  NAND3_X1 U4548 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A3(INSTADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n3613) );
  OAI21_X1 U4549 ( .B1(n5485), .B2(n3613), .A(n5532), .ZN(n3614) );
  NAND2_X1 U4550 ( .A1(n3615), .A2(n3614), .ZN(n5452) );
  INV_X1 U4551 ( .A(n5452), .ZN(n4102) );
  NAND3_X1 U4552 ( .A1(n4102), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5532), .ZN(n3616) );
  INV_X1 U4553 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U4554 ( .A1(n5441), .A2(n3616), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4224), .ZN(n3617) );
  INV_X1 U4555 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4232) );
  XNOR2_X1 U4556 ( .A(n3617), .B(n4232), .ZN(n5651) );
  AOI21_X1 U4557 ( .B1(n3671), .B2(n7068), .A(n4698), .ZN(n3631) );
  XNOR2_X1 U4558 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3619) );
  NAND2_X1 U4559 ( .A1(n3618), .A2(n3619), .ZN(n3637) );
  OAI21_X1 U4560 ( .B1(n3619), .B2(n3618), .A(n3637), .ZN(n4110) );
  NAND2_X1 U4561 ( .A1(n3631), .A2(n4110), .ZN(n3624) );
  XNOR2_X1 U4562 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3623) );
  AOI21_X1 U4563 ( .B1(n3318), .B2(n3623), .A(n3620), .ZN(n3622) );
  NAND2_X1 U4564 ( .A1(n3292), .A2(n5385), .ZN(n3621) );
  NAND2_X1 U4565 ( .A1(n4421), .A2(n3621), .ZN(n3639) );
  OR2_X1 U4566 ( .A1(n3622), .A2(n3639), .ZN(n3626) );
  NAND4_X1 U4567 ( .A1(n3624), .A2(n3671), .A3(n3623), .A4(n3626), .ZN(n3625)
         );
  NAND2_X1 U4568 ( .A1(n3625), .A2(n3660), .ZN(n3630) );
  INV_X1 U4569 ( .A(n3626), .ZN(n3628) );
  INV_X1 U4570 ( .A(n3631), .ZN(n3632) );
  NAND3_X1 U4571 ( .A1(n3632), .A2(STATE2_REG_0__SCAN_IN), .A3(n3627), .ZN(
        n3633) );
  NAND2_X1 U4572 ( .A1(n4756), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U4573 ( .A1(n3637), .A2(n3636), .ZN(n3647) );
  XNOR2_X1 U4574 ( .A(n4568), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3646)
         );
  XNOR2_X1 U4575 ( .A(n3647), .B(n3646), .ZN(n4109) );
  INV_X1 U4576 ( .A(n4109), .ZN(n3640) );
  NAND2_X1 U4577 ( .A1(n3671), .A2(n3640), .ZN(n3642) );
  INV_X1 U4578 ( .A(n3639), .ZN(n3641) );
  OAI211_X1 U4579 ( .C1(n3640), .C2(n3657), .A(n3642), .B(n3641), .ZN(n3644)
         );
  NOR2_X1 U4580 ( .A1(n3642), .A2(n3641), .ZN(n3643) );
  NAND2_X1 U4581 ( .A1(n3647), .A2(n3646), .ZN(n3649) );
  NAND2_X1 U4582 ( .A1(n7026), .A2(n4568), .ZN(n3648) );
  NAND2_X1 U4583 ( .A1(n3649), .A2(n3648), .ZN(n3655) );
  XNOR2_X1 U4584 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3654) );
  XNOR2_X1 U4585 ( .A(n3655), .B(n3654), .ZN(n4111) );
  INV_X1 U4586 ( .A(n4111), .ZN(n3650) );
  OAI22_X1 U4587 ( .A1(n3652), .A2(n3651), .B1(n3650), .B2(n3660), .ZN(n3659)
         );
  NOR2_X1 U4588 ( .A1(n4566), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3653)
         );
  AOI21_X1 U4589 ( .B1(n3655), .B2(n3654), .A(n3653), .ZN(n3663) );
  INV_X1 U4590 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7008) );
  NOR2_X1 U4591 ( .A1(n7008), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3656)
         );
  AND2_X1 U4592 ( .A1(n3663), .A2(n3656), .ZN(n4108) );
  NAND2_X1 U4593 ( .A1(n3657), .A2(n4108), .ZN(n3658) );
  NAND2_X1 U4594 ( .A1(n3659), .A2(n3658), .ZN(n3662) );
  AOI22_X1 U4595 ( .A1(n3668), .A2(n4108), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4647), .ZN(n3661) );
  NAND2_X1 U4596 ( .A1(n3662), .A2(n3661), .ZN(n3670) );
  INV_X1 U4597 ( .A(n3663), .ZN(n3665) );
  AND2_X1 U4598 ( .A1(n7008), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3664)
         );
  INV_X1 U4599 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U4600 ( .A1(n6238), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U4601 ( .A1(n3668), .A2(n4113), .ZN(n3669) );
  NAND2_X1 U4602 ( .A1(n3671), .A2(n4113), .ZN(n3672) );
  NAND2_X1 U4603 ( .A1(n4503), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6646) );
  AOI21_X1 U4604 ( .B1(n4657), .B2(n3675), .A(n4245), .ZN(n3676) );
  NAND2_X1 U4605 ( .A1(n3674), .A2(n3676), .ZN(n4134) );
  OR2_X1 U4606 ( .A1(n4134), .A2(n3318), .ZN(n4597) );
  NAND2_X1 U4607 ( .A1(n4717), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3822) );
  NAND2_X1 U4608 ( .A1(n6782), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3957) );
  INV_X1 U4609 ( .A(n3957), .ZN(n4336) );
  AOI21_X1 U4610 ( .B1(n4639), .B2(n3849), .A(n4336), .ZN(n3690) );
  AOI22_X1 U4611 ( .A1(n4337), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6782), .ZN(n3681) );
  AND2_X1 U4612 ( .A1(n3094), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3684) );
  NAND2_X1 U4613 ( .A1(n3684), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3680) );
  AND2_X1 U4614 ( .A1(n3681), .A2(n3680), .ZN(n3682) );
  OAI21_X1 U4615 ( .B1(n3679), .B2(n3822), .A(n3682), .ZN(n4510) );
  NAND2_X1 U4616 ( .A1(n4511), .A2(n4510), .ZN(n4509) );
  INV_X1 U4617 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6245) );
  NAND2_X1 U4618 ( .A1(n6782), .A2(n6245), .ZN(n4342) );
  OR2_X1 U4619 ( .A1(n4510), .A2(n4342), .ZN(n3683) );
  NAND2_X1 U4620 ( .A1(n4509), .A2(n3683), .ZN(n4515) );
  INV_X1 U4621 ( .A(n3684), .ZN(n3719) );
  NAND2_X1 U4622 ( .A1(n4641), .A2(n3849), .ZN(n3686) );
  AOI22_X1 U4623 ( .A1(n4337), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6782), .ZN(n3685) );
  OAI211_X1 U4624 ( .C1(n3719), .C2(n3635), .A(n3686), .B(n3685), .ZN(n4514)
         );
  NAND2_X1 U4625 ( .A1(n4515), .A2(n4514), .ZN(n4517) );
  INV_X1 U4626 ( .A(n4568), .ZN(n4946) );
  OAI21_X1 U4627 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3696), .ZN(n6477) );
  AOI22_X1 U4628 ( .A1(n4334), .A2(n6477), .B1(n4336), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3689) );
  NAND2_X1 U4629 ( .A1(n4083), .A2(EAX_REG_2__SCAN_IN), .ZN(n3688) );
  OAI211_X1 U4630 ( .C1(n3719), .C2(n4946), .A(n3689), .B(n3688), .ZN(n4529)
         );
  NAND2_X1 U4631 ( .A1(n4530), .A2(n4529), .ZN(n3694) );
  INV_X1 U4632 ( .A(n4517), .ZN(n3692) );
  INV_X1 U4633 ( .A(n3690), .ZN(n3691) );
  NAND2_X1 U4634 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  NAND2_X1 U4635 ( .A1(n3695), .A2(n3849), .ZN(n3702) );
  OAI21_X1 U4636 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3697), .A(n3713), 
        .ZN(n5300) );
  AOI22_X1 U4637 ( .A1(n4334), .A2(n5300), .B1(n4336), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4638 ( .A1(n4083), .A2(EAX_REG_3__SCAN_IN), .ZN(n3698) );
  OAI211_X1 U4639 ( .C1(n3719), .C2(n4566), .A(n3699), .B(n3698), .ZN(n3700)
         );
  INV_X1 U4640 ( .A(n3700), .ZN(n3701) );
  AND2_X2 U4641 ( .A1(n4618), .A2(n4617), .ZN(n4624) );
  NOR2_X1 U4642 ( .A1(n3703), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3704)
         );
  NOR2_X1 U4643 ( .A1(n3726), .A2(n3704), .ZN(n6340) );
  AOI22_X1 U4644 ( .A1(n4083), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6782), .ZN(n3705) );
  MUX2_X1 U4645 ( .A(n6340), .B(n3705), .S(n4342), .Z(n3706) );
  INV_X1 U4646 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6347) );
  XNOR2_X1 U4647 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .B(n3714), .ZN(n6356) );
  NAND2_X1 U4648 ( .A1(n6356), .A2(n4334), .ZN(n3708) );
  OAI21_X1 U4649 ( .B1(n6347), .B2(n3957), .A(n3708), .ZN(n3709) );
  AOI21_X1 U4650 ( .B1(n4083), .B2(EAX_REG_5__SCAN_IN), .A(n3709), .ZN(n3710)
         );
  NAND2_X1 U4651 ( .A1(n3712), .A2(n3849), .ZN(n3722) );
  INV_X1 U4652 ( .A(n3713), .ZN(n3716) );
  INV_X1 U4653 ( .A(n3714), .ZN(n3715) );
  OAI21_X1 U4654 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3716), .A(n3715), 
        .ZN(n6369) );
  NAND2_X1 U4655 ( .A1(n4083), .A2(EAX_REG_4__SCAN_IN), .ZN(n3718) );
  OAI21_X1 U4656 ( .B1(n6245), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6782), 
        .ZN(n3717) );
  OAI211_X1 U4657 ( .C1(n3719), .C2(n6238), .A(n3718), .B(n3717), .ZN(n3720)
         );
  OAI21_X1 U4658 ( .B1(n4342), .B2(n6369), .A(n3720), .ZN(n3721) );
  NAND2_X1 U4659 ( .A1(n3722), .A2(n3721), .ZN(n4623) );
  INV_X1 U4660 ( .A(n3724), .ZN(n3725) );
  NOR2_X1 U4661 ( .A1(n3726), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3727)
         );
  NOR2_X1 U4662 ( .A1(n3771), .A2(n3727), .ZN(n6322) );
  INV_X1 U4663 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6882) );
  OAI22_X1 U4664 ( .A1(n6322), .A2(n4342), .B1(n3957), .B2(n6882), .ZN(n3728)
         );
  AOI21_X1 U4665 ( .B1(n4083), .B2(EAX_REG_7__SCAN_IN), .A(n3728), .ZN(n3729)
         );
  AOI22_X1 U4666 ( .A1(n4311), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4667 ( .A1(n3096), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4668 ( .A1(n4313), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4669 ( .A1(n3344), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4670 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3741)
         );
  AOI22_X1 U4671 ( .A1(n4312), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4672 ( .A1(n3095), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4673 ( .A1(n4070), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4674 ( .A1(n3467), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4675 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  NOR2_X1 U4676 ( .A1(n3741), .A2(n3740), .ZN(n3744) );
  INV_X1 U4677 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5266) );
  XNOR2_X1 U4678 ( .A(n3791), .B(n5266), .ZN(n5592) );
  NAND2_X1 U4679 ( .A1(n5592), .A2(n4334), .ZN(n3743) );
  AOI22_X1 U4680 ( .A1(n4083), .A2(EAX_REG_11__SCAN_IN), .B1(n4336), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3742) );
  OAI211_X1 U4681 ( .C1(n3744), .C2(n3822), .A(n3743), .B(n3742), .ZN(n5263)
         );
  XOR2_X1 U4682 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3745), .Z(n6296) );
  AOI22_X1 U4683 ( .A1(n4311), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4684 ( .A1(n4313), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4312), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4685 ( .A1(n3096), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4686 ( .A1(n3095), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3746) );
  NAND4_X1 U4687 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3755)
         );
  AOI22_X1 U4688 ( .A1(n3395), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4689 ( .A1(n3401), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4690 ( .A1(n4314), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4691 ( .A1(n3467), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4692 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3754)
         );
  NOR2_X1 U4693 ( .A1(n3755), .A2(n3754), .ZN(n3758) );
  NAND2_X1 U4694 ( .A1(n4083), .A2(EAX_REG_10__SCAN_IN), .ZN(n3757) );
  NAND2_X1 U4695 ( .A1(n4336), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3756)
         );
  OAI211_X1 U4696 ( .C1(n3822), .C2(n3758), .A(n3757), .B(n3756), .ZN(n3759)
         );
  INV_X1 U4697 ( .A(n3759), .ZN(n3760) );
  OAI21_X1 U4698 ( .B1(n6296), .B2(n4342), .A(n3760), .ZN(n5259) );
  AOI22_X1 U4699 ( .A1(n4313), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4700 ( .A1(n3096), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4701 ( .A1(n3467), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4702 ( .A1(n3344), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3761) );
  NAND4_X1 U4703 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3770)
         );
  AOI22_X1 U4704 ( .A1(n4311), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4705 ( .A1(n3095), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4706 ( .A1(n4312), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4707 ( .A1(n3097), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4708 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3769)
         );
  NOR2_X1 U4709 ( .A1(n3770), .A2(n3769), .ZN(n3774) );
  XOR2_X1 U4710 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3771), .Z(n6312) );
  INV_X1 U4711 ( .A(n6312), .ZN(n5622) );
  AOI22_X1 U4712 ( .A1(n4336), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4334), 
        .B2(n5622), .ZN(n3773) );
  NAND2_X1 U4713 ( .A1(n4083), .A2(EAX_REG_8__SCAN_IN), .ZN(n3772) );
  OAI211_X1 U4714 ( .C1(n3822), .C2(n3774), .A(n3773), .B(n3772), .ZN(n5258)
         );
  INV_X1 U4715 ( .A(EAX_REG_9__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4716 ( .A1(n4311), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4717 ( .A1(n4313), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4718 ( .A1(n3467), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4719 ( .A1(n3095), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4720 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3784)
         );
  AOI22_X1 U4721 ( .A1(n4312), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4722 ( .A1(n3344), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4723 ( .A1(n4291), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4724 ( .A1(n3360), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3779) );
  NAND4_X1 U4725 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3783)
         );
  OAI21_X1 U4726 ( .B1(n3784), .B2(n3783), .A(n3849), .ZN(n3788) );
  INV_X1 U4727 ( .A(n3785), .ZN(n3786) );
  XNOR2_X1 U4728 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3786), .ZN(n5614) );
  AOI22_X1 U4729 ( .A1(n4334), .A2(n5614), .B1(n4336), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3787) );
  OAI211_X1 U4730 ( .C1(n3687), .C2(n3789), .A(n3788), .B(n3787), .ZN(n5283)
         );
  NAND4_X1 U4731 ( .A1(n5263), .A2(n5259), .A3(n5258), .A4(n5283), .ZN(n3790)
         );
  XOR2_X1 U4732 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3805), .Z(n6289) );
  AOI22_X1 U4733 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3395), .B1(n4289), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4734 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3344), .B1(n3095), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4735 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3467), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4736 ( .A1(n3096), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4737 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3801)
         );
  AOI22_X1 U4738 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4311), .B1(n4312), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4739 ( .A1(n4313), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4740 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4070), .B1(n3097), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4741 ( .A1(n3401), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3796) );
  NAND4_X1 U4742 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3800)
         );
  OR2_X1 U4743 ( .A1(n3801), .A2(n3800), .ZN(n3802) );
  AOI22_X1 U4744 ( .A1(n3849), .A2(n3802), .B1(n4336), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3804) );
  NAND2_X1 U4745 ( .A1(n4083), .A2(EAX_REG_12__SCAN_IN), .ZN(n3803) );
  OAI211_X1 U4746 ( .C1(n6289), .C2(n4342), .A(n3804), .B(n3803), .ZN(n5360)
         );
  NAND2_X1 U4747 ( .A1(n5260), .A2(n5360), .ZN(n4990) );
  INV_X1 U4748 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U4749 ( .A1(n3806), .A2(n6959), .ZN(n3808) );
  INV_X1 U4750 ( .A(n3852), .ZN(n3807) );
  NAND2_X1 U4751 ( .A1(n3808), .A2(n3807), .ZN(n6278) );
  AOI22_X1 U4752 ( .A1(n4311), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4753 ( .A1(n3095), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4754 ( .A1(n4070), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4755 ( .A1(n4314), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4756 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3818)
         );
  AOI22_X1 U4757 ( .A1(n3255), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4758 ( .A1(n3467), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4759 ( .A1(n4290), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4760 ( .A1(n3096), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3813) );
  NAND4_X1 U4761 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3817)
         );
  NOR2_X1 U4762 ( .A1(n3818), .A2(n3817), .ZN(n3821) );
  NAND2_X1 U4763 ( .A1(n4083), .A2(EAX_REG_13__SCAN_IN), .ZN(n3820) );
  NAND2_X1 U4764 ( .A1(n4336), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3819)
         );
  OAI211_X1 U4765 ( .C1(n3822), .C2(n3821), .A(n3820), .B(n3819), .ZN(n3823)
         );
  AOI21_X1 U4766 ( .B1(n6278), .B2(n4334), .A(n3823), .ZN(n4991) );
  AOI22_X1 U4767 ( .A1(n4313), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4768 ( .A1(n3360), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4769 ( .A1(n3095), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4770 ( .A1(n3395), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3826) );
  NAND4_X1 U4771 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3835)
         );
  AOI22_X1 U4772 ( .A1(n4311), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4773 ( .A1(n3442), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4774 ( .A1(n4314), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4775 ( .A1(n4290), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4776 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3834)
         );
  OAI21_X1 U4777 ( .B1(n3835), .B2(n3834), .A(n3849), .ZN(n3838) );
  XNOR2_X1 U4778 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3852), .ZN(n6269)
         );
  AOI22_X1 U4779 ( .A1(n4334), .A2(n6269), .B1(n4336), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U4780 ( .A1(n4083), .A2(EAX_REG_14__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4781 ( .A1(n3358), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4782 ( .A1(n3442), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4783 ( .A1(n4319), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4784 ( .A1(n4069), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4785 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3851)
         );
  AOI22_X1 U4786 ( .A1(n4313), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4787 ( .A1(n3095), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4788 ( .A1(n4290), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4789 ( .A1(n4314), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3845) );
  NAND4_X1 U4790 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3850)
         );
  OAI21_X1 U4791 ( .B1(n3851), .B2(n3850), .A(n3849), .ZN(n3855) );
  AND2_X2 U4792 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n3852), .ZN(n3868)
         );
  XNOR2_X1 U4793 ( .A(n3868), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5568)
         );
  AOI22_X1 U4794 ( .A1(n5568), .A2(n4334), .B1(n4336), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3854) );
  NAND2_X1 U4795 ( .A1(n4083), .A2(EAX_REG_15__SCAN_IN), .ZN(n3853) );
  INV_X1 U4796 ( .A(n3856), .ZN(n4579) );
  NAND2_X1 U4797 ( .A1(n4579), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4331) );
  AOI22_X1 U4798 ( .A1(n3395), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4799 ( .A1(n4069), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4800 ( .A1(n3096), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4801 ( .A1(n3344), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4802 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3866)
         );
  AOI22_X1 U4803 ( .A1(n3358), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4290), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4804 ( .A1(n3095), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4805 ( .A1(n4313), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4806 ( .A1(n3442), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4807 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3865)
         );
  NOR2_X1 U4808 ( .A1(n3866), .A2(n3865), .ZN(n3867) );
  OR2_X1 U4809 ( .A1(n4331), .A2(n3867), .ZN(n3871) );
  XNOR2_X1 U4810 ( .A(n3872), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5562)
         );
  INV_X1 U4811 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5560) );
  OAI22_X1 U4812 ( .A1(n5562), .A2(n4342), .B1(n5560), .B2(n3957), .ZN(n3869)
         );
  AOI21_X1 U4813 ( .B1(n4083), .B2(EAX_REG_16__SCAN_IN), .A(n3869), .ZN(n3870)
         );
  NAND2_X1 U4814 ( .A1(n3871), .A2(n3870), .ZN(n5230) );
  INV_X1 U4815 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n7038) );
  OAI21_X1 U4816 ( .B1(n3872), .B2(n5560), .A(n7038), .ZN(n3875) );
  AND2_X1 U4817 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3873) );
  NAND2_X1 U4818 ( .A1(n3875), .A2(n4015), .ZN(n5550) );
  AOI22_X1 U4819 ( .A1(n4311), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4312), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4820 ( .A1(n3442), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4821 ( .A1(n3096), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4822 ( .A1(n4291), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4823 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3885)
         );
  AOI22_X1 U4824 ( .A1(n3395), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4825 ( .A1(n3401), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4826 ( .A1(n4313), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4827 ( .A1(n4314), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4828 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3884)
         );
  NOR2_X1 U4829 ( .A1(n3885), .A2(n3884), .ZN(n3887) );
  AOI22_X1 U4830 ( .A1(n4083), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6782), .ZN(n3886) );
  OAI21_X1 U4831 ( .B1(n4331), .B2(n3887), .A(n3886), .ZN(n3888) );
  MUX2_X1 U4832 ( .A(n5550), .B(n3888), .S(n4342), .Z(n5214) );
  AND2_X2 U4833 ( .A1(n5212), .A2(n5214), .ZN(n5093) );
  AOI22_X1 U4834 ( .A1(n4311), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4835 ( .A1(n4313), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4836 ( .A1(n4290), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4837 ( .A1(n4291), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4838 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3898)
         );
  AOI22_X1 U4839 ( .A1(n3467), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4840 ( .A1(n3095), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4841 ( .A1(n3360), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4842 ( .A1(n4314), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4843 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  OR2_X1 U4844 ( .A1(n3898), .A2(n3897), .ZN(n3955) );
  INV_X1 U4845 ( .A(n3955), .ZN(n3919) );
  AOI22_X1 U4846 ( .A1(n4311), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4847 ( .A1(n4288), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4848 ( .A1(n4290), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3900) );
  INV_X1 U4849 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6816) );
  AOI22_X1 U4850 ( .A1(n4291), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4851 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3908)
         );
  AOI22_X1 U4852 ( .A1(n3467), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4853 ( .A1(n3095), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4854 ( .A1(n3360), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4855 ( .A1(n3344), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4856 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3907)
         );
  OR2_X1 U4857 ( .A1(n3908), .A2(n3907), .ZN(n3965) );
  AOI22_X1 U4858 ( .A1(n4311), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4859 ( .A1(n4288), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4860 ( .A1(n4290), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4289), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4861 ( .A1(n4291), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3909) );
  NAND4_X1 U4862 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3918)
         );
  AOI22_X1 U4863 ( .A1(n3467), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4864 ( .A1(n3095), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4865 ( .A1(n3360), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4866 ( .A1(n3344), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4867 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3917)
         );
  OR2_X1 U4868 ( .A1(n3918), .A2(n3917), .ZN(n3964) );
  NAND2_X1 U4869 ( .A1(n3965), .A2(n3964), .ZN(n3956) );
  NOR2_X1 U4870 ( .A1(n3919), .A2(n3956), .ZN(n3947) );
  AOI22_X1 U4871 ( .A1(n4311), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4872 ( .A1(n4288), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4873 ( .A1(n4312), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4874 ( .A1(n4291), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4875 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3929)
         );
  AOI22_X1 U4876 ( .A1(n3467), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4877 ( .A1(n3095), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4878 ( .A1(n3360), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4879 ( .A1(n4314), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3924) );
  NAND4_X1 U4880 ( .A1(n3927), .A2(n3926), .A3(n3925), .A4(n3924), .ZN(n3928)
         );
  OR2_X1 U4881 ( .A1(n3929), .A2(n3928), .ZN(n3948) );
  NAND2_X1 U4882 ( .A1(n3947), .A2(n3948), .ZN(n4062) );
  AOI22_X1 U4883 ( .A1(n4069), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4884 ( .A1(n4289), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4885 ( .A1(n3096), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4886 ( .A1(n3344), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U4887 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3939)
         );
  AOI22_X1 U4888 ( .A1(n4311), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4889 ( .A1(n3467), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4890 ( .A1(n4288), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4891 ( .A1(n4312), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3934) );
  NAND4_X1 U4892 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(n3938)
         );
  NOR2_X1 U4893 ( .A1(n3939), .A2(n3938), .ZN(n4063) );
  XNOR2_X1 U4894 ( .A(n4062), .B(n4063), .ZN(n3941) );
  AOI22_X1 U4895 ( .A1(n4083), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6782), .ZN(n3940) );
  OAI21_X1 U4896 ( .B1(n3941), .B2(n4331), .A(n3940), .ZN(n3946) );
  INV_X1 U4897 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5540) );
  OR2_X2 U4898 ( .A1(n4015), .A2(n5540), .ZN(n4017) );
  NAND2_X1 U4899 ( .A1(n3942), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4032)
         );
  INV_X1 U4900 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n7007) );
  INV_X1 U4901 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6955) );
  INV_X1 U4902 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5116) );
  INV_X1 U4903 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5457) );
  INV_X1 U4904 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5080) );
  OR2_X2 U4905 ( .A1(n3944), .A2(n5080), .ZN(n4086) );
  NAND2_X1 U4906 ( .A1(n3944), .A2(n5080), .ZN(n3945) );
  NAND2_X1 U4907 ( .A1(n4086), .A2(n3945), .ZN(n5450) );
  MUX2_X1 U4908 ( .A(n3946), .B(n5450), .S(n4334), .Z(n5079) );
  INV_X1 U4909 ( .A(n4331), .ZN(n4305) );
  XOR2_X1 U4910 ( .A(n3948), .B(n3947), .Z(n3951) );
  INV_X1 U4911 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3949) );
  OAI22_X1 U4912 ( .A1(n3687), .A2(n3949), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5457), .ZN(n3950) );
  AOI21_X1 U4913 ( .B1(n4305), .B2(n3951), .A(n3950), .ZN(n3953) );
  XNOR2_X1 U4914 ( .A(n3952), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5459)
         );
  MUX2_X1 U4915 ( .A(n3953), .B(n5459), .S(n4334), .Z(n5096) );
  XNOR2_X1 U4916 ( .A(n3954), .B(n5116), .ZN(n5478) );
  NAND2_X1 U4917 ( .A1(n5478), .A2(n4334), .ZN(n3962) );
  XNOR2_X1 U4918 ( .A(n3956), .B(n3955), .ZN(n3960) );
  INV_X1 U4919 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3958) );
  OAI22_X1 U4920 ( .A1(n3687), .A2(n3958), .B1(n3957), .B2(n5116), .ZN(n3959)
         );
  AOI21_X1 U4921 ( .B1(n4305), .B2(n3960), .A(n3959), .ZN(n3961) );
  AND2_X1 U4922 ( .A1(n3962), .A2(n3961), .ZN(n5112) );
  INV_X1 U4923 ( .A(n5112), .ZN(n3985) );
  INV_X1 U4924 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5125) );
  XNOR2_X1 U4925 ( .A(n3971), .B(n5125), .ZN(n5489) );
  XNOR2_X1 U4926 ( .A(n3965), .B(n3964), .ZN(n3967) );
  AOI22_X1 U4927 ( .A1(n4083), .A2(EAX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6782), .ZN(n3966) );
  OAI21_X1 U4928 ( .B1(n4331), .B2(n3967), .A(n3966), .ZN(n3968) );
  MUX2_X1 U4929 ( .A(n5489), .B(n3968), .S(n4342), .Z(n5124) );
  NAND2_X1 U4930 ( .A1(n3969), .A2(n6955), .ZN(n3970) );
  NAND2_X1 U4931 ( .A1(n3971), .A2(n3970), .ZN(n5498) );
  AOI22_X1 U4932 ( .A1(n4311), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4933 ( .A1(n4313), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4934 ( .A1(n3095), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4935 ( .A1(n3360), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U4936 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3981)
         );
  AOI22_X1 U4937 ( .A1(n3395), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4290), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4938 ( .A1(n3096), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4939 ( .A1(n4291), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4940 ( .A1(n4314), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4941 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3980)
         );
  NOR2_X1 U4942 ( .A1(n3981), .A2(n3980), .ZN(n3983) );
  AOI22_X1 U4943 ( .A1(n4083), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6782), .ZN(n3982) );
  OAI21_X1 U4944 ( .B1(n4331), .B2(n3983), .A(n3982), .ZN(n3984) );
  MUX2_X1 U4945 ( .A(n5498), .B(n3984), .S(n4342), .Z(n5138) );
  AND2_X1 U4946 ( .A1(n5124), .A2(n5138), .ZN(n5111) );
  NAND2_X1 U4947 ( .A1(n3985), .A2(n5111), .ZN(n4050) );
  AOI22_X1 U4948 ( .A1(n4311), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4949 ( .A1(n4313), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4950 ( .A1(n4312), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4289), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4951 ( .A1(n4291), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3986) );
  NAND4_X1 U4952 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3995)
         );
  AOI22_X1 U4953 ( .A1(n3467), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4954 ( .A1(n3095), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4955 ( .A1(n3360), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4956 ( .A1(n4314), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3990) );
  NAND4_X1 U4957 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n3994)
         );
  NOR2_X1 U4958 ( .A1(n3995), .A2(n3994), .ZN(n3998) );
  INV_X1 U4959 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5505) );
  AOI21_X1 U4960 ( .B1(n5505), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3996) );
  AOI21_X1 U4961 ( .B1(n4083), .B2(EAX_REG_21__SCAN_IN), .A(n3996), .ZN(n3997)
         );
  OAI21_X1 U4962 ( .B1(n4331), .B2(n3998), .A(n3997), .ZN(n4000) );
  XNOR2_X1 U4963 ( .A(n4034), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5507)
         );
  NAND2_X1 U4964 ( .A1(n5507), .A2(n4334), .ZN(n3999) );
  INV_X1 U4965 ( .A(n5153), .ZN(n4049) );
  XNOR2_X1 U4966 ( .A(n4017), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5526)
         );
  AOI22_X1 U4967 ( .A1(n3395), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4290), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4968 ( .A1(n4313), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4969 ( .A1(n3467), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4970 ( .A1(n4069), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4971 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4010)
         );
  AOI22_X1 U4972 ( .A1(n4311), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4973 ( .A1(n3095), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4974 ( .A1(n4291), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4975 ( .A1(n3344), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4976 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4009)
         );
  OR2_X1 U4977 ( .A1(n4010), .A2(n4009), .ZN(n4013) );
  INV_X1 U4978 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4011) );
  INV_X1 U4979 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5522) );
  OAI22_X1 U4980 ( .A1(n3687), .A2(n4011), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5522), .ZN(n4012) );
  AOI21_X1 U4981 ( .B1(n4305), .B2(n4013), .A(n4012), .ZN(n4014) );
  MUX2_X1 U4982 ( .A(n5526), .B(n4014), .S(n4342), .Z(n5180) );
  NAND2_X1 U4983 ( .A1(n4015), .A2(n5540), .ZN(n4016) );
  AND2_X1 U4984 ( .A1(n4017), .A2(n4016), .ZN(n5538) );
  AOI22_X1 U4985 ( .A1(n3395), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4986 ( .A1(n3096), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4987 ( .A1(n4290), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4988 ( .A1(n3095), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4018) );
  NAND4_X1 U4989 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4027)
         );
  AOI22_X1 U4990 ( .A1(n4313), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4991 ( .A1(n4314), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4992 ( .A1(n4311), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4993 ( .A1(n3467), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4022) );
  NAND4_X1 U4994 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4026)
         );
  OR2_X1 U4995 ( .A1(n4027), .A2(n4026), .ZN(n4030) );
  INV_X1 U4996 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4028) );
  OAI22_X1 U4997 ( .A1(n3687), .A2(n4028), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5540), .ZN(n4029) );
  AOI21_X1 U4998 ( .B1(n4305), .B2(n4030), .A(n4029), .ZN(n4031) );
  MUX2_X1 U4999 ( .A(n5538), .B(n4031), .S(n4342), .Z(n5199) );
  OR2_X1 U5000 ( .A1(n5180), .A2(n5199), .ZN(n5163) );
  NAND2_X1 U5001 ( .A1(n4032), .A2(n7007), .ZN(n4033) );
  AND2_X1 U5002 ( .A1(n4034), .A2(n4033), .ZN(n5515) );
  AOI22_X1 U5003 ( .A1(n4311), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5004 ( .A1(n4313), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5005 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4070), .B1(n3360), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5006 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3095), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4035) );
  NAND4_X1 U5007 ( .A1(n4038), .A2(n4037), .A3(n4036), .A4(n4035), .ZN(n4044)
         );
  AOI22_X1 U5008 ( .A1(n3395), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4290), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5009 ( .A1(n3467), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5010 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4314), .B1(n4296), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5011 ( .A1(n4291), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U5012 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4043)
         );
  OR2_X1 U5013 ( .A1(n4044), .A2(n4043), .ZN(n4047) );
  INV_X1 U5014 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4045) );
  OAI22_X1 U5015 ( .A1(n3687), .A2(n4045), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7007), .ZN(n4046) );
  AOI21_X1 U5016 ( .B1(n4305), .B2(n4047), .A(n4046), .ZN(n4048) );
  MUX2_X1 U5017 ( .A(n5515), .B(n4048), .S(n4342), .Z(n5164) );
  NOR2_X1 U5018 ( .A1(n5096), .A2(n5094), .ZN(n5078) );
  AOI22_X1 U5019 ( .A1(n4311), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5020 ( .A1(n4288), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5021 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4312), .B1(n4289), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5022 ( .A1(n4291), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4052) );
  NAND4_X1 U5023 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(n4061)
         );
  AOI22_X1 U5024 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3467), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5025 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3095), .B1(n4069), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5026 ( .A1(n3360), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5027 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3344), .B1(n4296), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4056) );
  NAND4_X1 U5028 ( .A1(n4059), .A2(n4058), .A3(n4057), .A4(n4056), .ZN(n4060)
         );
  OR2_X1 U5029 ( .A1(n4061), .A2(n4060), .ZN(n4081) );
  NOR2_X1 U5030 ( .A1(n4063), .A2(n4062), .ZN(n4082) );
  XOR2_X1 U5031 ( .A(n4081), .B(n4082), .Z(n4066) );
  INV_X1 U5032 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4064) );
  INV_X1 U5033 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5445) );
  OAI22_X1 U5034 ( .A1(n3687), .A2(n4064), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5445), .ZN(n4065) );
  AOI21_X1 U5035 ( .B1(n4066), .B2(n4305), .A(n4065), .ZN(n4068) );
  INV_X1 U5036 ( .A(n4086), .ZN(n4067) );
  XOR2_X1 U5037 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .B(n4067), .Z(n5443) );
  MUX2_X1 U5038 ( .A(n4068), .B(n5443), .S(n4334), .Z(n5067) );
  AOI22_X1 U5039 ( .A1(n4311), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5040 ( .A1(n4312), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5041 ( .A1(n4069), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5042 ( .A1(n4070), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4071) );
  NAND4_X1 U5043 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4080)
         );
  AOI22_X1 U5044 ( .A1(n3442), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5045 ( .A1(n3255), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5046 ( .A1(n4314), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5047 ( .A1(n4288), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U5048 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4079)
         );
  NOR2_X1 U5049 ( .A1(n4080), .A2(n4079), .ZN(n4287) );
  NAND2_X1 U5050 ( .A1(n4082), .A2(n4081), .ZN(n4286) );
  XNOR2_X1 U5051 ( .A(n4287), .B(n4286), .ZN(n4085) );
  AOI22_X1 U5052 ( .A1(n4083), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6782), .ZN(n4084) );
  OAI21_X1 U5053 ( .B1(n4085), .B2(n4331), .A(n4084), .ZN(n4090) );
  NOR2_X2 U5054 ( .A1(n4086), .A2(n5445), .ZN(n4087) );
  INV_X1 U5055 ( .A(n4087), .ZN(n4088) );
  INV_X1 U5056 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U5057 ( .A1(n4088), .A2(n5055), .ZN(n4089) );
  NAND2_X1 U5058 ( .A1(n4333), .A2(n4089), .ZN(n5054) );
  MUX2_X1 U5059 ( .A(n4090), .B(n5054), .S(n4334), .Z(n4091) );
  OAI21_X1 U5060 ( .B1(n3090), .B2(n4091), .A(n4308), .ZN(n5395) );
  AND3_X1 U5061 ( .A1(n4647), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U5062 ( .A1(n6864), .A2(n6782), .ZN(n5998) );
  NAND2_X1 U5063 ( .A1(n4406), .A2(n6186), .ZN(n6178) );
  NAND2_X1 U5064 ( .A1(n4092), .A2(n5998), .ZN(n6736) );
  NAND2_X1 U5065 ( .A1(n6736), .A2(n4647), .ZN(n4093) );
  NAND2_X1 U5066 ( .A1(n4094), .A2(n6782), .ZN(n6498) );
  INV_X1 U5067 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7046) );
  NOR2_X1 U5068 ( .A1(n6498), .A2(n7046), .ZN(n5655) );
  NAND2_X1 U5069 ( .A1(n4647), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4096) );
  NAND2_X1 U5070 ( .A1(n6245), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4095) );
  NAND2_X1 U5071 ( .A1(n4096), .A2(n4095), .ZN(n5647) );
  NOR2_X1 U5072 ( .A1(n6478), .A2(n5054), .ZN(n4097) );
  AOI211_X1 U5073 ( .C1(PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n6466), .A(n5655), 
        .B(n4097), .ZN(n4098) );
  NAND2_X1 U5074 ( .A1(n4101), .A2(n4100), .ZN(U2958) );
  NOR2_X1 U5075 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5652) );
  NAND3_X1 U5076 ( .A1(n3597), .A2(n5652), .A3(n4224), .ZN(n4997) );
  OR2_X1 U5078 ( .A1(n5452), .A2(n3141), .ZN(n5440) );
  INV_X1 U5080 ( .A(n4105), .ZN(n4107) );
  INV_X1 U5081 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4106) );
  NAND2_X1 U5082 ( .A1(n4107), .A2(n4106), .ZN(n4462) );
  NAND2_X1 U5083 ( .A1(n7068), .A2(n4462), .ZN(n4114) );
  NOR4_X1 U5084 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4112)
         );
  OR2_X1 U5085 ( .A1(n4113), .A2(n4112), .ZN(n4430) );
  NOR2_X1 U5086 ( .A1(READY_N), .A2(n4430), .ZN(n4452) );
  NAND2_X1 U5087 ( .A1(n4114), .A2(n4452), .ZN(n4117) );
  NAND3_X1 U5088 ( .A1(n4420), .A2(n4115), .A3(n7068), .ZN(n4116) );
  MUX2_X1 U5089 ( .A(n4117), .B(n4116), .S(n4724), .Z(n4124) );
  INV_X1 U5090 ( .A(n4134), .ZN(n4122) );
  OR2_X1 U5091 ( .A1(n4118), .A2(n4115), .ZN(n4121) );
  NAND2_X1 U5092 ( .A1(n4119), .A2(n4717), .ZN(n4259) );
  AND2_X1 U5093 ( .A1(n4259), .A2(n5023), .ZN(n4120) );
  NAND2_X1 U5094 ( .A1(n4121), .A2(n4120), .ZN(n4246) );
  NAND2_X1 U5095 ( .A1(n4122), .A2(n4246), .ZN(n4123) );
  NAND2_X1 U5096 ( .A1(n4123), .A2(n4340), .ZN(n4258) );
  NAND2_X1 U5097 ( .A1(n4124), .A2(n4258), .ZN(n4125) );
  INV_X1 U5098 ( .A(n6646), .ZN(n4636) );
  NAND2_X1 U5099 ( .A1(n4125), .A2(n4636), .ZN(n4132) );
  AOI21_X1 U5100 ( .B1(n3292), .B2(n4462), .A(READY_N), .ZN(n4129) );
  NAND2_X1 U5101 ( .A1(n5043), .A2(n5023), .ZN(n4128) );
  AOI21_X1 U5102 ( .B1(n4126), .B2(n4129), .A(n4128), .ZN(n4130) );
  INV_X1 U5103 ( .A(n4145), .ZN(n4519) );
  NAND2_X1 U5104 ( .A1(n4126), .A2(n4519), .ZN(n4468) );
  OAI21_X1 U5105 ( .B1(n4685), .B2(n4240), .A(n4597), .ZN(n4133) );
  INV_X1 U5106 ( .A(n4133), .ZN(n4135) );
  OR2_X1 U5107 ( .A1(n4134), .A2(n4421), .ZN(n4555) );
  NOR2_X1 U5108 ( .A1(n4340), .A2(n7068), .ZN(n6235) );
  INV_X1 U5109 ( .A(n6235), .ZN(n4593) );
  AND4_X1 U5110 ( .A1(n4468), .A2(n4135), .A3(n4555), .A4(n4593), .ZN(n4136)
         );
  NAND2_X1 U5111 ( .A1(n4392), .A2(n6502), .ZN(n4285) );
  NAND2_X1 U5112 ( .A1(n3122), .A2(EBX_REG_0__SCAN_IN), .ZN(n4138) );
  INV_X1 U5113 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4542) );
  NAND2_X1 U5114 ( .A1(n3122), .A2(n4542), .ZN(n4139) );
  OAI211_X1 U5115 ( .C1(n3123), .C2(EBX_REG_1__SCAN_IN), .A(n4139), .B(n4147), 
        .ZN(n4141) );
  NAND2_X1 U5116 ( .A1(n4141), .A2(n4140), .ZN(n4142) );
  XNOR2_X1 U5117 ( .A(n4499), .B(n4142), .ZN(n4520) );
  INV_X1 U5118 ( .A(n4142), .ZN(n4143) );
  NAND2_X1 U5119 ( .A1(n4143), .A2(n4499), .ZN(n4144) );
  NAND2_X1 U5120 ( .A1(n4518), .A2(n4144), .ZN(n4534) );
  INV_X1 U5121 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4146) );
  NAND2_X1 U5122 ( .A1(n4210), .A2(n4146), .ZN(n4148) );
  OAI211_X1 U5123 ( .C1(n4145), .C2(EBX_REG_2__SCAN_IN), .A(n4148), .B(n4349), 
        .ZN(n4150) );
  INV_X1 U5124 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4536) );
  NAND2_X1 U5125 ( .A1(n5169), .A2(n4536), .ZN(n4149) );
  INV_X1 U5126 ( .A(n4533), .ZN(n4151) );
  INV_X1 U5127 ( .A(n4153), .ZN(n4155) );
  NAND2_X1 U5128 ( .A1(n4498), .A2(n6837), .ZN(n4154) );
  NAND2_X1 U5129 ( .A1(n4155), .A2(n4154), .ZN(n4621) );
  MUX2_X1 U5130 ( .A(n5169), .B(n4220), .S(EBX_REG_4__SCAN_IN), .Z(n4156) );
  INV_X1 U5131 ( .A(n4156), .ZN(n4158) );
  NAND2_X1 U5132 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4157)
         );
  NAND2_X1 U5133 ( .A1(n4158), .A2(n4157), .ZN(n4674) );
  NAND2_X1 U5134 ( .A1(n3121), .A2(n3119), .ZN(n4668) );
  INV_X1 U5135 ( .A(n4668), .ZN(n4163) );
  MUX2_X1 U5136 ( .A(n4228), .B(n3131), .S(EBX_REG_5__SCAN_IN), .Z(n4159) );
  INV_X1 U5137 ( .A(n4159), .ZN(n4161) );
  NAND2_X1 U5138 ( .A1(n4498), .A2(n4893), .ZN(n4160) );
  NAND2_X1 U5139 ( .A1(n4161), .A2(n4160), .ZN(n4672) );
  NAND2_X1 U5140 ( .A1(n4163), .A2(n4162), .ZN(n4670) );
  NAND2_X1 U5141 ( .A1(n4210), .A2(n4164), .ZN(n4165) );
  OAI211_X1 U5142 ( .C1(n4145), .C2(EBX_REG_6__SCAN_IN), .A(n4165), .B(n4349), 
        .ZN(n4167) );
  INV_X1 U5143 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4795) );
  NAND2_X1 U5144 ( .A1(n3131), .A2(n4795), .ZN(n4166) );
  MUX2_X1 U5145 ( .A(n4228), .B(n5169), .S(EBX_REG_7__SCAN_IN), .Z(n4169) );
  NOR2_X1 U5146 ( .A1(n4356), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4168)
         );
  NOR2_X1 U5147 ( .A1(n4169), .A2(n4168), .ZN(n4839) );
  NAND2_X1 U5148 ( .A1(n4210), .A2(n5815), .ZN(n4170) );
  OAI211_X1 U5149 ( .C1(n4145), .C2(EBX_REG_8__SCAN_IN), .A(n4170), .B(n4349), 
        .ZN(n4172) );
  INV_X1 U5150 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U5151 ( .A1(n3131), .A2(n6829), .ZN(n4171) );
  NAND2_X1 U5152 ( .A1(n4172), .A2(n4171), .ZN(n5379) );
  MUX2_X1 U5153 ( .A(n4228), .B(n3131), .S(EBX_REG_9__SCAN_IN), .Z(n4173) );
  INV_X1 U5154 ( .A(n4173), .ZN(n4175) );
  NAND2_X1 U5155 ( .A1(n4498), .A2(n5808), .ZN(n4174) );
  NAND2_X1 U5156 ( .A1(n4175), .A2(n4174), .ZN(n5280) );
  MUX2_X1 U5157 ( .A(n5169), .B(n4220), .S(EBX_REG_10__SCAN_IN), .Z(n4177) );
  AND2_X1 U5158 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4176)
         );
  NOR2_X1 U5159 ( .A1(n4177), .A2(n4176), .ZN(n5366) );
  INV_X1 U5160 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U5161 ( .A1(n4228), .A2(n5363), .ZN(n4180) );
  NAND2_X1 U5162 ( .A1(n4349), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4178) );
  OAI211_X1 U5163 ( .C1(n4145), .C2(EBX_REG_11__SCAN_IN), .A(n4178), .B(n4210), 
        .ZN(n4179) );
  AND2_X1 U5164 ( .A1(n4180), .A2(n4179), .ZN(n5264) );
  INV_X1 U5165 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U5166 ( .A1(n4228), .A2(n6382), .ZN(n4183) );
  NAND2_X1 U5167 ( .A1(n4349), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4181) );
  OAI211_X1 U5168 ( .C1(n4145), .C2(EBX_REG_13__SCAN_IN), .A(n4181), .B(n4210), 
        .ZN(n4182) );
  AND2_X1 U5169 ( .A1(n4183), .A2(n4182), .ZN(n4982) );
  MUX2_X1 U5170 ( .A(n3131), .B(n4220), .S(EBX_REG_12__SCAN_IN), .Z(n4184) );
  INV_X1 U5171 ( .A(n4184), .ZN(n4186) );
  NAND2_X1 U5172 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4185) );
  NAND2_X1 U5173 ( .A1(n4186), .A2(n4185), .ZN(n5359) );
  MUX2_X1 U5174 ( .A(n5169), .B(n4220), .S(EBX_REG_14__SCAN_IN), .Z(n4189) );
  AND2_X1 U5175 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4188)
         );
  NOR2_X1 U5176 ( .A1(n4189), .A2(n4188), .ZN(n5356) );
  NOR2_X2 U5177 ( .A1(n4981), .A2(n5356), .ZN(n5250) );
  NAND2_X1 U5178 ( .A1(n4356), .A2(EBX_REG_15__SCAN_IN), .ZN(n4191) );
  NAND2_X1 U5179 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4190) );
  NAND2_X1 U5180 ( .A1(n4191), .A2(n4190), .ZN(n4192) );
  XNOR2_X1 U5181 ( .A(n4192), .B(n4349), .ZN(n5249) );
  NAND2_X1 U5182 ( .A1(n5250), .A2(n5249), .ZN(n5238) );
  MUX2_X1 U5183 ( .A(n3131), .B(n4220), .S(EBX_REG_16__SCAN_IN), .Z(n4194) );
  AND2_X1 U5184 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4193)
         );
  NOR2_X1 U5185 ( .A1(n4194), .A2(n4193), .ZN(n5240) );
  INV_X1 U5186 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U5187 ( .A1(n4228), .A2(n5348), .ZN(n4199) );
  NAND2_X1 U5188 ( .A1(n4349), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4197) );
  OAI211_X1 U5189 ( .C1(n4145), .C2(EBX_REG_17__SCAN_IN), .A(n4197), .B(n4210), 
        .ZN(n4198) );
  NAND2_X1 U5190 ( .A1(n4199), .A2(n4198), .ZN(n5216) );
  NAND2_X1 U5191 ( .A1(n3118), .A2(n4200), .ZN(n5184) );
  NAND2_X1 U5192 ( .A1(n4210), .A2(n5743), .ZN(n4201) );
  OAI211_X1 U5193 ( .C1(n4145), .C2(EBX_REG_19__SCAN_IN), .A(n4201), .B(n4349), 
        .ZN(n4203) );
  INV_X1 U5194 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6879) );
  NAND2_X1 U5195 ( .A1(n5169), .A2(n6879), .ZN(n4202) );
  AND2_X1 U5196 ( .A1(n4203), .A2(n4202), .ZN(n5188) );
  NAND2_X1 U5197 ( .A1(n4356), .A2(EBX_REG_18__SCAN_IN), .ZN(n4205) );
  NAND2_X1 U5198 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4204) );
  NAND2_X1 U5199 ( .A1(n4205), .A2(n4204), .ZN(n5168) );
  AND2_X1 U5200 ( .A1(n5168), .A2(n4349), .ZN(n5186) );
  NOR2_X1 U5201 ( .A1(n5168), .A2(n4349), .ZN(n5185) );
  OAI22_X1 U5202 ( .A1(n4356), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4145), .ZN(n5170) );
  MUX2_X1 U5203 ( .A(n5186), .B(n5185), .S(n5170), .Z(n4206) );
  NAND2_X1 U5204 ( .A1(n5167), .A2(n4206), .ZN(n5155) );
  MUX2_X1 U5205 ( .A(n4228), .B(n3131), .S(EBX_REG_21__SCAN_IN), .Z(n4207) );
  INV_X1 U5206 ( .A(n4207), .ZN(n4209) );
  NAND2_X1 U5207 ( .A1(n4498), .A2(n6925), .ZN(n4208) );
  NAND2_X1 U5208 ( .A1(n4209), .A2(n4208), .ZN(n5154) );
  INV_X1 U5209 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U5210 ( .A1(n4228), .A2(n5342), .ZN(n4213) );
  NAND2_X1 U5211 ( .A1(n4349), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4211) );
  OAI211_X1 U5212 ( .C1(EBX_REG_23__SCAN_IN), .C2(n4145), .A(n4211), .B(n4210), 
        .ZN(n4212) );
  AND2_X1 U5213 ( .A1(n4213), .A2(n4212), .ZN(n5128) );
  MUX2_X1 U5214 ( .A(n5169), .B(n4220), .S(EBX_REG_22__SCAN_IN), .Z(n4214) );
  INV_X1 U5215 ( .A(n4214), .ZN(n4216) );
  NAND2_X1 U5216 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4215) );
  NAND2_X1 U5217 ( .A1(n4216), .A2(n4215), .ZN(n5143) );
  AND2_X2 U5218 ( .A1(n5126), .A2(n3135), .ZN(n5099) );
  MUX2_X1 U5219 ( .A(n4228), .B(n5169), .S(EBX_REG_25__SCAN_IN), .Z(n4217) );
  INV_X1 U5220 ( .A(n4217), .ZN(n4219) );
  INV_X1 U5221 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U5222 ( .A1(n4498), .A2(n6866), .ZN(n4218) );
  NAND2_X1 U5223 ( .A1(n4219), .A2(n4218), .ZN(n5100) );
  MUX2_X1 U5224 ( .A(n3131), .B(n4220), .S(EBX_REG_24__SCAN_IN), .Z(n4222) );
  AND2_X1 U5225 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4221)
         );
  NOR2_X1 U5226 ( .A1(n4222), .A2(n4221), .ZN(n5115) );
  NOR2_X1 U5227 ( .A1(n5100), .A2(n5115), .ZN(n4223) );
  NAND2_X1 U5228 ( .A1(n4210), .A2(n4224), .ZN(n4225) );
  OAI211_X1 U5229 ( .C1(n4145), .C2(EBX_REG_26__SCAN_IN), .A(n4225), .B(n4349), 
        .ZN(n4227) );
  INV_X1 U5230 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U5231 ( .A1(n5169), .A2(n6827), .ZN(n4226) );
  NAND2_X1 U5232 ( .A1(n4227), .A2(n4226), .ZN(n5082) );
  NAND2_X1 U5233 ( .A1(n5081), .A2(n5082), .ZN(n5068) );
  MUX2_X1 U5234 ( .A(n4228), .B(n3131), .S(EBX_REG_27__SCAN_IN), .Z(n4229) );
  INV_X1 U5235 ( .A(n4229), .ZN(n4231) );
  INV_X1 U5236 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U5237 ( .A1(n4498), .A2(n5667), .ZN(n4230) );
  NAND2_X1 U5238 ( .A1(n4231), .A2(n4230), .ZN(n5069) );
  OR2_X2 U5239 ( .A1(n5068), .A2(n5069), .ZN(n5071) );
  NAND2_X1 U5240 ( .A1(n4210), .A2(n4232), .ZN(n4233) );
  OAI211_X1 U5241 ( .C1(n4145), .C2(EBX_REG_28__SCAN_IN), .A(n4233), .B(n4349), 
        .ZN(n4235) );
  INV_X1 U5242 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U5243 ( .A1(n3131), .A2(n5338), .ZN(n4234) );
  AND2_X1 U5244 ( .A1(n4235), .A2(n4234), .ZN(n5056) );
  NOR2_X4 U5245 ( .A1(n5071), .A2(n5056), .ZN(n5058) );
  OAI22_X1 U5246 ( .A1(n4356), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4145), .ZN(n4350) );
  AOI22_X1 U5247 ( .A1(n4356), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n4145), .ZN(n4354) );
  NAND2_X1 U5248 ( .A1(n4126), .A2(n4467), .ZN(n4614) );
  OR2_X1 U5249 ( .A1(n4240), .A2(n4239), .ZN(n4241) );
  AND2_X1 U5250 ( .A1(n4614), .A2(n4241), .ZN(n4242) );
  INV_X1 U5251 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6797) );
  NOR2_X1 U5252 ( .A1(n6498), .A2(n6797), .ZN(n4397) );
  INV_X1 U5253 ( .A(n4397), .ZN(n4265) );
  NAND2_X1 U5254 ( .A1(n4661), .A2(n7068), .ZN(n4243) );
  AOI21_X1 U5255 ( .B1(n3094), .B2(n4256), .A(n4243), .ZN(n4244) );
  AOI21_X1 U5256 ( .B1(n4356), .B2(n4245), .A(n4244), .ZN(n4247) );
  OAI211_X1 U5257 ( .C1(n3674), .C2(n4349), .A(n4247), .B(n4246), .ZN(n4248)
         );
  INV_X1 U5258 ( .A(n4248), .ZN(n4249) );
  NAND2_X1 U5259 ( .A1(n4250), .A2(n4249), .ZN(n4439) );
  OAI21_X1 U5260 ( .B1(n4251), .B2(n3510), .A(n4569), .ZN(n4252) );
  NOR2_X1 U5261 ( .A1(n4439), .A2(n4252), .ZN(n4253) );
  INV_X1 U5262 ( .A(n4340), .ZN(n4431) );
  NAND2_X1 U5263 ( .A1(n4431), .A2(n7068), .ZN(n4571) );
  NAND2_X2 U5264 ( .A1(n4976), .A2(n6521), .ZN(n4969) );
  INV_X1 U5265 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U5266 ( .A1(n6523), .A2(n6521), .ZN(n4543) );
  NAND2_X1 U5267 ( .A1(n4969), .A2(n4543), .ZN(n4279) );
  INV_X2 U5268 ( .A(n4279), .ZN(n6495) );
  NOR2_X1 U5269 ( .A1(n4146), .A2(n4542), .ZN(n6497) );
  NOR2_X1 U5270 ( .A1(n6837), .A2(n4255), .ZN(n4260) );
  NAND4_X1 U5271 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6497), .A4(n4260), .ZN(n4968) );
  NOR2_X1 U5272 ( .A1(n5822), .A2(n5815), .ZN(n5813) );
  NAND3_X1 U5273 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5813), .ZN(n4970) );
  NOR2_X1 U5274 ( .A1(n4968), .A2(n4970), .ZN(n4984) );
  OR2_X1 U5275 ( .A1(n5297), .A2(n4256), .ZN(n4257) );
  NAND2_X1 U5276 ( .A1(n4258), .A2(n4257), .ZN(n4453) );
  AOI21_X1 U5277 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4739) );
  INV_X1 U5278 ( .A(n4260), .ZN(n4891) );
  NOR2_X1 U5279 ( .A1(n4739), .A2(n4891), .ZN(n4889) );
  NAND3_X1 U5280 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4889), .ZN(n5806) );
  NOR2_X1 U5281 ( .A1(n4970), .A2(n5806), .ZN(n4268) );
  NAND2_X1 U5282 ( .A1(n6496), .A2(n4268), .ZN(n4978) );
  NAND2_X2 U5283 ( .A1(n5795), .A2(n4978), .ZN(n6482) );
  NAND3_X1 U5284 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n4971) );
  INV_X1 U5285 ( .A(n4971), .ZN(n5767) );
  AND2_X1 U5286 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5767), .ZN(n5763)
         );
  AND2_X1 U5287 ( .A1(n5763), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5769)
         );
  NAND2_X1 U5288 ( .A1(n5769), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5757) );
  NOR2_X1 U5289 ( .A1(n5757), .A2(n6942), .ZN(n4261) );
  NAND2_X1 U5290 ( .A1(n6482), .A2(n4261), .ZN(n5749) );
  NOR2_X2 U5291 ( .A1(n5749), .A2(n5728), .ZN(n5744) );
  NAND2_X1 U5292 ( .A1(n5744), .A2(n5723), .ZN(n5722) );
  INV_X1 U5293 ( .A(n5467), .ZN(n5469) );
  OR2_X2 U5294 ( .A1(n3132), .A2(n5473), .ZN(n5687) );
  NAND2_X1 U5295 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5678) );
  INV_X1 U5296 ( .A(n5653), .ZN(n4262) );
  NAND2_X1 U5297 ( .A1(n5666), .A2(n4262), .ZN(n5005) );
  INV_X1 U5298 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6843) );
  INV_X1 U5299 ( .A(n4263), .ZN(n4264) );
  OAI211_X1 U5300 ( .C1(n4960), .C2(n6500), .A(n4265), .B(n4264), .ZN(n4266)
         );
  INV_X1 U5301 ( .A(n4266), .ZN(n4283) );
  NAND2_X1 U5302 ( .A1(n5796), .A2(n4976), .ZN(n4973) );
  INV_X1 U5303 ( .A(n6521), .ZN(n4972) );
  OR2_X1 U5304 ( .A1(n5722), .A2(n5467), .ZN(n4278) );
  NAND2_X1 U5305 ( .A1(n4267), .A2(n6498), .ZN(n6522) );
  OAI21_X1 U5306 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n4976), .A(n6522), 
        .ZN(n4966) );
  INV_X1 U5307 ( .A(n4969), .ZN(n4270) );
  OAI22_X1 U5308 ( .A1(n5796), .A2(n4268), .B1(n4270), .B2(n4984), .ZN(n4272)
         );
  INV_X1 U5309 ( .A(n5757), .ZN(n4269) );
  AOI21_X1 U5310 ( .B1(n5796), .B2(n4270), .A(n4269), .ZN(n4271) );
  OR2_X1 U5311 ( .A1(n4272), .A2(n4271), .ZN(n4273) );
  OR2_X1 U5312 ( .A1(n4966), .A2(n4273), .ZN(n5760) );
  INV_X1 U5313 ( .A(n4274), .ZN(n4275) );
  NAND2_X1 U5314 ( .A1(n4275), .A2(n5723), .ZN(n4276) );
  AND2_X1 U5315 ( .A1(n5765), .A2(n4276), .ZN(n4277) );
  NOR2_X1 U5316 ( .A1(n5760), .A2(n4277), .ZN(n5715) );
  NAND2_X1 U5317 ( .A1(n4278), .A2(n5715), .ZN(n5710) );
  NAND2_X1 U5318 ( .A1(n5796), .A2(n4279), .ZN(n5725) );
  AND2_X1 U5319 ( .A1(n5725), .A2(n5473), .ZN(n4280) );
  AND2_X1 U5320 ( .A1(n5765), .A2(n5678), .ZN(n4281) );
  NOR2_X1 U5321 ( .A1(n5697), .A2(n4281), .ZN(n5668) );
  NAND2_X1 U5322 ( .A1(n5765), .A2(n5653), .ZN(n4282) );
  NAND2_X1 U5323 ( .A1(n5668), .A2(n4282), .ZN(n4389) );
  AOI21_X1 U5324 ( .B1(n5765), .B2(n6843), .A(n4389), .ZN(n5008) );
  NAND2_X1 U5325 ( .A1(n4285), .A2(n4284), .ZN(U2988) );
  NOR2_X1 U5326 ( .A1(n4287), .A2(n4286), .ZN(n4310) );
  AOI22_X1 U5327 ( .A1(n3358), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U5328 ( .A1(n4288), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3096), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4294) );
  AOI22_X1 U5329 ( .A1(n4290), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4289), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U5330 ( .A1(n4291), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4292) );
  NAND4_X1 U5331 ( .A1(n4295), .A2(n4294), .A3(n4293), .A4(n4292), .ZN(n4302)
         );
  AOI22_X1 U5332 ( .A1(n3442), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4300) );
  AOI22_X1 U5333 ( .A1(n3095), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U5334 ( .A1(n3360), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4298) );
  AOI22_X1 U5335 ( .A1(n4314), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4297) );
  NAND4_X1 U5336 ( .A1(n4300), .A2(n4299), .A3(n4298), .A4(n4297), .ZN(n4301)
         );
  OR2_X1 U5337 ( .A1(n4302), .A2(n4301), .ZN(n4309) );
  XOR2_X1 U5338 ( .A(n4310), .B(n4309), .Z(n4306) );
  INV_X1 U5339 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4303) );
  INV_X1 U5340 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5014) );
  OAI22_X1 U5341 ( .A1(n3687), .A2(n4303), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5014), .ZN(n4304) );
  AOI21_X1 U5342 ( .B1(n4306), .B2(n4305), .A(n4304), .ZN(n4307) );
  XNOR2_X1 U5343 ( .A(n4333), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5047)
         );
  MUX2_X1 U5344 ( .A(n4307), .B(n5047), .S(n4334), .Z(n5012) );
  NAND2_X1 U5345 ( .A1(n4310), .A2(n4309), .ZN(n4329) );
  AOI22_X1 U5346 ( .A1(n4311), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4318) );
  AOI22_X1 U5347 ( .A1(n4313), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4312), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4317) );
  AOI22_X1 U5348 ( .A1(n4314), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4316) );
  AOI22_X1 U5349 ( .A1(n3096), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4315) );
  NAND4_X1 U5350 ( .A1(n4318), .A2(n4317), .A3(n4316), .A4(n4315), .ZN(n4327)
         );
  AOI22_X1 U5351 ( .A1(n4319), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4291), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U5352 ( .A1(n3442), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U5353 ( .A1(n4069), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4296), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U5354 ( .A1(n4070), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4321), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4322) );
  NAND4_X1 U5355 ( .A1(n4325), .A2(n4324), .A3(n4323), .A4(n4322), .ZN(n4326)
         );
  NOR2_X1 U5356 ( .A1(n4327), .A2(n4326), .ZN(n4328) );
  XNOR2_X1 U5357 ( .A(n4329), .B(n4328), .ZN(n4332) );
  AOI22_X1 U5358 ( .A1(n4337), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6782), .ZN(n4330) );
  OAI21_X1 U5359 ( .B1(n4332), .B2(n4331), .A(n4330), .ZN(n4335) );
  XNOR2_X1 U5360 ( .A(n4345), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5028)
         );
  MUX2_X1 U5361 ( .A(n4335), .B(n5028), .S(n4334), .Z(n4395) );
  AOI22_X1 U5362 ( .A1(n4337), .A2(EAX_REG_31__SCAN_IN), .B1(n4336), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4338) );
  INV_X1 U5363 ( .A(n4338), .ZN(n4339) );
  NAND2_X1 U5364 ( .A1(n4126), .A2(n5023), .ZN(n4426) );
  NOR2_X1 U5365 ( .A1(n4340), .A2(n4430), .ZN(n4422) );
  NAND2_X1 U5366 ( .A1(n4422), .A2(n4636), .ZN(n6230) );
  NAND2_X1 U5367 ( .A1(n4647), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4341) );
  OR2_X1 U5368 ( .A1(n4342), .A2(n4341), .ZN(n6648) );
  NOR2_X1 U5369 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6741) );
  AND2_X1 U5370 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n4343) );
  NAND2_X1 U5371 ( .A1(n6741), .A2(n4343), .ZN(n4633) );
  NAND2_X1 U5372 ( .A1(n6648), .A2(n4633), .ZN(n4344) );
  INV_X1 U5373 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4346) );
  XNOR2_X2 U5374 ( .A(n4347), .B(n4346), .ZN(n5039) );
  AND2_X1 U5375 ( .A1(n5169), .A2(EBX_REG_29__SCAN_IN), .ZN(n4351) );
  AOI21_X1 U5376 ( .B1(n4350), .B2(n4349), .A(n4351), .ZN(n4385) );
  NAND2_X1 U5377 ( .A1(n5058), .A2(n4385), .ZN(n4387) );
  INV_X1 U5378 ( .A(n5058), .ZN(n4352) );
  AOI21_X1 U5379 ( .B1(n4352), .B2(n5169), .A(n4351), .ZN(n4353) );
  OAI21_X1 U5380 ( .B1(n4387), .B2(n4354), .A(n4353), .ZN(n4355) );
  OAI22_X1 U5381 ( .A1(n4356), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4145), .ZN(n4357) );
  INV_X1 U5382 ( .A(n5299), .ZN(n4361) );
  NOR2_X1 U5383 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5022) );
  INV_X1 U5384 ( .A(n5022), .ZN(n4375) );
  NAND3_X1 U5385 ( .A1(n4519), .A2(EBX_REG_31__SCAN_IN), .A3(n4375), .ZN(n4360) );
  NOR2_X2 U5386 ( .A1(n4361), .A2(n4360), .ZN(n6366) );
  OR2_X1 U5387 ( .A1(n4657), .A2(n4462), .ZN(n4362) );
  AOI21_X1 U5388 ( .B1(n4145), .B2(n4362), .A(n4375), .ZN(n4364) );
  INV_X1 U5389 ( .A(REIP_REG_14__SCAN_IN), .ZN(n7025) );
  INV_X1 U5390 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6971) );
  INV_X1 U5391 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5272) );
  INV_X1 U5392 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6675) );
  INV_X1 U5393 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6665) );
  NAND3_X1 U5394 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6359) );
  NOR2_X1 U5395 ( .A1(n6665), .A2(n6359), .ZN(n6328) );
  NAND2_X1 U5396 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6328), .ZN(n6318) );
  NAND2_X1 U5397 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n6330) );
  NOR2_X1 U5398 ( .A1(n6318), .A2(n6330), .ZN(n6307) );
  NAND2_X1 U5399 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6307), .ZN(n5284) );
  NOR2_X1 U5400 ( .A1(n6675), .A2(n5284), .ZN(n6299) );
  NAND2_X1 U5401 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6299), .ZN(n5271) );
  NOR2_X1 U5402 ( .A1(n5272), .A2(n5271), .ZN(n5269) );
  NAND2_X1 U5403 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5269), .ZN(n6275) );
  OR2_X1 U5404 ( .A1(n6971), .A2(n6275), .ZN(n6263) );
  NOR2_X1 U5405 ( .A1(n7025), .A2(n6263), .ZN(n4365) );
  NAND4_X1 U5406 ( .A1(n5237), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(REIP_REG_17__SCAN_IN), .ZN(n5204) );
  INV_X1 U5407 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6685) );
  AND2_X1 U5408 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n4367) );
  NAND3_X1 U5409 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4371) );
  INV_X1 U5410 ( .A(n4371), .ZN(n5098) );
  NAND2_X1 U5411 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5088) );
  INV_X1 U5412 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5449) );
  NOR2_X1 U5413 ( .A1(n5088), .A2(n5449), .ZN(n4370) );
  NAND2_X1 U5414 ( .A1(n5087), .A2(n4370), .ZN(n5074) );
  NAND2_X1 U5415 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4374) );
  INV_X1 U5416 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6703) );
  NAND3_X1 U5417 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_17__SCAN_IN), .ZN(n4366) );
  NAND2_X1 U5418 ( .A1(n4365), .A2(n5293), .ZN(n5235) );
  NOR2_X1 U5419 ( .A1(n4366), .A2(n5235), .ZN(n5223) );
  INV_X1 U5420 ( .A(n4367), .ZN(n4368) );
  NOR2_X1 U5421 ( .A1(n4368), .A2(n6685), .ZN(n4369) );
  AND2_X1 U5422 ( .A1(n5223), .A2(n4369), .ZN(n5142) );
  INV_X1 U5423 ( .A(n4370), .ZN(n4372) );
  NOR2_X1 U5424 ( .A1(n4372), .A2(n4371), .ZN(n4373) );
  NAND2_X1 U5425 ( .A1(n6360), .A2(n5293), .ZN(n5236) );
  AOI21_X1 U5426 ( .B1(n5142), .B2(n4373), .A(n5326), .ZN(n5089) );
  AOI21_X1 U5427 ( .B1(n6329), .B2(n4374), .A(n5089), .ZN(n5062) );
  OAI21_X1 U5428 ( .B1(REIP_REG_29__SCAN_IN), .B2(n6360), .A(n5062), .ZN(n5034) );
  AOI21_X1 U5429 ( .B1(n6329), .B2(n6797), .A(n5034), .ZN(n4378) );
  INV_X1 U5430 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6707) );
  NOR2_X1 U5431 ( .A1(n4462), .A2(n4375), .ZN(n4610) );
  NOR2_X1 U5432 ( .A1(n6740), .A2(n4610), .ZN(n4376) );
  AND2_X1 U5433 ( .A1(n5299), .A2(n4376), .ZN(n5021) );
  AOI22_X1 U5434 ( .A1(n5021), .A2(EBX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n6363), .ZN(n4377) );
  OAI21_X1 U5435 ( .B1(n4378), .B2(n6707), .A(n4377), .ZN(n4379) );
  AOI21_X1 U5436 ( .B1(n5333), .B2(n6366), .A(n4381), .ZN(n4382) );
  OR2_X1 U5437 ( .A1(n5058), .A2(n4385), .ZN(n4386) );
  NAND2_X1 U5438 ( .A1(n4387), .A2(n4386), .ZN(n5336) );
  OR2_X1 U5439 ( .A1(n5336), .A2(n6500), .ZN(n4388) );
  NAND2_X1 U5440 ( .A1(n6465), .A2(REIP_REG_29__SCAN_IN), .ZN(n5013) );
  OAI211_X1 U5441 ( .C1(n5005), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4388), .B(n5013), .ZN(n4391) );
  NAND2_X1 U5442 ( .A1(n4392), .A2(n6474), .ZN(n4401) );
  NOR2_X1 U5443 ( .A1(n6478), .A2(n5028), .ZN(n4396) );
  AOI211_X1 U5444 ( .C1(n6466), .C2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n4397), 
        .B(n4396), .ZN(n4398) );
  INV_X1 U5445 ( .A(n4399), .ZN(n4400) );
  NAND2_X1 U5446 ( .A1(n4401), .A2(n4400), .ZN(U2956) );
  NAND2_X1 U5447 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n4410) );
  INV_X1 U5448 ( .A(n4410), .ZN(n4402) );
  AOI21_X1 U5449 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n4402), .ZN(n4404) );
  NAND2_X1 U5450 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4409) );
  INV_X1 U5451 ( .A(n4409), .ZN(n4403) );
  INV_X1 U5452 ( .A(READY_N), .ZN(n6868) );
  INV_X1 U5453 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6975) );
  NOR2_X1 U5454 ( .A1(n6868), .A2(n6975), .ZN(n6656) );
  INV_X1 U5455 ( .A(n6656), .ZN(n4408) );
  OAI211_X1 U5456 ( .C1(n4404), .C2(n4403), .A(n4408), .B(n4462), .ZN(U3182)
         );
  AND2_X1 U5457 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n4644) );
  NAND2_X1 U5458 ( .A1(n4644), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5841) );
  INV_X1 U5459 ( .A(n5841), .ZN(n4456) );
  AOI21_X1 U5460 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6868), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4405) );
  NOR3_X1 U5461 ( .A1(n4456), .A2(n6741), .A3(n4405), .ZN(n4407) );
  OR2_X1 U5462 ( .A1(n4407), .A2(n4406), .ZN(U3150) );
  NAND2_X1 U5463 ( .A1(n4409), .A2(n4408), .ZN(n4413) );
  NAND2_X1 U5464 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n4412) );
  NOR2_X2 U5465 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6975), .ZN(n6746) );
  AOI21_X1 U5466 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(n4410), .A(n6746), 
        .ZN(n4411) );
  INV_X1 U5467 ( .A(NA_N), .ZN(n6815) );
  AOI221_X1 U5468 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6815), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6659) );
  AOI211_X1 U5469 ( .C1(n4413), .C2(n4412), .A(n4411), .B(n6659), .ZN(n4414)
         );
  INV_X1 U5470 ( .A(n4414), .ZN(U3181) );
  NOR2_X1 U5471 ( .A1(n5998), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5189) );
  INV_X1 U5472 ( .A(n5189), .ZN(n4415) );
  NAND2_X1 U5473 ( .A1(n4465), .A2(n4415), .ZN(n6229) );
  INV_X1 U5474 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n4416) );
  NAND2_X1 U5475 ( .A1(n6230), .A2(n4416), .ZN(n4418) );
  NAND2_X1 U5476 ( .A1(n6740), .A2(n5297), .ZN(n4425) );
  NAND2_X1 U5477 ( .A1(n6738), .A2(n4425), .ZN(n4417) );
  OAI21_X1 U5478 ( .B1(n6229), .B2(n4418), .A(n4417), .ZN(n4419) );
  INV_X1 U5479 ( .A(n4419), .ZN(U3474) );
  INV_X1 U5480 ( .A(n4420), .ZN(n4424) );
  INV_X1 U5481 ( .A(n4421), .ZN(n5291) );
  INV_X1 U5482 ( .A(n4426), .ZN(n4423) );
  OAI22_X1 U5483 ( .A1(n4424), .A2(n5291), .B1(n4423), .B2(n4422), .ZN(n6240)
         );
  AOI21_X1 U5484 ( .B1(n4425), .B2(n4462), .A(READY_N), .ZN(n6739) );
  NOR2_X1 U5485 ( .A1(n6240), .A2(n6739), .ZN(n4595) );
  NOR2_X1 U5486 ( .A1(n4595), .A2(n6646), .ZN(n6247) );
  INV_X1 U5487 ( .A(MORE_REG_SCAN_IN), .ZN(n4434) );
  INV_X1 U5488 ( .A(n4556), .ZN(n4428) );
  NAND3_X1 U5489 ( .A1(n4426), .A2(n4597), .A3(n4555), .ZN(n4427) );
  MUX2_X1 U5490 ( .A(n4428), .B(n4427), .S(n4420), .Z(n4429) );
  AOI21_X1 U5491 ( .B1(n4431), .B2(n4430), .A(n4429), .ZN(n4598) );
  INV_X1 U5492 ( .A(n4598), .ZN(n4432) );
  NAND2_X1 U5493 ( .A1(n6247), .A2(n4432), .ZN(n4433) );
  OAI21_X1 U5494 ( .B1(n6247), .B2(n4434), .A(n4433), .ZN(U3471) );
  INV_X1 U5495 ( .A(n4436), .ZN(n4799) );
  INV_X1 U5496 ( .A(n4126), .ZN(n4438) );
  NAND3_X1 U5497 ( .A1(n4698), .A2(n4661), .A3(n4724), .ZN(n4505) );
  NAND4_X1 U5498 ( .A1(n4438), .A2(n4437), .A3(n4593), .A4(n4505), .ZN(n4440)
         );
  OR2_X1 U5499 ( .A1(n4440), .A2(n4439), .ZN(n4580) );
  NAND2_X1 U5500 ( .A1(n4799), .A2(n4580), .ZN(n4444) );
  OAI21_X1 U5501 ( .B1(n4441), .B2(n4442), .A(n4579), .ZN(n4443) );
  OAI211_X1 U5502 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4571), .A(n4444), .B(n4443), .ZN(n4582) );
  INV_X1 U5503 ( .A(n6722), .ZN(n6234) );
  NAND2_X1 U5504 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4941) );
  INV_X1 U5505 ( .A(n4941), .ZN(n4446) );
  INV_X1 U5506 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U5507 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4445), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4542), .ZN(n4940) );
  INV_X1 U5508 ( .A(n6712), .ZN(n4937) );
  AOI222_X1 U5509 ( .A1(n4582), .A2(n6234), .B1(n4446), .B2(n4940), .C1(n4442), 
        .C2(n4937), .ZN(n4461) );
  INV_X1 U5510 ( .A(n4571), .ZN(n4581) );
  INV_X1 U5511 ( .A(n4462), .ZN(n4447) );
  OAI21_X1 U5512 ( .B1(n4581), .B2(n4126), .A(n4447), .ZN(n4448) );
  NAND2_X1 U5513 ( .A1(n4448), .A2(n4468), .ZN(n4450) );
  INV_X1 U5514 ( .A(n4555), .ZN(n4449) );
  AOI21_X1 U5515 ( .B1(n4450), .B2(n6868), .A(n4449), .ZN(n4451) );
  MUX2_X1 U5516 ( .A(n4451), .B(n4556), .S(n4420), .Z(n4455) );
  AND2_X1 U5517 ( .A1(n6235), .A2(n4452), .ZN(n4523) );
  NOR2_X1 U5518 ( .A1(n4453), .A2(n4523), .ZN(n4454) );
  NAND2_X1 U5519 ( .A1(n4455), .A2(n4454), .ZN(n4592) );
  NAND2_X1 U5520 ( .A1(n4592), .A2(n4636), .ZN(n6232) );
  NAND2_X1 U5521 ( .A1(n4456), .A2(FLUSH_REG_SCAN_IN), .ZN(n4458) );
  NAND2_X1 U5522 ( .A1(n4647), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4457) );
  AND2_X1 U5523 ( .A1(n4458), .A2(n4457), .ZN(n4459) );
  NAND2_X1 U5524 ( .A1(n6232), .A2(n4459), .ZN(n6720) );
  INV_X1 U5525 ( .A(n6720), .ZN(n6715) );
  OAI21_X1 U5526 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6712), .A(n6720), 
        .ZN(n6718) );
  INV_X1 U5527 ( .A(n6718), .ZN(n4460) );
  OAI22_X1 U5528 ( .A1(n4461), .A2(n6715), .B1(n3635), .B2(n4460), .ZN(U3460)
         );
  AND2_X1 U5529 ( .A1(n4614), .A2(n4571), .ZN(n4463) );
  NOR2_X1 U5530 ( .A1(n6418), .A2(n4657), .ZN(n6394) );
  NAND2_X1 U5531 ( .A1(n4644), .A2(n4647), .ZN(n6735) );
  INV_X1 U5532 ( .A(n6735), .ZN(n6411) );
  AOI222_X1 U5533 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6394), .B1(n6413), .B2(
        DATAO_REG_30__SCAN_IN), .C1(n6411), .C2(UWORD_REG_14__SCAN_IN), .ZN(
        n4464) );
  INV_X1 U5534 ( .A(n4464), .ZN(U2893) );
  INV_X1 U5535 ( .A(n4465), .ZN(n4466) );
  INV_X1 U5536 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6834) );
  OR2_X1 U5537 ( .A1(n4525), .A2(n4614), .ZN(n6464) );
  INV_X2 U5538 ( .A(n6464), .ZN(n7061) );
  INV_X1 U5539 ( .A(DATAI_12_), .ZN(n4469) );
  NOR2_X1 U5540 ( .A1(n7065), .A2(n4469), .ZN(n6455) );
  AOI21_X1 U5541 ( .B1(n7061), .B2(EAX_REG_28__SCAN_IN), .A(n6455), .ZN(n4470)
         );
  OAI21_X1 U5542 ( .B1(n6420), .B2(n6834), .A(n4470), .ZN(U2936) );
  INV_X1 U5543 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n7010) );
  INV_X1 U5544 ( .A(DATAI_10_), .ZN(n4471) );
  NOR2_X1 U5545 ( .A1(n7065), .A2(n4471), .ZN(n6451) );
  AOI21_X1 U5546 ( .B1(n7061), .B2(EAX_REG_26__SCAN_IN), .A(n6451), .ZN(n4472)
         );
  OAI21_X1 U5547 ( .B1(n7010), .B2(n6420), .A(n4472), .ZN(U2934) );
  INV_X1 U5548 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6862) );
  INV_X1 U5549 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4473) );
  OAI222_X1 U5550 ( .A1(n6419), .A2(n6862), .B1(n4496), .B2(n4473), .C1(n6735), 
        .C2(n7010), .ZN(U2897) );
  INV_X1 U5551 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4476) );
  INV_X1 U5552 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4475) );
  INV_X1 U5553 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4474) );
  OAI222_X1 U5554 ( .A1(n4476), .A2(n6419), .B1(n4496), .B2(n4475), .C1(n6735), 
        .C2(n4474), .ZN(U2901) );
  INV_X1 U5555 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4479) );
  INV_X1 U5556 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4478) );
  INV_X1 U5557 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4477) );
  OAI222_X1 U5558 ( .A1(n4479), .A2(n6419), .B1(n4496), .B2(n4478), .C1(n6735), 
        .C2(n4477), .ZN(U2907) );
  INV_X1 U5559 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4482) );
  INV_X1 U5560 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4481) );
  INV_X1 U5561 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4480) );
  OAI222_X1 U5562 ( .A1(n4482), .A2(n6419), .B1(n4496), .B2(n4481), .C1(n6735), 
        .C2(n4480), .ZN(U2900) );
  INV_X1 U5563 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4484) );
  INV_X1 U5564 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n4483) );
  OAI222_X1 U5565 ( .A1(n4484), .A2(n6419), .B1(n4496), .B2(n4303), .C1(n6735), 
        .C2(n4483), .ZN(U2894) );
  INV_X1 U5566 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4486) );
  INV_X1 U5567 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n4485) );
  OAI222_X1 U5568 ( .A1(n4486), .A2(n6419), .B1(n4496), .B2(n4064), .C1(n6735), 
        .C2(n4485), .ZN(U2896) );
  INV_X1 U5569 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4488) );
  INV_X1 U5570 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4487) );
  OAI222_X1 U5571 ( .A1(n4488), .A2(n6419), .B1(n4496), .B2(n3958), .C1(n6735), 
        .C2(n4487), .ZN(U2899) );
  INV_X1 U5572 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4491) );
  INV_X1 U5573 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4490) );
  INV_X1 U5574 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4489) );
  OAI222_X1 U5575 ( .A1(n4491), .A2(n6419), .B1(n4496), .B2(n4490), .C1(n6735), 
        .C2(n4489), .ZN(U2906) );
  INV_X1 U5576 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4493) );
  INV_X1 U5577 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4492) );
  OAI222_X1 U5578 ( .A1(n4493), .A2(n6419), .B1(n4496), .B2(n4011), .C1(n6735), 
        .C2(n4492), .ZN(U2904) );
  INV_X1 U5579 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4497) );
  INV_X1 U5580 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4495) );
  INV_X1 U5581 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4494) );
  OAI222_X1 U5582 ( .A1(n4497), .A2(n6419), .B1(n4496), .B2(n4495), .C1(n6735), 
        .C2(n4494), .ZN(U2902) );
  NAND2_X1 U5583 ( .A1(n4498), .A2(n6523), .ZN(n4500) );
  AND2_X1 U5584 ( .A1(n4500), .A2(n4499), .ZN(n6519) );
  INV_X1 U5585 ( .A(n6519), .ZN(n4513) );
  NOR2_X1 U5586 ( .A1(n4556), .A2(n6646), .ZN(n4501) );
  NAND2_X1 U5587 ( .A1(n4420), .A2(n4501), .ZN(n4508) );
  INV_X1 U5588 ( .A(n4512), .ZN(n5386) );
  NAND4_X1 U5589 ( .A1(n4504), .A2(n5386), .A3(n4503), .A4(n4502), .ZN(n4506)
         );
  NOR2_X1 U5590 ( .A1(n4506), .A2(n4505), .ZN(n4522) );
  NAND2_X1 U5591 ( .A1(n4522), .A2(n4519), .ZN(n4507) );
  NAND2_X2 U5592 ( .A1(n5381), .A2(n5386), .ZN(n5382) );
  INV_X2 U5593 ( .A(n5373), .ZN(n5381) );
  INV_X1 U5594 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6981) );
  OAI21_X1 U5595 ( .B1(n4511), .B2(n4510), .A(n4509), .ZN(n5644) );
  INV_X2 U5596 ( .A(n6379), .ZN(n5375) );
  OAI222_X1 U5597 ( .A1(n4513), .A2(n5382), .B1(n5381), .B2(n6981), .C1(n5644), 
        .C2(n5375), .ZN(U2859) );
  OR2_X1 U5598 ( .A1(n4515), .A2(n4514), .ZN(n4516) );
  NAND2_X1 U5599 ( .A1(n3113), .A2(n4516), .ZN(n5325) );
  INV_X1 U5600 ( .A(n5382), .ZN(n6378) );
  OAI21_X1 U5601 ( .B1(n4520), .B2(n4519), .A(n4518), .ZN(n5320) );
  AOI22_X1 U5602 ( .A1(n6378), .A2(n5320), .B1(n5373), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4521) );
  OAI21_X1 U5603 ( .B1(n5325), .B2(n5375), .A(n4521), .ZN(U2858) );
  AOI22_X1 U5604 ( .A1(n4523), .A2(n4636), .B1(n5291), .B2(n4522), .ZN(n4524)
         );
  OR2_X1 U5605 ( .A1(n4115), .A2(n5386), .ZN(n4526) );
  INV_X1 U5606 ( .A(n4526), .ZN(n4527) );
  INV_X1 U5607 ( .A(DATAI_1_), .ZN(n6438) );
  INV_X1 U5608 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4528) );
  OAI222_X1 U5609 ( .A1(n5325), .A2(n5438), .B1(n5437), .B2(n6438), .C1(n5436), 
        .C2(n4528), .ZN(U2890) );
  INV_X1 U5610 ( .A(DATAI_0_), .ZN(n6436) );
  INV_X1 U5611 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6417) );
  OAI222_X1 U5612 ( .A1(n5644), .A2(n5438), .B1(n5437), .B2(n6436), .C1(n5436), 
        .C2(n6417), .ZN(U2891) );
  NOR2_X1 U5613 ( .A1(n4530), .A2(n4529), .ZN(n4531) );
  NOR2_X1 U5614 ( .A1(n4618), .A2(n4531), .ZN(n6473) );
  NAND2_X1 U5615 ( .A1(n4534), .A2(n4533), .ZN(n4535) );
  NAND2_X1 U5616 ( .A1(n4532), .A2(n4535), .ZN(n6499) );
  OAI22_X1 U5617 ( .A1(n5382), .A2(n6499), .B1(n4536), .B2(n5381), .ZN(n4537)
         );
  AOI21_X1 U5618 ( .B1(n6473), .B2(n6379), .A(n4537), .ZN(n4538) );
  INV_X1 U5619 ( .A(n4538), .ZN(U2857) );
  NAND2_X1 U5620 ( .A1(n6523), .A2(n4973), .ZN(n6511) );
  AOI21_X1 U5621 ( .B1(n6522), .B2(n6511), .A(n4542), .ZN(n4548) );
  OAI21_X1 U5622 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n4749) );
  NAND3_X1 U5623 ( .A1(n5765), .A2(n4543), .A3(n4542), .ZN(n4546) );
  INV_X1 U5624 ( .A(REIP_REG_1__SCAN_IN), .ZN(n4544) );
  NOR2_X1 U5625 ( .A1(n6498), .A2(n4544), .ZN(n4745) );
  AOI21_X1 U5626 ( .B1(n6518), .B2(n5320), .A(n4745), .ZN(n4545) );
  OAI211_X1 U5627 ( .C1(n4749), .C2(n6515), .A(n4546), .B(n4545), .ZN(n4547)
         );
  OR2_X1 U5628 ( .A1(n4548), .A2(n4547), .ZN(U3017) );
  INV_X1 U5629 ( .A(n6473), .ZN(n5317) );
  INV_X1 U5630 ( .A(DATAI_2_), .ZN(n6440) );
  INV_X1 U5631 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4549) );
  OAI222_X1 U5632 ( .A1(n5317), .A2(n5438), .B1(n5437), .B2(n6440), .C1(n5436), 
        .C2(n4549), .ZN(U2889) );
  CLKBUF_X1 U5633 ( .A(n4553), .Z(n4939) );
  MUX2_X1 U5634 ( .A(n4554), .B(n4566), .S(n4939), .Z(n4557) );
  NAND2_X1 U5635 ( .A1(n4556), .A2(n4555), .ZN(n4574) );
  OAI21_X1 U5636 ( .B1(n4552), .B2(n4557), .A(n4574), .ZN(n4564) );
  NAND2_X1 U5637 ( .A1(n4568), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4558) );
  AND2_X1 U5638 ( .A1(n4558), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4559)
         );
  OAI22_X1 U5639 ( .A1(n4552), .A2(n4559), .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4561) );
  AOI21_X1 U5640 ( .B1(n4939), .B2(n4568), .A(n4566), .ZN(n4560) );
  NOR2_X1 U5641 ( .A1(n3096), .A2(n4560), .ZN(n6713) );
  OAI22_X1 U5642 ( .A1(n4571), .A2(n4561), .B1(n6713), .B2(n4569), .ZN(n4562)
         );
  INV_X1 U5643 ( .A(n4562), .ZN(n4563) );
  NAND2_X1 U5644 ( .A1(n4564), .A2(n4563), .ZN(n4565) );
  AOI21_X1 U5645 ( .B1(n4551), .B2(n4580), .A(n4565), .ZN(n6714) );
  MUX2_X1 U5646 ( .A(n4566), .B(n6714), .S(n4592), .Z(n4605) );
  AOI21_X1 U5647 ( .B1(n4605), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U5648 ( .A1(n5848), .A2(n4580), .ZN(n4576) );
  XNOR2_X1 U5649 ( .A(n4939), .B(n4568), .ZN(n4573) );
  XNOR2_X1 U5650 ( .A(n4568), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4570)
         );
  OAI22_X1 U5651 ( .A1(n4571), .A2(n4570), .B1(n4569), .B2(n4573), .ZN(n4572)
         );
  AOI21_X1 U5652 ( .B1(n4574), .B2(n4573), .A(n4572), .ZN(n4575) );
  AND2_X1 U5653 ( .A1(n4576), .A2(n4575), .ZN(n4938) );
  MUX2_X1 U5654 ( .A(n4946), .B(n4938), .S(n4592), .Z(n4586) );
  INV_X1 U5655 ( .A(n4586), .ZN(n4600) );
  CLKBUF_X1 U5656 ( .A(n4577), .Z(n4578) );
  AOI22_X1 U5657 ( .A1(n5952), .A2(n4580), .B1(n4579), .B2(n4578), .ZN(n6717)
         );
  NAND2_X1 U5658 ( .A1(n4581), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6723) );
  NAND3_X1 U5659 ( .A1(n6717), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6723), .ZN(n4583) );
  NAND2_X1 U5660 ( .A1(n4583), .A2(n4756), .ZN(n4585) );
  OAI211_X1 U5661 ( .C1(n4756), .C2(n4583), .A(n4592), .B(n4582), .ZN(n4584)
         );
  OAI211_X1 U5662 ( .C1(n4586), .C2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n4585), .B(n4584), .ZN(n4587) );
  OAI21_X1 U5663 ( .B1(n4600), .B2(n7026), .A(n4587), .ZN(n4588) );
  OAI21_X1 U5664 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4605), .A(n4588), 
        .ZN(n4608) );
  INV_X1 U5665 ( .A(n4590), .ZN(n5951) );
  NOR2_X1 U5666 ( .A1(n4589), .A2(n5951), .ZN(n4591) );
  XNOR2_X1 U5667 ( .A(n4591), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6233)
         );
  OAI22_X1 U5668 ( .A1(n6233), .A2(n4593), .B1(n4592), .B2(n6238), .ZN(n4594)
         );
  NOR2_X1 U5669 ( .A1(n4599), .A2(FLUSH_REG_SCAN_IN), .ZN(n4602) );
  AOI22_X1 U5670 ( .A1(n4594), .A2(n4599), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4602), .ZN(n4631) );
  OAI21_X1 U5671 ( .B1(MORE_REG_SCAN_IN), .B2(FLUSH_REG_SCAN_IN), .A(n4595), 
        .ZN(n4596) );
  NAND4_X1 U5672 ( .A1(n4631), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4607)
         );
  NAND2_X1 U5673 ( .A1(n4600), .A2(n4599), .ZN(n4606) );
  INV_X1 U5674 ( .A(n4601), .ZN(n4604) );
  INV_X1 U5675 ( .A(n4602), .ZN(n4603) );
  OAI22_X1 U5676 ( .A1(n4606), .A2(n4605), .B1(n4604), .B2(n4603), .ZN(n4629)
         );
  AOI211_X1 U5677 ( .C1(n4609), .C2(n4608), .A(n4607), .B(n4629), .ZN(n4628)
         );
  AOI21_X1 U5678 ( .B1(n4628), .B2(n4599), .A(n4647), .ZN(n4615) );
  INV_X1 U5679 ( .A(n4610), .ZN(n4613) );
  AOI21_X1 U5680 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n4611) );
  INV_X1 U5681 ( .A(n4611), .ZN(n4612) );
  OAI211_X1 U5682 ( .C1(n4614), .C2(n4613), .A(STATE2_REG_2__SCAN_IN), .B(
        n4612), .ZN(n4626) );
  NOR2_X1 U5683 ( .A1(n4615), .A2(n4626), .ZN(n6645) );
  OAI21_X1 U5684 ( .B1(n6645), .B2(n4647), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4616) );
  NAND2_X1 U5685 ( .A1(n4616), .A2(n5841), .ZN(U3453) );
  NOR2_X1 U5686 ( .A1(n4618), .A2(n4617), .ZN(n4619) );
  OR2_X1 U5687 ( .A1(n4624), .A2(n4619), .ZN(n5308) );
  AOI21_X1 U5688 ( .B1(n4532), .B2(n4621), .A(n4620), .ZN(n5302) );
  AOI22_X1 U5689 ( .A1(n6378), .A2(n5302), .B1(n5373), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4622) );
  OAI21_X1 U5690 ( .B1(n5308), .B2(n5375), .A(n4622), .ZN(U2856) );
  INV_X1 U5691 ( .A(DATAI_3_), .ZN(n6442) );
  INV_X1 U5692 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6410) );
  OAI222_X1 U5693 ( .A1(n5308), .A2(n5438), .B1(n5437), .B2(n6442), .C1(n5436), 
        .C2(n6410), .ZN(U2888) );
  AND2_X1 U5694 ( .A1(n4624), .A2(n4623), .ZN(n4667) );
  NOR2_X1 U5695 ( .A1(n4624), .A2(n4623), .ZN(n4625) );
  INV_X1 U5696 ( .A(DATAI_4_), .ZN(n6444) );
  INV_X1 U5697 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6912) );
  OAI222_X1 U5698 ( .A1(n6371), .A2(n5438), .B1(n5437), .B2(n6444), .C1(n5436), 
        .C2(n6912), .ZN(U2887) );
  INV_X1 U5699 ( .A(n6741), .ZN(n4645) );
  OAI21_X1 U5700 ( .B1(n6712), .B2(n4645), .A(n4626), .ZN(n4627) );
  AOI21_X1 U5701 ( .B1(n6782), .B2(READY_N), .A(n6645), .ZN(n6643) );
  MUX2_X1 U5702 ( .A(n4627), .B(n6643), .S(STATE2_REG_0__SCAN_IN), .Z(n4638)
         );
  INV_X1 U5703 ( .A(n4628), .ZN(n4635) );
  INV_X1 U5704 ( .A(n4629), .ZN(n4632) );
  OAI21_X1 U5705 ( .B1(n4632), .B2(n4630), .A(n4631), .ZN(n5839) );
  OAI21_X1 U5706 ( .B1(n5839), .B2(n5841), .A(n4633), .ZN(n4634) );
  AOI21_X1 U5707 ( .B1(n4636), .B2(n4635), .A(n4634), .ZN(n4637) );
  NAND2_X1 U5708 ( .A1(n4638), .A2(n4637), .ZN(U3148) );
  NAND2_X1 U5709 ( .A1(n5852), .A2(n4640), .ZN(n5907) );
  NAND2_X1 U5710 ( .A1(n5906), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5847) );
  NOR2_X1 U5711 ( .A1(n5907), .A2(n5847), .ZN(n5854) );
  NAND2_X1 U5712 ( .A1(n5848), .A2(n4799), .ZN(n6528) );
  INV_X1 U5713 ( .A(n6528), .ZN(n6124) );
  NAND3_X1 U5714 ( .A1(n6070), .A2(n6124), .A3(n5952), .ZN(n4642) );
  NAND2_X1 U5715 ( .A1(n4642), .A2(n6595), .ZN(n4653) );
  INV_X1 U5716 ( .A(n4653), .ZN(n4643) );
  OAI22_X1 U5717 ( .A1(n4654), .A2(n4643), .B1(n6530), .B2(n6782), .ZN(n6598)
         );
  INV_X1 U5718 ( .A(n6598), .ZN(n4665) );
  INV_X1 U5719 ( .A(n4644), .ZN(n5838) );
  NAND2_X1 U5720 ( .A1(n4645), .A2(n5838), .ZN(n4646) );
  INV_X1 U5721 ( .A(DATAI_7_), .ZN(n6448) );
  OR2_X1 U5722 ( .A1(n5840), .A2(n6448), .ZN(n6114) );
  INV_X1 U5723 ( .A(n5907), .ZN(n4649) );
  NAND2_X1 U5724 ( .A1(n6472), .A2(DATAI_31_), .ZN(n6642) );
  INV_X1 U5725 ( .A(n6642), .ZN(n6571) );
  NAND2_X1 U5726 ( .A1(n5906), .A2(n5956), .ZN(n4650) );
  NAND2_X1 U5727 ( .A1(n6472), .A2(DATAI_23_), .ZN(n6633) );
  OAI22_X1 U5728 ( .A1(n6596), .A2(n6633), .B1(n6595), .B2(n6632), .ZN(n4651)
         );
  AOI21_X1 U5729 ( .B1(n6534), .B2(n6571), .A(n4651), .ZN(n4656) );
  NAND2_X1 U5730 ( .A1(n5998), .A2(n6530), .ZN(n4652) );
  OAI211_X1 U5731 ( .C1(n4654), .C2(n4653), .A(n6182), .B(n4652), .ZN(n6599)
         );
  NAND2_X1 U5732 ( .A1(n6599), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4655) );
  OAI211_X1 U5733 ( .C1(n4665), .C2(n6114), .A(n4656), .B(n4655), .ZN(U3083)
         );
  OR2_X1 U5734 ( .A1(n5840), .A2(n6436), .ZN(n6084) );
  NAND2_X1 U5735 ( .A1(n6472), .A2(DATAI_24_), .ZN(n6133) );
  INV_X1 U5736 ( .A(n6133), .ZN(n6539) );
  NAND2_X1 U5737 ( .A1(n6472), .A2(DATAI_16_), .ZN(n6542) );
  OR2_X1 U5738 ( .A1(n4725), .A2(n4657), .ZN(n6083) );
  OAI22_X1 U5739 ( .A1(n6596), .A2(n6542), .B1(n6595), .B2(n6083), .ZN(n4658)
         );
  AOI21_X1 U5740 ( .B1(n6534), .B2(n6539), .A(n4658), .ZN(n4660) );
  NAND2_X1 U5741 ( .A1(n6599), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4659) );
  OAI211_X1 U5742 ( .C1(n4665), .C2(n6084), .A(n4660), .B(n4659), .ZN(U3076)
         );
  OR2_X1 U5743 ( .A1(n5840), .A2(n6442), .ZN(n6096) );
  NAND2_X1 U5744 ( .A1(n6472), .A2(DATAI_27_), .ZN(n6616) );
  INV_X1 U5745 ( .A(n6616), .ZN(n6552) );
  NAND2_X1 U5746 ( .A1(n6472), .A2(DATAI_19_), .ZN(n6611) );
  OR2_X1 U5747 ( .A1(n4725), .A2(n4661), .ZN(n6610) );
  OAI22_X1 U5748 ( .A1(n6596), .A2(n6611), .B1(n6595), .B2(n6610), .ZN(n4662)
         );
  AOI21_X1 U5749 ( .B1(n6534), .B2(n6552), .A(n4662), .ZN(n4664) );
  NAND2_X1 U5750 ( .A1(n6599), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4663) );
  OAI211_X1 U5751 ( .C1(n4665), .C2(n6096), .A(n4664), .B(n4663), .ZN(U3079)
         );
  NAND2_X1 U5752 ( .A1(n4667), .A2(n4666), .ZN(n4790) );
  OAI21_X1 U5753 ( .B1(n4667), .B2(n4666), .A(n4790), .ZN(n6352) );
  CLKBUF_X1 U5754 ( .A(n4668), .Z(n4669) );
  INV_X1 U5755 ( .A(n4670), .ZN(n4671) );
  AOI21_X1 U5756 ( .B1(n4672), .B2(n4669), .A(n4671), .ZN(n6350) );
  AOI22_X1 U5757 ( .A1(n6378), .A2(n6350), .B1(EBX_REG_5__SCAN_IN), .B2(n5373), 
        .ZN(n4673) );
  OAI21_X1 U5758 ( .B1(n6352), .B2(n5375), .A(n4673), .ZN(U2854) );
  OR2_X1 U5759 ( .A1(n4620), .A2(n4674), .ZN(n4675) );
  NAND2_X1 U5760 ( .A1(n4669), .A2(n4675), .ZN(n6364) );
  INV_X1 U5761 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6932) );
  OAI222_X1 U5762 ( .A1(n6364), .A2(n5382), .B1(n5381), .B2(n6932), .C1(n5375), 
        .C2(n6371), .ZN(U2855) );
  NAND2_X1 U5763 ( .A1(n6472), .A2(DATAI_20_), .ZN(n6618) );
  NOR2_X1 U5764 ( .A1(n4683), .A2(n6120), .ZN(n4689) );
  INV_X1 U5765 ( .A(n5855), .ZN(n5859) );
  AND2_X1 U5766 ( .A1(n4689), .A2(n5859), .ZN(n5905) );
  NOR2_X1 U5767 ( .A1(n5852), .A2(n5847), .ZN(n5846) );
  NAND2_X1 U5768 ( .A1(n6070), .A2(n3140), .ZN(n4903) );
  OR2_X1 U5769 ( .A1(n4903), .A2(n3679), .ZN(n4678) );
  NOR2_X1 U5770 ( .A1(n6072), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4677)
         );
  NAND2_X1 U5771 ( .A1(n6784), .A2(n4677), .ZN(n4731) );
  NAND2_X1 U5772 ( .A1(n4678), .A2(n4731), .ZN(n4680) );
  INV_X1 U5773 ( .A(n6784), .ZN(n4681) );
  INV_X1 U5774 ( .A(n6182), .ZN(n4679) );
  AOI21_X1 U5775 ( .B1(n4681), .B2(n5998), .A(n4679), .ZN(n4691) );
  OAI211_X1 U5776 ( .C1(n4695), .C2(n4680), .A(n4691), .B(n6535), .ZN(n4730)
         );
  INV_X1 U5777 ( .A(n4680), .ZN(n4682) );
  AND2_X1 U5778 ( .A1(n6535), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6037) );
  INV_X1 U5779 ( .A(n6037), .ZN(n6126) );
  OAI22_X1 U5780 ( .A1(n4695), .A2(n4682), .B1(n4681), .B2(n6126), .ZN(n4729)
         );
  OR2_X1 U5781 ( .A1(n5840), .A2(n6444), .ZN(n6100) );
  INV_X1 U5782 ( .A(n6100), .ZN(n6620) );
  AOI22_X1 U5783 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4730), .B1(n4729), 
        .B2(n6620), .ZN(n4688) );
  NOR2_X1 U5784 ( .A1(n5855), .A2(n5956), .ZN(n4684) );
  NAND2_X1 U5785 ( .A1(n6472), .A2(DATAI_28_), .ZN(n6623) );
  INV_X1 U5786 ( .A(n6623), .ZN(n6556) );
  OR2_X1 U5787 ( .A1(n4725), .A2(n4685), .ZN(n6617) );
  NOR2_X1 U5788 ( .A1(n6617), .A2(n4731), .ZN(n4686) );
  AOI21_X1 U5789 ( .B1(n4932), .B2(n6556), .A(n4686), .ZN(n4687) );
  OAI211_X1 U5790 ( .C1(n6618), .C2(n5947), .A(n4688), .B(n4687), .ZN(U3048)
         );
  NAND2_X1 U5791 ( .A1(n6472), .A2(DATAI_21_), .ZN(n6589) );
  NAND2_X1 U5792 ( .A1(n6039), .A2(n5952), .ZN(n4690) );
  AND2_X1 U5793 ( .A1(n6784), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6036)
         );
  NAND2_X1 U5794 ( .A1(n6036), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U5795 ( .A1(n4690), .A2(n6631), .ZN(n4692) );
  OAI211_X1 U5796 ( .C1(n4695), .C2(n4692), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n4691), .ZN(n6638) );
  INV_X1 U5797 ( .A(n4692), .ZN(n4694) );
  INV_X1 U5798 ( .A(n6036), .ZN(n4693) );
  OAI22_X1 U5799 ( .A1(n4695), .A2(n4694), .B1(n6782), .B2(n4693), .ZN(n6637)
         );
  INV_X1 U5800 ( .A(DATAI_5_), .ZN(n6446) );
  OR2_X1 U5801 ( .A1(n5840), .A2(n6446), .ZN(n6104) );
  AOI22_X1 U5802 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6638), .B1(n6637), 
        .B2(n6591), .ZN(n4701) );
  AND2_X1 U5803 ( .A1(n5855), .A2(n6120), .ZN(n4697) );
  NAND2_X1 U5804 ( .A1(n6472), .A2(DATAI_29_), .ZN(n6594) );
  OR2_X1 U5805 ( .A1(n4725), .A2(n4698), .ZN(n6588) );
  OAI22_X1 U5806 ( .A1(n6641), .A2(n6594), .B1(n6588), .B2(n6631), .ZN(n4699)
         );
  INV_X1 U5807 ( .A(n4699), .ZN(n4700) );
  OAI211_X1 U5808 ( .C1(n6589), .C2(n6634), .A(n4701), .B(n4700), .ZN(U3113)
         );
  INV_X1 U5809 ( .A(n6084), .ZN(n6532) );
  AOI22_X1 U5810 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n4730), .B1(n4729), 
        .B2(n6532), .ZN(n4704) );
  NOR2_X1 U5811 ( .A1(n6083), .A2(n4731), .ZN(n4702) );
  AOI21_X1 U5812 ( .B1(n4932), .B2(n6539), .A(n4702), .ZN(n4703) );
  OAI211_X1 U5813 ( .C1(n6542), .C2(n5947), .A(n4704), .B(n4703), .ZN(U3044)
         );
  AOI22_X1 U5814 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n4730), .B1(n4729), 
        .B2(n6591), .ZN(n4707) );
  INV_X1 U5815 ( .A(n6594), .ZN(n6560) );
  NOR2_X1 U5816 ( .A1(n6588), .A2(n4731), .ZN(n4705) );
  AOI21_X1 U5817 ( .B1(n4932), .B2(n6560), .A(n4705), .ZN(n4706) );
  OAI211_X1 U5818 ( .C1(n6589), .C2(n5947), .A(n4707), .B(n4706), .ZN(U3049)
         );
  NAND2_X1 U5819 ( .A1(n6472), .A2(DATAI_17_), .ZN(n6576) );
  OR2_X1 U5820 ( .A1(n5840), .A2(n6438), .ZN(n6088) );
  AOI22_X1 U5821 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4730), .B1(n4729), 
        .B2(n6578), .ZN(n4710) );
  NAND2_X1 U5822 ( .A1(n6472), .A2(DATAI_25_), .ZN(n6581) );
  INV_X1 U5823 ( .A(n6581), .ZN(n6544) );
  OR2_X1 U5824 ( .A1(n4725), .A2(n3292), .ZN(n6575) );
  NOR2_X1 U5825 ( .A1(n6575), .A2(n4731), .ZN(n4708) );
  AOI21_X1 U5826 ( .B1(n4932), .B2(n6544), .A(n4708), .ZN(n4709) );
  OAI211_X1 U5827 ( .C1(n6576), .C2(n5947), .A(n4710), .B(n4709), .ZN(U3045)
         );
  AOI22_X1 U5828 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6638), .B1(n6637), 
        .B2(n6578), .ZN(n4713) );
  OAI22_X1 U5829 ( .A1(n6641), .A2(n6581), .B1(n6575), .B2(n6631), .ZN(n4711)
         );
  INV_X1 U5830 ( .A(n4711), .ZN(n4712) );
  OAI211_X1 U5831 ( .C1(n6576), .C2(n6634), .A(n4713), .B(n4712), .ZN(U3109)
         );
  AOI22_X1 U5832 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6638), .B1(n6637), 
        .B2(n6532), .ZN(n4716) );
  OAI22_X1 U5833 ( .A1(n6641), .A2(n6133), .B1(n6083), .B2(n6631), .ZN(n4714)
         );
  INV_X1 U5834 ( .A(n4714), .ZN(n4715) );
  OAI211_X1 U5835 ( .C1(n6542), .C2(n6634), .A(n4716), .B(n4715), .ZN(U3108)
         );
  NAND2_X1 U5836 ( .A1(n6472), .A2(DATAI_22_), .ZN(n6625) );
  INV_X1 U5837 ( .A(DATAI_6_), .ZN(n7064) );
  OR2_X1 U5838 ( .A1(n5840), .A2(n7064), .ZN(n6108) );
  AOI22_X1 U5839 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n4730), .B1(n4729), 
        .B2(n6627), .ZN(n4720) );
  NAND2_X1 U5840 ( .A1(n6472), .A2(DATAI_30_), .ZN(n6630) );
  INV_X1 U5841 ( .A(n6630), .ZN(n6564) );
  OR2_X1 U5842 ( .A1(n4725), .A2(n4717), .ZN(n6624) );
  NOR2_X1 U5843 ( .A1(n6624), .A2(n4731), .ZN(n4718) );
  AOI21_X1 U5844 ( .B1(n4932), .B2(n6564), .A(n4718), .ZN(n4719) );
  OAI211_X1 U5845 ( .C1(n6625), .C2(n5947), .A(n4720), .B(n4719), .ZN(U3050)
         );
  INV_X1 U5846 ( .A(n6096), .ZN(n6613) );
  AOI22_X1 U5847 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n4730), .B1(n4729), 
        .B2(n6613), .ZN(n4723) );
  NOR2_X1 U5848 ( .A1(n6610), .A2(n4731), .ZN(n4721) );
  AOI21_X1 U5849 ( .B1(n4932), .B2(n6552), .A(n4721), .ZN(n4722) );
  OAI211_X1 U5850 ( .C1(n6611), .C2(n5947), .A(n4723), .B(n4722), .ZN(U3047)
         );
  NAND2_X1 U5851 ( .A1(n6472), .A2(DATAI_18_), .ZN(n6604) );
  OR2_X1 U5852 ( .A1(n5840), .A2(n6440), .ZN(n6092) );
  AOI22_X1 U5853 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n4730), .B1(n4729), 
        .B2(n6606), .ZN(n4728) );
  NAND2_X1 U5854 ( .A1(n6472), .A2(DATAI_26_), .ZN(n6609) );
  INV_X1 U5855 ( .A(n6609), .ZN(n6548) );
  OR2_X1 U5856 ( .A1(n4725), .A2(n4724), .ZN(n6603) );
  NOR2_X1 U5857 ( .A1(n6603), .A2(n4731), .ZN(n4726) );
  AOI21_X1 U5858 ( .B1(n4932), .B2(n6548), .A(n4726), .ZN(n4727) );
  OAI211_X1 U5859 ( .C1(n6604), .C2(n5947), .A(n4728), .B(n4727), .ZN(U3046)
         );
  INV_X1 U5860 ( .A(n6114), .ZN(n6636) );
  AOI22_X1 U5861 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n4730), .B1(n4729), 
        .B2(n6636), .ZN(n4734) );
  NOR2_X1 U5862 ( .A1(n6632), .A2(n4731), .ZN(n4732) );
  AOI21_X1 U5863 ( .B1(n4932), .B2(n6571), .A(n4732), .ZN(n4733) );
  OAI211_X1 U5864 ( .C1(n6633), .C2(n5947), .A(n4734), .B(n4733), .ZN(U3051)
         );
  INV_X1 U5865 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6978) );
  OAI222_X1 U5866 ( .A1(n6352), .A2(n5438), .B1(n5437), .B2(n6446), .C1(n5436), 
        .C2(n6978), .ZN(U2886) );
  CLKBUF_X1 U5867 ( .A(n4735), .Z(n4736) );
  XNOR2_X1 U5868 ( .A(n4737), .B(n4736), .ZN(n4754) );
  AOI21_X1 U5869 ( .B1(n6497), .B2(n6495), .A(n6496), .ZN(n5832) );
  NOR2_X1 U5870 ( .A1(n4739), .A2(n5832), .ZN(n4950) );
  OAI211_X1 U5871 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4950), .B(n4891), .ZN(n4742) );
  INV_X1 U5872 ( .A(n6497), .ZN(n4738) );
  AOI21_X1 U5873 ( .B1(n4969), .B2(n4738), .A(n4966), .ZN(n6509) );
  NAND2_X1 U5874 ( .A1(n6496), .A2(n4739), .ZN(n6507) );
  NAND2_X1 U5875 ( .A1(n6509), .A2(n6507), .ZN(n4951) );
  OAI22_X1 U5876 ( .A1(n6500), .A2(n6364), .B1(n6665), .B2(n6498), .ZN(n4740)
         );
  AOI21_X1 U5877 ( .B1(n4951), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4740), 
        .ZN(n4741) );
  OAI211_X1 U5878 ( .C1(n6515), .C2(n4754), .A(n4742), .B(n4741), .ZN(U3014)
         );
  INV_X1 U5879 ( .A(n5325), .ZN(n4743) );
  NAND2_X1 U5880 ( .A1(n4743), .A2(n6472), .ZN(n4748) );
  INV_X1 U5881 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4746) );
  AND2_X1 U5882 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4744)
         );
  AOI211_X1 U5883 ( .C1(n5632), .C2(n4746), .A(n4745), .B(n4744), .ZN(n4747)
         );
  OAI211_X1 U5884 ( .C1(n4749), .C2(n5625), .A(n4748), .B(n4747), .ZN(U2985)
         );
  INV_X1 U5885 ( .A(n6371), .ZN(n4752) );
  AOI22_X1 U5886 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6465), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4750) );
  OAI21_X1 U5887 ( .B1(n6369), .B2(n6478), .A(n4750), .ZN(n4751) );
  AOI21_X1 U5888 ( .B1(n4752), .B2(n6472), .A(n4751), .ZN(n4753) );
  OAI21_X1 U5889 ( .B1(n5625), .B2(n4754), .A(n4753), .ZN(U2982) );
  INV_X1 U5890 ( .A(n5861), .ZN(n4757) );
  NOR3_X1 U5891 ( .A1(n4757), .A2(n5906), .A3(n6120), .ZN(n6121) );
  AND3_X1 U5892 ( .A1(n4756), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6073) );
  NOR3_X1 U5893 ( .A1(n4757), .A2(n5906), .A3(n6245), .ZN(n5853) );
  AND2_X1 U5894 ( .A1(n5848), .A2(n4436), .ZN(n6082) );
  INV_X1 U5895 ( .A(n6082), .ZN(n6071) );
  NAND2_X1 U5896 ( .A1(n4551), .A2(n5952), .ZN(n6180) );
  NAND2_X1 U5897 ( .A1(n6073), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4783) );
  OAI21_X1 U5898 ( .B1(n6071), .B2(n6180), .A(n4783), .ZN(n4760) );
  OR3_X1 U5899 ( .A1(n5853), .A2(n5998), .A3(n4760), .ZN(n4758) );
  NAND2_X1 U5900 ( .A1(n4782), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4763)
         );
  NAND3_X1 U5901 ( .A1(n5861), .A2(n4759), .A3(n6120), .ZN(n6069) );
  AOI22_X1 U5902 ( .A1(n4760), .A2(n6186), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6073), .ZN(n4784) );
  OAI22_X1 U5903 ( .A1(n4784), .A2(n6104), .B1(n6588), .B2(n4783), .ZN(n4761)
         );
  AOI21_X1 U5904 ( .B1(n6560), .B2(n6117), .A(n4761), .ZN(n4762) );
  OAI211_X1 U5905 ( .C1(n6171), .C2(n6589), .A(n4763), .B(n4762), .ZN(U3129)
         );
  NAND2_X1 U5906 ( .A1(n4782), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4766)
         );
  OAI22_X1 U5907 ( .A1(n4784), .A2(n6108), .B1(n6624), .B2(n4783), .ZN(n4764)
         );
  AOI21_X1 U5908 ( .B1(n6564), .B2(n6117), .A(n4764), .ZN(n4765) );
  OAI211_X1 U5909 ( .C1(n6171), .C2(n6625), .A(n4766), .B(n4765), .ZN(U3130)
         );
  NAND2_X1 U5910 ( .A1(n4782), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4769)
         );
  OAI22_X1 U5911 ( .A1(n4784), .A2(n6100), .B1(n6617), .B2(n4783), .ZN(n4767)
         );
  AOI21_X1 U5912 ( .B1(n6556), .B2(n6117), .A(n4767), .ZN(n4768) );
  OAI211_X1 U5913 ( .C1(n6171), .C2(n6618), .A(n4769), .B(n4768), .ZN(U3128)
         );
  NAND2_X1 U5914 ( .A1(n4782), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4772)
         );
  OAI22_X1 U5915 ( .A1(n4784), .A2(n6092), .B1(n6603), .B2(n4783), .ZN(n4770)
         );
  AOI21_X1 U5916 ( .B1(n6548), .B2(n6117), .A(n4770), .ZN(n4771) );
  OAI211_X1 U5917 ( .C1(n6171), .C2(n6604), .A(n4772), .B(n4771), .ZN(U3126)
         );
  NAND2_X1 U5918 ( .A1(n4782), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4775)
         );
  OAI22_X1 U5919 ( .A1(n4784), .A2(n6088), .B1(n6575), .B2(n4783), .ZN(n4773)
         );
  AOI21_X1 U5920 ( .B1(n6544), .B2(n6117), .A(n4773), .ZN(n4774) );
  OAI211_X1 U5921 ( .C1(n6171), .C2(n6576), .A(n4775), .B(n4774), .ZN(U3125)
         );
  NAND2_X1 U5922 ( .A1(n4782), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4778)
         );
  OAI22_X1 U5923 ( .A1(n4784), .A2(n6096), .B1(n6610), .B2(n4783), .ZN(n4776)
         );
  AOI21_X1 U5924 ( .B1(n6552), .B2(n6117), .A(n4776), .ZN(n4777) );
  OAI211_X1 U5925 ( .C1(n6171), .C2(n6611), .A(n4778), .B(n4777), .ZN(U3127)
         );
  NAND2_X1 U5926 ( .A1(n4782), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4781)
         );
  OAI22_X1 U5927 ( .A1(n4784), .A2(n6114), .B1(n6632), .B2(n4783), .ZN(n4779)
         );
  AOI21_X1 U5928 ( .B1(n6571), .B2(n6117), .A(n4779), .ZN(n4780) );
  OAI211_X1 U5929 ( .C1(n6171), .C2(n6633), .A(n4781), .B(n4780), .ZN(U3131)
         );
  NAND2_X1 U5930 ( .A1(n4782), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4787)
         );
  OAI22_X1 U5931 ( .A1(n4784), .A2(n6084), .B1(n6083), .B2(n4783), .ZN(n4785)
         );
  AOI21_X1 U5932 ( .B1(n6539), .B2(n6117), .A(n4785), .ZN(n4786) );
  OAI211_X1 U5933 ( .C1(n6171), .C2(n6542), .A(n4787), .B(n4786), .ZN(U3124)
         );
  INV_X1 U5934 ( .A(n4788), .ZN(n4791) );
  INV_X1 U5935 ( .A(n4789), .ZN(n4836) );
  AOI21_X1 U5936 ( .B1(n4791), .B2(n4790), .A(n4836), .ZN(n6341) );
  AND2_X1 U5937 ( .A1(n4670), .A2(n4792), .ZN(n4794) );
  OR2_X1 U5938 ( .A1(n4794), .A2(n4793), .ZN(n6336) );
  OAI22_X1 U5939 ( .A1(n5382), .A2(n6336), .B1(n4795), .B2(n5381), .ZN(n4796)
         );
  AOI21_X1 U5940 ( .B1(n6341), .B2(n6379), .A(n4796), .ZN(n4797) );
  INV_X1 U5941 ( .A(n4797), .ZN(U2853) );
  NAND2_X1 U5942 ( .A1(n5859), .A2(n4842), .ZN(n4802) );
  INV_X1 U5943 ( .A(n4802), .ZN(n4798) );
  AOI21_X1 U5944 ( .B1(n4798), .B2(STATEBS16_REG_SCAN_IN), .A(n5998), .ZN(
        n4805) );
  NOR2_X1 U5945 ( .A1(n4551), .A2(n5992), .ZN(n5862) );
  NOR2_X1 U5946 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4843) );
  AND2_X1 U5947 ( .A1(n4843), .A2(n6535), .ZN(n5865) );
  NAND2_X1 U5948 ( .A1(n5865), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4827) );
  INV_X1 U5949 ( .A(n4827), .ZN(n4800) );
  AOI21_X1 U5950 ( .B1(n5862), .B2(n5952), .A(n4800), .ZN(n4804) );
  INV_X1 U5951 ( .A(n4804), .ZN(n4801) );
  AOI22_X1 U5952 ( .A1(n4805), .A2(n4801), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5865), .ZN(n4833) );
  NOR2_X1 U5953 ( .A1(n4802), .A2(n6120), .ZN(n4899) );
  OAI22_X1 U5954 ( .A1(n4935), .A2(n6611), .B1(n6610), .B2(n4827), .ZN(n4803)
         );
  AOI21_X1 U5955 ( .B1(n6552), .B2(n4829), .A(n4803), .ZN(n4808) );
  NAND2_X1 U5956 ( .A1(n4805), .A2(n4804), .ZN(n4806) );
  NAND2_X1 U5957 ( .A1(n4830), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4807) );
  OAI211_X1 U5958 ( .C1(n4833), .C2(n6096), .A(n4808), .B(n4807), .ZN(U3031)
         );
  OAI22_X1 U5959 ( .A1(n4935), .A2(n6604), .B1(n6603), .B2(n4827), .ZN(n4809)
         );
  AOI21_X1 U5960 ( .B1(n6548), .B2(n4829), .A(n4809), .ZN(n4811) );
  NAND2_X1 U5961 ( .A1(n4830), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4810) );
  OAI211_X1 U5962 ( .C1(n4833), .C2(n6092), .A(n4811), .B(n4810), .ZN(U3030)
         );
  OAI22_X1 U5963 ( .A1(n4935), .A2(n6542), .B1(n6083), .B2(n4827), .ZN(n4812)
         );
  AOI21_X1 U5964 ( .B1(n6539), .B2(n4829), .A(n4812), .ZN(n4814) );
  NAND2_X1 U5965 ( .A1(n4830), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4813) );
  OAI211_X1 U5966 ( .C1(n4833), .C2(n6084), .A(n4814), .B(n4813), .ZN(U3028)
         );
  OAI22_X1 U5967 ( .A1(n4935), .A2(n6633), .B1(n6632), .B2(n4827), .ZN(n4815)
         );
  AOI21_X1 U5968 ( .B1(n6571), .B2(n4829), .A(n4815), .ZN(n4817) );
  NAND2_X1 U5969 ( .A1(n4830), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4816) );
  OAI211_X1 U5970 ( .C1(n4833), .C2(n6114), .A(n4817), .B(n4816), .ZN(U3035)
         );
  OAI22_X1 U5971 ( .A1(n4935), .A2(n6589), .B1(n6588), .B2(n4827), .ZN(n4818)
         );
  AOI21_X1 U5972 ( .B1(n6560), .B2(n4829), .A(n4818), .ZN(n4820) );
  NAND2_X1 U5973 ( .A1(n4830), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4819) );
  OAI211_X1 U5974 ( .C1(n4833), .C2(n6104), .A(n4820), .B(n4819), .ZN(U3033)
         );
  OAI22_X1 U5975 ( .A1(n4935), .A2(n6576), .B1(n6575), .B2(n4827), .ZN(n4821)
         );
  AOI21_X1 U5976 ( .B1(n6544), .B2(n4829), .A(n4821), .ZN(n4823) );
  NAND2_X1 U5977 ( .A1(n4830), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4822) );
  OAI211_X1 U5978 ( .C1(n4833), .C2(n6088), .A(n4823), .B(n4822), .ZN(U3029)
         );
  OAI22_X1 U5979 ( .A1(n4935), .A2(n6625), .B1(n6624), .B2(n4827), .ZN(n4824)
         );
  AOI21_X1 U5980 ( .B1(n6564), .B2(n4829), .A(n4824), .ZN(n4826) );
  NAND2_X1 U5981 ( .A1(n4830), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4825) );
  OAI211_X1 U5982 ( .C1(n4833), .C2(n6108), .A(n4826), .B(n4825), .ZN(U3034)
         );
  OAI22_X1 U5983 ( .A1(n4935), .A2(n6618), .B1(n6617), .B2(n4827), .ZN(n4828)
         );
  AOI21_X1 U5984 ( .B1(n6556), .B2(n4829), .A(n4828), .ZN(n4832) );
  NAND2_X1 U5985 ( .A1(n4830), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4831) );
  OAI211_X1 U5986 ( .C1(n4833), .C2(n6100), .A(n4832), .B(n4831), .ZN(U3032)
         );
  OAI21_X1 U5987 ( .B1(n4836), .B2(n4835), .A(n5377), .ZN(n6325) );
  INV_X1 U5988 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6896) );
  OAI222_X1 U5989 ( .A1(n6325), .A2(n5438), .B1(n5437), .B2(n6448), .C1(n5436), 
        .C2(n6896), .ZN(U2884) );
  INV_X1 U5990 ( .A(n6341), .ZN(n4837) );
  INV_X1 U5991 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6407) );
  OAI222_X1 U5992 ( .A1(n4837), .A2(n5438), .B1(n5437), .B2(n7064), .C1(n5436), 
        .C2(n6407), .ZN(U2885) );
  NOR2_X1 U5993 ( .A1(n4793), .A2(n4839), .ZN(n4840) );
  OR2_X1 U5994 ( .A1(n4838), .A2(n4840), .ZN(n6319) );
  INV_X1 U5995 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4841) );
  OAI222_X1 U5996 ( .A1(n6319), .A2(n5382), .B1(n4841), .B2(n5381), .C1(n6325), 
        .C2(n5375), .ZN(U2852) );
  NAND2_X1 U5997 ( .A1(n4842), .A2(n5855), .ZN(n5995) );
  OR2_X1 U5998 ( .A1(n5998), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6177) );
  INV_X1 U5999 ( .A(n6177), .ZN(n4846) );
  NAND2_X1 U6000 ( .A1(n4843), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5999) );
  NOR2_X1 U6001 ( .A1(n5999), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4853)
         );
  NAND2_X1 U6002 ( .A1(n4850), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6080) );
  OAI21_X1 U6003 ( .B1(n4853), .B2(n6864), .A(n6080), .ZN(n4845) );
  INV_X1 U6004 ( .A(n6079), .ZN(n4844) );
  INV_X1 U6005 ( .A(n6033), .ZN(n6525) );
  AOI21_X1 U6006 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6525), .A(n5840), .ZN(
        n5864) );
  OAI21_X1 U6007 ( .B1(n4844), .B2(n6782), .A(n5864), .ZN(n6074) );
  AOI211_X1 U6008 ( .C1(n4846), .C2(n5992), .A(n4845), .B(n6074), .ZN(n4849)
         );
  INV_X1 U6009 ( .A(n5992), .ZN(n4852) );
  OAI21_X1 U6010 ( .B1(n4852), .B2(n5998), .A(n6529), .ZN(n4847) );
  NAND3_X1 U6011 ( .A1(n5994), .A2(n6596), .A3(n4847), .ZN(n4848) );
  NAND2_X1 U6012 ( .A1(n4849), .A2(n4848), .ZN(n4875) );
  NAND2_X1 U6013 ( .A1(n4875), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4856) );
  NOR2_X1 U6014 ( .A1(n6070), .A2(n5998), .ZN(n6129) );
  NOR2_X1 U6015 ( .A1(n4850), .A2(n6782), .ZN(n6075) );
  INV_X1 U6016 ( .A(n6075), .ZN(n6122) );
  NOR3_X1 U6017 ( .A1(n6122), .A2(n6525), .A3(n6079), .ZN(n4851) );
  AOI21_X1 U6018 ( .B1(n6129), .B2(n4852), .A(n4851), .ZN(n4877) );
  INV_X1 U6019 ( .A(n4853), .ZN(n4876) );
  OAI22_X1 U6020 ( .A1(n4877), .A2(n6092), .B1(n6603), .B2(n4876), .ZN(n4854)
         );
  AOI21_X1 U6021 ( .B1(n6548), .B2(n4879), .A(n4854), .ZN(n4855) );
  OAI211_X1 U6022 ( .C1(n5994), .C2(n6604), .A(n4856), .B(n4855), .ZN(U3086)
         );
  NAND2_X1 U6023 ( .A1(n4875), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4859) );
  OAI22_X1 U6024 ( .A1(n4877), .A2(n6100), .B1(n6617), .B2(n4876), .ZN(n4857)
         );
  AOI21_X1 U6025 ( .B1(n6556), .B2(n4879), .A(n4857), .ZN(n4858) );
  OAI211_X1 U6026 ( .C1(n5994), .C2(n6618), .A(n4859), .B(n4858), .ZN(U3088)
         );
  NAND2_X1 U6027 ( .A1(n4875), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4862) );
  OAI22_X1 U6028 ( .A1(n4877), .A2(n6084), .B1(n6083), .B2(n4876), .ZN(n4860)
         );
  AOI21_X1 U6029 ( .B1(n6539), .B2(n4879), .A(n4860), .ZN(n4861) );
  OAI211_X1 U6030 ( .C1(n5994), .C2(n6542), .A(n4862), .B(n4861), .ZN(U3084)
         );
  NAND2_X1 U6031 ( .A1(n4875), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4865) );
  OAI22_X1 U6032 ( .A1(n4877), .A2(n6088), .B1(n6575), .B2(n4876), .ZN(n4863)
         );
  AOI21_X1 U6033 ( .B1(n6544), .B2(n4879), .A(n4863), .ZN(n4864) );
  OAI211_X1 U6034 ( .C1(n5994), .C2(n6576), .A(n4865), .B(n4864), .ZN(U3085)
         );
  NAND2_X1 U6035 ( .A1(n4875), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4868) );
  OAI22_X1 U6036 ( .A1(n4877), .A2(n6104), .B1(n6588), .B2(n4876), .ZN(n4866)
         );
  AOI21_X1 U6037 ( .B1(n6560), .B2(n4879), .A(n4866), .ZN(n4867) );
  OAI211_X1 U6038 ( .C1(n5994), .C2(n6589), .A(n4868), .B(n4867), .ZN(U3089)
         );
  NAND2_X1 U6039 ( .A1(n4875), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4871) );
  OAI22_X1 U6040 ( .A1(n4877), .A2(n6096), .B1(n6610), .B2(n4876), .ZN(n4869)
         );
  AOI21_X1 U6041 ( .B1(n6552), .B2(n4879), .A(n4869), .ZN(n4870) );
  OAI211_X1 U6042 ( .C1(n5994), .C2(n6611), .A(n4871), .B(n4870), .ZN(U3087)
         );
  NAND2_X1 U6043 ( .A1(n4875), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4874) );
  OAI22_X1 U6044 ( .A1(n4877), .A2(n6114), .B1(n6632), .B2(n4876), .ZN(n4872)
         );
  AOI21_X1 U6045 ( .B1(n6571), .B2(n4879), .A(n4872), .ZN(n4873) );
  OAI211_X1 U6046 ( .C1(n5994), .C2(n6633), .A(n4874), .B(n4873), .ZN(U3091)
         );
  NAND2_X1 U6047 ( .A1(n4875), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4881) );
  OAI22_X1 U6048 ( .A1(n4877), .A2(n6108), .B1(n6624), .B2(n4876), .ZN(n4878)
         );
  AOI21_X1 U6049 ( .B1(n6564), .B2(n4879), .A(n4878), .ZN(n4880) );
  OAI211_X1 U6050 ( .C1(n5994), .C2(n6625), .A(n4881), .B(n4880), .ZN(U3090)
         );
  CLKBUF_X1 U6051 ( .A(n4882), .Z(n4884) );
  XNOR2_X1 U6052 ( .A(n4884), .B(n4883), .ZN(n4898) );
  INV_X1 U6053 ( .A(n6352), .ZN(n4887) );
  INV_X1 U6054 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6667) );
  NOR2_X1 U6055 ( .A1(n6498), .A2(n6667), .ZN(n4895) );
  AOI21_X1 U6056 ( .B1(n6466), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4895), 
        .ZN(n4885) );
  OAI21_X1 U6057 ( .B1(n6356), .B2(n6478), .A(n4885), .ZN(n4886) );
  AOI21_X1 U6058 ( .B1(n4887), .B2(n6472), .A(n4886), .ZN(n4888) );
  OAI21_X1 U6059 ( .B1(n5625), .B2(n4898), .A(n4888), .ZN(U2981) );
  NAND2_X1 U6060 ( .A1(n6497), .A2(n6495), .ZN(n4890) );
  INV_X1 U6061 ( .A(n4889), .ZN(n4892) );
  OAI22_X1 U6062 ( .A1(n4891), .A2(n4890), .B1(n5796), .B2(n4892), .ZN(n4894)
         );
  INV_X1 U6063 ( .A(n5765), .ZN(n5805) );
  NOR2_X1 U6064 ( .A1(n4893), .A2(n4892), .ZN(n5830) );
  OAI21_X1 U6065 ( .B1(n5805), .B2(n5830), .A(n6509), .ZN(n5835) );
  OAI21_X1 U6066 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4894), .A(n5835), 
        .ZN(n4897) );
  AOI21_X1 U6067 ( .B1(n6518), .B2(n6350), .A(n4895), .ZN(n4896) );
  OAI211_X1 U6068 ( .C1(n6515), .C2(n4898), .A(n4897), .B(n4896), .ZN(U3013)
         );
  OAI21_X1 U6069 ( .B1(n4899), .B2(n4932), .A(n6177), .ZN(n4900) );
  AOI21_X1 U6070 ( .B1(n4900), .B2(n4903), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4902) );
  NOR2_X1 U6071 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4901) );
  AND2_X1 U6072 ( .A1(n6784), .A2(n4901), .ZN(n4906) );
  AOI21_X1 U6073 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6033), .A(n5840), .ZN(
        n6123) );
  NAND2_X1 U6074 ( .A1(n4928), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4909) );
  INV_X1 U6075 ( .A(n6576), .ZN(n6140) );
  OR2_X1 U6076 ( .A1(n4903), .A2(n5998), .ZN(n4905) );
  NAND3_X1 U6077 ( .A1(n6075), .A2(n6525), .A3(n6535), .ZN(n4904) );
  INV_X1 U6078 ( .A(n4906), .ZN(n4929) );
  OAI22_X1 U6079 ( .A1(n4930), .A2(n6088), .B1(n6575), .B2(n4929), .ZN(n4907)
         );
  AOI21_X1 U6080 ( .B1(n4932), .B2(n6140), .A(n4907), .ZN(n4908) );
  OAI211_X1 U6081 ( .C1(n4935), .C2(n6581), .A(n4909), .B(n4908), .ZN(U3037)
         );
  NAND2_X1 U6082 ( .A1(n4928), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4912) );
  INV_X1 U6083 ( .A(n6604), .ZN(n6145) );
  OAI22_X1 U6084 ( .A1(n4930), .A2(n6092), .B1(n6603), .B2(n4929), .ZN(n4910)
         );
  AOI21_X1 U6085 ( .B1(n4932), .B2(n6145), .A(n4910), .ZN(n4911) );
  OAI211_X1 U6086 ( .C1(n4935), .C2(n6609), .A(n4912), .B(n4911), .ZN(U3038)
         );
  NAND2_X1 U6087 ( .A1(n4928), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4915) );
  INV_X1 U6088 ( .A(n6611), .ZN(n6150) );
  OAI22_X1 U6089 ( .A1(n4930), .A2(n6096), .B1(n6610), .B2(n4929), .ZN(n4913)
         );
  AOI21_X1 U6090 ( .B1(n4932), .B2(n6150), .A(n4913), .ZN(n4914) );
  OAI211_X1 U6091 ( .C1(n4935), .C2(n6616), .A(n4915), .B(n4914), .ZN(U3039)
         );
  NAND2_X1 U6092 ( .A1(n4928), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4918) );
  INV_X1 U6093 ( .A(n6542), .ZN(n6135) );
  OAI22_X1 U6094 ( .A1(n4930), .A2(n6084), .B1(n6083), .B2(n4929), .ZN(n4916)
         );
  AOI21_X1 U6095 ( .B1(n4932), .B2(n6135), .A(n4916), .ZN(n4917) );
  OAI211_X1 U6096 ( .C1(n4935), .C2(n6133), .A(n4918), .B(n4917), .ZN(U3036)
         );
  NAND2_X1 U6097 ( .A1(n4928), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4921) );
  INV_X1 U6098 ( .A(n6589), .ZN(n6160) );
  OAI22_X1 U6099 ( .A1(n4930), .A2(n6104), .B1(n6588), .B2(n4929), .ZN(n4919)
         );
  AOI21_X1 U6100 ( .B1(n4932), .B2(n6160), .A(n4919), .ZN(n4920) );
  OAI211_X1 U6101 ( .C1(n4935), .C2(n6594), .A(n4921), .B(n4920), .ZN(U3041)
         );
  NAND2_X1 U6102 ( .A1(n4928), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4924) );
  INV_X1 U6103 ( .A(n6625), .ZN(n6165) );
  OAI22_X1 U6104 ( .A1(n4930), .A2(n6108), .B1(n6624), .B2(n4929), .ZN(n4922)
         );
  AOI21_X1 U6105 ( .B1(n4932), .B2(n6165), .A(n4922), .ZN(n4923) );
  OAI211_X1 U6106 ( .C1(n4935), .C2(n6630), .A(n4924), .B(n4923), .ZN(U3042)
         );
  NAND2_X1 U6107 ( .A1(n4928), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4927) );
  INV_X1 U6108 ( .A(n6633), .ZN(n6173) );
  OAI22_X1 U6109 ( .A1(n4930), .A2(n6114), .B1(n6632), .B2(n4929), .ZN(n4925)
         );
  AOI21_X1 U6110 ( .B1(n4932), .B2(n6173), .A(n4925), .ZN(n4926) );
  OAI211_X1 U6111 ( .C1(n4935), .C2(n6642), .A(n4927), .B(n4926), .ZN(U3043)
         );
  NAND2_X1 U6112 ( .A1(n4928), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4934) );
  INV_X1 U6113 ( .A(n6618), .ZN(n6155) );
  OAI22_X1 U6114 ( .A1(n4930), .A2(n6100), .B1(n6617), .B2(n4929), .ZN(n4931)
         );
  AOI21_X1 U6115 ( .B1(n4932), .B2(n6155), .A(n4931), .ZN(n4933) );
  OAI211_X1 U6116 ( .C1(n4935), .C2(n6623), .A(n4934), .B(n4933), .ZN(U3040)
         );
  INV_X1 U6117 ( .A(n4939), .ZN(n4936) );
  AOI21_X1 U6118 ( .B1(n4937), .B2(n4936), .A(n6715), .ZN(n4947) );
  INV_X1 U6119 ( .A(n4938), .ZN(n4944) );
  NAND2_X1 U6120 ( .A1(n4939), .A2(n4946), .ZN(n4942) );
  OAI22_X1 U6121 ( .A1(n6712), .A2(n4942), .B1(n4941), .B2(n4940), .ZN(n4943)
         );
  AOI21_X1 U6122 ( .B1(n4944), .B2(n6234), .A(n4943), .ZN(n4945) );
  OAI22_X1 U6123 ( .A1(n4947), .A2(n4946), .B1(n6715), .B2(n4945), .ZN(U3459)
         );
  XNOR2_X1 U6124 ( .A(n4948), .B(n4949), .ZN(n4959) );
  AOI22_X1 U6125 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4951), .B1(n4950), 
        .B2(n6837), .ZN(n4953) );
  INV_X1 U6126 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6884) );
  NOR2_X1 U6127 ( .A1(n6498), .A2(n6884), .ZN(n4954) );
  AOI21_X1 U6128 ( .B1(n6518), .B2(n5302), .A(n4954), .ZN(n4952) );
  OAI211_X1 U6129 ( .C1(n4959), .C2(n6515), .A(n4953), .B(n4952), .ZN(U3015)
         );
  INV_X1 U6130 ( .A(n5308), .ZN(n4957) );
  AOI21_X1 U6131 ( .B1(n6466), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4954), 
        .ZN(n4955) );
  OAI21_X1 U6132 ( .B1(n5300), .B2(n6478), .A(n4955), .ZN(n4956) );
  AOI21_X1 U6133 ( .B1(n4957), .B2(n6472), .A(n4956), .ZN(n4958) );
  OAI21_X1 U6134 ( .B1(n4959), .B2(n5625), .A(n4958), .ZN(U2983) );
  INV_X1 U6135 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5031) );
  OAI222_X1 U6136 ( .A1(n5375), .A2(n5019), .B1(n5382), .B2(n4960), .C1(n5031), 
        .C2(n5381), .ZN(U2829) );
  CLKBUF_X1 U6137 ( .A(n4961), .Z(n4965) );
  INV_X1 U6139 ( .A(n5529), .ZN(n4963) );
  AOI21_X1 U6140 ( .B1(n4965), .B2(n4964), .A(n4963), .ZN(n4996) );
  AND2_X1 U6141 ( .A1(n5806), .A2(n6496), .ZN(n4967) );
  AOI211_X1 U6142 ( .C1(n4969), .C2(n4968), .A(n4967), .B(n4966), .ZN(n5816)
         );
  INV_X1 U6143 ( .A(n5816), .ZN(n5824) );
  AOI21_X1 U6144 ( .B1(n4970), .B2(n5765), .A(n5824), .ZN(n6487) );
  NAND2_X1 U6145 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4974) );
  AOI22_X1 U6146 ( .A1(n4974), .A2(n4973), .B1(n4972), .B2(n4971), .ZN(n4975)
         );
  NAND2_X1 U6147 ( .A1(n6487), .A2(n4975), .ZN(n5791) );
  INV_X1 U6148 ( .A(n4976), .ZN(n4977) );
  NAND3_X1 U6149 ( .A1(n4977), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n4984), 
        .ZN(n4979) );
  NAND3_X1 U6150 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n6948), .ZN(n4985) );
  AOI21_X1 U6151 ( .B1(n4979), .B2(n4978), .A(n4985), .ZN(n5790) );
  NAND2_X1 U6152 ( .A1(n4980), .A2(n5359), .ZN(n5358) );
  INV_X1 U6153 ( .A(n5358), .ZN(n4983) );
  OAI21_X1 U6154 ( .B1(n4983), .B2(n4982), .A(n4981), .ZN(n6277) );
  NAND2_X1 U6155 ( .A1(n6465), .A2(REIP_REG_13__SCAN_IN), .ZN(n4993) );
  INV_X1 U6156 ( .A(n4984), .ZN(n4986) );
  OR3_X1 U6157 ( .A1(n6521), .A2(n4986), .A3(n4985), .ZN(n4987) );
  OAI211_X1 U6158 ( .C1(n6277), .C2(n6500), .A(n4993), .B(n4987), .ZN(n4988)
         );
  AOI211_X1 U6159 ( .C1(n5791), .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5790), .B(n4988), .ZN(n4989) );
  OAI21_X1 U6160 ( .B1(n4996), .B2(n6515), .A(n4989), .ZN(U3005) );
  XNOR2_X1 U6161 ( .A(n5362), .B(n3824), .ZN(n6380) );
  NAND2_X1 U6162 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4992)
         );
  OAI211_X1 U6163 ( .C1(n6478), .C2(n6278), .A(n4993), .B(n4992), .ZN(n4994)
         );
  AOI21_X1 U6164 ( .B1(n6380), .B2(n6472), .A(n4994), .ZN(n4995) );
  OAI21_X1 U6165 ( .B1(n4996), .B2(n5625), .A(n4995), .ZN(U2973) );
  AND2_X1 U6166 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6779) );
  XNOR2_X1 U6167 ( .A(n5532), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5461)
         );
  INV_X1 U6168 ( .A(n4997), .ZN(n4999) );
  NOR2_X1 U6169 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U6170 ( .A1(n4999), .A2(n4998), .ZN(n5000) );
  INV_X1 U6171 ( .A(n6779), .ZN(n5004) );
  NOR3_X1 U6172 ( .A1(n5005), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5004), 
        .ZN(n5006) );
  NOR2_X1 U6173 ( .A1(n6498), .A2(n6707), .ZN(n5037) );
  OAI21_X1 U6174 ( .B1(n5805), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5008), 
        .ZN(n5009) );
  NAND2_X1 U6175 ( .A1(n5009), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5010) );
  OAI211_X1 U6176 ( .C1(n3145), .C2(n6515), .A(n5011), .B(n5010), .ZN(U2987)
         );
  AOI21_X1 U6177 ( .B1(n5012), .B2(n4308), .A(n4393), .ZN(n5046) );
  NAND2_X1 U6178 ( .A1(n5046), .A2(n6472), .ZN(n5017) );
  OAI21_X1 U6179 ( .B1(n5630), .B2(n5014), .A(n5013), .ZN(n5015) );
  AOI21_X1 U6180 ( .B1(n5632), .B2(n5047), .A(n5015), .ZN(n5016) );
  OAI211_X1 U6181 ( .C1(n5018), .C2(n5625), .A(n5017), .B(n5016), .ZN(U2957)
         );
  INV_X1 U6182 ( .A(n5019), .ZN(n5020) );
  NAND2_X1 U6183 ( .A1(n5020), .A2(n3093), .ZN(n5036) );
  INV_X1 U6184 ( .A(n5021), .ZN(n5026) );
  NOR2_X1 U6185 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5022), .ZN(n5024) );
  NAND3_X1 U6186 ( .A1(n5299), .A2(n5024), .A3(n5023), .ZN(n5025) );
  INV_X1 U6187 ( .A(n5028), .ZN(n5029) );
  AOI22_X1 U6188 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5029), .ZN(n5030) );
  OAI21_X1 U6189 ( .B1(n6310), .B2(n5031), .A(n5030), .ZN(n5033) );
  NOR3_X1 U6190 ( .A1(n5051), .A2(REIP_REG_30__SCAN_IN), .A3(n6703), .ZN(n5032) );
  AOI211_X1 U6191 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5034), .A(n5033), .B(n5032), .ZN(n5035) );
  OAI211_X1 U6192 ( .C1(n4960), .C2(n6335), .A(n5036), .B(n5035), .ZN(U2797)
         );
  AOI21_X1 U6193 ( .B1(n6466), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5037), 
        .ZN(n5038) );
  OAI21_X1 U6194 ( .B1(n6478), .B2(n5039), .A(n5038), .ZN(n5040) );
  OAI21_X1 U6195 ( .B1(n3145), .B2(n5625), .A(n5041), .ZN(U2955) );
  NAND3_X1 U6196 ( .A1(n5042), .A2(n5386), .A3(n5436), .ZN(n5045) );
  NOR2_X2 U6197 ( .A1(n6387), .A2(n5043), .ZN(n6384) );
  AOI22_X1 U6198 ( .A1(n6384), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6387), .ZN(n5044) );
  NAND2_X1 U6199 ( .A1(n5045), .A2(n5044), .ZN(U2860) );
  INV_X1 U6200 ( .A(n5046), .ZN(n5392) );
  INV_X1 U6201 ( .A(n5336), .ZN(n5050) );
  INV_X1 U6202 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5337) );
  AOI22_X1 U6203 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5047), .ZN(n5048) );
  OAI21_X1 U6204 ( .B1(n6310), .B2(n5337), .A(n5048), .ZN(n5049) );
  AOI21_X1 U6205 ( .B1(n5050), .B2(n6366), .A(n5049), .ZN(n5053) );
  MUX2_X1 U6206 ( .A(n5051), .B(n5062), .S(REIP_REG_29__SCAN_IN), .Z(n5052) );
  OAI211_X1 U6207 ( .C1(n5392), .C2(n3130), .A(n5053), .B(n5052), .ZN(U2798)
         );
  OAI22_X1 U6208 ( .A1(n5055), .A2(n6348), .B1(n5027), .B2(n5054), .ZN(n5060)
         );
  AND2_X1 U6209 ( .A1(n5071), .A2(n5056), .ZN(n5057) );
  OR2_X1 U6210 ( .A1(n5058), .A2(n5057), .ZN(n5658) );
  NOR2_X1 U6211 ( .A1(n5658), .A2(n6335), .ZN(n5059) );
  AOI211_X1 U6212 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6358), .A(n5060), .B(n5059), 
        .ZN(n5065) );
  INV_X1 U6213 ( .A(n5074), .ZN(n5061) );
  NAND2_X1 U6214 ( .A1(n5061), .A2(REIP_REG_27__SCAN_IN), .ZN(n5063) );
  MUX2_X1 U6215 ( .A(n5063), .B(n5062), .S(REIP_REG_28__SCAN_IN), .Z(n5064) );
  OAI211_X1 U6216 ( .C1(n5395), .C2(n3130), .A(n5065), .B(n5064), .ZN(U2799)
         );
  AOI21_X1 U6217 ( .B1(n5067), .B2(n5066), .A(n3090), .ZN(n5447) );
  INV_X1 U6218 ( .A(n5447), .ZN(n5398) );
  NAND2_X1 U6219 ( .A1(n5084), .A2(n5069), .ZN(n5070) );
  NAND2_X1 U6220 ( .A1(n5071), .A2(n5070), .ZN(n5664) );
  AOI22_X1 U6221 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5443), .ZN(n5073) );
  NAND2_X1 U6222 ( .A1(n6358), .A2(EBX_REG_27__SCAN_IN), .ZN(n5072) );
  OAI211_X1 U6223 ( .C1(n5664), .C2(n6335), .A(n5073), .B(n5072), .ZN(n5076)
         );
  NOR2_X1 U6224 ( .A1(n5074), .A2(REIP_REG_27__SCAN_IN), .ZN(n5075) );
  OAI21_X1 U6225 ( .B1(n5398), .B2(n3130), .A(n5077), .ZN(U2800) );
  AND2_X1 U6226 ( .A1(n5093), .A2(n5078), .ZN(n5095) );
  OAI21_X1 U6227 ( .B1(n5095), .B2(n5079), .A(n5066), .ZN(n5456) );
  OAI22_X1 U6228 ( .A1(n5080), .A2(n6348), .B1(n5027), .B2(n5450), .ZN(n5086)
         );
  OR2_X1 U6229 ( .A1(n5081), .A2(n5082), .ZN(n5083) );
  NAND2_X1 U6230 ( .A1(n5084), .A2(n5083), .ZN(n5673) );
  NOR2_X1 U6231 ( .A1(n5673), .A2(n6335), .ZN(n5085) );
  AOI211_X1 U6232 ( .C1(EBX_REG_26__SCAN_IN), .C2(n6358), .A(n5086), .B(n5085), 
        .ZN(n5092) );
  INV_X1 U6233 ( .A(n5087), .ZN(n5119) );
  NOR2_X1 U6234 ( .A1(n5119), .A2(n5088), .ZN(n5090) );
  OAI21_X1 U6235 ( .B1(n5090), .B2(REIP_REG_26__SCAN_IN), .A(n5089), .ZN(n5091) );
  OAI211_X1 U6236 ( .C1(n5456), .C2(n3130), .A(n5092), .B(n5091), .ZN(U2801)
         );
  INV_X1 U6237 ( .A(n5093), .ZN(n5213) );
  AOI21_X1 U6238 ( .B1(n5096), .B2(n5114), .A(n5095), .ZN(n5097) );
  INV_X1 U6239 ( .A(n5097), .ZN(n5465) );
  AOI21_X1 U6240 ( .B1(n5142), .B2(n5098), .A(n5326), .ZN(n5134) );
  INV_X1 U6241 ( .A(n5115), .ZN(n5102) );
  INV_X1 U6242 ( .A(n5100), .ZN(n5101) );
  AOI21_X1 U6243 ( .B1(n5129), .B2(n5102), .A(n5101), .ZN(n5103) );
  OR2_X1 U6244 ( .A1(n5081), .A2(n5103), .ZN(n5686) );
  AOI22_X1 U6245 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5459), .ZN(n5105) );
  NAND2_X1 U6246 ( .A1(n6358), .A2(EBX_REG_25__SCAN_IN), .ZN(n5104) );
  OAI211_X1 U6247 ( .C1(n5686), .C2(n6335), .A(n5105), .B(n5104), .ZN(n5108)
         );
  XNOR2_X1 U6248 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5106) );
  NOR2_X1 U6249 ( .A1(n5119), .A2(n5106), .ZN(n5107) );
  OAI21_X1 U6250 ( .B1(n5465), .B2(n3130), .A(n5109), .ZN(U2802) );
  NOR2_X2 U6251 ( .A1(n5213), .A2(n5110), .ZN(n5139) );
  NAND2_X1 U6252 ( .A1(n5139), .A2(n5111), .ZN(n5123) );
  NAND2_X1 U6253 ( .A1(n5123), .A2(n5112), .ZN(n5113) );
  XOR2_X1 U6254 ( .A(n5115), .B(n5129), .Z(n5694) );
  OAI22_X1 U6255 ( .A1(n5116), .A2(n6348), .B1(n5027), .B2(n5478), .ZN(n5117)
         );
  AOI21_X1 U6256 ( .B1(EBX_REG_24__SCAN_IN), .B2(n6358), .A(n5117), .ZN(n5118)
         );
  OAI21_X1 U6257 ( .B1(n5694), .B2(n6335), .A(n5118), .ZN(n5121) );
  NOR2_X1 U6258 ( .A1(n5119), .A2(REIP_REG_24__SCAN_IN), .ZN(n5120) );
  OAI21_X1 U6259 ( .B1(n5405), .B2(n3130), .A(n5122), .ZN(U2803) );
  OAI22_X1 U6260 ( .A1(n5125), .A2(n6348), .B1(n5027), .B2(n5489), .ZN(n5132)
         );
  INV_X1 U6261 ( .A(n5126), .ZN(n5127) );
  AOI21_X1 U6262 ( .B1(n5126), .B2(n5143), .A(n5128), .ZN(n5130) );
  OR2_X1 U6263 ( .A1(n5130), .A2(n5129), .ZN(n5701) );
  NOR2_X1 U6264 ( .A1(n5701), .A2(n6335), .ZN(n5131) );
  AOI211_X1 U6265 ( .C1(EBX_REG_23__SCAN_IN), .C2(n6358), .A(n5132), .B(n5131), 
        .ZN(n5137) );
  INV_X1 U6266 ( .A(n5133), .ZN(n5159) );
  NAND2_X1 U6267 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5147) );
  NOR2_X1 U6268 ( .A1(n5159), .A2(n5147), .ZN(n5135) );
  OAI21_X1 U6269 ( .B1(n5135), .B2(REIP_REG_23__SCAN_IN), .A(n5134), .ZN(n5136) );
  OAI211_X1 U6270 ( .C1(n5487), .C2(n3130), .A(n5137), .B(n5136), .ZN(U2804)
         );
  NOR2_X1 U6271 ( .A1(n5139), .A2(n5138), .ZN(n5140) );
  NOR2_X1 U6272 ( .A1(n5141), .A2(n5140), .ZN(n5500) );
  INV_X1 U6273 ( .A(n5500), .ZN(n5410) );
  NOR2_X1 U6274 ( .A1(n5142), .A2(n5326), .ZN(n5174) );
  INV_X1 U6275 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6910) );
  XNOR2_X1 U6276 ( .A(n5127), .B(n5143), .ZN(n5707) );
  NAND2_X1 U6277 ( .A1(n5707), .A2(n6366), .ZN(n5146) );
  INV_X1 U6278 ( .A(n5498), .ZN(n5144) );
  AOI22_X1 U6279 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5144), .ZN(n5145) );
  OAI211_X1 U6280 ( .C1(n6310), .C2(n6910), .A(n5146), .B(n5145), .ZN(n5150)
         );
  INV_X1 U6281 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7043) );
  INV_X1 U6282 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6691) );
  INV_X1 U6283 ( .A(n5147), .ZN(n5148) );
  AOI211_X1 U6284 ( .C1(n7043), .C2(n6691), .A(n5148), .B(n5159), .ZN(n5149)
         );
  AOI211_X1 U6285 ( .C1(n5174), .C2(REIP_REG_22__SCAN_IN), .A(n5150), .B(n5149), .ZN(n5151) );
  OAI21_X1 U6286 ( .B1(n5410), .B2(n3130), .A(n5151), .ZN(U2805) );
  XNOR2_X1 U6287 ( .A(n5166), .B(n5153), .ZN(n5510) );
  NAND2_X1 U6288 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  NAND2_X1 U6289 ( .A1(n5127), .A2(n5156), .ZN(n5717) );
  AOI22_X1 U6290 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5507), .ZN(n5158) );
  NAND2_X1 U6291 ( .A1(n6358), .A2(EBX_REG_21__SCAN_IN), .ZN(n5157) );
  OAI211_X1 U6292 ( .C1(n5717), .C2(n6335), .A(n5158), .B(n5157), .ZN(n5161)
         );
  NOR2_X1 U6293 ( .A1(n5159), .A2(REIP_REG_21__SCAN_IN), .ZN(n5160) );
  OAI21_X1 U6294 ( .B1(n5510), .B2(n3130), .A(n5162), .ZN(U2806) );
  OR2_X2 U6295 ( .A1(n5213), .A2(n5163), .ZN(n5182) );
  AND2_X1 U6296 ( .A1(n5182), .A2(n5164), .ZN(n5165) );
  NOR2_X1 U6297 ( .A1(n5166), .A2(n5165), .ZN(n5516) );
  INV_X1 U6298 ( .A(n5516), .ZN(n5415) );
  MUX2_X1 U6299 ( .A(n3131), .B(n5168), .S(n5167), .Z(n5171) );
  XNOR2_X1 U6300 ( .A(n5171), .B(n5170), .ZN(n5730) );
  INV_X1 U6301 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5173) );
  AOI22_X1 U6302 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5515), .ZN(n5172) );
  OAI21_X1 U6303 ( .B1(n6310), .B2(n5173), .A(n5172), .ZN(n5178) );
  AOI21_X1 U6304 ( .B1(n5183), .B2(REIP_REG_19__SCAN_IN), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5176) );
  INV_X1 U6305 ( .A(n5174), .ZN(n5175) );
  NOR2_X1 U6306 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  AOI211_X1 U6307 ( .C1(n6366), .C2(n5730), .A(n5178), .B(n5177), .ZN(n5179)
         );
  OAI21_X1 U6308 ( .B1(n5415), .B2(n3130), .A(n5179), .ZN(U2807) );
  NAND2_X1 U6309 ( .A1(n5197), .A2(n5180), .ZN(n5181) );
  NAND2_X2 U6310 ( .A1(n5182), .A2(n5181), .ZN(n5523) );
  INV_X1 U6311 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6688) );
  AOI22_X1 U6312 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6358), .B1(n5183), .B2(n6688), .ZN(n5196) );
  INV_X1 U6313 ( .A(n5218), .ZN(n5187) );
  OR2_X1 U6314 ( .A1(n5186), .A2(n5185), .ZN(n5200) );
  NAND2_X1 U6315 ( .A1(n5187), .A2(n5200), .ZN(n5203) );
  XNOR2_X1 U6316 ( .A(n5203), .B(n5188), .ZN(n5739) );
  NAND2_X1 U6317 ( .A1(n5293), .A2(n5189), .ZN(n6346) );
  OAI22_X1 U6318 ( .A1(n5326), .A2(n5223), .B1(REIP_REG_18__SCAN_IN), .B2(
        n5204), .ZN(n5190) );
  NAND2_X1 U6319 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5190), .ZN(n5191) );
  AND2_X1 U6320 ( .A1(n6346), .A2(n5191), .ZN(n5193) );
  AOI22_X1 U6321 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5526), .ZN(n5192) );
  OAI211_X1 U6322 ( .C1(n5739), .C2(n6335), .A(n5193), .B(n5192), .ZN(n5194)
         );
  INV_X1 U6323 ( .A(n5194), .ZN(n5195) );
  OAI211_X1 U6324 ( .C1(n5523), .C2(n3130), .A(n5196), .B(n5195), .ZN(U2808)
         );
  INV_X1 U6325 ( .A(n5197), .ZN(n5198) );
  AOI21_X1 U6326 ( .B1(n5199), .B2(n5213), .A(n5198), .ZN(n5542) );
  INV_X1 U6327 ( .A(n5542), .ZN(n5420) );
  INV_X1 U6328 ( .A(n5200), .ZN(n5201) );
  NAND2_X1 U6329 ( .A1(n5218), .A2(n5201), .ZN(n5202) );
  NAND2_X1 U6330 ( .A1(n5203), .A2(n5202), .ZN(n5748) );
  INV_X1 U6331 ( .A(n5748), .ZN(n5210) );
  INV_X1 U6332 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5347) );
  NOR2_X1 U6333 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5204), .ZN(n5205) );
  NOR2_X1 U6334 ( .A1(n6362), .A2(n5205), .ZN(n5207) );
  AOI22_X1 U6335 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5538), .ZN(n5206) );
  OAI211_X1 U6336 ( .C1(n6310), .C2(n5347), .A(n5207), .B(n5206), .ZN(n5209)
         );
  NOR3_X1 U6337 ( .A1(n5223), .A2(n5326), .A3(n6685), .ZN(n5208) );
  AOI211_X1 U6338 ( .C1(n6366), .C2(n5210), .A(n5209), .B(n5208), .ZN(n5211)
         );
  OAI21_X1 U6339 ( .B1(n5420), .B2(n3130), .A(n5211), .ZN(U2809) );
  OAI21_X1 U6340 ( .B1(n5232), .B2(n5214), .A(n5213), .ZN(n5548) );
  NAND2_X1 U6341 ( .A1(n5215), .A2(n5216), .ZN(n5217) );
  NAND2_X1 U6342 ( .A1(n5218), .A2(n5217), .ZN(n5756) );
  NOR2_X1 U6343 ( .A1(n5756), .A2(n6335), .ZN(n5221) );
  NOR2_X1 U6344 ( .A1(n5027), .A2(n5550), .ZN(n5220) );
  OAI22_X1 U6345 ( .A1(n6310), .A2(n5348), .B1(n7038), .B2(n6348), .ZN(n5219)
         );
  NOR4_X1 U6346 ( .A1(n5221), .A2(n6362), .A3(n5220), .A4(n5219), .ZN(n5227)
         );
  INV_X1 U6347 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U6348 ( .A1(n5237), .A2(REIP_REG_15__SCAN_IN), .ZN(n5234) );
  INV_X1 U6349 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5222) );
  OAI21_X1 U6350 ( .B1(n6998), .B2(n5234), .A(n5222), .ZN(n5225) );
  INV_X1 U6351 ( .A(n5223), .ZN(n5224) );
  NAND3_X1 U6352 ( .A1(n5225), .A2(n5236), .A3(n5224), .ZN(n5226) );
  OAI211_X1 U6353 ( .C1(n5548), .C2(n3130), .A(n5227), .B(n5226), .ZN(U2810)
         );
  NOR2_X1 U6354 ( .A1(n5229), .A2(n5230), .ZN(n5231) );
  OR2_X1 U6355 ( .A1(n5232), .A2(n5231), .ZN(n6383) );
  AOI22_X1 U6356 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n6363), .B1(n5562), 
        .B2(n3129), .ZN(n5233) );
  OAI21_X1 U6357 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5234), .A(n5233), .ZN(n5245) );
  NAND2_X1 U6358 ( .A1(n5236), .A2(n5235), .ZN(n6262) );
  INV_X1 U6359 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7023) );
  NAND2_X1 U6360 ( .A1(n5237), .A2(n7023), .ZN(n5254) );
  AOI21_X1 U6361 ( .B1(n6262), .B2(n5254), .A(n6998), .ZN(n5244) );
  CLKBUF_X1 U6362 ( .A(n5238), .Z(n5239) );
  NAND2_X1 U6363 ( .A1(n5239), .A2(n5240), .ZN(n5241) );
  NAND2_X1 U6364 ( .A1(n5215), .A2(n5241), .ZN(n5772) );
  AOI21_X1 U6365 ( .B1(n6358), .B2(EBX_REG_16__SCAN_IN), .A(n6362), .ZN(n5242)
         );
  OAI21_X1 U6366 ( .B1(n5772), .B2(n6335), .A(n5242), .ZN(n5243) );
  NOR3_X1 U6367 ( .A1(n5245), .A2(n5244), .A3(n5243), .ZN(n5246) );
  OAI21_X1 U6368 ( .B1(n6383), .B2(n3130), .A(n5246), .ZN(U2811) );
  AOI21_X1 U6369 ( .B1(n5248), .B2(n5247), .A(n5229), .ZN(n5570) );
  INV_X1 U6370 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5352) );
  OAI22_X1 U6371 ( .A1(n6310), .A2(n5352), .B1(n7023), .B2(n6262), .ZN(n5256)
         );
  OR2_X1 U6372 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  NAND2_X1 U6373 ( .A1(n5239), .A2(n5251), .ZN(n5781) );
  OAI21_X1 U6374 ( .B1(n5027), .B2(n5568), .A(n6346), .ZN(n5252) );
  AOI21_X1 U6375 ( .B1(PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n6363), .A(n5252), 
        .ZN(n5253) );
  OAI211_X1 U6376 ( .C1(n6335), .C2(n5781), .A(n5254), .B(n5253), .ZN(n5255)
         );
  AOI211_X1 U6377 ( .C1(n5570), .C2(n3093), .A(n5256), .B(n5255), .ZN(n5257)
         );
  INV_X1 U6378 ( .A(n5257), .ZN(U2812) );
  INV_X1 U6379 ( .A(n5258), .ZN(n5378) );
  NAND2_X1 U6380 ( .A1(n5376), .A2(n5283), .ZN(n5371) );
  INV_X1 U6381 ( .A(n5259), .ZN(n5372) );
  NOR2_X1 U6382 ( .A1(n5371), .A2(n5372), .ZN(n5370) );
  INV_X1 U6383 ( .A(n5261), .ZN(n5262) );
  OAI21_X1 U6384 ( .B1(n5370), .B2(n5263), .A(n5262), .ZN(n5596) );
  INV_X1 U6385 ( .A(n5592), .ZN(n5276) );
  NOR2_X1 U6386 ( .A1(n5368), .A2(n5264), .ZN(n5265) );
  OR2_X1 U6387 ( .A1(n4980), .A2(n5265), .ZN(n6479) );
  OAI22_X1 U6388 ( .A1(n6479), .A2(n6335), .B1(n5266), .B2(n6348), .ZN(n5267)
         );
  INV_X1 U6389 ( .A(n5267), .ZN(n5268) );
  OAI211_X1 U6390 ( .C1(n6310), .C2(n5363), .A(n5268), .B(n6346), .ZN(n5275)
         );
  OAI21_X1 U6391 ( .B1(n5269), .B2(n6360), .A(n5293), .ZN(n6285) );
  INV_X1 U6392 ( .A(n6285), .ZN(n5273) );
  INV_X1 U6393 ( .A(n5269), .ZN(n6280) );
  NAND2_X1 U6394 ( .A1(n6329), .A2(n6280), .ZN(n5270) );
  OAI22_X1 U6395 ( .A1(n5273), .A2(n5272), .B1(n5271), .B2(n5270), .ZN(n5274)
         );
  AOI211_X1 U6396 ( .C1(n3129), .C2(n5276), .A(n5275), .B(n5274), .ZN(n5277)
         );
  OAI21_X1 U6397 ( .B1(n3130), .B2(n5596), .A(n5277), .ZN(U2816) );
  NAND2_X1 U6398 ( .A1(n6329), .A2(n5284), .ZN(n6308) );
  NAND2_X1 U6399 ( .A1(n6308), .A2(n5293), .ZN(n6306) );
  INV_X1 U6400 ( .A(n5367), .ZN(n5279) );
  AOI21_X1 U6401 ( .B1(n5280), .B2(n5278), .A(n5279), .ZN(n6489) );
  AOI22_X1 U6402 ( .A1(n6306), .A2(REIP_REG_9__SCAN_IN), .B1(n6366), .B2(n6489), .ZN(n5281) );
  OAI211_X1 U6403 ( .C1(n6348), .C2(n5282), .A(n5281), .B(n6346), .ZN(n5290)
         );
  OAI21_X1 U6404 ( .B1(n5376), .B2(n5283), .A(n5371), .ZN(n5618) );
  INV_X1 U6405 ( .A(n5614), .ZN(n5286) );
  NOR2_X1 U6406 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6360), .ZN(n6298) );
  INV_X1 U6407 ( .A(n5284), .ZN(n5285) );
  AOI22_X1 U6408 ( .A1(n3129), .A2(n5286), .B1(n6298), .B2(n5285), .ZN(n5288)
         );
  NAND2_X1 U6409 ( .A1(n6358), .A2(EBX_REG_9__SCAN_IN), .ZN(n5287) );
  OAI211_X1 U6410 ( .C1(n5618), .C2(n3130), .A(n5288), .B(n5287), .ZN(n5289)
         );
  OR2_X1 U6411 ( .A1(n5290), .A2(n5289), .ZN(U2818) );
  NAND2_X1 U6412 ( .A1(n5299), .A2(n5291), .ZN(n5292) );
  INV_X1 U6413 ( .A(n5293), .ZN(n6317) );
  INV_X1 U6414 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6662) );
  NOR2_X1 U6415 ( .A1(n6317), .A2(n6662), .ZN(n5295) );
  OAI21_X1 U6416 ( .B1(n6360), .B2(REIP_REG_1__SCAN_IN), .A(n5295), .ZN(n5294)
         );
  INV_X1 U6417 ( .A(n5294), .ZN(n5309) );
  NOR2_X1 U6418 ( .A1(n6884), .A2(n4544), .ZN(n5296) );
  AOI21_X1 U6419 ( .B1(n5296), .B2(n5295), .A(n5326), .ZN(n6357) );
  OAI21_X1 U6420 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5309), .A(n6357), .ZN(n5307)
         );
  INV_X1 U6421 ( .A(n5297), .ZN(n5298) );
  NAND2_X1 U6422 ( .A1(n5299), .A2(n5298), .ZN(n5329) );
  INV_X1 U6423 ( .A(n5300), .ZN(n5301) );
  AOI22_X1 U6424 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6363), .B1(n3129), 
        .B2(n5301), .ZN(n5304) );
  NAND2_X1 U6425 ( .A1(n6366), .A2(n5302), .ZN(n5303) );
  OAI211_X1 U6426 ( .C1(n6070), .C2(n5329), .A(n5304), .B(n5303), .ZN(n5305)
         );
  AOI21_X1 U6427 ( .B1(EBX_REG_3__SCAN_IN), .B2(n6358), .A(n5305), .ZN(n5306)
         );
  OAI211_X1 U6428 ( .C1(n6370), .C2(n5308), .A(n5307), .B(n5306), .ZN(U2824)
         );
  NAND2_X1 U6429 ( .A1(n6358), .A2(EBX_REG_2__SCAN_IN), .ZN(n5316) );
  AOI221_X1 U6430 ( .B1(n6360), .B2(n6662), .C1(n4544), .C2(n6662), .A(n5309), 
        .ZN(n5310) );
  AOI21_X1 U6431 ( .B1(n6363), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n5310), 
        .ZN(n5315) );
  INV_X1 U6432 ( .A(n5329), .ZN(n6368) );
  INV_X1 U6433 ( .A(n6499), .ZN(n5311) );
  AOI22_X1 U6434 ( .A1(n6368), .A2(n5848), .B1(n6366), .B2(n5311), .ZN(n5314)
         );
  INV_X1 U6435 ( .A(n6477), .ZN(n5312) );
  NAND2_X1 U6436 ( .A1(n3129), .A2(n5312), .ZN(n5313) );
  OAI21_X1 U6437 ( .B1(n5317), .B2(n6370), .A(n3136), .ZN(U2825) );
  NAND2_X1 U6438 ( .A1(n6329), .A2(n4544), .ZN(n5319) );
  AOI22_X1 U6439 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6317), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5318) );
  OAI211_X1 U6440 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n5027), .A(n5319), 
        .B(n5318), .ZN(n5323) );
  INV_X1 U6441 ( .A(n5320), .ZN(n5321) );
  OAI22_X1 U6442 ( .A1(n6335), .A2(n5321), .B1(n4436), .B2(n5329), .ZN(n5322)
         );
  AOI211_X1 U6443 ( .C1(EBX_REG_1__SCAN_IN), .C2(n6358), .A(n5323), .B(n5322), 
        .ZN(n5324) );
  OAI21_X1 U6444 ( .B1(n6370), .B2(n5325), .A(n5324), .ZN(U2826) );
  INV_X1 U6445 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6846) );
  OAI22_X1 U6446 ( .A1(n5326), .A2(n6846), .B1(n6310), .B2(n6981), .ZN(n5327)
         );
  INV_X1 U6447 ( .A(n5327), .ZN(n5332) );
  OAI21_X1 U6448 ( .B1(n6363), .B2(n3129), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5328) );
  OAI21_X1 U6449 ( .B1(n5329), .B2(n3679), .A(n5328), .ZN(n5330) );
  AOI21_X1 U6450 ( .B1(n6366), .B2(n6519), .A(n5330), .ZN(n5331) );
  OAI211_X1 U6451 ( .C1(n6370), .C2(n5644), .A(n5332), .B(n5331), .ZN(U2827)
         );
  INV_X1 U6452 ( .A(n5333), .ZN(n5335) );
  INV_X1 U6453 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5334) );
  OAI22_X1 U6454 ( .A1(n5335), .A2(n5382), .B1(n5381), .B2(n5334), .ZN(U2828)
         );
  OAI222_X1 U6455 ( .A1(n5375), .A2(n5392), .B1(n5381), .B2(n5337), .C1(n5336), 
        .C2(n5382), .ZN(U2830) );
  OAI222_X1 U6456 ( .A1(n5338), .A2(n5381), .B1(n5382), .B2(n5658), .C1(n5395), 
        .C2(n5375), .ZN(U2831) );
  INV_X1 U6457 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5339) );
  OAI222_X1 U6458 ( .A1(n5339), .A2(n5381), .B1(n5382), .B2(n5664), .C1(n5398), 
        .C2(n5375), .ZN(U2832) );
  OAI222_X1 U6459 ( .A1(n6827), .A2(n5381), .B1(n5382), .B2(n5673), .C1(n5456), 
        .C2(n5375), .ZN(U2833) );
  INV_X1 U6460 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5340) );
  OAI222_X1 U6461 ( .A1(n5340), .A2(n5381), .B1(n5382), .B2(n5686), .C1(n5465), 
        .C2(n5375), .ZN(U2834) );
  INV_X1 U6462 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5341) );
  OAI222_X1 U6463 ( .A1(n5341), .A2(n5381), .B1(n5382), .B2(n5694), .C1(n5375), 
        .C2(n5405), .ZN(U2835) );
  OAI222_X1 U6464 ( .A1(n5342), .A2(n5381), .B1(n5382), .B2(n5701), .C1(n5487), 
        .C2(n5375), .ZN(U2836) );
  INV_X1 U6465 ( .A(n5707), .ZN(n5343) );
  OAI222_X1 U6466 ( .A1(n6910), .A2(n5381), .B1(n5382), .B2(n5343), .C1(n5375), 
        .C2(n5410), .ZN(U2837) );
  INV_X1 U6467 ( .A(EBX_REG_21__SCAN_IN), .ZN(n7016) );
  OAI222_X1 U6468 ( .A1(n7016), .A2(n5381), .B1(n5382), .B2(n5717), .C1(n5510), 
        .C2(n5375), .ZN(U2838) );
  AOI22_X1 U6469 ( .A1(n5730), .A2(n6378), .B1(EBX_REG_20__SCAN_IN), .B2(n5373), .ZN(n5344) );
  OAI21_X1 U6470 ( .B1(n5415), .B2(n5375), .A(n5344), .ZN(U2839) );
  OAI22_X1 U6471 ( .A1(n5739), .A2(n5382), .B1(n6879), .B2(n5381), .ZN(n5345)
         );
  INV_X1 U6472 ( .A(n5345), .ZN(n5346) );
  OAI21_X1 U6473 ( .B1(n5523), .B2(n5375), .A(n5346), .ZN(U2840) );
  OAI222_X1 U6474 ( .A1(n5375), .A2(n5420), .B1(n5381), .B2(n5347), .C1(n5748), 
        .C2(n5382), .ZN(U2841) );
  OAI22_X1 U6475 ( .A1(n5756), .A2(n5382), .B1(n5348), .B2(n5381), .ZN(n5349)
         );
  INV_X1 U6476 ( .A(n5349), .ZN(n5350) );
  OAI21_X1 U6477 ( .B1(n5548), .B2(n5375), .A(n5350), .ZN(U2842) );
  INV_X1 U6478 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5351) );
  OAI222_X1 U6479 ( .A1(n5351), .A2(n5381), .B1(n5382), .B2(n5772), .C1(n6383), 
        .C2(n5375), .ZN(U2843) );
  INV_X1 U6480 ( .A(n5570), .ZN(n5424) );
  OAI222_X1 U6481 ( .A1(n5382), .A2(n5781), .B1(n5381), .B2(n5352), .C1(n5424), 
        .C2(n5375), .ZN(U2844) );
  INV_X1 U6482 ( .A(n5247), .ZN(n5353) );
  AOI21_X1 U6483 ( .B1(n5355), .B2(n5354), .A(n5353), .ZN(n6271) );
  INV_X1 U6484 ( .A(n6271), .ZN(n5426) );
  XNOR2_X1 U6485 ( .A(n4981), .B(n5356), .ZN(n6267) );
  INV_X1 U6486 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5357) );
  OAI222_X1 U6487 ( .A1(n5426), .A2(n5375), .B1(n5382), .B2(n6267), .C1(n5357), 
        .C2(n5381), .ZN(U2845) );
  OAI21_X1 U6488 ( .B1(n4980), .B2(n5359), .A(n5358), .ZN(n6286) );
  INV_X1 U6489 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6869) );
  OR2_X1 U6490 ( .A1(n5261), .A2(n5360), .ZN(n5361) );
  AND2_X1 U6491 ( .A1(n5362), .A2(n5361), .ZN(n6290) );
  INV_X1 U6492 ( .A(n6290), .ZN(n5430) );
  OAI222_X1 U6493 ( .A1(n6286), .A2(n5382), .B1(n5381), .B2(n6869), .C1(n5375), 
        .C2(n5430), .ZN(U2847) );
  OAI22_X1 U6494 ( .A1(n6479), .A2(n5382), .B1(n5363), .B2(n5381), .ZN(n5364)
         );
  INV_X1 U6495 ( .A(n5364), .ZN(n5365) );
  OAI21_X1 U6496 ( .B1(n5596), .B2(n5375), .A(n5365), .ZN(U2848) );
  AND2_X1 U6497 ( .A1(n5367), .A2(n5366), .ZN(n5369) );
  OR2_X1 U6498 ( .A1(n5369), .A2(n5368), .ZN(n6294) );
  INV_X1 U6499 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6958) );
  AOI21_X1 U6500 ( .B1(n5372), .B2(n5371), .A(n5370), .ZN(n6297) );
  INV_X1 U6501 ( .A(n6297), .ZN(n5433) );
  OAI222_X1 U6502 ( .A1(n6294), .A2(n5382), .B1(n5381), .B2(n6958), .C1(n5375), 
        .C2(n5433), .ZN(U2849) );
  AOI22_X1 U6503 ( .A1(n6489), .A2(n6378), .B1(n5373), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5374) );
  OAI21_X1 U6504 ( .B1(n5618), .B2(n5375), .A(n5374), .ZN(U2850) );
  AOI21_X1 U6505 ( .B1(n5378), .B2(n5377), .A(n5376), .ZN(n6313) );
  OR2_X1 U6506 ( .A1(n4838), .A2(n5379), .ZN(n5380) );
  NAND2_X1 U6507 ( .A1(n5278), .A2(n5380), .ZN(n6304) );
  OAI22_X1 U6508 ( .A1(n6304), .A2(n5382), .B1(n6829), .B2(n5381), .ZN(n5383)
         );
  AOI21_X1 U6509 ( .B1(n6313), .B2(n6379), .A(n5383), .ZN(n5384) );
  INV_X1 U6510 ( .A(n5384), .ZN(U2851) );
  AOI22_X1 U6511 ( .A1(n6384), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6387), .ZN(n5389) );
  NOR3_X1 U6512 ( .A1(n6387), .A2(n5386), .A3(n5385), .ZN(n5387) );
  NAND2_X1 U6513 ( .A1(n6388), .A2(DATAI_14_), .ZN(n5388) );
  OAI211_X1 U6514 ( .C1(n5019), .C2(n5438), .A(n5389), .B(n5388), .ZN(U2861)
         );
  AOI22_X1 U6515 ( .A1(n6384), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6387), .ZN(n5391) );
  NAND2_X1 U6516 ( .A1(n6388), .A2(DATAI_13_), .ZN(n5390) );
  OAI211_X1 U6517 ( .C1(n5392), .C2(n5438), .A(n5391), .B(n5390), .ZN(U2862)
         );
  AOI22_X1 U6518 ( .A1(n6384), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6387), .ZN(n5394) );
  NAND2_X1 U6519 ( .A1(n6388), .A2(DATAI_12_), .ZN(n5393) );
  OAI211_X1 U6520 ( .C1(n5395), .C2(n5438), .A(n5394), .B(n5393), .ZN(U2863)
         );
  AOI22_X1 U6521 ( .A1(n6384), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6387), .ZN(n5397) );
  NAND2_X1 U6522 ( .A1(n6388), .A2(DATAI_11_), .ZN(n5396) );
  OAI211_X1 U6523 ( .C1(n5398), .C2(n5438), .A(n5397), .B(n5396), .ZN(U2864)
         );
  AOI22_X1 U6524 ( .A1(n6384), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6387), .ZN(n5400) );
  NAND2_X1 U6525 ( .A1(n6388), .A2(DATAI_10_), .ZN(n5399) );
  OAI211_X1 U6526 ( .C1(n5456), .C2(n5438), .A(n5400), .B(n5399), .ZN(U2865)
         );
  AOI22_X1 U6527 ( .A1(n6384), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6387), .ZN(n5402) );
  NAND2_X1 U6528 ( .A1(n6388), .A2(DATAI_9_), .ZN(n5401) );
  OAI211_X1 U6529 ( .C1(n5465), .C2(n5438), .A(n5402), .B(n5401), .ZN(U2866)
         );
  AOI22_X1 U6530 ( .A1(n6384), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6387), .ZN(n5404) );
  NAND2_X1 U6531 ( .A1(n6388), .A2(DATAI_8_), .ZN(n5403) );
  OAI211_X1 U6532 ( .C1(n5405), .C2(n5438), .A(n5404), .B(n5403), .ZN(U2867)
         );
  AOI22_X1 U6533 ( .A1(n6384), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6387), .ZN(n5407) );
  NAND2_X1 U6534 ( .A1(n6388), .A2(DATAI_7_), .ZN(n5406) );
  OAI211_X1 U6535 ( .C1(n5487), .C2(n5438), .A(n5407), .B(n5406), .ZN(U2868)
         );
  AOI22_X1 U6536 ( .A1(n6384), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6387), .ZN(n5409) );
  NAND2_X1 U6537 ( .A1(n6388), .A2(DATAI_6_), .ZN(n5408) );
  OAI211_X1 U6538 ( .C1(n5410), .C2(n5438), .A(n5409), .B(n5408), .ZN(U2869)
         );
  AOI22_X1 U6539 ( .A1(n6384), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6387), .ZN(n5412) );
  NAND2_X1 U6540 ( .A1(n6388), .A2(DATAI_5_), .ZN(n5411) );
  OAI211_X1 U6541 ( .C1(n5510), .C2(n5438), .A(n5412), .B(n5411), .ZN(U2870)
         );
  AOI22_X1 U6542 ( .A1(n6384), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6387), .ZN(n5414) );
  NAND2_X1 U6543 ( .A1(n6388), .A2(DATAI_4_), .ZN(n5413) );
  OAI211_X1 U6544 ( .C1(n5415), .C2(n5438), .A(n5414), .B(n5413), .ZN(U2871)
         );
  AOI22_X1 U6545 ( .A1(n6384), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6387), .ZN(n5417) );
  NAND2_X1 U6546 ( .A1(n6388), .A2(DATAI_3_), .ZN(n5416) );
  OAI211_X1 U6547 ( .C1(n5523), .C2(n5438), .A(n5417), .B(n5416), .ZN(U2872)
         );
  AOI22_X1 U6548 ( .A1(n6384), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6387), .ZN(n5419) );
  NAND2_X1 U6549 ( .A1(n6388), .A2(DATAI_2_), .ZN(n5418) );
  OAI211_X1 U6550 ( .C1(n5420), .C2(n5438), .A(n5419), .B(n5418), .ZN(U2873)
         );
  AOI22_X1 U6551 ( .A1(n6384), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6387), .ZN(n5422) );
  NAND2_X1 U6552 ( .A1(n6388), .A2(DATAI_1_), .ZN(n5421) );
  OAI211_X1 U6553 ( .C1(n5548), .C2(n5438), .A(n5422), .B(n5421), .ZN(U2874)
         );
  AOI22_X1 U6554 ( .A1(n5434), .A2(DATAI_15_), .B1(n6387), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5423) );
  OAI21_X1 U6555 ( .B1(n5424), .B2(n5438), .A(n5423), .ZN(U2876) );
  AOI22_X1 U6556 ( .A1(n5434), .A2(DATAI_14_), .B1(n6387), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5425) );
  OAI21_X1 U6557 ( .B1(n5426), .B2(n5438), .A(n5425), .ZN(U2877) );
  INV_X1 U6558 ( .A(n6380), .ZN(n5428) );
  AOI22_X1 U6559 ( .A1(n5434), .A2(DATAI_13_), .B1(n6387), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5427) );
  OAI21_X1 U6560 ( .B1(n5428), .B2(n5438), .A(n5427), .ZN(U2878) );
  AOI22_X1 U6561 ( .A1(n5434), .A2(DATAI_12_), .B1(n6387), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5429) );
  OAI21_X1 U6562 ( .B1(n5430), .B2(n5438), .A(n5429), .ZN(U2879) );
  AOI22_X1 U6563 ( .A1(n5434), .A2(DATAI_11_), .B1(n6387), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5431) );
  OAI21_X1 U6564 ( .B1(n5596), .B2(n5438), .A(n5431), .ZN(U2880) );
  AOI22_X1 U6565 ( .A1(n5434), .A2(DATAI_10_), .B1(n6387), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5432) );
  OAI21_X1 U6566 ( .B1(n5433), .B2(n5438), .A(n5432), .ZN(U2881) );
  AOI22_X1 U6567 ( .A1(n5434), .A2(DATAI_9_), .B1(n6387), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5435) );
  OAI21_X1 U6568 ( .B1(n5618), .B2(n5438), .A(n5435), .ZN(U2882) );
  INV_X1 U6569 ( .A(n6313), .ZN(n5439) );
  INV_X1 U6570 ( .A(DATAI_8_), .ZN(n6943) );
  INV_X1 U6571 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6849) );
  OAI222_X1 U6572 ( .A1(n5439), .A2(n5438), .B1(n5437), .B2(n6943), .C1(n5436), 
        .C2(n6849), .ZN(U2883) );
  NAND2_X1 U6573 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  XNOR2_X1 U6574 ( .A(n5442), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5671)
         );
  NAND2_X1 U6575 ( .A1(n5632), .A2(n5443), .ZN(n5444) );
  NAND2_X1 U6576 ( .A1(n6465), .A2(REIP_REG_27__SCAN_IN), .ZN(n5663) );
  OAI211_X1 U6577 ( .C1(n5445), .C2(n5630), .A(n5444), .B(n5663), .ZN(n5446)
         );
  AOI21_X1 U6578 ( .B1(n5447), .B2(n6472), .A(n5446), .ZN(n5448) );
  OAI21_X1 U6579 ( .B1(n5671), .B2(n5625), .A(n5448), .ZN(U2959) );
  NOR2_X1 U6580 ( .A1(n6498), .A2(n5449), .ZN(n5674) );
  NOR2_X1 U6581 ( .A1(n6478), .A2(n5450), .ZN(n5451) );
  AOI211_X1 U6582 ( .C1(PHYADDRPOINTER_REG_26__SCAN_IN), .C2(n6466), .A(n5674), 
        .B(n5451), .ZN(n5455) );
  XNOR2_X1 U6583 ( .A(n3573), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5453)
         );
  XNOR2_X1 U6584 ( .A(n5452), .B(n5453), .ZN(n5672) );
  NAND2_X1 U6585 ( .A1(n5672), .A2(n6474), .ZN(n5454) );
  OAI211_X1 U6586 ( .C1(n5456), .C2(n6178), .A(n5455), .B(n5454), .ZN(U2960)
         );
  NAND2_X1 U6587 ( .A1(n6465), .A2(REIP_REG_25__SCAN_IN), .ZN(n5685) );
  OAI21_X1 U6588 ( .B1(n5630), .B2(n5457), .A(n5685), .ZN(n5458) );
  AOI21_X1 U6589 ( .B1(n5632), .B2(n5459), .A(n5458), .ZN(n5464) );
  OAI21_X1 U6590 ( .B1(n5462), .B2(n5461), .A(n5460), .ZN(n5684) );
  NAND2_X1 U6591 ( .A1(n5684), .A2(n6474), .ZN(n5463) );
  OAI211_X1 U6592 ( .C1(n5465), .C2(n6178), .A(n5464), .B(n5463), .ZN(U2961)
         );
  XNOR2_X1 U6593 ( .A(n5532), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5521)
         );
  AOI21_X2 U6594 ( .B1(n5519), .B2(n5521), .A(n5466), .ZN(n5513) );
  NOR2_X1 U6595 ( .A1(n5532), .A2(n5733), .ZN(n5483) );
  NAND2_X1 U6596 ( .A1(n5532), .A2(n5733), .ZN(n5482) );
  XNOR2_X1 U6597 ( .A(n3573), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5503)
         );
  NAND4_X1 U6599 ( .A1(n5532), .A2(n5467), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n5692), .ZN(n5468) );
  OAI21_X1 U6600 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5692), .A(n5468), 
        .ZN(n5476) );
  NAND2_X1 U6601 ( .A1(n3597), .A2(n5708), .ZN(n5493) );
  NOR2_X1 U6602 ( .A1(n5493), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5471)
         );
  NOR3_X1 U6603 ( .A1(n3597), .A2(n5469), .A3(n6999), .ZN(n5470) );
  NOR3_X1 U6604 ( .A1(n5471), .A2(n5470), .A3(n5692), .ZN(n5475) );
  NAND2_X1 U6605 ( .A1(n5471), .A2(n5692), .ZN(n5472) );
  AOI21_X1 U6606 ( .B1(n5473), .B2(n5472), .A(n5502), .ZN(n5474) );
  NAND2_X1 U6607 ( .A1(n6465), .A2(REIP_REG_24__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U6608 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5477)
         );
  OAI211_X1 U6609 ( .C1(n6478), .C2(n5478), .A(n5693), .B(n5477), .ZN(n5479)
         );
  AOI21_X1 U6610 ( .B1(n5480), .B2(n6472), .A(n5479), .ZN(n5481) );
  OAI21_X1 U6611 ( .B1(n5699), .B2(n5625), .A(n5481), .ZN(U2962) );
  INV_X1 U6612 ( .A(n5482), .ZN(n5484) );
  NOR2_X1 U6613 ( .A1(n5484), .A2(n5483), .ZN(n5512) );
  NAND2_X1 U6614 ( .A1(n5513), .A2(n5512), .ZN(n5511) );
  OAI22_X1 U6615 ( .A1(n5502), .A2(n5493), .B1(n5485), .B2(n5511), .ZN(n5486)
         );
  XNOR2_X1 U6616 ( .A(n5486), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5705)
         );
  INV_X1 U6617 ( .A(n5487), .ZN(n5491) );
  NAND2_X1 U6618 ( .A1(n6465), .A2(REIP_REG_23__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U6619 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5488)
         );
  OAI211_X1 U6620 ( .C1(n6478), .C2(n5489), .A(n5700), .B(n5488), .ZN(n5490)
         );
  AOI21_X1 U6621 ( .B1(n5491), .B2(n6472), .A(n5490), .ZN(n5492) );
  OAI21_X1 U6622 ( .B1(n5705), .B2(n5625), .A(n5492), .ZN(U2963) );
  OAI21_X1 U6623 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n3597), .A(n5502), 
        .ZN(n5496) );
  INV_X1 U6624 ( .A(n5493), .ZN(n5494) );
  AOI21_X1 U6625 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5532), .A(n5494), 
        .ZN(n5495) );
  XNOR2_X1 U6626 ( .A(n5496), .B(n5495), .ZN(n5713) );
  NOR2_X1 U6627 ( .A1(n6498), .A2(n7043), .ZN(n5706) );
  AOI21_X1 U6628 ( .B1(n6466), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5706), 
        .ZN(n5497) );
  OAI21_X1 U6629 ( .B1(n5498), .B2(n6478), .A(n5497), .ZN(n5499) );
  AOI21_X1 U6630 ( .B1(n5500), .B2(n6472), .A(n5499), .ZN(n5501) );
  OAI21_X1 U6631 ( .B1(n5713), .B2(n5625), .A(n5501), .ZN(U2964) );
  OAI21_X1 U6632 ( .B1(n3099), .B2(n5503), .A(n5502), .ZN(n5714) );
  NAND2_X1 U6633 ( .A1(n5714), .A2(n6474), .ZN(n5509) );
  NAND2_X1 U6634 ( .A1(n6465), .A2(REIP_REG_21__SCAN_IN), .ZN(n5716) );
  OAI21_X1 U6635 ( .B1(n5630), .B2(n5505), .A(n5716), .ZN(n5506) );
  AOI21_X1 U6636 ( .B1(n5632), .B2(n5507), .A(n5506), .ZN(n5508) );
  OAI211_X1 U6637 ( .C1(n6178), .C2(n5510), .A(n5509), .B(n5508), .ZN(U2965)
         );
  OAI21_X1 U6638 ( .B1(n5513), .B2(n5512), .A(n5511), .ZN(n5737) );
  NAND2_X1 U6639 ( .A1(n6465), .A2(REIP_REG_20__SCAN_IN), .ZN(n5731) );
  OAI21_X1 U6640 ( .B1(n5630), .B2(n7007), .A(n5731), .ZN(n5514) );
  AOI21_X1 U6641 ( .B1(n5632), .B2(n5515), .A(n5514), .ZN(n5518) );
  NAND2_X1 U6642 ( .A1(n5516), .A2(n6472), .ZN(n5517) );
  OAI211_X1 U6643 ( .C1(n5737), .C2(n5625), .A(n5518), .B(n5517), .ZN(U2966)
         );
  XOR2_X1 U6644 ( .A(n5521), .B(n5520), .Z(n5746) );
  NAND2_X1 U6645 ( .A1(n6465), .A2(REIP_REG_19__SCAN_IN), .ZN(n5738) );
  OAI21_X1 U6646 ( .B1(n5630), .B2(n5522), .A(n5738), .ZN(n5525) );
  NOR2_X1 U6647 ( .A1(n5523), .A2(n6178), .ZN(n5524) );
  OAI21_X1 U6648 ( .B1(n5746), .B2(n5625), .A(n5527), .ZN(U2967) );
  AOI21_X2 U6650 ( .B1(n5572), .B2(n5531), .A(n5530), .ZN(n5565) );
  XNOR2_X1 U6651 ( .A(n5532), .B(n6928), .ZN(n5566) );
  INV_X2 U6652 ( .A(n5535), .ZN(n5555) );
  NAND2_X1 U6653 ( .A1(n5532), .A2(n5768), .ZN(n5556) );
  NAND2_X2 U6654 ( .A1(n5555), .A2(n5556), .ZN(n5554) );
  INV_X1 U6655 ( .A(n5536), .ZN(n5534) );
  XNOR2_X1 U6656 ( .A(n5537), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5754)
         );
  NAND2_X1 U6657 ( .A1(n5632), .A2(n5538), .ZN(n5539) );
  NAND2_X1 U6658 ( .A1(n6465), .A2(REIP_REG_18__SCAN_IN), .ZN(n5747) );
  OAI211_X1 U6659 ( .C1(n5630), .C2(n5540), .A(n5539), .B(n5747), .ZN(n5541)
         );
  AOI21_X1 U6660 ( .B1(n5542), .B2(n6472), .A(n5541), .ZN(n5543) );
  OAI21_X1 U6661 ( .B1(n5754), .B2(n5625), .A(n5543), .ZN(U2968) );
  INV_X1 U6662 ( .A(n5544), .ZN(n5547) );
  OR2_X1 U6663 ( .A1(n5532), .A2(n5768), .ZN(n5558) );
  XNOR2_X1 U6664 ( .A(n3573), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5545)
         );
  AOI21_X1 U6665 ( .B1(n5554), .B2(n5558), .A(n5545), .ZN(n5546) );
  AOI21_X1 U6666 ( .B1(n5547), .B2(n5554), .A(n5546), .ZN(n5762) );
  INV_X1 U6667 ( .A(n5548), .ZN(n5552) );
  NAND2_X1 U6668 ( .A1(n6465), .A2(REIP_REG_17__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U6669 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5549)
         );
  OAI211_X1 U6670 ( .C1(n6478), .C2(n5550), .A(n5755), .B(n5549), .ZN(n5551)
         );
  AOI21_X1 U6671 ( .B1(n5552), .B2(n6472), .A(n5551), .ZN(n5553) );
  OAI21_X1 U6672 ( .B1(n5762), .B2(n5625), .A(n5553), .ZN(U2969) );
  INV_X1 U6673 ( .A(n5554), .ZN(n5559) );
  AOI21_X1 U6674 ( .B1(n5556), .B2(n5558), .A(n5555), .ZN(n5557) );
  AOI21_X1 U6675 ( .B1(n5559), .B2(n5558), .A(n5557), .ZN(n5775) );
  NAND2_X1 U6676 ( .A1(n5775), .A2(n6474), .ZN(n5564) );
  NAND2_X1 U6677 ( .A1(n6465), .A2(REIP_REG_16__SCAN_IN), .ZN(n5770) );
  OAI21_X1 U6678 ( .B1(n5630), .B2(n5560), .A(n5770), .ZN(n5561) );
  AOI21_X1 U6679 ( .B1(n5632), .B2(n5562), .A(n5561), .ZN(n5563) );
  OAI211_X1 U6680 ( .C1(n6178), .C2(n6383), .A(n5564), .B(n5563), .ZN(U2970)
         );
  XOR2_X1 U6681 ( .A(n5566), .B(n3100), .Z(n5785) );
  NOR2_X1 U6682 ( .A1(n6498), .A2(n7023), .ZN(n5778) );
  AOI21_X1 U6683 ( .B1(n6466), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5778), 
        .ZN(n5567) );
  OAI21_X1 U6684 ( .B1(n5568), .B2(n6478), .A(n5567), .ZN(n5569) );
  AOI21_X1 U6685 ( .B1(n5570), .B2(n6472), .A(n5569), .ZN(n5571) );
  OAI21_X1 U6686 ( .B1(n5785), .B2(n5625), .A(n5571), .ZN(U2971) );
  XNOR2_X1 U6687 ( .A(n3573), .B(n5788), .ZN(n5573) );
  XNOR2_X1 U6688 ( .A(n5572), .B(n5573), .ZN(n5794) );
  NAND2_X1 U6689 ( .A1(n6465), .A2(REIP_REG_14__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U6690 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5574)
         );
  OAI211_X1 U6691 ( .C1(n6478), .C2(n6269), .A(n5786), .B(n5574), .ZN(n5575)
         );
  AOI21_X1 U6692 ( .B1(n6271), .B2(n6472), .A(n5575), .ZN(n5576) );
  OAI21_X1 U6693 ( .B1(n5794), .B2(n5625), .A(n5576), .ZN(U2972) );
  INV_X1 U6694 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U6695 ( .A1(n5578), .A2(n5597), .ZN(n5590) );
  NOR2_X1 U6696 ( .A1(n3573), .A2(n6486), .ZN(n5589) );
  AOI21_X1 U6697 ( .B1(n5590), .B2(n5587), .A(n5589), .ZN(n5582) );
  OAI21_X1 U6698 ( .B1(n5532), .B2(n5580), .A(n5579), .ZN(n5581) );
  XNOR2_X1 U6699 ( .A(n5582), .B(n5581), .ZN(n5804) );
  INV_X1 U6700 ( .A(n6289), .ZN(n5584) );
  AOI22_X1 U6701 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6465), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5583) );
  OAI21_X1 U6702 ( .B1(n6478), .B2(n5584), .A(n5583), .ZN(n5585) );
  AOI21_X1 U6703 ( .B1(n6290), .B2(n6472), .A(n5585), .ZN(n5586) );
  OAI21_X1 U6704 ( .B1(n5804), .B2(n5625), .A(n5586), .ZN(U2974) );
  INV_X1 U6705 ( .A(n5587), .ZN(n5588) );
  NOR2_X1 U6706 ( .A1(n5589), .A2(n5588), .ZN(n5591) );
  XOR2_X1 U6707 ( .A(n5591), .B(n5590), .Z(n6483) );
  NAND2_X1 U6708 ( .A1(n6483), .A2(n6474), .ZN(n5595) );
  NOR2_X1 U6709 ( .A1(n6498), .A2(n5272), .ZN(n6480) );
  NOR2_X1 U6710 ( .A1(n6478), .A2(n5592), .ZN(n5593) );
  AOI211_X1 U6711 ( .C1(n6466), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6480), 
        .B(n5593), .ZN(n5594) );
  OAI211_X1 U6712 ( .C1(n6178), .C2(n5596), .A(n5595), .B(n5594), .ZN(U2975)
         );
  INV_X1 U6713 ( .A(n5597), .ZN(n5599) );
  NOR2_X1 U6714 ( .A1(n5599), .A2(n5598), .ZN(n5607) );
  NAND2_X1 U6715 ( .A1(n5619), .A2(n5620), .ZN(n5602) );
  NAND2_X1 U6716 ( .A1(n5602), .A2(n5601), .ZN(n5613) );
  OR2_X1 U6717 ( .A1(n5613), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U6718 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  XOR2_X1 U6719 ( .A(n5607), .B(n5606), .Z(n5812) );
  INV_X1 U6720 ( .A(n6296), .ZN(n5609) );
  AOI22_X1 U6721 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6465), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5608) );
  OAI21_X1 U6722 ( .B1(n6478), .B2(n5609), .A(n5608), .ZN(n5610) );
  AOI21_X1 U6723 ( .B1(n6297), .B2(n6472), .A(n5610), .ZN(n5611) );
  OAI21_X1 U6724 ( .B1(n5812), .B2(n5625), .A(n5611), .ZN(U2976) );
  XNOR2_X1 U6725 ( .A(n3573), .B(n5808), .ZN(n5612) );
  XNOR2_X1 U6726 ( .A(n5613), .B(n5612), .ZN(n6490) );
  NAND2_X1 U6727 ( .A1(n6490), .A2(n6474), .ZN(n5617) );
  NOR2_X1 U6728 ( .A1(n6498), .A2(n6675), .ZN(n6488) );
  NOR2_X1 U6729 ( .A1(n6478), .A2(n5614), .ZN(n5615) );
  AOI211_X1 U6730 ( .C1(n6466), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6488), 
        .B(n5615), .ZN(n5616) );
  OAI211_X1 U6731 ( .C1(n6178), .C2(n5618), .A(n5617), .B(n5616), .ZN(U2977)
         );
  XNOR2_X1 U6732 ( .A(n5620), .B(n5619), .ZN(n5821) );
  NAND2_X1 U6733 ( .A1(n6465), .A2(REIP_REG_8__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U6734 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5621)
         );
  OAI211_X1 U6735 ( .C1(n6478), .C2(n5622), .A(n5814), .B(n5621), .ZN(n5623)
         );
  AOI21_X1 U6736 ( .B1(n6313), .B2(n6472), .A(n5623), .ZN(n5624) );
  OAI21_X1 U6737 ( .B1(n5821), .B2(n5625), .A(n5624), .ZN(U2978) );
  AND2_X1 U6738 ( .A1(n5628), .A2(n5627), .ZN(n5629) );
  XOR2_X1 U6739 ( .A(n5626), .B(n5629), .Z(n5828) );
  NAND2_X1 U6740 ( .A1(n5828), .A2(n6474), .ZN(n5634) );
  NAND2_X1 U6741 ( .A1(n6465), .A2(REIP_REG_7__SCAN_IN), .ZN(n5825) );
  OAI21_X1 U6742 ( .B1(n5630), .B2(n6882), .A(n5825), .ZN(n5631) );
  AOI21_X1 U6743 ( .B1(n5632), .B2(n6322), .A(n5631), .ZN(n5633) );
  OAI211_X1 U6744 ( .C1(n6178), .C2(n6325), .A(n5634), .B(n5633), .ZN(U2979)
         );
  NAND2_X1 U6746 ( .A1(n3106), .A2(n5638), .ZN(n5639) );
  XNOR2_X1 U6747 ( .A(n5635), .B(n5639), .ZN(n5837) );
  INV_X1 U6748 ( .A(n6340), .ZN(n5641) );
  AOI22_X1 U6749 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6465), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n5640) );
  OAI21_X1 U6750 ( .B1(n5641), .B2(n6478), .A(n5640), .ZN(n5642) );
  AOI21_X1 U6751 ( .B1(n6341), .B2(n6472), .A(n5642), .ZN(n5643) );
  OAI21_X1 U6752 ( .B1(n5625), .B2(n5837), .A(n5643), .ZN(U2980) );
  INV_X1 U6753 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U6754 ( .A1(n5645), .A2(n6472), .ZN(n5650) );
  NAND2_X1 U6755 ( .A1(n6465), .A2(REIP_REG_0__SCAN_IN), .ZN(n6512) );
  NOR2_X1 U6756 ( .A1(n5646), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6514)
         );
  OR3_X1 U6757 ( .A1(n6513), .A2(n6514), .A3(n5625), .ZN(n5649) );
  OAI21_X1 U6758 ( .B1(n6466), .B2(n5647), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5648) );
  NAND4_X1 U6759 ( .A1(n5650), .A2(n6512), .A3(n5649), .A4(n5648), .ZN(U2986)
         );
  INV_X1 U6760 ( .A(n5651), .ZN(n5662) );
  INV_X1 U6761 ( .A(n5668), .ZN(n5660) );
  INV_X1 U6762 ( .A(n5652), .ZN(n5654) );
  NAND3_X1 U6763 ( .A1(n5666), .A2(n5654), .A3(n5653), .ZN(n5657) );
  INV_X1 U6764 ( .A(n5655), .ZN(n5656) );
  OAI211_X1 U6765 ( .C1(n6500), .C2(n5658), .A(n5657), .B(n5656), .ZN(n5659)
         );
  AOI21_X1 U6766 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5660), .A(n5659), 
        .ZN(n5661) );
  OAI21_X1 U6767 ( .B1(n5662), .B2(n6515), .A(n5661), .ZN(U2990) );
  OAI21_X1 U6768 ( .B1(n5664), .B2(n6500), .A(n5663), .ZN(n5665) );
  AOI21_X1 U6769 ( .B1(n5666), .B2(n5667), .A(n5665), .ZN(n5670) );
  OR2_X1 U6770 ( .A1(n5668), .A2(n5667), .ZN(n5669) );
  OAI211_X1 U6771 ( .C1(n5671), .C2(n6515), .A(n5670), .B(n5669), .ZN(U2991)
         );
  NAND2_X1 U6772 ( .A1(n5672), .A2(n6502), .ZN(n5683) );
  INV_X1 U6773 ( .A(n5673), .ZN(n5675) );
  AOI21_X1 U6774 ( .B1(n5675), .B2(n6518), .A(n5674), .ZN(n5682) );
  NAND2_X1 U6775 ( .A1(n5697), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5681) );
  INV_X1 U6776 ( .A(n5687), .ZN(n5679) );
  INV_X1 U6777 ( .A(n5676), .ZN(n5677) );
  NAND3_X1 U6778 ( .A1(n5679), .A2(n5678), .A3(n5677), .ZN(n5680) );
  NAND4_X1 U6779 ( .A1(n5683), .A2(n5682), .A3(n5681), .A4(n5680), .ZN(U2992)
         );
  INV_X1 U6780 ( .A(n5684), .ZN(n5691) );
  OAI21_X1 U6781 ( .B1(n5686), .B2(n6500), .A(n5685), .ZN(n5689) );
  NOR2_X1 U6782 ( .A1(n5687), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5688)
         );
  AOI211_X1 U6783 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5697), .A(n5689), .B(n5688), .ZN(n5690) );
  OAI21_X1 U6784 ( .B1(n5691), .B2(n6515), .A(n5690), .ZN(U2993) );
  OAI21_X1 U6785 ( .B1(n3132), .B2(n6999), .A(n5692), .ZN(n5696) );
  OAI21_X1 U6786 ( .B1(n5694), .B2(n6500), .A(n5693), .ZN(n5695) );
  AOI21_X1 U6787 ( .B1(n5697), .B2(n5696), .A(n5695), .ZN(n5698) );
  OAI21_X1 U6788 ( .B1(n5699), .B2(n6515), .A(n5698), .ZN(U2994) );
  OAI21_X1 U6789 ( .B1(n5701), .B2(n6500), .A(n5700), .ZN(n5703) );
  NOR2_X1 U6790 ( .A1(n3132), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5702)
         );
  AOI211_X1 U6791 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5710), .A(n5703), .B(n5702), .ZN(n5704) );
  OAI21_X1 U6792 ( .B1(n5705), .B2(n6515), .A(n5704), .ZN(U2995) );
  AOI21_X1 U6793 ( .B1(n5707), .B2(n6518), .A(n5706), .ZN(n5712) );
  OAI21_X1 U6794 ( .B1(n5722), .B2(n6925), .A(n5708), .ZN(n5709) );
  NAND2_X1 U6795 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  OAI211_X1 U6796 ( .C1(n5713), .C2(n6515), .A(n5712), .B(n5711), .ZN(U2996)
         );
  NAND2_X1 U6797 ( .A1(n5714), .A2(n6502), .ZN(n5721) );
  INV_X1 U6798 ( .A(n5715), .ZN(n5719) );
  OAI21_X1 U6799 ( .B1(n5717), .B2(n6500), .A(n5716), .ZN(n5718) );
  AOI21_X1 U6800 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5719), .A(n5718), 
        .ZN(n5720) );
  OAI211_X1 U6801 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5722), .A(n5721), .B(n5720), .ZN(U2997) );
  NOR2_X1 U6802 ( .A1(n5724), .A2(n5723), .ZN(n5735) );
  INV_X1 U6803 ( .A(n5760), .ZN(n5727) );
  NAND2_X1 U6804 ( .A1(n5725), .A2(n6942), .ZN(n5726) );
  NAND2_X1 U6805 ( .A1(n5727), .A2(n5726), .ZN(n5752) );
  AND2_X1 U6806 ( .A1(n5765), .A2(n5728), .ZN(n5729) );
  NOR2_X1 U6807 ( .A1(n5752), .A2(n5729), .ZN(n5740) );
  NAND2_X1 U6808 ( .A1(n5730), .A2(n6518), .ZN(n5732) );
  OAI211_X1 U6809 ( .C1(n5740), .C2(n5733), .A(n5732), .B(n5731), .ZN(n5734)
         );
  AOI21_X1 U6810 ( .B1(n5744), .B2(n5735), .A(n5734), .ZN(n5736) );
  OAI21_X1 U6811 ( .B1(n5737), .B2(n6515), .A(n5736), .ZN(U2998) );
  OAI21_X1 U6812 ( .B1(n5739), .B2(n6500), .A(n5738), .ZN(n5742) );
  NOR2_X1 U6813 ( .A1(n5740), .A2(n5743), .ZN(n5741) );
  AOI211_X1 U6814 ( .C1(n5744), .C2(n5743), .A(n5742), .B(n5741), .ZN(n5745)
         );
  OAI21_X1 U6815 ( .B1(n5746), .B2(n6515), .A(n5745), .ZN(U2999) );
  OAI21_X1 U6816 ( .B1(n5748), .B2(n6500), .A(n5747), .ZN(n5751) );
  NOR2_X1 U6817 ( .A1(n5749), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5750)
         );
  AOI211_X1 U6818 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n5752), .A(n5751), .B(n5750), .ZN(n5753) );
  OAI21_X1 U6819 ( .B1(n5754), .B2(n6515), .A(n5753), .ZN(U3000) );
  OAI21_X1 U6820 ( .B1(n5756), .B2(n6500), .A(n5755), .ZN(n5759) );
  INV_X1 U6821 ( .A(n6482), .ZN(n5797) );
  NOR3_X1 U6822 ( .A1(n5797), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5757), 
        .ZN(n5758) );
  AOI211_X1 U6823 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5760), .A(n5759), .B(n5758), .ZN(n5761) );
  OAI21_X1 U6824 ( .B1(n5762), .B2(n6515), .A(n5761), .ZN(U3001) );
  INV_X1 U6825 ( .A(n5763), .ZN(n5766) );
  INV_X1 U6826 ( .A(n6487), .ZN(n5764) );
  AOI21_X1 U6827 ( .B1(n5766), .B2(n5765), .A(n5764), .ZN(n5777) );
  AND2_X1 U6828 ( .A1(n6482), .A2(n5767), .ZN(n5789) );
  NAND3_X1 U6829 ( .A1(n5789), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n6928), .ZN(n5780) );
  AOI21_X1 U6830 ( .B1(n5777), .B2(n5780), .A(n5768), .ZN(n5774) );
  NAND3_X1 U6831 ( .A1(n6482), .A2(n5769), .A3(n5768), .ZN(n5771) );
  OAI211_X1 U6832 ( .C1(n6500), .C2(n5772), .A(n5771), .B(n5770), .ZN(n5773)
         );
  AOI211_X1 U6833 ( .C1(n5775), .C2(n6502), .A(n5774), .B(n5773), .ZN(n5776)
         );
  INV_X1 U6834 ( .A(n5776), .ZN(U3002) );
  INV_X1 U6835 ( .A(n5777), .ZN(n5783) );
  INV_X1 U6836 ( .A(n5778), .ZN(n5779) );
  OAI211_X1 U6837 ( .C1(n6500), .C2(n5781), .A(n5780), .B(n5779), .ZN(n5782)
         );
  AOI21_X1 U6838 ( .B1(n5783), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5782), 
        .ZN(n5784) );
  OAI21_X1 U6839 ( .B1(n5785), .B2(n6515), .A(n5784), .ZN(U3003) );
  OAI21_X1 U6840 ( .B1(n6267), .B2(n6500), .A(n5786), .ZN(n5787) );
  AOI21_X1 U6841 ( .B1(n5789), .B2(n5788), .A(n5787), .ZN(n5793) );
  OAI21_X1 U6842 ( .B1(n5791), .B2(n5790), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5792) );
  OAI211_X1 U6843 ( .C1(n5794), .C2(n6515), .A(n5793), .B(n5792), .ZN(U3004)
         );
  INV_X1 U6844 ( .A(n6286), .ZN(n5802) );
  INV_X1 U6845 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6679) );
  OAI221_X1 U6846 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5796), .C1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n5795), .A(n6487), .ZN(n5799) );
  NOR3_X1 U6847 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5797), .A3(n6486), 
        .ZN(n5798) );
  AOI21_X1 U6848 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n5799), .A(n5798), 
        .ZN(n5800) );
  OAI21_X1 U6849 ( .B1(n6498), .B2(n6679), .A(n5800), .ZN(n5801) );
  AOI21_X1 U6850 ( .B1(n5802), .B2(n6518), .A(n5801), .ZN(n5803) );
  OAI21_X1 U6851 ( .B1(n5804), .B2(n6515), .A(n5803), .ZN(U3006) );
  OAI21_X1 U6852 ( .B1(n5805), .B2(n5813), .A(n5816), .ZN(n6491) );
  INV_X1 U6853 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6677) );
  OAI22_X1 U6854 ( .A1(n6294), .A2(n6500), .B1(n6677), .B2(n6498), .ZN(n5810)
         );
  NOR2_X1 U6855 ( .A1(n5832), .A2(n5806), .ZN(n5823) );
  NAND2_X1 U6856 ( .A1(n5813), .A2(n5823), .ZN(n6494) );
  AOI221_X1 U6857 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5808), .C2(n5807), .A(n6494), 
        .ZN(n5809) );
  AOI211_X1 U6858 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6491), .A(n5810), .B(n5809), .ZN(n5811) );
  OAI21_X1 U6859 ( .B1(n6515), .B2(n5812), .A(n5811), .ZN(U3008) );
  AOI21_X1 U6860 ( .B1(n5822), .B2(n5815), .A(n5813), .ZN(n5819) );
  OAI21_X1 U6861 ( .B1(n6500), .B2(n6304), .A(n5814), .ZN(n5818) );
  NOR2_X1 U6862 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  AOI211_X1 U6863 ( .C1(n5819), .C2(n5823), .A(n5818), .B(n5817), .ZN(n5820)
         );
  OAI21_X1 U6864 ( .B1(n6515), .B2(n5821), .A(n5820), .ZN(U3010) );
  AOI22_X1 U6865 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n5824), .B1(n5823), 
        .B2(n5822), .ZN(n5826) );
  OAI211_X1 U6866 ( .C1(n6500), .C2(n6319), .A(n5826), .B(n5825), .ZN(n5827)
         );
  AOI21_X1 U6867 ( .B1(n5828), .B2(n6502), .A(n5827), .ZN(n5829) );
  INV_X1 U6868 ( .A(n5829), .ZN(U3011) );
  INV_X1 U6869 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6669) );
  OAI22_X1 U6870 ( .A1(n6500), .A2(n6336), .B1(n6669), .B2(n6498), .ZN(n5834)
         );
  INV_X1 U6871 ( .A(n5830), .ZN(n5831) );
  NOR3_X1 U6872 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5832), .A3(n5831), 
        .ZN(n5833) );
  AOI211_X1 U6873 ( .C1(INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n5835), .A(n5834), 
        .B(n5833), .ZN(n5836) );
  OAI21_X1 U6874 ( .B1(n6515), .B2(n5837), .A(n5836), .ZN(U3012) );
  NOR2_X1 U6875 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4599), .ZN(n5857) );
  OAI222_X1 U6876 ( .A1(n6120), .A2(n5998), .B1(n5857), .B2(n3679), .C1(n5839), 
        .C2(n5838), .ZN(n5843) );
  NOR2_X1 U6877 ( .A1(n5839), .A2(FLUSH_REG_SCAN_IN), .ZN(n5842) );
  OAI21_X1 U6878 ( .B1(n5842), .B2(n5841), .A(n5840), .ZN(n6524) );
  MUX2_X1 U6879 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n5843), .S(n6524), 
        .Z(U3465) );
  OAI211_X1 U6880 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5906), .A(n5847), .B(
        n6186), .ZN(n5844) );
  OAI21_X1 U6881 ( .B1(n4436), .B2(n5857), .A(n5844), .ZN(n5845) );
  MUX2_X1 U6882 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5845), .S(n6524), 
        .Z(U3464) );
  AOI21_X1 U6883 ( .B1(n5852), .B2(n5847), .A(n5846), .ZN(n5850) );
  INV_X1 U6884 ( .A(n5848), .ZN(n5849) );
  OAI22_X1 U6885 ( .A1(n5850), .A2(n5998), .B1(n5849), .B2(n5857), .ZN(n5851)
         );
  MUX2_X1 U6886 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5851), .S(n6524), 
        .Z(U3463) );
  INV_X1 U6887 ( .A(n5852), .ZN(n5856) );
  AOI211_X1 U6888 ( .C1(n5856), .C2(n5855), .A(n5854), .B(n5853), .ZN(n5858)
         );
  OAI222_X1 U6889 ( .A1(n6177), .A2(n5859), .B1(n5998), .B2(n5858), .C1(n5857), 
        .C2(n6070), .ZN(n5860) );
  MUX2_X1 U6890 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5860), .S(n6524), 
        .Z(U3462) );
  NAND3_X1 U6891 ( .A1(n5899), .A2(n6186), .A3(n6223), .ZN(n5863) );
  AOI21_X1 U6892 ( .B1(n5863), .B2(n6177), .A(n5862), .ZN(n5867) );
  OAI21_X1 U6893 ( .B1(n6782), .B2(n6079), .A(n5864), .ZN(n5910) );
  AND2_X1 U6894 ( .A1(n5865), .A2(n6072), .ZN(n5896) );
  OAI21_X1 U6895 ( .B1(n5896), .B2(n6864), .A(n6080), .ZN(n5866) );
  NOR3_X2 U6896 ( .A1(n5867), .A2(n5910), .A3(n5866), .ZN(n5904) );
  INV_X1 U6897 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5872) );
  NAND3_X1 U6898 ( .A1(n6075), .A2(n6033), .A3(n6079), .ZN(n5868) );
  OAI21_X1 U6899 ( .B1(n6529), .B2(n5992), .A(n5868), .ZN(n5897) );
  INV_X1 U6900 ( .A(n6083), .ZN(n6531) );
  AOI22_X1 U6901 ( .A1(n6532), .A2(n5897), .B1(n6531), .B2(n5896), .ZN(n5869)
         );
  OAI21_X1 U6902 ( .B1(n5899), .B2(n6542), .A(n5869), .ZN(n5870) );
  AOI21_X1 U6903 ( .B1(n6539), .B2(n5901), .A(n5870), .ZN(n5871) );
  OAI21_X1 U6904 ( .B1(n5904), .B2(n5872), .A(n5871), .ZN(U3020) );
  INV_X1 U6905 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5876) );
  INV_X1 U6906 ( .A(n6575), .ZN(n6543) );
  AOI22_X1 U6907 ( .A1(n6578), .A2(n5897), .B1(n6543), .B2(n5896), .ZN(n5873)
         );
  OAI21_X1 U6908 ( .B1(n5899), .B2(n6576), .A(n5873), .ZN(n5874) );
  AOI21_X1 U6909 ( .B1(n6544), .B2(n5901), .A(n5874), .ZN(n5875) );
  OAI21_X1 U6910 ( .B1(n5904), .B2(n5876), .A(n5875), .ZN(U3021) );
  INV_X1 U6911 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5880) );
  INV_X1 U6912 ( .A(n6603), .ZN(n6547) );
  AOI22_X1 U6913 ( .A1(n6606), .A2(n5897), .B1(n6547), .B2(n5896), .ZN(n5877)
         );
  OAI21_X1 U6914 ( .B1(n5899), .B2(n6604), .A(n5877), .ZN(n5878) );
  AOI21_X1 U6915 ( .B1(n6548), .B2(n5901), .A(n5878), .ZN(n5879) );
  OAI21_X1 U6916 ( .B1(n5904), .B2(n5880), .A(n5879), .ZN(U3022) );
  INV_X1 U6917 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5884) );
  INV_X1 U6918 ( .A(n6610), .ZN(n6551) );
  AOI22_X1 U6919 ( .A1(n6613), .A2(n5897), .B1(n6551), .B2(n5896), .ZN(n5881)
         );
  OAI21_X1 U6920 ( .B1(n5899), .B2(n6611), .A(n5881), .ZN(n5882) );
  AOI21_X1 U6921 ( .B1(n6552), .B2(n5901), .A(n5882), .ZN(n5883) );
  OAI21_X1 U6922 ( .B1(n5904), .B2(n5884), .A(n5883), .ZN(U3023) );
  INV_X1 U6923 ( .A(n6617), .ZN(n6555) );
  AOI22_X1 U6924 ( .A1(n6620), .A2(n5897), .B1(n6555), .B2(n5896), .ZN(n5885)
         );
  OAI21_X1 U6925 ( .B1(n5899), .B2(n6618), .A(n5885), .ZN(n5886) );
  AOI21_X1 U6926 ( .B1(n6556), .B2(n5901), .A(n5886), .ZN(n5887) );
  OAI21_X1 U6927 ( .B1(n5904), .B2(n7014), .A(n5887), .ZN(U3024) );
  INV_X1 U6928 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5891) );
  INV_X1 U6929 ( .A(n6588), .ZN(n6559) );
  AOI22_X1 U6930 ( .A1(n6591), .A2(n5897), .B1(n6559), .B2(n5896), .ZN(n5888)
         );
  OAI21_X1 U6931 ( .B1(n5899), .B2(n6589), .A(n5888), .ZN(n5889) );
  AOI21_X1 U6932 ( .B1(n6560), .B2(n5901), .A(n5889), .ZN(n5890) );
  OAI21_X1 U6933 ( .B1(n5904), .B2(n5891), .A(n5890), .ZN(U3025) );
  INV_X1 U6934 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5895) );
  INV_X1 U6935 ( .A(n6624), .ZN(n6563) );
  AOI22_X1 U6936 ( .A1(n6627), .A2(n5897), .B1(n6563), .B2(n5896), .ZN(n5892)
         );
  OAI21_X1 U6937 ( .B1(n5899), .B2(n6625), .A(n5892), .ZN(n5893) );
  AOI21_X1 U6938 ( .B1(n6564), .B2(n5901), .A(n5893), .ZN(n5894) );
  OAI21_X1 U6939 ( .B1(n5904), .B2(n5895), .A(n5894), .ZN(U3026) );
  INV_X1 U6940 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5903) );
  INV_X1 U6941 ( .A(n6632), .ZN(n6568) );
  AOI22_X1 U6942 ( .A1(n6636), .A2(n5897), .B1(n6568), .B2(n5896), .ZN(n5898)
         );
  OAI21_X1 U6943 ( .B1(n5899), .B2(n6633), .A(n5898), .ZN(n5900) );
  AOI21_X1 U6944 ( .B1(n6571), .B2(n5901), .A(n5900), .ZN(n5902) );
  OAI21_X1 U6945 ( .B1(n5904), .B2(n5903), .A(n5902), .ZN(U3027) );
  AOI22_X1 U6946 ( .A1(n5905), .A2(n6177), .B1(n5951), .B2(n6082), .ZN(n5911)
         );
  AOI21_X1 U6947 ( .B1(n5957), .B2(STATEBS16_REG_SCAN_IN), .A(n5998), .ZN(
        n5961) );
  NOR2_X1 U6948 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5908) );
  AND2_X1 U6949 ( .A1(n5908), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5963)
         );
  AND2_X1 U6950 ( .A1(n5963), .A2(n6072), .ZN(n5943) );
  OAI21_X1 U6951 ( .B1(n5943), .B2(n6864), .A(n6122), .ZN(n5909) );
  AOI211_X1 U6952 ( .C1(n5911), .C2(n5961), .A(n5910), .B(n5909), .ZN(n5918)
         );
  INV_X1 U6953 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5917) );
  INV_X1 U6954 ( .A(n5957), .ZN(n5912) );
  INV_X1 U6955 ( .A(n6080), .ZN(n6526) );
  NAND3_X1 U6956 ( .A1(n6526), .A2(n6033), .A3(n6079), .ZN(n5913) );
  OAI21_X1 U6957 ( .B1(n6529), .B2(n6071), .A(n5913), .ZN(n5944) );
  AOI22_X1 U6958 ( .A1(n6532), .A2(n5944), .B1(n6531), .B2(n5943), .ZN(n5914)
         );
  OAI21_X1 U6959 ( .B1(n5947), .B2(n6133), .A(n5914), .ZN(n5915) );
  AOI21_X1 U6960 ( .B1(n6135), .B2(n5958), .A(n5915), .ZN(n5916) );
  OAI21_X1 U6961 ( .B1(n5918), .B2(n5917), .A(n5916), .ZN(U3052) );
  INV_X1 U6962 ( .A(n5918), .ZN(n5949) );
  AOI22_X1 U6963 ( .A1(n6578), .A2(n5944), .B1(n6543), .B2(n5943), .ZN(n5920)
         );
  NAND2_X1 U6964 ( .A1(n5958), .A2(n6140), .ZN(n5919) );
  OAI211_X1 U6965 ( .C1(n5947), .C2(n6581), .A(n5920), .B(n5919), .ZN(n5921)
         );
  AOI21_X1 U6966 ( .B1(n5949), .B2(INSTQUEUE_REG_4__1__SCAN_IN), .A(n5921), 
        .ZN(n5922) );
  INV_X1 U6967 ( .A(n5922), .ZN(U3053) );
  AOI22_X1 U6968 ( .A1(n6606), .A2(n5944), .B1(n6547), .B2(n5943), .ZN(n5924)
         );
  NAND2_X1 U6969 ( .A1(n5958), .A2(n6145), .ZN(n5923) );
  OAI211_X1 U6970 ( .C1(n5947), .C2(n6609), .A(n5924), .B(n5923), .ZN(n5925)
         );
  AOI21_X1 U6971 ( .B1(n5949), .B2(INSTQUEUE_REG_4__2__SCAN_IN), .A(n5925), 
        .ZN(n5926) );
  INV_X1 U6972 ( .A(n5926), .ZN(U3054) );
  AOI22_X1 U6973 ( .A1(n6613), .A2(n5944), .B1(n6551), .B2(n5943), .ZN(n5928)
         );
  NAND2_X1 U6974 ( .A1(n5958), .A2(n6150), .ZN(n5927) );
  OAI211_X1 U6975 ( .C1(n5947), .C2(n6616), .A(n5928), .B(n5927), .ZN(n5929)
         );
  AOI21_X1 U6976 ( .B1(n5949), .B2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n5929), 
        .ZN(n5930) );
  INV_X1 U6977 ( .A(n5930), .ZN(U3055) );
  AOI22_X1 U6978 ( .A1(n6620), .A2(n5944), .B1(n6555), .B2(n5943), .ZN(n5932)
         );
  NAND2_X1 U6979 ( .A1(n5958), .A2(n6155), .ZN(n5931) );
  OAI211_X1 U6980 ( .C1(n5947), .C2(n6623), .A(n5932), .B(n5931), .ZN(n5933)
         );
  AOI21_X1 U6981 ( .B1(n5949), .B2(INSTQUEUE_REG_4__4__SCAN_IN), .A(n5933), 
        .ZN(n5934) );
  INV_X1 U6982 ( .A(n5934), .ZN(U3056) );
  AOI22_X1 U6983 ( .A1(n6591), .A2(n5944), .B1(n6559), .B2(n5943), .ZN(n5936)
         );
  NAND2_X1 U6984 ( .A1(n5958), .A2(n6160), .ZN(n5935) );
  OAI211_X1 U6985 ( .C1(n5947), .C2(n6594), .A(n5936), .B(n5935), .ZN(n5937)
         );
  AOI21_X1 U6986 ( .B1(n5949), .B2(INSTQUEUE_REG_4__5__SCAN_IN), .A(n5937), 
        .ZN(n5938) );
  INV_X1 U6987 ( .A(n5938), .ZN(U3057) );
  AOI22_X1 U6988 ( .A1(n6627), .A2(n5944), .B1(n6563), .B2(n5943), .ZN(n5940)
         );
  NAND2_X1 U6989 ( .A1(n5958), .A2(n6165), .ZN(n5939) );
  OAI211_X1 U6990 ( .C1(n5947), .C2(n6630), .A(n5940), .B(n5939), .ZN(n5941)
         );
  AOI21_X1 U6991 ( .B1(n5949), .B2(INSTQUEUE_REG_4__6__SCAN_IN), .A(n5941), 
        .ZN(n5942) );
  INV_X1 U6992 ( .A(n5942), .ZN(U3058) );
  AOI22_X1 U6993 ( .A1(n6636), .A2(n5944), .B1(n6568), .B2(n5943), .ZN(n5946)
         );
  NAND2_X1 U6994 ( .A1(n5958), .A2(n6173), .ZN(n5945) );
  OAI211_X1 U6995 ( .C1(n5947), .C2(n6642), .A(n5946), .B(n5945), .ZN(n5948)
         );
  AOI21_X1 U6996 ( .B1(n5949), .B2(INSTQUEUE_REG_4__7__SCAN_IN), .A(n5948), 
        .ZN(n5950) );
  INV_X1 U6997 ( .A(n5950), .ZN(U3059) );
  AND2_X1 U6998 ( .A1(n5952), .A2(n5951), .ZN(n5954) );
  NAND2_X1 U6999 ( .A1(n5963), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5984) );
  INV_X1 U7000 ( .A(n5984), .ZN(n5953) );
  AOI21_X1 U7001 ( .B1(n6082), .B2(n5954), .A(n5953), .ZN(n5960) );
  INV_X1 U7002 ( .A(n5960), .ZN(n5955) );
  AOI22_X1 U7003 ( .A1(n5961), .A2(n5955), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5963), .ZN(n5990) );
  OAI22_X1 U7004 ( .A1(n5985), .A2(n6133), .B1(n6083), .B2(n5984), .ZN(n5959)
         );
  AOI21_X1 U7005 ( .B1(n6135), .B2(n6570), .A(n5959), .ZN(n5965) );
  NAND2_X1 U7006 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  NAND2_X1 U7007 ( .A1(n5987), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5964) );
  OAI211_X1 U7008 ( .C1(n5990), .C2(n6084), .A(n5965), .B(n5964), .ZN(U3060)
         );
  OAI22_X1 U7009 ( .A1(n5985), .A2(n6581), .B1(n6575), .B2(n5984), .ZN(n5966)
         );
  AOI21_X1 U7010 ( .B1(n6140), .B2(n6570), .A(n5966), .ZN(n5968) );
  NAND2_X1 U7011 ( .A1(n5987), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5967) );
  OAI211_X1 U7012 ( .C1(n5990), .C2(n6088), .A(n5968), .B(n5967), .ZN(U3061)
         );
  OAI22_X1 U7013 ( .A1(n5985), .A2(n6609), .B1(n6603), .B2(n5984), .ZN(n5969)
         );
  AOI21_X1 U7014 ( .B1(n6145), .B2(n6570), .A(n5969), .ZN(n5971) );
  NAND2_X1 U7015 ( .A1(n5987), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5970) );
  OAI211_X1 U7016 ( .C1(n5990), .C2(n6092), .A(n5971), .B(n5970), .ZN(U3062)
         );
  OAI22_X1 U7017 ( .A1(n5985), .A2(n6616), .B1(n6610), .B2(n5984), .ZN(n5972)
         );
  AOI21_X1 U7018 ( .B1(n6150), .B2(n6570), .A(n5972), .ZN(n5974) );
  NAND2_X1 U7019 ( .A1(n5987), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5973) );
  OAI211_X1 U7020 ( .C1(n5990), .C2(n6096), .A(n5974), .B(n5973), .ZN(U3063)
         );
  OAI22_X1 U7021 ( .A1(n5985), .A2(n6623), .B1(n6617), .B2(n5984), .ZN(n5975)
         );
  AOI21_X1 U7022 ( .B1(n6155), .B2(n6570), .A(n5975), .ZN(n5977) );
  NAND2_X1 U7023 ( .A1(n5987), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5976) );
  OAI211_X1 U7024 ( .C1(n5990), .C2(n6100), .A(n5977), .B(n5976), .ZN(U3064)
         );
  OAI22_X1 U7025 ( .A1(n5985), .A2(n6594), .B1(n6588), .B2(n5984), .ZN(n5978)
         );
  AOI21_X1 U7026 ( .B1(n6160), .B2(n6570), .A(n5978), .ZN(n5980) );
  NAND2_X1 U7027 ( .A1(n5987), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5979) );
  OAI211_X1 U7028 ( .C1(n5990), .C2(n6104), .A(n5980), .B(n5979), .ZN(U3065)
         );
  OAI22_X1 U7029 ( .A1(n5985), .A2(n6630), .B1(n6624), .B2(n5984), .ZN(n5981)
         );
  AOI21_X1 U7030 ( .B1(n6165), .B2(n6570), .A(n5981), .ZN(n5983) );
  NAND2_X1 U7031 ( .A1(n5987), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5982) );
  OAI211_X1 U7032 ( .C1(n5990), .C2(n6108), .A(n5983), .B(n5982), .ZN(U3066)
         );
  OAI22_X1 U7033 ( .A1(n5985), .A2(n6642), .B1(n6632), .B2(n5984), .ZN(n5986)
         );
  AOI21_X1 U7034 ( .B1(n6173), .B2(n6570), .A(n5986), .ZN(n5989) );
  NAND2_X1 U7035 ( .A1(n5987), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5988) );
  OAI211_X1 U7036 ( .C1(n5990), .C2(n6114), .A(n5989), .B(n5988), .ZN(U3067)
         );
  INV_X1 U7037 ( .A(n5995), .ZN(n5991) );
  AOI21_X1 U7038 ( .B1(n5991), .B2(STATEBS16_REG_SCAN_IN), .A(n5998), .ZN(
        n5997) );
  OR2_X1 U7039 ( .A1(n5999), .A2(n6072), .ZN(n6023) );
  OAI21_X1 U7040 ( .B1(n6180), .B2(n5992), .A(n6023), .ZN(n6001) );
  INV_X1 U7041 ( .A(n5999), .ZN(n5993) );
  AOI22_X1 U7042 ( .A1(n5997), .A2(n6001), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5993), .ZN(n6030) );
  INV_X1 U7043 ( .A(n6065), .ZN(n6024) );
  OAI22_X1 U7044 ( .A1(n6024), .A2(n6542), .B1(n6083), .B2(n6023), .ZN(n5996)
         );
  AOI21_X1 U7045 ( .B1(n6539), .B2(n6026), .A(n5996), .ZN(n6004) );
  INV_X1 U7046 ( .A(n5997), .ZN(n6002) );
  NAND2_X1 U7047 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  NAND2_X1 U7048 ( .A1(n6027), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6003) );
  OAI211_X1 U7049 ( .C1(n6030), .C2(n6084), .A(n6004), .B(n6003), .ZN(U3092)
         );
  OAI22_X1 U7050 ( .A1(n6024), .A2(n6576), .B1(n6575), .B2(n6023), .ZN(n6005)
         );
  AOI21_X1 U7051 ( .B1(n6544), .B2(n6026), .A(n6005), .ZN(n6007) );
  NAND2_X1 U7052 ( .A1(n6027), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6006) );
  OAI211_X1 U7053 ( .C1(n6030), .C2(n6088), .A(n6007), .B(n6006), .ZN(U3093)
         );
  OAI22_X1 U7054 ( .A1(n6024), .A2(n6604), .B1(n6603), .B2(n6023), .ZN(n6008)
         );
  AOI21_X1 U7055 ( .B1(n6548), .B2(n6026), .A(n6008), .ZN(n6010) );
  NAND2_X1 U7056 ( .A1(n6027), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6009) );
  OAI211_X1 U7057 ( .C1(n6030), .C2(n6092), .A(n6010), .B(n6009), .ZN(U3094)
         );
  OAI22_X1 U7058 ( .A1(n6024), .A2(n6611), .B1(n6610), .B2(n6023), .ZN(n6011)
         );
  AOI21_X1 U7059 ( .B1(n6552), .B2(n6026), .A(n6011), .ZN(n6013) );
  NAND2_X1 U7060 ( .A1(n6027), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6012) );
  OAI211_X1 U7061 ( .C1(n6030), .C2(n6096), .A(n6013), .B(n6012), .ZN(U3095)
         );
  OAI22_X1 U7062 ( .A1(n6024), .A2(n6618), .B1(n6617), .B2(n6023), .ZN(n6014)
         );
  AOI21_X1 U7063 ( .B1(n6556), .B2(n6026), .A(n6014), .ZN(n6016) );
  NAND2_X1 U7064 ( .A1(n6027), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6015) );
  OAI211_X1 U7065 ( .C1(n6030), .C2(n6100), .A(n6016), .B(n6015), .ZN(U3096)
         );
  OAI22_X1 U7066 ( .A1(n6024), .A2(n6589), .B1(n6588), .B2(n6023), .ZN(n6017)
         );
  AOI21_X1 U7067 ( .B1(n6560), .B2(n6026), .A(n6017), .ZN(n6019) );
  NAND2_X1 U7068 ( .A1(n6027), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6018) );
  OAI211_X1 U7069 ( .C1(n6030), .C2(n6104), .A(n6019), .B(n6018), .ZN(U3097)
         );
  OAI22_X1 U7070 ( .A1(n6024), .A2(n6625), .B1(n6624), .B2(n6023), .ZN(n6020)
         );
  AOI21_X1 U7071 ( .B1(n6564), .B2(n6026), .A(n6020), .ZN(n6022) );
  NAND2_X1 U7072 ( .A1(n6027), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6021) );
  OAI211_X1 U7073 ( .C1(n6030), .C2(n6108), .A(n6022), .B(n6021), .ZN(U3098)
         );
  OAI22_X1 U7074 ( .A1(n6024), .A2(n6633), .B1(n6632), .B2(n6023), .ZN(n6025)
         );
  AOI21_X1 U7075 ( .B1(n6571), .B2(n6026), .A(n6025), .ZN(n6029) );
  NAND2_X1 U7076 ( .A1(n6027), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n6028) );
  OAI211_X1 U7077 ( .C1(n6030), .C2(n6114), .A(n6029), .B(n6028), .ZN(U3099)
         );
  INV_X1 U7078 ( .A(n6641), .ZN(n6031) );
  OAI21_X1 U7079 ( .B1(n6065), .B2(n6031), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6032) );
  NAND2_X1 U7080 ( .A1(n6032), .A2(n6186), .ZN(n6040) );
  INV_X1 U7081 ( .A(n6040), .ZN(n6035) );
  NOR3_X1 U7082 ( .A1(n6122), .A2(n6033), .A3(n6535), .ZN(n6034) );
  NAND2_X1 U7083 ( .A1(n6036), .A2(n6072), .ZN(n6063) );
  AOI211_X1 U7084 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6063), .A(n6037), .B(
        n6526), .ZN(n6038) );
  NAND2_X1 U7085 ( .A1(n6062), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6043)
         );
  OAI22_X1 U7086 ( .A1(n6641), .A2(n6542), .B1(n6063), .B2(n6083), .ZN(n6041)
         );
  AOI21_X1 U7087 ( .B1(n6065), .B2(n6539), .A(n6041), .ZN(n6042) );
  OAI211_X1 U7088 ( .C1(n6068), .C2(n6084), .A(n6043), .B(n6042), .ZN(U3100)
         );
  NAND2_X1 U7089 ( .A1(n6062), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6046)
         );
  OAI22_X1 U7090 ( .A1(n6641), .A2(n6576), .B1(n6063), .B2(n6575), .ZN(n6044)
         );
  AOI21_X1 U7091 ( .B1(n6065), .B2(n6544), .A(n6044), .ZN(n6045) );
  OAI211_X1 U7092 ( .C1(n6068), .C2(n6088), .A(n6046), .B(n6045), .ZN(U3101)
         );
  NAND2_X1 U7093 ( .A1(n6062), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6049)
         );
  OAI22_X1 U7094 ( .A1(n6641), .A2(n6604), .B1(n6063), .B2(n6603), .ZN(n6047)
         );
  AOI21_X1 U7095 ( .B1(n6065), .B2(n6548), .A(n6047), .ZN(n6048) );
  OAI211_X1 U7096 ( .C1(n6068), .C2(n6092), .A(n6049), .B(n6048), .ZN(U3102)
         );
  NAND2_X1 U7097 ( .A1(n6062), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6052)
         );
  OAI22_X1 U7098 ( .A1(n6641), .A2(n6611), .B1(n6063), .B2(n6610), .ZN(n6050)
         );
  AOI21_X1 U7099 ( .B1(n6065), .B2(n6552), .A(n6050), .ZN(n6051) );
  OAI211_X1 U7100 ( .C1(n6068), .C2(n6096), .A(n6052), .B(n6051), .ZN(U3103)
         );
  NAND2_X1 U7101 ( .A1(n6062), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6055)
         );
  OAI22_X1 U7102 ( .A1(n6641), .A2(n6618), .B1(n6063), .B2(n6617), .ZN(n6053)
         );
  AOI21_X1 U7103 ( .B1(n6065), .B2(n6556), .A(n6053), .ZN(n6054) );
  OAI211_X1 U7104 ( .C1(n6068), .C2(n6100), .A(n6055), .B(n6054), .ZN(U3104)
         );
  NAND2_X1 U7105 ( .A1(n6062), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6058)
         );
  OAI22_X1 U7106 ( .A1(n6641), .A2(n6589), .B1(n6063), .B2(n6588), .ZN(n6056)
         );
  AOI21_X1 U7107 ( .B1(n6065), .B2(n6560), .A(n6056), .ZN(n6057) );
  OAI211_X1 U7108 ( .C1(n6068), .C2(n6104), .A(n6058), .B(n6057), .ZN(U3105)
         );
  NAND2_X1 U7109 ( .A1(n6062), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6061)
         );
  OAI22_X1 U7110 ( .A1(n6641), .A2(n6625), .B1(n6063), .B2(n6624), .ZN(n6059)
         );
  AOI21_X1 U7111 ( .B1(n6065), .B2(n6564), .A(n6059), .ZN(n6060) );
  OAI211_X1 U7112 ( .C1(n6068), .C2(n6108), .A(n6061), .B(n6060), .ZN(U3106)
         );
  NAND2_X1 U7113 ( .A1(n6062), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6067)
         );
  OAI22_X1 U7114 ( .A1(n6641), .A2(n6633), .B1(n6063), .B2(n6632), .ZN(n6064)
         );
  AOI21_X1 U7115 ( .B1(n6065), .B2(n6571), .A(n6064), .ZN(n6066) );
  OAI211_X1 U7116 ( .C1(n6068), .C2(n6114), .A(n6067), .B(n6066), .ZN(U3107)
         );
  AOI21_X1 U7117 ( .B1(n6634), .B2(n6069), .A(n6245), .ZN(n6078) );
  OAI21_X1 U7118 ( .B1(n6071), .B2(n6070), .A(n6186), .ZN(n6077) );
  NAND2_X1 U7119 ( .A1(n6073), .A2(n6072), .ZN(n6113) );
  AOI211_X1 U7120 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6113), .A(n6075), .B(
        n6074), .ZN(n6076) );
  NAND2_X1 U7121 ( .A1(n6112), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6087)
         );
  NOR3_X1 U7122 ( .A1(n6080), .A2(n6525), .A3(n6079), .ZN(n6081) );
  AOI21_X1 U7123 ( .B1(n6129), .B2(n6082), .A(n6081), .ZN(n6115) );
  OAI22_X1 U7124 ( .A1(n6115), .A2(n6084), .B1(n6083), .B2(n6113), .ZN(n6085)
         );
  AOI21_X1 U7125 ( .B1(n6117), .B2(n6135), .A(n6085), .ZN(n6086) );
  OAI211_X1 U7126 ( .C1(n6634), .C2(n6133), .A(n6087), .B(n6086), .ZN(U3116)
         );
  NAND2_X1 U7127 ( .A1(n6112), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6091)
         );
  OAI22_X1 U7128 ( .A1(n6115), .A2(n6088), .B1(n6575), .B2(n6113), .ZN(n6089)
         );
  AOI21_X1 U7129 ( .B1(n6140), .B2(n6117), .A(n6089), .ZN(n6090) );
  OAI211_X1 U7130 ( .C1(n6634), .C2(n6581), .A(n6091), .B(n6090), .ZN(U3117)
         );
  NAND2_X1 U7131 ( .A1(n6112), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6095)
         );
  OAI22_X1 U7132 ( .A1(n6115), .A2(n6092), .B1(n6603), .B2(n6113), .ZN(n6093)
         );
  AOI21_X1 U7133 ( .B1(n6145), .B2(n6117), .A(n6093), .ZN(n6094) );
  OAI211_X1 U7134 ( .C1(n6634), .C2(n6609), .A(n6095), .B(n6094), .ZN(U3118)
         );
  NAND2_X1 U7135 ( .A1(n6112), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6099)
         );
  OAI22_X1 U7136 ( .A1(n6115), .A2(n6096), .B1(n6610), .B2(n6113), .ZN(n6097)
         );
  AOI21_X1 U7137 ( .B1(n6150), .B2(n6117), .A(n6097), .ZN(n6098) );
  OAI211_X1 U7138 ( .C1(n6634), .C2(n6616), .A(n6099), .B(n6098), .ZN(U3119)
         );
  NAND2_X1 U7139 ( .A1(n6112), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6103)
         );
  OAI22_X1 U7140 ( .A1(n6115), .A2(n6100), .B1(n6617), .B2(n6113), .ZN(n6101)
         );
  AOI21_X1 U7141 ( .B1(n6155), .B2(n6117), .A(n6101), .ZN(n6102) );
  OAI211_X1 U7142 ( .C1(n6634), .C2(n6623), .A(n6103), .B(n6102), .ZN(U3120)
         );
  NAND2_X1 U7143 ( .A1(n6112), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6107)
         );
  OAI22_X1 U7144 ( .A1(n6115), .A2(n6104), .B1(n6588), .B2(n6113), .ZN(n6105)
         );
  AOI21_X1 U7145 ( .B1(n6160), .B2(n6117), .A(n6105), .ZN(n6106) );
  OAI211_X1 U7146 ( .C1(n6634), .C2(n6594), .A(n6107), .B(n6106), .ZN(U3121)
         );
  NAND2_X1 U7147 ( .A1(n6112), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6111)
         );
  OAI22_X1 U7148 ( .A1(n6115), .A2(n6108), .B1(n6624), .B2(n6113), .ZN(n6109)
         );
  AOI21_X1 U7149 ( .B1(n6165), .B2(n6117), .A(n6109), .ZN(n6110) );
  OAI211_X1 U7150 ( .C1(n6634), .C2(n6630), .A(n6111), .B(n6110), .ZN(U3122)
         );
  NAND2_X1 U7151 ( .A1(n6112), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6119)
         );
  OAI22_X1 U7152 ( .A1(n6115), .A2(n6114), .B1(n6632), .B2(n6113), .ZN(n6116)
         );
  AOI21_X1 U7153 ( .B1(n6173), .B2(n6117), .A(n6116), .ZN(n6118) );
  OAI211_X1 U7154 ( .C1(n6634), .C2(n6642), .A(n6119), .B(n6118), .ZN(U3123)
         );
  NAND2_X1 U7155 ( .A1(n6528), .A2(n6186), .ZN(n6533) );
  AOI211_X1 U7156 ( .C1(n6529), .C2(n6533), .A(n6225), .B(n6121), .ZN(n6128)
         );
  OAI211_X1 U7157 ( .C1(n6124), .C2(n6177), .A(n6123), .B(n6122), .ZN(n6537)
         );
  NOR2_X1 U7158 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6125), .ZN(n6168)
         );
  OAI21_X1 U7159 ( .B1(n6168), .B2(n6864), .A(n6126), .ZN(n6127) );
  NOR3_X2 U7160 ( .A1(n6128), .A2(n6537), .A3(n6127), .ZN(n6176) );
  INV_X1 U7161 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6137) );
  INV_X1 U7162 ( .A(n6129), .ZN(n6131) );
  NAND3_X1 U7163 ( .A1(n6526), .A2(n6525), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6130) );
  OAI21_X1 U7164 ( .B1(n6131), .B2(n6528), .A(n6130), .ZN(n6169) );
  AOI22_X1 U7165 ( .A1(n6169), .A2(n6532), .B1(n6531), .B2(n6168), .ZN(n6132)
         );
  OAI21_X1 U7166 ( .B1(n6133), .B2(n6171), .A(n6132), .ZN(n6134) );
  AOI21_X1 U7167 ( .B1(n6135), .B2(n6225), .A(n6134), .ZN(n6136) );
  OAI21_X1 U7168 ( .B1(n6176), .B2(n6137), .A(n6136), .ZN(U3132) );
  INV_X1 U7169 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6142) );
  AOI22_X1 U7170 ( .A1(n6169), .A2(n6578), .B1(n6543), .B2(n6168), .ZN(n6138)
         );
  OAI21_X1 U7171 ( .B1(n6171), .B2(n6581), .A(n6138), .ZN(n6139) );
  AOI21_X1 U7172 ( .B1(n6140), .B2(n6225), .A(n6139), .ZN(n6141) );
  OAI21_X1 U7173 ( .B1(n6176), .B2(n6142), .A(n6141), .ZN(U3133) );
  INV_X1 U7174 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6147) );
  AOI22_X1 U7175 ( .A1(n6169), .A2(n6606), .B1(n6547), .B2(n6168), .ZN(n6143)
         );
  OAI21_X1 U7176 ( .B1(n6171), .B2(n6609), .A(n6143), .ZN(n6144) );
  AOI21_X1 U7177 ( .B1(n6145), .B2(n6225), .A(n6144), .ZN(n6146) );
  OAI21_X1 U7178 ( .B1(n6176), .B2(n6147), .A(n6146), .ZN(U3134) );
  INV_X1 U7179 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6152) );
  AOI22_X1 U7180 ( .A1(n6169), .A2(n6613), .B1(n6551), .B2(n6168), .ZN(n6148)
         );
  OAI21_X1 U7181 ( .B1(n6171), .B2(n6616), .A(n6148), .ZN(n6149) );
  AOI21_X1 U7182 ( .B1(n6150), .B2(n6225), .A(n6149), .ZN(n6151) );
  OAI21_X1 U7183 ( .B1(n6176), .B2(n6152), .A(n6151), .ZN(U3135) );
  INV_X1 U7184 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6157) );
  AOI22_X1 U7185 ( .A1(n6169), .A2(n6620), .B1(n6555), .B2(n6168), .ZN(n6153)
         );
  OAI21_X1 U7186 ( .B1(n6171), .B2(n6623), .A(n6153), .ZN(n6154) );
  AOI21_X1 U7187 ( .B1(n6155), .B2(n6225), .A(n6154), .ZN(n6156) );
  OAI21_X1 U7188 ( .B1(n6176), .B2(n6157), .A(n6156), .ZN(U3136) );
  INV_X1 U7189 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6162) );
  AOI22_X1 U7190 ( .A1(n6169), .A2(n6591), .B1(n6559), .B2(n6168), .ZN(n6158)
         );
  OAI21_X1 U7191 ( .B1(n6171), .B2(n6594), .A(n6158), .ZN(n6159) );
  AOI21_X1 U7192 ( .B1(n6160), .B2(n6225), .A(n6159), .ZN(n6161) );
  OAI21_X1 U7193 ( .B1(n6176), .B2(n6162), .A(n6161), .ZN(U3137) );
  INV_X1 U7194 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6167) );
  AOI22_X1 U7195 ( .A1(n6169), .A2(n6627), .B1(n6563), .B2(n6168), .ZN(n6163)
         );
  OAI21_X1 U7196 ( .B1(n6171), .B2(n6630), .A(n6163), .ZN(n6164) );
  AOI21_X1 U7197 ( .B1(n6165), .B2(n6225), .A(n6164), .ZN(n6166) );
  OAI21_X1 U7198 ( .B1(n6176), .B2(n6167), .A(n6166), .ZN(U3138) );
  INV_X1 U7199 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6175) );
  AOI22_X1 U7200 ( .A1(n6169), .A2(n6636), .B1(n6568), .B2(n6168), .ZN(n6170)
         );
  OAI21_X1 U7201 ( .B1(n6171), .B2(n6642), .A(n6170), .ZN(n6172) );
  AOI21_X1 U7202 ( .B1(n6173), .B2(n6225), .A(n6172), .ZN(n6174) );
  OAI21_X1 U7203 ( .B1(n6176), .B2(n6175), .A(n6174), .ZN(U3139) );
  OAI21_X1 U7204 ( .B1(n6179), .B2(n6178), .A(n6177), .ZN(n6185) );
  OR2_X1 U7205 ( .A1(n6180), .A2(n6528), .ZN(n6181) );
  NAND2_X1 U7206 ( .A1(n6181), .A2(n6191), .ZN(n6187) );
  INV_X1 U7207 ( .A(n6187), .ZN(n6184) );
  OAI21_X1 U7208 ( .B1(n6186), .B2(n6188), .A(n6182), .ZN(n6183) );
  INV_X1 U7209 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7210 ( .A1(n6187), .A2(n6186), .ZN(n6190) );
  NAND2_X1 U7211 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6188), .ZN(n6189) );
  NAND2_X1 U7212 ( .A1(n6190), .A2(n6189), .ZN(n6221) );
  INV_X1 U7213 ( .A(n6191), .ZN(n6220) );
  AOI22_X1 U7214 ( .A1(n6221), .A2(n6532), .B1(n6220), .B2(n6531), .ZN(n6192)
         );
  OAI21_X1 U7215 ( .B1(n6223), .B2(n6542), .A(n6192), .ZN(n6193) );
  AOI21_X1 U7216 ( .B1(n6539), .B2(n6225), .A(n6193), .ZN(n6194) );
  OAI21_X1 U7217 ( .B1(n6228), .B2(n6195), .A(n6194), .ZN(U3140) );
  INV_X1 U7218 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6199) );
  AOI22_X1 U7219 ( .A1(n6221), .A2(n6578), .B1(n6220), .B2(n6543), .ZN(n6196)
         );
  OAI21_X1 U7220 ( .B1(n6223), .B2(n6576), .A(n6196), .ZN(n6197) );
  AOI21_X1 U7221 ( .B1(n6544), .B2(n6225), .A(n6197), .ZN(n6198) );
  OAI21_X1 U7222 ( .B1(n6228), .B2(n6199), .A(n6198), .ZN(U3141) );
  INV_X1 U7223 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6203) );
  AOI22_X1 U7224 ( .A1(n6221), .A2(n6606), .B1(n6220), .B2(n6547), .ZN(n6200)
         );
  OAI21_X1 U7225 ( .B1(n6223), .B2(n6604), .A(n6200), .ZN(n6201) );
  AOI21_X1 U7226 ( .B1(n6548), .B2(n6225), .A(n6201), .ZN(n6202) );
  OAI21_X1 U7227 ( .B1(n6228), .B2(n6203), .A(n6202), .ZN(U3142) );
  INV_X1 U7228 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6207) );
  AOI22_X1 U7229 ( .A1(n6221), .A2(n6613), .B1(n6220), .B2(n6551), .ZN(n6204)
         );
  OAI21_X1 U7230 ( .B1(n6223), .B2(n6611), .A(n6204), .ZN(n6205) );
  AOI21_X1 U7231 ( .B1(n6552), .B2(n6225), .A(n6205), .ZN(n6206) );
  OAI21_X1 U7232 ( .B1(n6228), .B2(n6207), .A(n6206), .ZN(U3143) );
  INV_X1 U7233 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6211) );
  AOI22_X1 U7234 ( .A1(n6221), .A2(n6620), .B1(n6220), .B2(n6555), .ZN(n6208)
         );
  OAI21_X1 U7235 ( .B1(n6223), .B2(n6618), .A(n6208), .ZN(n6209) );
  AOI21_X1 U7236 ( .B1(n6556), .B2(n6225), .A(n6209), .ZN(n6210) );
  OAI21_X1 U7237 ( .B1(n6228), .B2(n6211), .A(n6210), .ZN(U3144) );
  INV_X1 U7238 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6215) );
  AOI22_X1 U7239 ( .A1(n6221), .A2(n6591), .B1(n6220), .B2(n6559), .ZN(n6212)
         );
  OAI21_X1 U7240 ( .B1(n6223), .B2(n6589), .A(n6212), .ZN(n6213) );
  AOI21_X1 U7241 ( .B1(n6560), .B2(n6225), .A(n6213), .ZN(n6214) );
  OAI21_X1 U7242 ( .B1(n6228), .B2(n6215), .A(n6214), .ZN(U3145) );
  INV_X1 U7243 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6219) );
  AOI22_X1 U7244 ( .A1(n6221), .A2(n6627), .B1(n6220), .B2(n6563), .ZN(n6216)
         );
  OAI21_X1 U7245 ( .B1(n6223), .B2(n6625), .A(n6216), .ZN(n6217) );
  AOI21_X1 U7246 ( .B1(n6564), .B2(n6225), .A(n6217), .ZN(n6218) );
  OAI21_X1 U7247 ( .B1(n6228), .B2(n6219), .A(n6218), .ZN(U3146) );
  INV_X1 U7248 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n6227) );
  AOI22_X1 U7249 ( .A1(n6221), .A2(n6636), .B1(n6220), .B2(n6568), .ZN(n6222)
         );
  OAI21_X1 U7250 ( .B1(n6223), .B2(n6633), .A(n6222), .ZN(n6224) );
  AOI21_X1 U7251 ( .B1(n6571), .B2(n6225), .A(n6224), .ZN(n6226) );
  OAI21_X1 U7252 ( .B1(n6228), .B2(n6227), .A(n6226), .ZN(U3147) );
  INV_X1 U7253 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n6876) );
  NOR2_X1 U7254 ( .A1(n6876), .A2(n6419), .ZN(U2892) );
  AOI21_X1 U7255 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n6230), .A(n6229), .ZN(
        n6231) );
  INV_X1 U7256 ( .A(n6231), .ZN(U2788) );
  INV_X1 U7257 ( .A(n6232), .ZN(n6236) );
  INV_X1 U7258 ( .A(n6233), .ZN(n6367) );
  NAND4_X1 U7259 ( .A1(n6236), .A2(n6367), .A3(n6235), .A4(n6234), .ZN(n6237)
         );
  OAI21_X1 U7260 ( .B1(n6720), .B2(n6238), .A(n6237), .ZN(U3455) );
  INV_X1 U7261 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6992) );
  AOI21_X1 U7262 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6992), .A(n4106), .ZN(n6243) );
  INV_X1 U7263 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6239) );
  AOI21_X1 U7264 ( .B1(n6243), .B2(n6239), .A(n6746), .ZN(U2789) );
  OAI21_X1 U7265 ( .B1(n6240), .B2(n6646), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6241) );
  OAI21_X1 U7266 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6647), .A(n6241), .ZN(
        U2790) );
  NOR2_X1 U7267 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6244) );
  OAI21_X1 U7268 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6244), .A(n6734), .ZN(n6242)
         );
  OAI21_X1 U7269 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6734), .A(n6242), .ZN(
        U2791) );
  NOR2_X1 U7270 ( .A1(n6746), .A2(n6243), .ZN(n6711) );
  OAI21_X1 U7271 ( .B1(n6244), .B2(BS16_N), .A(n6711), .ZN(n6709) );
  OAI21_X1 U7272 ( .B1(n6711), .B2(n6245), .A(n6709), .ZN(U2792) );
  INV_X1 U7273 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6246) );
  OAI21_X1 U7274 ( .B1(n6247), .B2(n6246), .A(n5625), .ZN(U2793) );
  NOR2_X1 U7275 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n6791) );
  AOI211_X1 U7276 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_13__SCAN_IN), .B(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n6248) );
  INV_X1 U7277 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6964) );
  INV_X1 U7278 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6934) );
  NAND4_X1 U7279 ( .A1(n6791), .A2(n6248), .A3(n6964), .A4(n6934), .ZN(n6256)
         );
  OR4_X1 U7280 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6255) );
  OR4_X1 U7281 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(
        n6254) );
  NOR4_X1 U7282 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n6252) );
  NOR4_X1 U7283 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6251) );
  NOR4_X1 U7284 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6250) );
  NOR4_X1 U7285 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6249) );
  NAND4_X1 U7286 ( .A1(n6252), .A2(n6251), .A3(n6250), .A4(n6249), .ZN(n6253)
         );
  NOR4_X2 U7287 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n6732)
         );
  INV_X1 U7288 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6258) );
  NOR3_X1 U7289 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7290 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6259), .A(n6732), .ZN(n6257)
         );
  OAI21_X1 U7291 ( .B1(n6732), .B2(n6258), .A(n6257), .ZN(U2794) );
  INV_X1 U7292 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6261) );
  NOR2_X1 U7293 ( .A1(REIP_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n6726) );
  OAI21_X1 U7294 ( .B1(n6259), .B2(n6726), .A(n6732), .ZN(n6260) );
  OAI21_X1 U7295 ( .B1(n6732), .B2(n6261), .A(n6260), .ZN(U2795) );
  INV_X1 U7296 ( .A(n6262), .ZN(n6265) );
  OAI21_X1 U7297 ( .B1(n6360), .B2(n6263), .A(n7025), .ZN(n6264) );
  AOI22_X1 U7298 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6358), .B1(n6265), .B2(n6264), .ZN(n6274) );
  INV_X1 U7299 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6266) );
  OAI22_X1 U7300 ( .A1(n6267), .A2(n6335), .B1(n6266), .B2(n6348), .ZN(n6268)
         );
  INV_X1 U7301 ( .A(n6268), .ZN(n6273) );
  INV_X1 U7302 ( .A(n6269), .ZN(n6270) );
  AOI22_X1 U7303 ( .A1(n6271), .A2(n3093), .B1(n6270), .B2(n3129), .ZN(n6272)
         );
  NAND4_X1 U7304 ( .A1(n6274), .A2(n6273), .A3(n6272), .A4(n6346), .ZN(U2813)
         );
  NOR3_X1 U7305 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6360), .A3(n6275), .ZN(n6276) );
  AOI211_X1 U7306 ( .C1(n6363), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6362), 
        .B(n6276), .ZN(n6284) );
  INV_X1 U7307 ( .A(n6277), .ZN(n6377) );
  AOI22_X1 U7308 ( .A1(n6377), .A2(n6366), .B1(EBX_REG_13__SCAN_IN), .B2(n6358), .ZN(n6283) );
  INV_X1 U7309 ( .A(n6278), .ZN(n6279) );
  AOI22_X1 U7310 ( .A1(n6380), .A2(n3093), .B1(n6279), .B2(n3129), .ZN(n6282)
         );
  NOR3_X1 U7311 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6360), .A3(n6280), .ZN(n6288) );
  OAI21_X1 U7312 ( .B1(n6288), .B2(n6285), .A(REIP_REG_13__SCAN_IN), .ZN(n6281) );
  NAND4_X1 U7313 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(U2814)
         );
  AOI22_X1 U7314 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6358), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6285), .ZN(n6293) );
  OAI21_X1 U7315 ( .B1(n6286), .B2(n6335), .A(n6346), .ZN(n6287) );
  AOI211_X1 U7316 ( .C1(n6363), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6288), 
        .B(n6287), .ZN(n6292) );
  AOI22_X1 U7317 ( .A1(n6290), .A2(n3093), .B1(n3129), .B2(n6289), .ZN(n6291)
         );
  NAND3_X1 U7318 ( .A1(n6293), .A2(n6292), .A3(n6291), .ZN(U2815) );
  OAI22_X1 U7319 ( .A1(n6310), .A2(n6958), .B1(n6335), .B2(n6294), .ZN(n6295)
         );
  AOI211_X1 U7320 ( .C1(n6363), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6362), 
        .B(n6295), .ZN(n6303) );
  AOI22_X1 U7321 ( .A1(n6297), .A2(n3093), .B1(n3129), .B2(n6296), .ZN(n6302)
         );
  OAI21_X1 U7322 ( .B1(n6298), .B2(n6306), .A(REIP_REG_10__SCAN_IN), .ZN(n6301) );
  NAND3_X1 U7323 ( .A1(n6329), .A2(n6299), .A3(n6677), .ZN(n6300) );
  NAND4_X1 U7324 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .ZN(U2817)
         );
  INV_X1 U7325 ( .A(n6304), .ZN(n6305) );
  AOI22_X1 U7326 ( .A1(n6306), .A2(REIP_REG_8__SCAN_IN), .B1(n6366), .B2(n6305), .ZN(n6316) );
  INV_X1 U7327 ( .A(n6307), .ZN(n6309) );
  OAI22_X1 U7328 ( .A1(n6310), .A2(n6829), .B1(n6309), .B2(n6308), .ZN(n6311)
         );
  AOI211_X1 U7329 ( .C1(n6363), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6362), 
        .B(n6311), .ZN(n6315) );
  AOI22_X1 U7330 ( .A1(n6313), .A2(n3093), .B1(n3129), .B2(n6312), .ZN(n6314)
         );
  NAND3_X1 U7331 ( .A1(n6316), .A2(n6315), .A3(n6314), .ZN(U2819) );
  INV_X1 U7332 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6672) );
  AOI21_X1 U7333 ( .B1(n6329), .B2(n6318), .A(n6317), .ZN(n6344) );
  INV_X1 U7334 ( .A(n6319), .ZN(n6320) );
  AOI22_X1 U7335 ( .A1(n6358), .A2(EBX_REG_7__SCAN_IN), .B1(n6366), .B2(n6320), 
        .ZN(n6321) );
  OAI211_X1 U7336 ( .C1(n6348), .C2(n6882), .A(n6321), .B(n6346), .ZN(n6327)
         );
  INV_X1 U7337 ( .A(n6322), .ZN(n6323) );
  OAI22_X1 U7338 ( .A1(n6325), .A2(n3130), .B1(n6323), .B2(n5027), .ZN(n6326)
         );
  NOR2_X1 U7339 ( .A1(n6327), .A2(n6326), .ZN(n6332) );
  NAND2_X1 U7340 ( .A1(n6329), .A2(n6328), .ZN(n6345) );
  NOR2_X1 U7341 ( .A1(n6667), .A2(n6345), .ZN(n6338) );
  OAI211_X1 U7342 ( .C1(REIP_REG_7__SCAN_IN), .C2(REIP_REG_6__SCAN_IN), .A(
        n6338), .B(n6330), .ZN(n6331) );
  OAI211_X1 U7343 ( .C1(n6672), .C2(n6344), .A(n6332), .B(n6331), .ZN(U2820)
         );
  INV_X1 U7344 ( .A(n6344), .ZN(n6339) );
  NAND2_X1 U7345 ( .A1(n6358), .A2(EBX_REG_6__SCAN_IN), .ZN(n6334) );
  AOI21_X1 U7346 ( .B1(n6363), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6362), 
        .ZN(n6333) );
  OAI211_X1 U7347 ( .C1(n6336), .C2(n6335), .A(n6334), .B(n6333), .ZN(n6337)
         );
  AOI221_X1 U7348 ( .B1(n6339), .B2(REIP_REG_6__SCAN_IN), .C1(n6338), .C2(
        n6669), .A(n6337), .ZN(n6343) );
  AOI22_X1 U7349 ( .A1(n6341), .A2(n3093), .B1(n6340), .B2(n3129), .ZN(n6342)
         );
  NAND2_X1 U7350 ( .A1(n6343), .A2(n6342), .ZN(U2821) );
  AOI21_X1 U7351 ( .B1(n6667), .B2(n6345), .A(n6344), .ZN(n6354) );
  OAI21_X1 U7352 ( .B1(n6348), .B2(n6347), .A(n6346), .ZN(n6349) );
  AOI21_X1 U7353 ( .B1(n6366), .B2(n6350), .A(n6349), .ZN(n6351) );
  OAI21_X1 U7354 ( .B1(n6352), .B2(n6370), .A(n6351), .ZN(n6353) );
  OAI21_X1 U7355 ( .B1(n6356), .B2(n5027), .A(n6355), .ZN(U2822) );
  AOI22_X1 U7356 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6358), .B1(
        REIP_REG_4__SCAN_IN), .B2(n6357), .ZN(n6376) );
  NOR3_X1 U7357 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6360), .A3(n6359), .ZN(n6361)
         );
  AOI211_X1 U7358 ( .C1(n6363), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6362), 
        .B(n6361), .ZN(n6375) );
  INV_X1 U7359 ( .A(n6364), .ZN(n6365) );
  AOI22_X1 U7360 ( .A1(n6368), .A2(n6367), .B1(n6366), .B2(n6365), .ZN(n6374)
         );
  OAI22_X1 U7361 ( .A1(n6371), .A2(n6370), .B1(n6369), .B2(n5027), .ZN(n6372)
         );
  INV_X1 U7362 ( .A(n6372), .ZN(n6373) );
  NAND4_X1 U7363 ( .A1(n6376), .A2(n6375), .A3(n6374), .A4(n6373), .ZN(U2823)
         );
  AOI22_X1 U7364 ( .A1(n6380), .A2(n6379), .B1(n6378), .B2(n6377), .ZN(n6381)
         );
  OAI21_X1 U7365 ( .B1(n6382), .B2(n5381), .A(n6381), .ZN(U2846) );
  INV_X1 U7366 ( .A(n6383), .ZN(n6386) );
  AOI22_X1 U7367 ( .A1(n6386), .A2(n6385), .B1(n6384), .B2(DATAI_16_), .ZN(
        n6390) );
  AOI22_X1 U7368 ( .A1(n6388), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6387), .ZN(n6389) );
  NAND2_X1 U7369 ( .A1(n6390), .A2(n6389), .ZN(U2875) );
  AOI22_X1 U7370 ( .A1(n6394), .A2(EAX_REG_28__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n6391) );
  OAI21_X1 U7371 ( .B1(n6834), .B2(n6735), .A(n6391), .ZN(U2895) );
  INV_X1 U7372 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n6914) );
  AOI22_X1 U7373 ( .A1(n6394), .A2(EAX_REG_25__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U7374 ( .B1(n6914), .B2(n6735), .A(n6392), .ZN(U2898) );
  INV_X1 U7375 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6812) );
  AOI22_X1 U7376 ( .A1(n6394), .A2(EAX_REG_20__SCAN_IN), .B1(n6411), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n6393) );
  OAI21_X1 U7377 ( .B1(n6812), .B2(n6419), .A(n6393), .ZN(U2903) );
  INV_X1 U7378 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n7042) );
  AOI22_X1 U7379 ( .A1(n6394), .A2(EAX_REG_18__SCAN_IN), .B1(n6411), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n6395) );
  OAI21_X1 U7380 ( .B1(n7042), .B2(n6419), .A(n6395), .ZN(U2905) );
  INV_X1 U7381 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6946) );
  AOI22_X1 U7382 ( .A1(n6411), .A2(LWORD_REG_15__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6396) );
  OAI21_X1 U7383 ( .B1(n6946), .B2(n6418), .A(n6396), .ZN(U2908) );
  INV_X1 U7384 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6878) );
  AOI22_X1 U7385 ( .A1(n6411), .A2(LWORD_REG_14__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6397) );
  OAI21_X1 U7386 ( .B1(n6878), .B2(n6418), .A(n6397), .ZN(U2909) );
  INV_X1 U7387 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6399) );
  AOI22_X1 U7388 ( .A1(n6411), .A2(LWORD_REG_13__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6398) );
  OAI21_X1 U7389 ( .B1(n6399), .B2(n6418), .A(n6398), .ZN(U2910) );
  INV_X1 U7390 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6457) );
  AOI22_X1 U7391 ( .A1(n6411), .A2(LWORD_REG_12__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6400) );
  OAI21_X1 U7392 ( .B1(n6457), .B2(n6418), .A(n6400), .ZN(U2911) );
  INV_X1 U7393 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6402) );
  AOI22_X1 U7394 ( .A1(n6411), .A2(LWORD_REG_11__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6401) );
  OAI21_X1 U7395 ( .B1(n6402), .B2(n6418), .A(n6401), .ZN(U2912) );
  INV_X1 U7396 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6453) );
  AOI22_X1 U7397 ( .A1(n6411), .A2(LWORD_REG_10__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6403) );
  OAI21_X1 U7398 ( .B1(n6453), .B2(n6418), .A(n6403), .ZN(U2913) );
  AOI22_X1 U7399 ( .A1(n6411), .A2(LWORD_REG_9__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6404) );
  OAI21_X1 U7400 ( .B1(n3789), .B2(n6418), .A(n6404), .ZN(U2914) );
  INV_X1 U7401 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6956) );
  INV_X1 U7402 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n6405) );
  OAI222_X1 U7403 ( .A1(n6419), .A2(n6956), .B1(n6418), .B2(n6849), .C1(n6735), 
        .C2(n6405), .ZN(U2915) );
  INV_X1 U7404 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n6875) );
  INV_X1 U7405 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6931) );
  OAI222_X1 U7406 ( .A1(n6419), .A2(n6875), .B1(n6418), .B2(n6896), .C1(n6735), 
        .C2(n6931), .ZN(U2916) );
  AOI22_X1 U7407 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6411), .B1(n6413), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6406) );
  OAI21_X1 U7408 ( .B1(n6407), .B2(n6418), .A(n6406), .ZN(U2917) );
  AOI22_X1 U7409 ( .A1(n6411), .A2(LWORD_REG_5__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6408) );
  OAI21_X1 U7410 ( .B1(n6978), .B2(n6418), .A(n6408), .ZN(U2918) );
  AOI22_X1 U7411 ( .A1(n6411), .A2(LWORD_REG_4__SCAN_IN), .B1(n6413), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6409) );
  OAI21_X1 U7412 ( .B1(n6912), .B2(n6418), .A(n6409), .ZN(U2919) );
  INV_X1 U7413 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n6926) );
  INV_X1 U7414 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n7011) );
  OAI222_X1 U7415 ( .A1(n6419), .A2(n6926), .B1(n6418), .B2(n6410), .C1(n6735), 
        .C2(n7011), .ZN(U2920) );
  INV_X1 U7416 ( .A(n6418), .ZN(n6414) );
  AOI222_X1 U7417 ( .A1(n6413), .A2(DATAO_REG_2__SCAN_IN), .B1(n6414), .B2(
        EAX_REG_2__SCAN_IN), .C1(n6411), .C2(LWORD_REG_2__SCAN_IN), .ZN(n6412)
         );
  INV_X1 U7418 ( .A(n6412), .ZN(U2921) );
  INV_X1 U7419 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6847) );
  AOI22_X1 U7420 ( .A1(EAX_REG_1__SCAN_IN), .A2(n6414), .B1(n6413), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6415) );
  OAI21_X1 U7421 ( .B1(n6847), .B2(n6735), .A(n6415), .ZN(U2922) );
  INV_X1 U7422 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n6962) );
  INV_X1 U7423 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6416) );
  OAI222_X1 U7424 ( .A1(n6419), .A2(n6962), .B1(n6418), .B2(n6417), .C1(n6735), 
        .C2(n6416), .ZN(U2923) );
  AOI22_X1 U7425 ( .A1(n7062), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n7061), .ZN(n6421) );
  OAI21_X1 U7426 ( .B1(n7065), .B2(n6436), .A(n6421), .ZN(U2924) );
  AOI22_X1 U7427 ( .A1(n7062), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n7061), .ZN(n6422) );
  OAI21_X1 U7428 ( .B1(n7065), .B2(n6438), .A(n6422), .ZN(U2925) );
  AOI22_X1 U7429 ( .A1(n7062), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n7061), .ZN(n6423) );
  OAI21_X1 U7430 ( .B1(n7065), .B2(n6440), .A(n6423), .ZN(U2926) );
  AOI22_X1 U7431 ( .A1(n7062), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n7061), .ZN(n6424) );
  OAI21_X1 U7432 ( .B1(n7065), .B2(n6442), .A(n6424), .ZN(U2927) );
  AOI22_X1 U7433 ( .A1(n7062), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n7061), .ZN(n6425) );
  OAI21_X1 U7434 ( .B1(n7065), .B2(n6444), .A(n6425), .ZN(U2928) );
  AOI22_X1 U7435 ( .A1(n7062), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n7061), .ZN(n6426) );
  OAI21_X1 U7436 ( .B1(n7065), .B2(n6446), .A(n6426), .ZN(U2929) );
  AOI22_X1 U7437 ( .A1(n7062), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n7061), .ZN(n6427) );
  OAI21_X1 U7438 ( .B1(n7065), .B2(n7064), .A(n6427), .ZN(U2930) );
  AOI22_X1 U7439 ( .A1(n7062), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n7061), .ZN(n6428) );
  OAI21_X1 U7440 ( .B1(n7065), .B2(n6448), .A(n6428), .ZN(U2931) );
  AOI22_X1 U7441 ( .A1(n7062), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n7061), .ZN(n6429) );
  OAI21_X1 U7442 ( .B1(n7065), .B2(n6943), .A(n6429), .ZN(U2932) );
  INV_X1 U7443 ( .A(DATAI_9_), .ZN(n7040) );
  AOI22_X1 U7444 ( .A1(n7062), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n7061), .ZN(n6430) );
  OAI21_X1 U7445 ( .B1(n7065), .B2(n7040), .A(n6430), .ZN(U2933) );
  INV_X1 U7446 ( .A(DATAI_11_), .ZN(n6929) );
  AOI22_X1 U7447 ( .A1(n7062), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n7061), .ZN(n6431) );
  OAI21_X1 U7448 ( .B1(n7065), .B2(n6929), .A(n6431), .ZN(U2935) );
  INV_X1 U7449 ( .A(DATAI_13_), .ZN(n6796) );
  AOI22_X1 U7450 ( .A1(n7062), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n7061), .ZN(n6432) );
  OAI21_X1 U7451 ( .B1(n7065), .B2(n6796), .A(n6432), .ZN(U2937) );
  INV_X1 U7452 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6803) );
  INV_X1 U7453 ( .A(DATAI_14_), .ZN(n6433) );
  NOR2_X1 U7454 ( .A1(n7065), .A2(n6433), .ZN(n6459) );
  AOI21_X1 U7455 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6462), .A(n6459), .ZN(
        n6434) );
  OAI21_X1 U7456 ( .B1(n6803), .B2(n6464), .A(n6434), .ZN(U2938) );
  AOI22_X1 U7457 ( .A1(n7062), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n7061), .ZN(n6435) );
  OAI21_X1 U7458 ( .B1(n7065), .B2(n6436), .A(n6435), .ZN(U2939) );
  AOI22_X1 U7459 ( .A1(n7062), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n7061), .ZN(n6437) );
  OAI21_X1 U7460 ( .B1(n7065), .B2(n6438), .A(n6437), .ZN(U2940) );
  AOI22_X1 U7461 ( .A1(n7062), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n7061), .ZN(n6439) );
  OAI21_X1 U7462 ( .B1(n7065), .B2(n6440), .A(n6439), .ZN(U2941) );
  AOI22_X1 U7463 ( .A1(n7062), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n7061), .ZN(n6441) );
  OAI21_X1 U7464 ( .B1(n7065), .B2(n6442), .A(n6441), .ZN(U2942) );
  AOI22_X1 U7465 ( .A1(n7062), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n7061), .ZN(n6443) );
  OAI21_X1 U7466 ( .B1(n7065), .B2(n6444), .A(n6443), .ZN(U2943) );
  AOI22_X1 U7467 ( .A1(n7062), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n7061), .ZN(n6445) );
  OAI21_X1 U7468 ( .B1(n7065), .B2(n6446), .A(n6445), .ZN(U2944) );
  AOI22_X1 U7469 ( .A1(n7062), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n7061), .ZN(n6447) );
  OAI21_X1 U7470 ( .B1(n7065), .B2(n6448), .A(n6447), .ZN(U2946) );
  AOI22_X1 U7471 ( .A1(n7062), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n7061), .ZN(n6449) );
  OAI21_X1 U7472 ( .B1(n7065), .B2(n6943), .A(n6449), .ZN(U2947) );
  AOI22_X1 U7473 ( .A1(n7062), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n7061), .ZN(n6450) );
  OAI21_X1 U7474 ( .B1(n7065), .B2(n7040), .A(n6450), .ZN(U2948) );
  AOI21_X1 U7475 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6462), .A(n6451), .ZN(
        n6452) );
  OAI21_X1 U7476 ( .B1(n6453), .B2(n6464), .A(n6452), .ZN(U2949) );
  AOI22_X1 U7477 ( .A1(n6462), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n7061), .ZN(n6454) );
  OAI21_X1 U7478 ( .B1(n7065), .B2(n6929), .A(n6454), .ZN(U2950) );
  AOI21_X1 U7479 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n7062), .A(n6455), .ZN(
        n6456) );
  OAI21_X1 U7480 ( .B1(n6457), .B2(n6464), .A(n6456), .ZN(U2951) );
  AOI22_X1 U7481 ( .A1(n6462), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n7061), .ZN(n6458) );
  OAI21_X1 U7482 ( .B1(n7065), .B2(n6796), .A(n6458), .ZN(U2952) );
  AOI21_X1 U7483 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6462), .A(n6459), .ZN(
        n6460) );
  OAI21_X1 U7484 ( .B1(n6878), .B2(n6464), .A(n6460), .ZN(U2953) );
  INV_X1 U7485 ( .A(n7065), .ZN(n6461) );
  AOI22_X1 U7486 ( .A1(n6462), .A2(LWORD_REG_15__SCAN_IN), .B1(n6461), .B2(
        DATAI_15_), .ZN(n6463) );
  OAI21_X1 U7487 ( .B1(n6946), .B2(n6464), .A(n6463), .ZN(U2954) );
  AOI22_X1 U7488 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6465), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6476) );
  INV_X1 U7489 ( .A(n6467), .ZN(n6469) );
  NAND2_X1 U7490 ( .A1(n6469), .A2(n6468), .ZN(n6471) );
  XNOR2_X1 U7491 ( .A(n6471), .B(n6470), .ZN(n6503) );
  AOI22_X1 U7492 ( .A1(n6474), .A2(n6503), .B1(n6473), .B2(n6472), .ZN(n6475)
         );
  OAI211_X1 U7493 ( .C1(n6478), .C2(n6477), .A(n6476), .B(n6475), .ZN(U2984)
         );
  INV_X1 U7494 ( .A(n6479), .ZN(n6481) );
  AOI21_X1 U7495 ( .B1(n6481), .B2(n6518), .A(n6480), .ZN(n6485) );
  AOI22_X1 U7496 ( .A1(n6502), .A2(n6483), .B1(n6486), .B2(n6482), .ZN(n6484)
         );
  OAI211_X1 U7497 ( .C1(n6487), .C2(n6486), .A(n6485), .B(n6484), .ZN(U3007)
         );
  AOI21_X1 U7498 ( .B1(n6489), .B2(n6518), .A(n6488), .ZN(n6493) );
  AOI22_X1 U7499 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n6491), .B1(n6490), 
        .B2(n6502), .ZN(n6492) );
  OAI211_X1 U7500 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6494), .A(n6493), 
        .B(n6492), .ZN(U3009) );
  NAND2_X1 U7501 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6495), .ZN(n6510)
         );
  NAND3_X1 U7502 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n6497), .A3(n6496), 
        .ZN(n6506) );
  OAI22_X1 U7503 ( .A1(n6500), .A2(n6499), .B1(n6662), .B2(n6498), .ZN(n6501)
         );
  INV_X1 U7504 ( .A(n6501), .ZN(n6505) );
  NAND2_X1 U7505 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  AND4_X1 U7506 ( .A1(n6507), .A2(n6506), .A3(n6505), .A4(n6504), .ZN(n6508)
         );
  OAI221_X1 U7507 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6510), .C1(n4146), .C2(n6509), .A(n6508), .ZN(U3016) );
  NAND2_X1 U7508 ( .A1(n6512), .A2(n6511), .ZN(n6517) );
  NOR3_X1 U7509 ( .A1(n6515), .A2(n6514), .A3(n6513), .ZN(n6516) );
  AOI211_X1 U7510 ( .C1(n6519), .C2(n6518), .A(n6517), .B(n6516), .ZN(n6520)
         );
  OAI221_X1 U7511 ( .B1(n6523), .B2(n6522), .C1(n6523), .C2(n6521), .A(n6520), 
        .ZN(U3018) );
  NOR2_X1 U7512 ( .A1(n7008), .A2(n6524), .ZN(U3019) );
  NAND3_X1 U7513 ( .A1(n6526), .A2(n6525), .A3(n6535), .ZN(n6527) );
  OAI21_X1 U7514 ( .B1(n6529), .B2(n6528), .A(n6527), .ZN(n6569) );
  NOR2_X1 U7515 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6530), .ZN(n6567)
         );
  AOI22_X1 U7516 ( .A1(n6532), .A2(n6569), .B1(n6531), .B2(n6567), .ZN(n6541)
         );
  NOR3_X1 U7517 ( .A1(n6534), .A2(n6570), .A3(n6533), .ZN(n6538) );
  OAI21_X1 U7518 ( .B1(n6864), .B2(n6567), .A(n6535), .ZN(n6536) );
  AOI22_X1 U7519 ( .A1(n6572), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6539), 
        .B2(n6570), .ZN(n6540) );
  OAI211_X1 U7520 ( .C1(n6542), .C2(n6602), .A(n6541), .B(n6540), .ZN(U3068)
         );
  AOI22_X1 U7521 ( .A1(n6578), .A2(n6569), .B1(n6543), .B2(n6567), .ZN(n6546)
         );
  AOI22_X1 U7522 ( .A1(n6572), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6544), 
        .B2(n6570), .ZN(n6545) );
  OAI211_X1 U7523 ( .C1(n6576), .C2(n6602), .A(n6546), .B(n6545), .ZN(U3069)
         );
  AOI22_X1 U7524 ( .A1(n6606), .A2(n6569), .B1(n6547), .B2(n6567), .ZN(n6550)
         );
  AOI22_X1 U7525 ( .A1(n6572), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6548), 
        .B2(n6570), .ZN(n6549) );
  OAI211_X1 U7526 ( .C1(n6604), .C2(n6602), .A(n6550), .B(n6549), .ZN(U3070)
         );
  AOI22_X1 U7527 ( .A1(n6613), .A2(n6569), .B1(n6551), .B2(n6567), .ZN(n6554)
         );
  AOI22_X1 U7528 ( .A1(n6572), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6552), 
        .B2(n6570), .ZN(n6553) );
  OAI211_X1 U7529 ( .C1(n6611), .C2(n6602), .A(n6554), .B(n6553), .ZN(U3071)
         );
  AOI22_X1 U7530 ( .A1(n6620), .A2(n6569), .B1(n6555), .B2(n6567), .ZN(n6558)
         );
  AOI22_X1 U7531 ( .A1(n6572), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6556), 
        .B2(n6570), .ZN(n6557) );
  OAI211_X1 U7532 ( .C1(n6618), .C2(n6602), .A(n6558), .B(n6557), .ZN(U3072)
         );
  AOI22_X1 U7533 ( .A1(n6591), .A2(n6569), .B1(n6559), .B2(n6567), .ZN(n6562)
         );
  AOI22_X1 U7534 ( .A1(n6572), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6560), 
        .B2(n6570), .ZN(n6561) );
  OAI211_X1 U7535 ( .C1(n6589), .C2(n6602), .A(n6562), .B(n6561), .ZN(U3073)
         );
  AOI22_X1 U7536 ( .A1(n6627), .A2(n6569), .B1(n6563), .B2(n6567), .ZN(n6566)
         );
  AOI22_X1 U7537 ( .A1(n6572), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6564), 
        .B2(n6570), .ZN(n6565) );
  OAI211_X1 U7538 ( .C1(n6625), .C2(n6602), .A(n6566), .B(n6565), .ZN(U3074)
         );
  AOI22_X1 U7539 ( .A1(n6636), .A2(n6569), .B1(n6568), .B2(n6567), .ZN(n6574)
         );
  AOI22_X1 U7540 ( .A1(n6572), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6571), 
        .B2(n6570), .ZN(n6573) );
  OAI211_X1 U7541 ( .C1(n6633), .C2(n6602), .A(n6574), .B(n6573), .ZN(U3075)
         );
  OAI22_X1 U7542 ( .A1(n6596), .A2(n6576), .B1(n6595), .B2(n6575), .ZN(n6577)
         );
  INV_X1 U7543 ( .A(n6577), .ZN(n6580) );
  AOI22_X1 U7544 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6599), .B1(n6598), 
        .B2(n6578), .ZN(n6579) );
  OAI211_X1 U7545 ( .C1(n6581), .C2(n6602), .A(n6580), .B(n6579), .ZN(U3077)
         );
  OAI22_X1 U7546 ( .A1(n6596), .A2(n6604), .B1(n6595), .B2(n6603), .ZN(n6582)
         );
  INV_X1 U7547 ( .A(n6582), .ZN(n6584) );
  AOI22_X1 U7548 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6599), .B1(n6598), 
        .B2(n6606), .ZN(n6583) );
  OAI211_X1 U7549 ( .C1(n6609), .C2(n6602), .A(n6584), .B(n6583), .ZN(U3078)
         );
  OAI22_X1 U7550 ( .A1(n6596), .A2(n6618), .B1(n6595), .B2(n6617), .ZN(n6585)
         );
  INV_X1 U7551 ( .A(n6585), .ZN(n6587) );
  AOI22_X1 U7552 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6599), .B1(n6598), 
        .B2(n6620), .ZN(n6586) );
  OAI211_X1 U7553 ( .C1(n6623), .C2(n6602), .A(n6587), .B(n6586), .ZN(U3080)
         );
  OAI22_X1 U7554 ( .A1(n6596), .A2(n6589), .B1(n6595), .B2(n6588), .ZN(n6590)
         );
  INV_X1 U7555 ( .A(n6590), .ZN(n6593) );
  AOI22_X1 U7556 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6599), .B1(n6598), 
        .B2(n6591), .ZN(n6592) );
  OAI211_X1 U7557 ( .C1(n6594), .C2(n6602), .A(n6593), .B(n6592), .ZN(U3081)
         );
  OAI22_X1 U7558 ( .A1(n6596), .A2(n6625), .B1(n6595), .B2(n6624), .ZN(n6597)
         );
  INV_X1 U7559 ( .A(n6597), .ZN(n6601) );
  AOI22_X1 U7560 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6599), .B1(n6598), 
        .B2(n6627), .ZN(n6600) );
  OAI211_X1 U7561 ( .C1(n6630), .C2(n6602), .A(n6601), .B(n6600), .ZN(U3082)
         );
  OAI22_X1 U7562 ( .A1(n6634), .A2(n6604), .B1(n6603), .B2(n6631), .ZN(n6605)
         );
  INV_X1 U7563 ( .A(n6605), .ZN(n6608) );
  AOI22_X1 U7564 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6638), .B1(n6637), 
        .B2(n6606), .ZN(n6607) );
  OAI211_X1 U7565 ( .C1(n6609), .C2(n6641), .A(n6608), .B(n6607), .ZN(U3110)
         );
  OAI22_X1 U7566 ( .A1(n6634), .A2(n6611), .B1(n6610), .B2(n6631), .ZN(n6612)
         );
  INV_X1 U7567 ( .A(n6612), .ZN(n6615) );
  AOI22_X1 U7568 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6638), .B1(n6637), 
        .B2(n6613), .ZN(n6614) );
  OAI211_X1 U7569 ( .C1(n6616), .C2(n6641), .A(n6615), .B(n6614), .ZN(U3111)
         );
  OAI22_X1 U7570 ( .A1(n6634), .A2(n6618), .B1(n6617), .B2(n6631), .ZN(n6619)
         );
  INV_X1 U7571 ( .A(n6619), .ZN(n6622) );
  AOI22_X1 U7572 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6638), .B1(n6637), 
        .B2(n6620), .ZN(n6621) );
  OAI211_X1 U7573 ( .C1(n6623), .C2(n6641), .A(n6622), .B(n6621), .ZN(U3112)
         );
  OAI22_X1 U7574 ( .A1(n6634), .A2(n6625), .B1(n6624), .B2(n6631), .ZN(n6626)
         );
  INV_X1 U7575 ( .A(n6626), .ZN(n6629) );
  AOI22_X1 U7576 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6638), .B1(n6637), 
        .B2(n6627), .ZN(n6628) );
  OAI211_X1 U7577 ( .C1(n6630), .C2(n6641), .A(n6629), .B(n6628), .ZN(U3114)
         );
  OAI22_X1 U7578 ( .A1(n6634), .A2(n6633), .B1(n6632), .B2(n6631), .ZN(n6635)
         );
  INV_X1 U7579 ( .A(n6635), .ZN(n6640) );
  AOI22_X1 U7580 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6638), .B1(n6637), 
        .B2(n6636), .ZN(n6639) );
  OAI211_X1 U7581 ( .C1(n6642), .C2(n6641), .A(n6640), .B(n6639), .ZN(U3115)
         );
  INV_X1 U7582 ( .A(n6643), .ZN(n6644) );
  OAI211_X1 U7583 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(n6644), .B(STATE2_REG_1__SCAN_IN), .ZN(n6653) );
  INV_X1 U7584 ( .A(n6645), .ZN(n6651) );
  OAI21_X1 U7585 ( .B1(n6647), .B2(READY_N), .A(n6646), .ZN(n6650) );
  INV_X1 U7586 ( .A(n6648), .ZN(n6649) );
  AOI21_X1 U7587 ( .B1(n6651), .B2(n6650), .A(n6649), .ZN(n6652) );
  NAND2_X1 U7588 ( .A1(n6653), .A2(n6652), .ZN(U3149) );
  INV_X1 U7589 ( .A(n6711), .ZN(n6654) );
  AND2_X1 U7590 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6654), .ZN(U3151) );
  AND2_X1 U7591 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6654), .ZN(U3152) );
  AND2_X1 U7592 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6654), .ZN(U3153) );
  INV_X1 U7593 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n7045) );
  NOR2_X1 U7594 ( .A1(n6711), .A2(n7045), .ZN(U3154) );
  INV_X1 U7595 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6993) );
  NOR2_X1 U7596 ( .A1(n6711), .A2(n6993), .ZN(U3155) );
  AND2_X1 U7597 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6654), .ZN(U3156) );
  AND2_X1 U7598 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6654), .ZN(U3157) );
  AND2_X1 U7599 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6654), .ZN(U3158) );
  AND2_X1 U7600 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6654), .ZN(U3159) );
  AND2_X1 U7601 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6654), .ZN(U3160) );
  NOR2_X1 U7602 ( .A1(n6711), .A2(n6964), .ZN(U3161) );
  AND2_X1 U7603 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6654), .ZN(U3162) );
  AND2_X1 U7604 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6654), .ZN(U3163) );
  AND2_X1 U7605 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6654), .ZN(U3164) );
  AND2_X1 U7606 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6654), .ZN(U3165) );
  AND2_X1 U7607 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6654), .ZN(U3166) );
  AND2_X1 U7608 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6654), .ZN(U3167) );
  AND2_X1 U7609 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6654), .ZN(U3168) );
  INV_X1 U7610 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6800) );
  NOR2_X1 U7611 ( .A1(n6711), .A2(n6800), .ZN(U3169) );
  AND2_X1 U7612 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6654), .ZN(U3170) );
  AND2_X1 U7613 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6654), .ZN(U3171) );
  AND2_X1 U7614 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6654), .ZN(U3172) );
  INV_X1 U7615 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6819) );
  NOR2_X1 U7616 ( .A1(n6711), .A2(n6819), .ZN(U3173) );
  AND2_X1 U7617 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6654), .ZN(U3174) );
  AND2_X1 U7618 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6654), .ZN(U3175) );
  NOR2_X1 U7619 ( .A1(n6711), .A2(n6934), .ZN(U3176) );
  INV_X1 U7620 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6894) );
  NOR2_X1 U7621 ( .A1(n6711), .A2(n6894), .ZN(U3177) );
  AND2_X1 U7622 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6654), .ZN(U3178) );
  AND2_X1 U7623 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6654), .ZN(U3179) );
  AND2_X1 U7624 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6654), .ZN(U3180) );
  AOI221_X1 U7625 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6868), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6655) );
  AOI221_X1 U7626 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6655), .C2(HOLD), .A(n4106), .ZN(n6660) );
  NAND3_X1 U7627 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .A3(
        STATE_REG_2__SCAN_IN), .ZN(n6658) );
  NAND4_X1 U7628 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .A3(n6656), .A4(n6815), .ZN(n6657) );
  OAI211_X1 U7629 ( .C1(n6660), .C2(n6659), .A(n6658), .B(n6657), .ZN(U3183)
         );
  NAND2_X1 U7630 ( .A1(n6746), .A2(n6992), .ZN(n6706) );
  NOR2_X2 U7631 ( .A1(n6992), .A2(n6734), .ZN(n6704) );
  AOI22_X1 U7632 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6734), .ZN(n6661) );
  OAI21_X1 U7633 ( .B1(n6662), .B2(n6706), .A(n6661), .ZN(U3184) );
  AOI22_X1 U7634 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6734), .ZN(n6663) );
  OAI21_X1 U7635 ( .B1(n6884), .B2(n6706), .A(n6663), .ZN(U3185) );
  AOI22_X1 U7636 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6734), .ZN(n6664) );
  OAI21_X1 U7637 ( .B1(n6665), .B2(n6706), .A(n6664), .ZN(U3186) );
  AOI22_X1 U7638 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6734), .ZN(n6666) );
  OAI21_X1 U7639 ( .B1(n6667), .B2(n6706), .A(n6666), .ZN(U3187) );
  AOI22_X1 U7640 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6734), .ZN(n6668) );
  OAI21_X1 U7641 ( .B1(n6669), .B2(n6706), .A(n6668), .ZN(U3188) );
  AOI22_X1 U7642 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6734), .ZN(n6670) );
  OAI21_X1 U7643 ( .B1(n6672), .B2(n6706), .A(n6670), .ZN(U3189) );
  INV_X1 U7644 ( .A(n6704), .ZN(n6702) );
  INV_X1 U7645 ( .A(n6706), .ZN(n6700) );
  AOI22_X1 U7646 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6734), .ZN(n6671) );
  OAI21_X1 U7647 ( .B1(n6672), .B2(n6702), .A(n6671), .ZN(U3190) );
  AOI22_X1 U7648 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6734), .ZN(n6673) );
  OAI21_X1 U7649 ( .B1(n6675), .B2(n6706), .A(n6673), .ZN(U3191) );
  AOI22_X1 U7650 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6734), .ZN(n6674) );
  OAI21_X1 U7651 ( .B1(n6675), .B2(n6702), .A(n6674), .ZN(U3192) );
  AOI22_X1 U7652 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6734), .ZN(n6676) );
  OAI21_X1 U7653 ( .B1(n6677), .B2(n6702), .A(n6676), .ZN(U3193) );
  AOI22_X1 U7654 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6734), .ZN(n6678) );
  OAI21_X1 U7655 ( .B1(n6679), .B2(n6706), .A(n6678), .ZN(U3194) );
  AOI22_X1 U7656 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6734), .ZN(n6680) );
  OAI21_X1 U7657 ( .B1(n6971), .B2(n6706), .A(n6680), .ZN(U3195) );
  AOI22_X1 U7658 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6734), .ZN(n6681) );
  OAI21_X1 U7659 ( .B1(n6971), .B2(n6702), .A(n6681), .ZN(U3196) );
  AOI22_X1 U7660 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6734), .ZN(n6682) );
  OAI21_X1 U7661 ( .B1(n7023), .B2(n6706), .A(n6682), .ZN(U3197) );
  INV_X1 U7662 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6972) );
  OAI222_X1 U7663 ( .A1(n6702), .A2(n7023), .B1(n6972), .B2(n6746), .C1(n6998), 
        .C2(n6706), .ZN(U3198) );
  AOI22_X1 U7664 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6734), .ZN(n6683) );
  OAI21_X1 U7665 ( .B1(n6998), .B2(n6702), .A(n6683), .ZN(U3199) );
  AOI22_X1 U7666 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6734), .ZN(n6684) );
  OAI21_X1 U7667 ( .B1(n6685), .B2(n6706), .A(n6684), .ZN(U3200) );
  AOI22_X1 U7668 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6734), .ZN(n6686) );
  OAI21_X1 U7669 ( .B1(n6688), .B2(n6706), .A(n6686), .ZN(U3201) );
  INV_X1 U7670 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6828) );
  INV_X1 U7671 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6687) );
  OAI222_X1 U7672 ( .A1(n6702), .A2(n6688), .B1(n6828), .B2(n6746), .C1(n6687), 
        .C2(n6706), .ZN(U3202) );
  AOI22_X1 U7673 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6734), .ZN(n6689) );
  OAI21_X1 U7674 ( .B1(n6691), .B2(n6706), .A(n6689), .ZN(U3203) );
  AOI22_X1 U7675 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6734), .ZN(n6690) );
  OAI21_X1 U7676 ( .B1(n6691), .B2(n6702), .A(n6690), .ZN(U3204) );
  AOI22_X1 U7677 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6734), .ZN(n6692) );
  OAI21_X1 U7678 ( .B1(n7043), .B2(n6702), .A(n6692), .ZN(U3205) );
  INV_X1 U7679 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6694) );
  AOI22_X1 U7680 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6734), .ZN(n6693) );
  OAI21_X1 U7681 ( .B1(n6694), .B2(n6706), .A(n6693), .ZN(U3206) );
  INV_X1 U7682 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6977) );
  AOI22_X1 U7683 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6734), .ZN(n6695) );
  OAI21_X1 U7684 ( .B1(n6977), .B2(n6706), .A(n6695), .ZN(U3207) );
  AOI22_X1 U7685 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6734), .ZN(n6696) );
  OAI21_X1 U7686 ( .B1(n6977), .B2(n6702), .A(n6696), .ZN(U3208) );
  INV_X1 U7687 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6945) );
  AOI22_X1 U7688 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6734), .ZN(n6697) );
  OAI21_X1 U7689 ( .B1(n6945), .B2(n6706), .A(n6697), .ZN(U3209) );
  AOI22_X1 U7690 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6734), .ZN(n6698) );
  OAI21_X1 U7691 ( .B1(n6945), .B2(n6702), .A(n6698), .ZN(U3210) );
  AOI22_X1 U7692 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6734), .ZN(n6699) );
  OAI21_X1 U7693 ( .B1(n7046), .B2(n6702), .A(n6699), .ZN(U3211) );
  AOI22_X1 U7694 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6734), .ZN(n6701) );
  OAI21_X1 U7695 ( .B1(n6703), .B2(n6702), .A(n6701), .ZN(U3212) );
  AOI22_X1 U7696 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6734), .ZN(n6705) );
  OAI21_X1 U7697 ( .B1(n6707), .B2(n6706), .A(n6705), .ZN(U3213) );
  MUX2_X1 U7698 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6746), .Z(U3445) );
  MUX2_X1 U7699 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6746), .Z(U3446) );
  MUX2_X1 U7700 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6746), .Z(U3447) );
  INV_X1 U7701 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6730) );
  INV_X1 U7702 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U7703 ( .A1(n6746), .A2(n6730), .B1(n6838), .B2(n6734), .ZN(U3448)
         );
  OAI21_X1 U7704 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6711), .A(n6709), .ZN(
        n6708) );
  INV_X1 U7705 ( .A(n6708), .ZN(U3451) );
  INV_X1 U7706 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6710) );
  OAI21_X1 U7707 ( .B1(n6711), .B2(n6710), .A(n6709), .ZN(U3452) );
  OAI22_X1 U7708 ( .A1(n6714), .A2(n6722), .B1(n6713), .B2(n6712), .ZN(n6716)
         );
  MUX2_X1 U7709 ( .A(n6716), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6715), 
        .Z(U3456) );
  OAI22_X1 U7710 ( .A1(n6717), .A2(n6722), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n4599), .ZN(n6719) );
  OAI22_X1 U7711 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6720), .B1(n6719), .B2(n6718), .ZN(n6721) );
  OAI21_X1 U7712 ( .B1(n6723), .B2(n6722), .A(n6721), .ZN(U3461) );
  INV_X1 U7713 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6725) );
  NOR3_X1 U7714 ( .A1(n6725), .A2(REIP_REG_0__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6724) );
  AOI221_X1 U7715 ( .B1(n6726), .B2(n6725), .C1(REIP_REG_1__SCAN_IN), .C2(
        REIP_REG_0__SCAN_IN), .A(n6724), .ZN(n6728) );
  INV_X1 U7716 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6727) );
  INV_X1 U7717 ( .A(n6732), .ZN(n6729) );
  AOI22_X1 U7718 ( .A1(n6732), .A2(n6728), .B1(n6727), .B2(n6729), .ZN(U3468)
         );
  NOR2_X1 U7719 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6731) );
  AOI22_X1 U7720 ( .A1(n6732), .A2(n6731), .B1(n6730), .B2(n6729), .ZN(U3469)
         );
  NAND2_X1 U7721 ( .A1(n6734), .A2(W_R_N_REG_SCAN_IN), .ZN(n6733) );
  OAI21_X1 U7722 ( .B1(n6734), .B2(READREQUEST_REG_SCAN_IN), .A(n6733), .ZN(
        U3470) );
  NOR2_X1 U7723 ( .A1(n6735), .A2(READY_N), .ZN(n6737) );
  NOR3_X1 U7724 ( .A1(n6738), .A2(n6737), .A3(n6736), .ZN(n6745) );
  OAI211_X1 U7725 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6740), .A(n6739), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6742) );
  AOI21_X1 U7726 ( .B1(n6742), .B2(STATE2_REG_0__SCAN_IN), .A(n6741), .ZN(
        n6744) );
  NAND2_X1 U7727 ( .A1(n6745), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6743) );
  OAI21_X1 U7728 ( .B1(n6745), .B2(n6744), .A(n6743), .ZN(U3472) );
  MUX2_X1 U7729 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6746), .Z(U3473) );
  NAND4_X1 U7730 ( .A1(EAX_REG_15__SCAN_IN), .A2(DATAI_11_), .A3(
        DATAO_REG_3__SCAN_IN), .A4(n6928), .ZN(n6778) );
  NAND4_X1 U7731 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(DATAI_8_), .A3(
        DATAI_23_), .A4(n6948), .ZN(n6777) );
  INV_X1 U7732 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6965) );
  NOR4_X1 U7733 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        DATAO_REG_0__SCAN_IN), .A3(n6965), .A4(n6964), .ZN(n6753) );
  NOR4_X1 U7734 ( .A1(REIP_REG_25__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .A3(DATAO_REG_8__SCAN_IN), .A4(n6958), 
        .ZN(n6752) );
  NAND4_X1 U7735 ( .A1(EAX_REG_5__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        ADDRESS_REG_14__SCAN_IN), .A4(n6981), .ZN(n6750) );
  NAND4_X1 U7736 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        LWORD_REG_7__SCAN_IN), .A3(n6934), .A4(n6932), .ZN(n6749) );
  INV_X1 U7737 ( .A(DATAI_22_), .ZN(n6805) );
  NAND4_X1 U7738 ( .A1(DATAI_30_), .A2(DATAWIDTH_REG_9__SCAN_IN), .A3(NA_N), 
        .A4(n6805), .ZN(n6748) );
  NAND4_X1 U7739 ( .A1(EAX_REG_30__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .A3(
        DATAWIDTH_REG_13__SCAN_IN), .A4(n6796), .ZN(n6747) );
  NOR4_X1 U7740 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n6751)
         );
  NAND3_X1 U7741 ( .A1(n6753), .A2(n6752), .A3(n6751), .ZN(n6776) );
  NAND4_X1 U7742 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        EBX_REG_21__SCAN_IN), .A3(PHYADDRPOINTER_REG_20__SCAN_IN), .A4(
        UWORD_REG_10__SCAN_IN), .ZN(n6757) );
  NAND4_X1 U7743 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n6850), .A3(n7064), 
        .A4(n7011), .ZN(n6756) );
  NAND4_X1 U7744 ( .A1(REIP_REG_22__SCAN_IN), .A2(DATAO_REG_18__SCAN_IN), .A3(
        n7023), .A4(n7025), .ZN(n6755) );
  NAND4_X1 U7745 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(DATAI_9_), .A3(
        n5055), .A4(n6998), .ZN(n6754) );
  NOR4_X1 U7746 ( .A1(n6757), .A2(n6756), .A3(n6755), .A4(n6754), .ZN(n6774)
         );
  INV_X1 U7747 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6980) );
  INV_X1 U7748 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6961) );
  INV_X1 U7749 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n7002) );
  NAND4_X1 U7750 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n6980), .A3(n6961), 
        .A4(n7002), .ZN(n6762) );
  INV_X1 U7751 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6761) );
  NAND4_X1 U7752 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(
        INSTQUEUE_REG_10__2__SCAN_IN), .A3(INSTQUEUE_REG_13__2__SCAN_IN), .A4(
        INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6759) );
  NAND4_X1 U7753 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(
        INSTQUEUE_REG_14__7__SCAN_IN), .A3(INSTQUEUE_REG_8__7__SCAN_IN), .A4(
        INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n6758) );
  OR4_X1 U7754 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(
        INSTQUEUE_REG_9__6__SCAN_IN), .A3(n6759), .A4(n6758), .ZN(n6760) );
  NOR4_X1 U7755 ( .A1(n6762), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .A3(n6761), 
        .A4(n6760), .ZN(n6773) );
  NAND4_X1 U7756 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(DATAI_29_), .A4(n6878), .ZN(n6766) );
  NAND4_X1 U7757 ( .A1(EBX_REG_12__SCAN_IN), .A2(DATAO_REG_31__SCAN_IN), .A3(
        DATAO_REG_7__SCAN_IN), .A4(n6879), .ZN(n6765) );
  NAND4_X1 U7758 ( .A1(EAX_REG_4__SCAN_IN), .A2(DATAO_REG_2__SCAN_IN), .A3(
        n5340), .A4(n6910), .ZN(n6764) );
  INV_X1 U7759 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6891) );
  INV_X1 U7760 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6906) );
  NAND4_X1 U7761 ( .A1(EAX_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(n6891), .A4(n6906), .ZN(n6763) );
  NOR4_X1 U7762 ( .A1(n6766), .A2(n6765), .A3(n6764), .A4(n6763), .ZN(n6772)
         );
  NAND4_X1 U7763 ( .A1(EBX_REG_26__SCAN_IN), .A2(EBX_REG_8__SCAN_IN), .A3(
        ADDRESS_REG_18__SCAN_IN), .A4(n6837), .ZN(n6770) );
  NAND4_X1 U7764 ( .A1(DATAO_REG_20__SCAN_IN), .A2(UWORD_REG_12__SCAN_IN), 
        .A3(n6835), .A4(n6838), .ZN(n6769) );
  INV_X1 U7765 ( .A(DATAI_19_), .ZN(n6861) );
  NAND4_X1 U7766 ( .A1(STATE2_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A3(DATAO_REG_26__SCAN_IN), .A4(
        n6861), .ZN(n6768) );
  NAND4_X1 U7767 ( .A1(EAX_REG_8__SCAN_IN), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n6846), .A4(n6847), .ZN(n6767) );
  NOR4_X1 U7768 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n6771)
         );
  NAND4_X1 U7769 ( .A1(n6774), .A2(n6773), .A3(n6772), .A4(n6771), .ZN(n6775)
         );
  NOR4_X1 U7770 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6794)
         );
  NOR4_X1 U7771 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(
        INSTQUEUE_REG_7__0__SCAN_IN), .A3(INSTQUEUE_REG_4__1__SCAN_IN), .A4(
        n5917), .ZN(n6792) );
  AND4_X1 U7772 ( .A1(n7046), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .A3(
        INSTQUEUE_REG_5__4__SCAN_IN), .A4(REIP_REG_27__SCAN_IN), .ZN(n6780) );
  NAND4_X1 U7773 ( .A1(n6780), .A2(n6779), .A3(UWORD_REG_9__SCAN_IN), .A4(
        STATE_REG_1__SCAN_IN), .ZN(n6786) );
  AND4_X1 U7774 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(
        INSTQUEUE_REG_1__5__SCAN_IN), .A3(INSTQUEUE_REG_11__1__SCAN_IN), .A4(
        n6868), .ZN(n6781) );
  INV_X1 U7775 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6991) );
  AND2_X1 U7776 ( .A1(n6781), .A2(n6991), .ZN(n6783) );
  NAND4_X1 U7777 ( .A1(n6784), .A2(STATE_REG_2__SCAN_IN), .A3(n6783), .A4(
        n6782), .ZN(n6785) );
  NOR2_X1 U7778 ( .A1(n6786), .A2(n6785), .ZN(n6790) );
  INV_X1 U7779 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6892) );
  INV_X1 U7780 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n7017) );
  NAND4_X1 U7781 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n7014), .A3(n6892), 
        .A4(n7017), .ZN(n6788) );
  INV_X1 U7782 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n7013) );
  INV_X1 U7783 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6885) );
  NAND4_X1 U7784 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6142), .A3(n7013), 
        .A4(n6885), .ZN(n6787) );
  NOR2_X1 U7785 ( .A1(n6788), .A2(n6787), .ZN(n6789) );
  AND4_X1 U7786 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n6793)
         );
  AOI21_X1 U7787 ( .B1(n6794), .B2(n6793), .A(keyinput124), .ZN(n7060) );
  AOI22_X1 U7788 ( .A1(n6797), .A2(keyinput65), .B1(keyinput17), .B2(n6796), 
        .ZN(n6795) );
  OAI221_X1 U7789 ( .B1(n6797), .B2(keyinput65), .C1(n6796), .C2(keyinput17), 
        .A(n6795), .ZN(n6810) );
  AOI22_X1 U7790 ( .A1(n6800), .A2(keyinput51), .B1(n6799), .B2(keyinput27), 
        .ZN(n6798) );
  OAI221_X1 U7791 ( .B1(n6800), .B2(keyinput51), .C1(n6799), .C2(keyinput27), 
        .A(n6798), .ZN(n6809) );
  INV_X1 U7792 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6802) );
  AOI22_X1 U7793 ( .A1(n6803), .A2(keyinput18), .B1(n6802), .B2(keyinput83), 
        .ZN(n6801) );
  OAI221_X1 U7794 ( .B1(n6803), .B2(keyinput18), .C1(n6802), .C2(keyinput83), 
        .A(n6801), .ZN(n6808) );
  INV_X1 U7795 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6806) );
  AOI22_X1 U7796 ( .A1(n6806), .A2(keyinput94), .B1(keyinput38), .B2(n6805), 
        .ZN(n6804) );
  OAI221_X1 U7797 ( .B1(n6806), .B2(keyinput94), .C1(n6805), .C2(keyinput38), 
        .A(n6804), .ZN(n6807) );
  NOR4_X1 U7798 ( .A1(n6810), .A2(n6809), .A3(n6808), .A4(n6807), .ZN(n6859)
         );
  INV_X1 U7799 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6813) );
  AOI22_X1 U7800 ( .A1(n6813), .A2(keyinput48), .B1(keyinput108), .B2(n6812), 
        .ZN(n6811) );
  OAI221_X1 U7801 ( .B1(n6813), .B2(keyinput48), .C1(n6812), .C2(keyinput108), 
        .A(n6811), .ZN(n6825) );
  AOI22_X1 U7802 ( .A1(n6816), .A2(keyinput7), .B1(keyinput99), .B2(n6815), 
        .ZN(n6814) );
  OAI221_X1 U7803 ( .B1(n6816), .B2(keyinput7), .C1(n6815), .C2(keyinput99), 
        .A(n6814), .ZN(n6824) );
  INV_X1 U7804 ( .A(DATAI_30_), .ZN(n6818) );
  AOI22_X1 U7805 ( .A1(n6819), .A2(keyinput62), .B1(n6818), .B2(keyinput110), 
        .ZN(n6817) );
  OAI221_X1 U7806 ( .B1(n6819), .B2(keyinput62), .C1(n6818), .C2(keyinput110), 
        .A(n6817), .ZN(n6823) );
  XNOR2_X1 U7807 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .B(keyinput116), .ZN(n6821) );
  XNOR2_X1 U7808 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .B(keyinput87), .ZN(n6820)
         );
  NAND2_X1 U7809 ( .A1(n6821), .A2(n6820), .ZN(n6822) );
  NOR4_X1 U7810 ( .A1(n6825), .A2(n6824), .A3(n6823), .A4(n6822), .ZN(n6858)
         );
  AOI22_X1 U7811 ( .A1(n6828), .A2(keyinput13), .B1(n6827), .B2(keyinput72), 
        .ZN(n6826) );
  OAI221_X1 U7812 ( .B1(n6828), .B2(keyinput13), .C1(n6827), .C2(keyinput72), 
        .A(n6826), .ZN(n6832) );
  XNOR2_X1 U7813 ( .A(n6829), .B(keyinput31), .ZN(n6831) );
  XOR2_X1 U7814 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .B(keyinput95), .Z(n6830)
         );
  OR3_X1 U7815 ( .A1(n6832), .A2(n6831), .A3(n6830), .ZN(n6841) );
  AOI22_X1 U7816 ( .A1(n6835), .A2(keyinput40), .B1(keyinput81), .B2(n6834), 
        .ZN(n6833) );
  OAI221_X1 U7817 ( .B1(n6835), .B2(keyinput40), .C1(n6834), .C2(keyinput81), 
        .A(n6833), .ZN(n6840) );
  AOI22_X1 U7818 ( .A1(n6838), .A2(keyinput22), .B1(n6837), .B2(keyinput77), 
        .ZN(n6836) );
  OAI221_X1 U7819 ( .B1(n6838), .B2(keyinput22), .C1(n6837), .C2(keyinput77), 
        .A(n6836), .ZN(n6839) );
  NOR3_X1 U7820 ( .A1(n6841), .A2(n6840), .A3(n6839), .ZN(n6857) );
  INV_X1 U7821 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6844) );
  AOI22_X1 U7822 ( .A1(n6844), .A2(keyinput52), .B1(keyinput26), .B2(n6843), 
        .ZN(n6842) );
  OAI221_X1 U7823 ( .B1(n6844), .B2(keyinput52), .C1(n6843), .C2(keyinput26), 
        .A(n6842), .ZN(n6855) );
  AOI22_X1 U7824 ( .A1(n6847), .A2(keyinput53), .B1(n6846), .B2(keyinput106), 
        .ZN(n6845) );
  OAI221_X1 U7825 ( .B1(n6847), .B2(keyinput53), .C1(n6846), .C2(keyinput106), 
        .A(n6845), .ZN(n6854) );
  AOI22_X1 U7826 ( .A1(n6850), .A2(keyinput10), .B1(keyinput97), .B2(n6849), 
        .ZN(n6848) );
  OAI221_X1 U7827 ( .B1(n6850), .B2(keyinput10), .C1(n6849), .C2(keyinput97), 
        .A(n6848), .ZN(n6853) );
  AOI22_X1 U7828 ( .A1(n4103), .A2(keyinput73), .B1(keyinput23), .B2(n4146), 
        .ZN(n6851) );
  OAI221_X1 U7829 ( .B1(n4103), .B2(keyinput73), .C1(n4146), .C2(keyinput23), 
        .A(n6851), .ZN(n6852) );
  NOR4_X1 U7830 ( .A1(n6855), .A2(n6854), .A3(n6853), .A4(n6852), .ZN(n6856)
         );
  NAND4_X1 U7831 ( .A1(n6859), .A2(n6858), .A3(n6857), .A4(n6856), .ZN(n7058)
         );
  AOI22_X1 U7832 ( .A1(n6862), .A2(keyinput111), .B1(n6861), .B2(keyinput29), 
        .ZN(n6860) );
  OAI221_X1 U7833 ( .B1(n6862), .B2(keyinput111), .C1(n6861), .C2(keyinput29), 
        .A(n6860), .ZN(n6873) );
  AOI22_X1 U7834 ( .A1(n6864), .A2(keyinput0), .B1(n5917), .B2(keyinput119), 
        .ZN(n6863) );
  OAI221_X1 U7835 ( .B1(n6864), .B2(keyinput0), .C1(n5917), .C2(keyinput119), 
        .A(n6863), .ZN(n6872) );
  AOI22_X1 U7836 ( .A1(n6866), .A2(keyinput91), .B1(n6761), .B2(keyinput12), 
        .ZN(n6865) );
  OAI221_X1 U7837 ( .B1(n6866), .B2(keyinput91), .C1(n6761), .C2(keyinput12), 
        .A(n6865), .ZN(n6871) );
  AOI22_X1 U7838 ( .A1(n6869), .A2(keyinput4), .B1(n6868), .B2(keyinput37), 
        .ZN(n6867) );
  OAI221_X1 U7839 ( .B1(n6869), .B2(keyinput4), .C1(n6868), .C2(keyinput37), 
        .A(n6867), .ZN(n6870) );
  NOR4_X1 U7840 ( .A1(n6873), .A2(n6872), .A3(n6871), .A4(n6870), .ZN(n6923)
         );
  AOI22_X1 U7841 ( .A1(n6876), .A2(keyinput21), .B1(keyinput47), .B2(n6875), 
        .ZN(n6874) );
  OAI221_X1 U7842 ( .B1(n6876), .B2(keyinput21), .C1(n6875), .C2(keyinput47), 
        .A(n6874), .ZN(n6889) );
  AOI22_X1 U7843 ( .A1(n6879), .A2(keyinput35), .B1(keyinput70), .B2(n6878), 
        .ZN(n6877) );
  OAI221_X1 U7844 ( .B1(n6879), .B2(keyinput35), .C1(n6878), .C2(keyinput70), 
        .A(n6877), .ZN(n6888) );
  INV_X1 U7845 ( .A(DATAI_29_), .ZN(n6881) );
  AOI22_X1 U7846 ( .A1(n6882), .A2(keyinput46), .B1(keyinput32), .B2(n6881), 
        .ZN(n6880) );
  OAI221_X1 U7847 ( .B1(n6882), .B2(keyinput46), .C1(n6881), .C2(keyinput32), 
        .A(n6880), .ZN(n6887) );
  AOI22_X1 U7848 ( .A1(n6885), .A2(keyinput2), .B1(keyinput58), .B2(n6884), 
        .ZN(n6883) );
  OAI221_X1 U7849 ( .B1(n6885), .B2(keyinput2), .C1(n6884), .C2(keyinput58), 
        .A(n6883), .ZN(n6886) );
  NOR4_X1 U7850 ( .A1(n6889), .A2(n6888), .A3(n6887), .A4(n6886), .ZN(n6922)
         );
  AOI22_X1 U7851 ( .A1(n6892), .A2(keyinput19), .B1(keyinput11), .B2(n6891), 
        .ZN(n6890) );
  OAI221_X1 U7852 ( .B1(n6892), .B2(keyinput19), .C1(n6891), .C2(keyinput11), 
        .A(n6890), .ZN(n6904) );
  INV_X1 U7853 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U7854 ( .A1(n6895), .A2(keyinput43), .B1(keyinput6), .B2(n6894), 
        .ZN(n6893) );
  OAI221_X1 U7855 ( .B1(n6895), .B2(keyinput43), .C1(n6894), .C2(keyinput6), 
        .A(n6893), .ZN(n6903) );
  XOR2_X1 U7856 ( .A(n6896), .B(keyinput14), .Z(n6901) );
  INV_X1 U7857 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6897) );
  XOR2_X1 U7858 ( .A(n6897), .B(keyinput1), .Z(n6900) );
  XNOR2_X1 U7859 ( .A(STATE2_REG_2__SCAN_IN), .B(keyinput90), .ZN(n6899) );
  XNOR2_X1 U7860 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(keyinput121), .ZN(
        n6898) );
  NAND4_X1 U7861 ( .A1(n6901), .A2(n6900), .A3(n6899), .A4(n6898), .ZN(n6902)
         );
  NOR3_X1 U7862 ( .A1(n6904), .A2(n6903), .A3(n6902), .ZN(n6921) );
  INV_X1 U7863 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6907) );
  AOI22_X1 U7864 ( .A1(n6907), .A2(keyinput42), .B1(keyinput79), .B2(n6906), 
        .ZN(n6905) );
  OAI221_X1 U7865 ( .B1(n6907), .B2(keyinput42), .C1(n6906), .C2(keyinput79), 
        .A(n6905), .ZN(n6919) );
  INV_X1 U7866 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U7867 ( .A1(n6910), .A2(keyinput30), .B1(n6909), .B2(keyinput67), 
        .ZN(n6908) );
  OAI221_X1 U7868 ( .B1(n6910), .B2(keyinput30), .C1(n6909), .C2(keyinput67), 
        .A(n6908), .ZN(n6918) );
  AOI22_X1 U7869 ( .A1(n6912), .A2(keyinput8), .B1(n5340), .B2(keyinput71), 
        .ZN(n6911) );
  OAI221_X1 U7870 ( .B1(n6912), .B2(keyinput8), .C1(n5340), .C2(keyinput71), 
        .A(n6911), .ZN(n6917) );
  INV_X1 U7871 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6915) );
  AOI22_X1 U7872 ( .A1(n6915), .A2(keyinput92), .B1(n6914), .B2(keyinput78), 
        .ZN(n6913) );
  OAI221_X1 U7873 ( .B1(n6915), .B2(keyinput92), .C1(n6914), .C2(keyinput78), 
        .A(n6913), .ZN(n6916) );
  NOR4_X1 U7874 ( .A1(n6919), .A2(n6918), .A3(n6917), .A4(n6916), .ZN(n6920)
         );
  NAND4_X1 U7875 ( .A1(n6923), .A2(n6922), .A3(n6921), .A4(n6920), .ZN(n7057)
         );
  AOI22_X1 U7876 ( .A1(n6926), .A2(keyinput36), .B1(n6925), .B2(keyinput107), 
        .ZN(n6924) );
  OAI221_X1 U7877 ( .B1(n6926), .B2(keyinput36), .C1(n6925), .C2(keyinput107), 
        .A(n6924), .ZN(n6938) );
  AOI22_X1 U7878 ( .A1(n6929), .A2(keyinput54), .B1(n6928), .B2(keyinput61), 
        .ZN(n6927) );
  OAI221_X1 U7879 ( .B1(n6929), .B2(keyinput54), .C1(n6928), .C2(keyinput61), 
        .A(n6927), .ZN(n6937) );
  AOI22_X1 U7880 ( .A1(n6932), .A2(keyinput63), .B1(keyinput103), .B2(n6931), 
        .ZN(n6930) );
  OAI221_X1 U7881 ( .B1(n6932), .B2(keyinput63), .C1(n6931), .C2(keyinput103), 
        .A(n6930), .ZN(n6936) );
  AOI22_X1 U7882 ( .A1(n6934), .A2(keyinput104), .B1(n6142), .B2(keyinput57), 
        .ZN(n6933) );
  OAI221_X1 U7883 ( .B1(n6934), .B2(keyinput104), .C1(n6142), .C2(keyinput57), 
        .A(n6933), .ZN(n6935) );
  NOR4_X1 U7884 ( .A1(n6938), .A2(n6937), .A3(n6936), .A4(n6935), .ZN(n6989)
         );
  INV_X1 U7885 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6940) );
  AOI22_X1 U7886 ( .A1(n6940), .A2(keyinput20), .B1(keyinput44), .B2(n6227), 
        .ZN(n6939) );
  OAI221_X1 U7887 ( .B1(n6940), .B2(keyinput20), .C1(n6227), .C2(keyinput44), 
        .A(n6939), .ZN(n6953) );
  AOI22_X1 U7888 ( .A1(n6943), .A2(keyinput60), .B1(n6942), .B2(keyinput75), 
        .ZN(n6941) );
  OAI221_X1 U7889 ( .B1(n6943), .B2(keyinput60), .C1(n6942), .C2(keyinput75), 
        .A(n6941), .ZN(n6952) );
  AOI22_X1 U7890 ( .A1(n6946), .A2(keyinput50), .B1(keyinput76), .B2(n6945), 
        .ZN(n6944) );
  OAI221_X1 U7891 ( .B1(n6946), .B2(keyinput50), .C1(n6945), .C2(keyinput76), 
        .A(n6944), .ZN(n6951) );
  INV_X1 U7892 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6949) );
  AOI22_X1 U7893 ( .A1(n6949), .A2(keyinput127), .B1(keyinput113), .B2(n6948), 
        .ZN(n6947) );
  OAI221_X1 U7894 ( .B1(n6949), .B2(keyinput127), .C1(n6948), .C2(keyinput113), 
        .A(n6947), .ZN(n6950) );
  NOR4_X1 U7895 ( .A1(n6953), .A2(n6952), .A3(n6951), .A4(n6950), .ZN(n6988)
         );
  AOI22_X1 U7896 ( .A1(n6956), .A2(keyinput3), .B1(n6955), .B2(keyinput49), 
        .ZN(n6954) );
  OAI221_X1 U7897 ( .B1(n6956), .B2(keyinput3), .C1(n6955), .C2(keyinput49), 
        .A(n6954), .ZN(n6969) );
  AOI22_X1 U7898 ( .A1(n6959), .A2(keyinput98), .B1(n6958), .B2(keyinput68), 
        .ZN(n6957) );
  OAI221_X1 U7899 ( .B1(n6959), .B2(keyinput98), .C1(n6958), .C2(keyinput68), 
        .A(n6957), .ZN(n6968) );
  AOI22_X1 U7900 ( .A1(n6962), .A2(keyinput74), .B1(n6961), .B2(keyinput39), 
        .ZN(n6960) );
  OAI221_X1 U7901 ( .B1(n6962), .B2(keyinput74), .C1(n6961), .C2(keyinput39), 
        .A(n6960), .ZN(n6967) );
  AOI22_X1 U7902 ( .A1(n6965), .A2(keyinput25), .B1(keyinput120), .B2(n6964), 
        .ZN(n6963) );
  OAI221_X1 U7903 ( .B1(n6965), .B2(keyinput25), .C1(n6964), .C2(keyinput120), 
        .A(n6963), .ZN(n6966) );
  NOR4_X1 U7904 ( .A1(n6969), .A2(n6968), .A3(n6967), .A4(n6966), .ZN(n6987)
         );
  AOI22_X1 U7905 ( .A1(n6972), .A2(keyinput56), .B1(n6971), .B2(keyinput80), 
        .ZN(n6970) );
  OAI221_X1 U7906 ( .B1(n6972), .B2(keyinput56), .C1(n6971), .C2(keyinput80), 
        .A(n6970), .ZN(n6985) );
  INV_X1 U7907 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6974) );
  AOI22_X1 U7908 ( .A1(n6975), .A2(keyinput28), .B1(n6974), .B2(keyinput115), 
        .ZN(n6973) );
  OAI221_X1 U7909 ( .B1(n6975), .B2(keyinput28), .C1(n6974), .C2(keyinput115), 
        .A(n6973), .ZN(n6984) );
  AOI22_X1 U7910 ( .A1(n6978), .A2(keyinput45), .B1(keyinput102), .B2(n6977), 
        .ZN(n6976) );
  OAI221_X1 U7911 ( .B1(n6978), .B2(keyinput45), .C1(n6977), .C2(keyinput102), 
        .A(n6976), .ZN(n6983) );
  AOI22_X1 U7912 ( .A1(n6981), .A2(keyinput86), .B1(n6980), .B2(keyinput105), 
        .ZN(n6979) );
  OAI221_X1 U7913 ( .B1(n6981), .B2(keyinput86), .C1(n6980), .C2(keyinput105), 
        .A(n6979), .ZN(n6982) );
  NOR4_X1 U7914 ( .A1(n6985), .A2(n6984), .A3(n6983), .A4(n6982), .ZN(n6986)
         );
  NAND4_X1 U7915 ( .A1(n6989), .A2(n6988), .A3(n6987), .A4(n6986), .ZN(n7056)
         );
  AOI22_X1 U7916 ( .A1(n6992), .A2(keyinput101), .B1(n6991), .B2(keyinput41), 
        .ZN(n6990) );
  OAI221_X1 U7917 ( .B1(n6992), .B2(keyinput101), .C1(n6991), .C2(keyinput41), 
        .A(n6990), .ZN(n6996) );
  XOR2_X1 U7918 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .B(keyinput69), .Z(n6995)
         );
  XNOR2_X1 U7919 ( .A(n6993), .B(keyinput55), .ZN(n6994) );
  OR3_X1 U7920 ( .A1(n6996), .A2(n6995), .A3(n6994), .ZN(n7005) );
  AOI22_X1 U7921 ( .A1(n6999), .A2(keyinput84), .B1(keyinput66), .B2(n6998), 
        .ZN(n6997) );
  OAI221_X1 U7922 ( .B1(n6999), .B2(keyinput84), .C1(n6998), .C2(keyinput66), 
        .A(n6997), .ZN(n7004) );
  INV_X1 U7923 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n7001) );
  AOI22_X1 U7924 ( .A1(n7002), .A2(keyinput59), .B1(keyinput16), .B2(n7001), 
        .ZN(n7000) );
  OAI221_X1 U7925 ( .B1(n7002), .B2(keyinput59), .C1(n7001), .C2(keyinput16), 
        .A(n7000), .ZN(n7003) );
  NOR3_X1 U7926 ( .A1(n7005), .A2(n7004), .A3(n7003), .ZN(n7054) );
  NAND2_X1 U7927 ( .A1(n7007), .A2(keyinput89), .ZN(n7006) );
  OAI221_X1 U7928 ( .B1(n7008), .B2(keyinput124), .C1(n7007), .C2(keyinput89), 
        .A(n7006), .ZN(n7021) );
  AOI22_X1 U7929 ( .A1(n7011), .A2(keyinput85), .B1(keyinput9), .B2(n7010), 
        .ZN(n7009) );
  OAI221_X1 U7930 ( .B1(n7011), .B2(keyinput85), .C1(n7010), .C2(keyinput9), 
        .A(n7009), .ZN(n7020) );
  AOI22_X1 U7931 ( .A1(n7014), .A2(keyinput117), .B1(keyinput82), .B2(n7013), 
        .ZN(n7012) );
  OAI221_X1 U7932 ( .B1(n7014), .B2(keyinput117), .C1(n7013), .C2(keyinput82), 
        .A(n7012), .ZN(n7019) );
  AOI22_X1 U7933 ( .A1(n7017), .A2(keyinput126), .B1(keyinput93), .B2(n7016), 
        .ZN(n7015) );
  OAI221_X1 U7934 ( .B1(n7017), .B2(keyinput126), .C1(n7016), .C2(keyinput93), 
        .A(n7015), .ZN(n7018) );
  NOR4_X1 U7935 ( .A1(n7021), .A2(n7020), .A3(n7019), .A4(n7018), .ZN(n7053)
         );
  AOI22_X1 U7936 ( .A1(n7064), .A2(keyinput34), .B1(n7023), .B2(keyinput114), 
        .ZN(n7022) );
  OAI221_X1 U7937 ( .B1(n7064), .B2(keyinput34), .C1(n7023), .C2(keyinput114), 
        .A(n7022), .ZN(n7035) );
  AOI22_X1 U7938 ( .A1(n7026), .A2(keyinput64), .B1(keyinput112), .B2(n7025), 
        .ZN(n7024) );
  OAI221_X1 U7939 ( .B1(n7026), .B2(keyinput64), .C1(n7025), .C2(keyinput112), 
        .A(n7024), .ZN(n7034) );
  INV_X1 U7940 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n7029) );
  INV_X1 U7941 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n7028) );
  AOI22_X1 U7942 ( .A1(n7029), .A2(keyinput24), .B1(n7028), .B2(keyinput122), 
        .ZN(n7027) );
  OAI221_X1 U7943 ( .B1(n7029), .B2(keyinput24), .C1(n7028), .C2(keyinput122), 
        .A(n7027), .ZN(n7033) );
  INV_X1 U7944 ( .A(DATAI_23_), .ZN(n7031) );
  AOI22_X1 U7945 ( .A1(n7031), .A2(keyinput96), .B1(n6175), .B2(keyinput100), 
        .ZN(n7030) );
  OAI221_X1 U7946 ( .B1(n7031), .B2(keyinput96), .C1(n6175), .C2(keyinput100), 
        .A(n7030), .ZN(n7032) );
  NOR4_X1 U7947 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n7052)
         );
  INV_X1 U7948 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n7037) );
  AOI22_X1 U7949 ( .A1(n7038), .A2(keyinput109), .B1(n7037), .B2(keyinput118), 
        .ZN(n7036) );
  OAI221_X1 U7950 ( .B1(n7038), .B2(keyinput109), .C1(n7037), .C2(keyinput118), 
        .A(n7036), .ZN(n7050) );
  AOI22_X1 U7951 ( .A1(n7040), .A2(keyinput125), .B1(n5055), .B2(keyinput88), 
        .ZN(n7039) );
  OAI221_X1 U7952 ( .B1(n7040), .B2(keyinput125), .C1(n5055), .C2(keyinput88), 
        .A(n7039), .ZN(n7049) );
  AOI22_X1 U7953 ( .A1(n7043), .A2(keyinput15), .B1(keyinput123), .B2(n7042), 
        .ZN(n7041) );
  OAI221_X1 U7954 ( .B1(n7043), .B2(keyinput15), .C1(n7042), .C2(keyinput123), 
        .A(n7041), .ZN(n7048) );
  AOI22_X1 U7955 ( .A1(n7046), .A2(keyinput33), .B1(keyinput5), .B2(n7045), 
        .ZN(n7044) );
  OAI221_X1 U7956 ( .B1(n7046), .B2(keyinput33), .C1(n7045), .C2(keyinput5), 
        .A(n7044), .ZN(n7047) );
  NOR4_X1 U7957 ( .A1(n7050), .A2(n7049), .A3(n7048), .A4(n7047), .ZN(n7051)
         );
  NAND4_X1 U7958 ( .A1(n7054), .A2(n7053), .A3(n7052), .A4(n7051), .ZN(n7055)
         );
  NOR4_X1 U7959 ( .A1(n7058), .A2(n7057), .A3(n7056), .A4(n7055), .ZN(n7059)
         );
  OAI21_X1 U7960 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n7060), .A(n7059), 
        .ZN(n7067) );
  AOI22_X1 U7961 ( .A1(n7062), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n7061), .ZN(n7063) );
  OAI21_X1 U7962 ( .B1(n7065), .B2(n7064), .A(n7063), .ZN(n7066) );
  XNOR2_X1 U7963 ( .A(n7067), .B(n7066), .ZN(U2945) );
  AND2_X2 U4089 ( .A1(n4442), .A2(n3154), .ZN(n3338) );
  AND4_X1 U4177 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3275)
         );
  AND4_X1 U4182 ( .A1(n3263), .A2(n3262), .A3(n3261), .A4(n3260), .ZN(n3274)
         );
  AND4_X1 U4187 ( .A1(n3267), .A2(n3266), .A3(n3265), .A4(n3264), .ZN(n3273)
         );
  AND2_X1 U3580 ( .A1(n3289), .A2(n3288), .ZN(n3311) );
  OAI22_X1 U4205 ( .A1(n4340), .A2(n3279), .B1(n4240), .B2(n4647), .ZN(n3280)
         );
  BUF_X1 U6138 ( .A(n4962), .Z(n5529) );
  NAND2_X1 U6598 ( .A1(n5504), .A2(n5503), .ZN(n5502) );
  XNOR2_X1 U5079 ( .A(n4104), .B(n4103), .ZN(n4392) );
  OR2_X2 U3718 ( .A1(n3292), .A2(n3127), .ZN(n4145) );
  NOR2_X1 U5077 ( .A1(n4102), .A2(n4997), .ZN(n4383) );
  BUF_X2 U3543 ( .A(n3312), .Z(n5385) );
  CLKBUF_X2 U3556 ( .A(n3442), .Z(n3467) );
  CLKBUF_X1 U3569 ( .A(n3324), .Z(n4289) );
  CLKBUF_X1 U3667 ( .A(n3387), .Z(n3388) );
  AND4_X1 U3668 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), .ZN(n3272)
         );
  CLKBUF_X1 U3674 ( .A(n3315), .Z(n4115) );
  NAND2_X1 U3679 ( .A1(n4657), .A2(n3292), .ZN(n4421) );
  CLKBUF_X1 U3680 ( .A(n5504), .Z(n3099) );
  CLKBUF_X1 U3682 ( .A(n4834), .Z(n5377) );
  NAND2_X1 U3737 ( .A1(n5529), .A2(n5528), .ZN(n5572) );
  AND2_X2 U3769 ( .A1(n3153), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4442)
         );
  AND4_X2 U3796 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3159)
         );
  INV_X1 U3860 ( .A(n3292), .ZN(n7068) );
  NAND4_X2 U3951 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n4254)
         );
  CLKBUF_X1 U4011 ( .A(n5565), .Z(n3100) );
endmodule

