

module b17_C_AntiSAT_k_256_4 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9793, n9795, n9796, n9797, n9798, n9799, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272;

  INV_X1 U11237 ( .A(n20086), .ZN(n20078) );
  INV_X1 U11238 ( .A(n14372), .ZN(n14376) );
  OAI21_X1 U11239 ( .B1(n10993), .B2(n10095), .A(n10996), .ZN(n10094) );
  NAND2_X1 U11240 ( .A1(n10843), .A2(n13630), .ZN(n10844) );
  XNOR2_X1 U11241 ( .A(n10804), .B(n10834), .ZN(n10978) );
  CLKBUF_X2 U11242 ( .A(n12766), .Z(n16013) );
  NAND2_X1 U11243 ( .A1(n13188), .A2(n13187), .ZN(n14065) );
  NOR2_X1 U11244 ( .A1(n13251), .A2(n10134), .ZN(n13587) );
  NOR2_X2 U11246 ( .A1(n15041), .A2(n15339), .ZN(n15043) );
  NAND2_X1 U11247 ( .A1(n10641), .A2(n10656), .ZN(n19731) );
  NAND2_X1 U11248 ( .A1(n10635), .A2(n10636), .ZN(n10712) );
  NAND2_X1 U11249 ( .A1(n11191), .A2(n10044), .ZN(n17333) );
  NAND2_X1 U11250 ( .A1(n9820), .A2(n10645), .ZN(n19770) );
  INV_X1 U11251 ( .A(n13140), .ZN(n13154) );
  NAND2_X1 U11252 ( .A1(n10618), .A2(n10617), .ZN(n13712) );
  INV_X1 U11253 ( .A(n17186), .ZN(n9806) );
  INV_X1 U11254 ( .A(n9842), .ZN(n17210) );
  CLKBUF_X2 U11255 ( .A(n10679), .Z(n14141) );
  AND2_X1 U11256 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10553), .ZN(
        n14151) );
  INV_X2 U11257 ( .A(n11055), .ZN(n13905) );
  OR2_X1 U11258 ( .A1(n11014), .A2(n11013), .ZN(n10244) );
  INV_X4 U11259 ( .A(n21272), .ZN(n9801) );
  CLKBUF_X2 U11260 ( .A(n10542), .Z(n14353) );
  CLKBUF_X2 U11261 ( .A(n10544), .Z(n14351) );
  CLKBUF_X2 U11262 ( .A(n10308), .Z(n14352) );
  CLKBUF_X2 U11264 ( .A(n11949), .Z(n12376) );
  CLKBUF_X2 U11265 ( .A(n11802), .Z(n9803) );
  CLKBUF_X2 U11266 ( .A(n11874), .Z(n12351) );
  CLKBUF_X2 U11267 ( .A(n11876), .Z(n9804) );
  NAND3_X1 U11268 ( .A1(n9911), .A2(n9827), .A3(n9910), .ZN(n12793) );
  CLKBUF_X1 U11269 ( .A(n11759), .Z(n20249) );
  NAND2_X1 U11270 ( .A1(n10315), .A2(n10314), .ZN(n10344) );
  AND2_X4 U11271 ( .A1(n13069), .A2(n11635), .ZN(n11729) );
  AND2_X2 U11272 ( .A1(n13215), .A2(n11634), .ZN(n11949) );
  NOR2_X2 U11273 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11635) );
  CLKBUF_X1 U11274 ( .A(n19691), .Z(n9793) );
  OAI221_X1 U11275 ( .B1(n13510), .B2(n16413), .C1(n19206), .C2(n16413), .A(
        n20977), .ZN(n19691) );
  INV_X1 U11277 ( .A(n21271), .ZN(n9795) );
  CLKBUF_X2 U11278 ( .A(n11785), .Z(n12447) );
  INV_X1 U11279 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9998) );
  NOR2_X1 U11280 ( .A1(n9972), .A2(n10645), .ZN(n10705) );
  XOR2_X1 U11282 ( .A(n21036), .B(keyinput171), .Z(n21038) );
  NAND2_X1 U11284 ( .A1(n10779), .A2(n9826), .ZN(n10804) );
  AOI21_X1 U11286 ( .B1(n11119), .B2(n11295), .A(n9931), .ZN(n9930) );
  NAND2_X1 U11287 ( .A1(n11772), .A2(n11771), .ZN(n11847) );
  XNOR2_X1 U11288 ( .A(n13085), .B(n12695), .ZN(n20166) );
  AND2_X1 U11289 ( .A1(n11673), .A2(n11672), .ZN(n11759) );
  NAND2_X1 U11290 ( .A1(n10885), .A2(n10941), .ZN(n10888) );
  NAND2_X1 U11291 ( .A1(n9989), .A2(n9822), .ZN(n13964) );
  NAND2_X1 U11292 ( .A1(n10635), .A2(n10648), .ZN(n13745) );
  NOR2_X1 U11293 ( .A1(n17747), .A2(n11270), .ZN(n11272) );
  OAI21_X1 U11294 ( .B1(n17858), .B2(n9932), .A(n9930), .ZN(n17850) );
  NOR2_X1 U11295 ( .A1(n11736), .A2(n11735), .ZN(n11752) );
  INV_X1 U11296 ( .A(n11759), .ZN(n13824) );
  NAND2_X1 U11297 ( .A1(n10945), .A2(n10941), .ZN(n14022) );
  NOR2_X1 U11298 ( .A1(n15147), .A2(n15146), .ZN(n15145) );
  NAND2_X1 U11299 ( .A1(n11375), .A2(n13515), .ZN(n11511) );
  NOR2_X1 U11300 ( .A1(n13621), .A2(n16323), .ZN(n13639) );
  NOR2_X1 U11301 ( .A1(n10978), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13598) );
  NAND2_X1 U11302 ( .A1(n10635), .A2(n10642), .ZN(n19456) );
  INV_X2 U11303 ( .A(n17163), .ZN(n11145) );
  INV_X1 U11304 ( .A(n9801), .ZN(n11038) );
  INV_X1 U11305 ( .A(n17699), .ZN(n17901) );
  NAND2_X1 U11306 ( .A1(n16485), .A2(n17820), .ZN(n16470) );
  NOR3_X1 U11307 ( .A1(n17607), .A2(n17615), .A3(n17973), .ZN(n17597) );
  INV_X1 U11308 ( .A(n20043), .ZN(n20081) );
  CLKBUF_X3 U11309 ( .A(n13635), .Z(n19075) );
  NOR2_X2 U11310 ( .A1(n17136), .A2(n16769), .ZN(n17112) );
  INV_X2 U11311 ( .A(n10244), .ZN(n17231) );
  NAND2_X1 U11312 ( .A1(n17832), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17831) );
  INV_X1 U11313 ( .A(n20050), .ZN(n15945) );
  INV_X1 U11314 ( .A(n20171), .ZN(n20163) );
  INV_X1 U11315 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19951) );
  OR2_X1 U11316 ( .A1(n11236), .A2(n11235), .ZN(n9796) );
  INV_X4 U11317 ( .A(n10227), .ZN(n17195) );
  XNOR2_X2 U11319 ( .A(n10972), .B(n11397), .ZN(n10974) );
  INV_X2 U11320 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15725) );
  NOR2_X4 U11321 ( .A1(n15886), .A2(n13840), .ZN(n17284) );
  NAND4_X1 U11322 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n9797) );
  INV_X4 U11323 ( .A(n11758), .ZN(n20238) );
  INV_X2 U11324 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9798) );
  INV_X2 U11325 ( .A(n13515), .ZN(n14024) );
  BUF_X4 U11326 ( .A(n13906), .Z(n9799) );
  AOI21_X2 U11327 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17620), .A(
        n18392), .ZN(n17747) );
  AOI21_X1 U11328 ( .B1(n15558), .B2(n10118), .A(n10110), .ZN(n10109) );
  NOR2_X2 U11329 ( .A1(n15406), .A2(n15578), .ZN(n15556) );
  XNOR2_X1 U11330 ( .A(n12637), .B(n12636), .ZN(n12800) );
  AOI21_X1 U11331 ( .B1(n12465), .B2(n12466), .A(n12637), .ZN(n14716) );
  AOI21_X1 U11332 ( .B1(n14425), .B2(n14424), .A(n14411), .ZN(n14737) );
  NAND3_X1 U11333 ( .A1(n12781), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14762), .ZN(n14739) );
  NOR2_X1 U11334 ( .A1(n15375), .A2(n15534), .ZN(n15361) );
  OAI21_X1 U11335 ( .B1(n13964), .B2(n11002), .A(n10955), .ZN(n10956) );
  OAI21_X1 U11336 ( .B1(n14411), .B2(n14412), .A(n12465), .ZN(n14725) );
  NAND2_X1 U11337 ( .A1(n10938), .A2(n9990), .ZN(n9989) );
  OAI21_X1 U11338 ( .B1(n11589), .B2(n10190), .A(n10187), .ZN(n15384) );
  INV_X1 U11340 ( .A(n14315), .ZN(n9802) );
  OAI21_X1 U11341 ( .B1(n15416), .B2(n11588), .A(n15413), .ZN(n15404) );
  XNOR2_X1 U11342 ( .A(n14259), .B(n10243), .ZN(n15147) );
  NAND2_X1 U11343 ( .A1(n15150), .A2(n14237), .ZN(n14259) );
  NOR2_X1 U11344 ( .A1(n15141), .A2(n15142), .ZN(n13995) );
  AOI21_X1 U11345 ( .B1(n13480), .B2(n13478), .A(n10801), .ZN(n13584) );
  AND2_X1 U11346 ( .A1(n10066), .A2(n16022), .ZN(n10065) );
  NAND2_X1 U11347 ( .A1(n10777), .A2(n19141), .ZN(n10802) );
  CLKBUF_X1 U11348 ( .A(n10988), .Z(n10990) );
  NAND2_X1 U11349 ( .A1(n10978), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13595) );
  NAND2_X1 U11350 ( .A1(n17295), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n17294) );
  NOR2_X1 U11351 ( .A1(n10958), .A2(n10957), .ZN(n13923) );
  AND2_X1 U11352 ( .A1(n14985), .A2(n9916), .ZN(n14988) );
  INV_X1 U11353 ( .A(n10804), .ZN(n10836) );
  AND2_X1 U11354 ( .A1(n10834), .A2(n10833), .ZN(n10835) );
  AND2_X1 U11355 ( .A1(n13813), .A2(n12775), .ZN(n14819) );
  NAND2_X1 U11356 ( .A1(n14022), .A2(n10944), .ZN(n10958) );
  AND2_X2 U11357 ( .A1(n20079), .A2(n13499), .ZN(n20086) );
  OAI21_X1 U11358 ( .B1(n16429), .B2(n11269), .A(n10041), .ZN(n10040) );
  NOR2_X2 U11359 ( .A1(n19697), .A2(n19577), .ZN(n19633) );
  AND2_X1 U11360 ( .A1(n10746), .A2(n10745), .ZN(n10834) );
  AND2_X1 U11362 ( .A1(n12739), .A2(n12738), .ZN(n16029) );
  NOR2_X2 U11363 ( .A1(n19720), .A2(n19719), .ZN(n19830) );
  NAND2_X2 U11365 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17849), .ZN(n17769) );
  INV_X1 U11366 ( .A(n12016), .ZN(n9918) );
  INV_X1 U11367 ( .A(n17911), .ZN(n17849) );
  AND2_X1 U11368 ( .A1(n13151), .A2(n13186), .ZN(n13152) );
  INV_X1 U11369 ( .A(n17753), .ZN(n17825) );
  NAND2_X1 U11370 ( .A1(n17916), .A2(n17744), .ZN(n17661) );
  OR2_X1 U11371 ( .A1(n13150), .A2(n13149), .ZN(n13151) );
  NAND2_X1 U11372 ( .A1(n18731), .A2(n18939), .ZN(n16583) );
  NAND2_X1 U11373 ( .A1(n9818), .A2(n10645), .ZN(n19686) );
  NAND2_X1 U11374 ( .A1(n11911), .A2(n13402), .ZN(n11970) );
  NAND2_X1 U11375 ( .A1(n10037), .A2(n9882), .ZN(n18731) );
  AND2_X1 U11377 ( .A1(n10655), .A2(n13712), .ZN(n10078) );
  CLKBUF_X1 U11378 ( .A(n12698), .Z(n20481) );
  AND2_X1 U11379 ( .A1(n11891), .A2(n11924), .ZN(n11911) );
  NOR2_X1 U11380 ( .A1(n17438), .A2(n18291), .ZN(n17363) );
  CLKBUF_X1 U11381 ( .A(n13242), .Z(n9817) );
  NAND2_X1 U11382 ( .A1(n18213), .A2(n18752), .ZN(n18149) );
  NAND2_X1 U11383 ( .A1(n12958), .A2(n12957), .ZN(n15698) );
  NAND2_X1 U11384 ( .A1(n11910), .A2(n11909), .ZN(n13402) );
  AND2_X1 U11385 ( .A1(n10624), .A2(n15695), .ZN(n10642) );
  NAND2_X1 U11386 ( .A1(n17850), .A2(n10246), .ZN(n11123) );
  NAND2_X1 U11387 ( .A1(n10871), .A2(n10941), .ZN(n10869) );
  XNOR2_X1 U11388 ( .A(n11892), .B(n20365), .ZN(n20476) );
  CLKBUF_X1 U11389 ( .A(n16287), .Z(n16310) );
  NAND2_X1 U11390 ( .A1(n10416), .A2(n10415), .ZN(n10622) );
  OR2_X1 U11391 ( .A1(n10858), .A2(n10006), .ZN(n10871) );
  CLKBUF_X1 U11392 ( .A(n17534), .Z(n17543) );
  OR2_X1 U11393 ( .A1(n10614), .A2(n10613), .ZN(n10628) );
  NAND2_X1 U11394 ( .A1(n10859), .A2(n10848), .ZN(n10858) );
  XNOR2_X1 U11395 ( .A(n10418), .B(n10419), .ZN(n10606) );
  NAND2_X1 U11396 ( .A1(n10859), .A2(n13515), .ZN(n10941) );
  NAND2_X1 U11397 ( .A1(n11849), .A2(n11848), .ZN(n20276) );
  NOR2_X2 U11398 ( .A1(n18272), .A2(n17542), .ZN(n17534) );
  OAI22_X1 U11399 ( .A1(n10413), .A2(n16379), .B1(n19980), .B2(n19935), .ZN(
        n10419) );
  NAND2_X1 U11400 ( .A1(n9938), .A2(n10048), .ZN(n11118) );
  INV_X1 U11401 ( .A(n10131), .ZN(n11390) );
  NOR2_X1 U11402 ( .A1(n11247), .A2(n11252), .ZN(n12834) );
  CLKBUF_X1 U11403 ( .A(n10406), .Z(n10424) );
  OR2_X1 U11404 ( .A1(n11867), .A2(n11868), .ZN(n11865) );
  OAI211_X1 U11405 ( .C1(n10406), .C2(n16365), .A(n10242), .B(n10395), .ZN(
        n10614) );
  AND2_X1 U11406 ( .A1(n10840), .A2(n10841), .ZN(n10853) );
  OAI211_X1 U11407 ( .C1(n10406), .C2(n16356), .A(n10412), .B(n10411), .ZN(
        n10418) );
  NAND2_X1 U11408 ( .A1(n17882), .A2(n11113), .ZN(n17871) );
  NAND2_X1 U11409 ( .A1(n17884), .A2(n17883), .ZN(n17882) );
  NAND2_X1 U11410 ( .A1(n11783), .A2(n9844), .ZN(n11846) );
  OR2_X1 U11411 ( .A1(n17870), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10049) );
  NAND2_X1 U11412 ( .A1(n10373), .A2(n11347), .ZN(n11557) );
  OAI211_X1 U11413 ( .C1(n10367), .C2(n10366), .A(n15796), .B(n11555), .ZN(
        n11553) );
  AND2_X1 U11414 ( .A1(n13013), .A2(n11780), .ZN(n13798) );
  OR2_X1 U11415 ( .A1(n10963), .A2(n14024), .ZN(n11380) );
  NAND2_X1 U11416 ( .A1(n13002), .A2(n20249), .ZN(n13001) );
  AND3_X1 U11417 ( .A1(n14371), .A2(n10317), .A3(n10316), .ZN(n16394) );
  INV_X1 U11418 ( .A(n18282), .ZN(n13836) );
  AND2_X1 U11419 ( .A1(n11777), .A2(n11763), .ZN(n13002) );
  AOI211_X1 U11420 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n11035), .B(n11034), .ZN(n17417) );
  AND2_X1 U11421 ( .A1(n14395), .A2(n12530), .ZN(n12985) );
  AND2_X1 U11422 ( .A1(n10346), .A2(n10364), .ZN(n11549) );
  OR2_X1 U11423 ( .A1(n12523), .A2(n11764), .ZN(n13015) );
  AND2_X1 U11424 ( .A1(n13784), .A2(n12690), .ZN(n12687) );
  AND3_X1 U11425 ( .A1(n10364), .A2(n10354), .A3(n10344), .ZN(n10360) );
  OR2_X1 U11426 ( .A1(n10571), .A2(n10570), .ZN(n11392) );
  INV_X1 U11427 ( .A(n10345), .ZN(n10343) );
  INV_X1 U11428 ( .A(n10364), .ZN(n11334) );
  INV_X1 U11429 ( .A(n12972), .ZN(n19340) );
  NAND2_X2 U11430 ( .A1(n10262), .A2(n10261), .ZN(n13570) );
  OR2_X1 U11431 ( .A1(n11813), .A2(n11812), .ZN(n12746) );
  INV_X2 U11432 ( .A(n13779), .ZN(n13784) );
  NAND2_X1 U11433 ( .A1(n10340), .A2(n10339), .ZN(n10368) );
  NAND2_X1 U11434 ( .A1(n11705), .A2(n11704), .ZN(n12690) );
  NAND4_X2 U11435 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n12524) );
  AND3_X1 U11436 ( .A1(n11721), .A2(n11720), .A3(n11719), .ZN(n11727) );
  NAND2_X1 U11437 ( .A1(n10239), .A2(n10300), .ZN(n10301) );
  NAND2_X2 U11438 ( .A1(n18945), .A2(n18822), .ZN(n18869) );
  AND4_X1 U11439 ( .A1(n11703), .A2(n11702), .A3(n11701), .A4(n11700), .ZN(
        n11704) );
  AND4_X1 U11440 ( .A1(n11699), .A2(n11698), .A3(n11697), .A4(n11696), .ZN(
        n11705) );
  AND4_X1 U11441 ( .A1(n11667), .A2(n11666), .A3(n11665), .A4(n11664), .ZN(
        n11673) );
  AND4_X1 U11442 ( .A1(n11671), .A2(n11670), .A3(n11669), .A4(n11668), .ZN(
        n11672) );
  INV_X8 U11443 ( .A(n11054), .ZN(n17237) );
  NOR2_X1 U11444 ( .A1(n11734), .A2(n11733), .ZN(n11735) );
  AND4_X1 U11445 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n11751) );
  AND4_X1 U11446 ( .A1(n11744), .A2(n11743), .A3(n11742), .A4(n11741), .ZN(
        n11750) );
  AND4_X1 U11447 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n11749) );
  AND4_X1 U11448 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(
        n11721) );
  AND4_X1 U11449 ( .A1(n11714), .A2(n11713), .A3(n11712), .A4(n11711), .ZN(
        n11720) );
  AND4_X1 U11450 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n11643) );
  AND4_X1 U11451 ( .A1(n11691), .A2(n11690), .A3(n11689), .A4(n11688), .ZN(
        n11692) );
  AND4_X1 U11452 ( .A1(n11687), .A2(n11686), .A3(n11685), .A4(n11684), .ZN(
        n11693) );
  AND4_X1 U11453 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n11694) );
  AND4_X1 U11454 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n11695) );
  AND3_X1 U11455 ( .A1(n11660), .A2(n11659), .A3(n11658), .ZN(n11661) );
  AND4_X1 U11456 ( .A1(n11640), .A2(n11639), .A3(n11638), .A4(n11637), .ZN(
        n11641) );
  AND4_X1 U11457 ( .A1(n11628), .A2(n11627), .A3(n11626), .A4(n11625), .ZN(
        n11642) );
  INV_X2 U11458 ( .A(n17246), .ZN(n17215) );
  NOR2_X2 U11459 ( .A1(n18514), .A2(n18513), .ZN(n18613) );
  AND3_X1 U11460 ( .A1(n10299), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10298), .ZN(n10300) );
  INV_X1 U11461 ( .A(n11011), .ZN(n17177) );
  OR2_X2 U11462 ( .A1(n18897), .A2(n11016), .ZN(n11054) );
  NAND2_X2 U11463 ( .A1(n19988), .A2(n19861), .ZN(n19915) );
  BUF_X2 U11464 ( .A(n11801), .Z(n12448) );
  BUF_X2 U11465 ( .A(n10545), .Z(n14354) );
  BUF_X2 U11466 ( .A(n11807), .Z(n12420) );
  NAND2_X2 U11467 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11006), .ZN(
        n17246) );
  INV_X2 U11468 ( .A(n16572), .ZN(n16574) );
  INV_X1 U11469 ( .A(n19840), .ZN(n19154) );
  OR3_X2 U11470 ( .A1(n18892), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n16718) );
  INV_X4 U11471 ( .A(n17151), .ZN(n11226) );
  OR2_X2 U11472 ( .A1(n11010), .A2(n11009), .ZN(n17186) );
  INV_X2 U11473 ( .A(n18946), .ZN(n18945) );
  AND2_X2 U11474 ( .A1(n11635), .A2(n11634), .ZN(n11874) );
  OR2_X2 U11475 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15793), .ZN(
        n11056) );
  AND2_X2 U11476 ( .A1(n11618), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13215) );
  AND2_X2 U11477 ( .A1(n11620), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11634) );
  NAND3_X1 U11478 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n18744), .ZN(n11076) );
  NAND2_X1 U11479 ( .A1(n18897), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11010) );
  NAND3_X1 U11480 ( .A1(n18744), .A2(n18897), .A3(n21179), .ZN(n17072) );
  CLKBUF_X1 U11481 ( .A(n10379), .Z(n15711) );
  NAND2_X1 U11482 ( .A1(n18916), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11012) );
  AND2_X2 U11483 ( .A1(n10201), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11629) );
  INV_X1 U11484 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18910) );
  INV_X1 U11485 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10379) );
  INV_X2 U11486 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16379) );
  AND2_X1 U11487 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18744) );
  INV_X2 U11488 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21179) );
  INV_X1 U11489 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11618) );
  AND2_X1 U11490 ( .A1(n11847), .A2(n11846), .ZN(n11850) );
  XNOR2_X1 U11491 ( .A(n11847), .B(n11784), .ZN(n11938) );
  AOI21_X1 U11492 ( .B1(n10380), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10381), 
        .ZN(n10382) );
  NOR2_X2 U11493 ( .A1(n18739), .A2(n18759), .ZN(n18213) );
  NOR2_X2 U11494 ( .A1(n17546), .A2(n17376), .ZN(n17368) );
  NAND2_X2 U11495 ( .A1(n16034), .A2(n12732), .ZN(n16031) );
  NAND2_X1 U11497 ( .A1(n11727), .A2(n11726), .ZN(n9805) );
  NAND2_X2 U11498 ( .A1(n17697), .A2(n11132), .ZN(n17659) );
  OR2_X1 U11499 ( .A1(n13085), .A2(n12696), .ZN(n12697) );
  NAND2_X2 U11500 ( .A1(n12778), .A2(n14858), .ZN(n14785) );
  NAND2_X2 U11501 ( .A1(n14786), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12780) );
  AOI21_X1 U11502 ( .B1(n14796), .B2(n10231), .A(n14858), .ZN(n12777) );
  OAI21_X2 U11503 ( .B1(n10196), .B2(n9984), .A(n9982), .ZN(n15423) );
  NAND2_X2 U11504 ( .A1(n9828), .A2(n10846), .ZN(n10196) );
  INV_X1 U11505 ( .A(n14272), .ZN(n9807) );
  OR3_X4 U11506 ( .A1(n15493), .A2(n10083), .A3(n10082), .ZN(n9840) );
  NOR2_X2 U11507 ( .A1(n13448), .A2(n13488), .ZN(n13487) );
  INV_X1 U11508 ( .A(n11312), .ZN(n16393) );
  NAND2_X4 U11509 ( .A1(n10302), .A2(n10301), .ZN(n10354) );
  INV_X2 U11510 ( .A(n10352), .ZN(n10328) );
  OAI21_X2 U11511 ( .B1(n12638), .B2(n12661), .A(n13825), .ZN(n11757) );
  AND2_X4 U11512 ( .A1(n12690), .A2(n9797), .ZN(n12529) );
  NAND2_X2 U11513 ( .A1(n10615), .A2(n10074), .ZN(n10617) );
  AND2_X2 U11514 ( .A1(n10405), .A2(n10387), .ZN(n10615) );
  NOR2_X2 U11515 ( .A1(n18933), .A2(n18149), .ZN(n18113) );
  NAND2_X2 U11516 ( .A1(n11312), .A2(n11582), .ZN(n11546) );
  NAND2_X1 U11517 ( .A1(n16397), .A2(n19970), .ZN(n11312) );
  NAND2_X1 U11518 ( .A1(n19971), .A2(n10368), .ZN(n11582) );
  NAND2_X2 U11519 ( .A1(n11844), .A2(n11769), .ZN(n11858) );
  NAND2_X1 U11520 ( .A1(n15440), .A2(n15439), .ZN(n15658) );
  NOR2_X2 U11521 ( .A1(n14807), .A2(n16045), .ZN(n14796) );
  NAND2_X1 U11522 ( .A1(n11359), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9809) );
  NAND2_X2 U11523 ( .A1(n11359), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10406) );
  XNOR2_X2 U11525 ( .A(n12713), .B(n12706), .ZN(n13289) );
  NAND2_X2 U11526 ( .A1(n20197), .A2(n12705), .ZN(n12713) );
  NOR2_X4 U11527 ( .A1(n13597), .A2(n13598), .ZN(n13596) );
  INV_X1 U11528 ( .A(n12766), .ZN(n9810) );
  OR2_X1 U11529 ( .A1(n18897), .A2(n11016), .ZN(n9811) );
  NOR2_X1 U11530 ( .A1(n11010), .A2(n11012), .ZN(n9812) );
  INV_X1 U11531 ( .A(n14159), .ZN(n9813) );
  INV_X1 U11532 ( .A(n14159), .ZN(n9814) );
  INV_X1 U11533 ( .A(n14159), .ZN(n10308) );
  NAND2_X2 U11534 ( .A1(n15710), .A2(n16370), .ZN(n14159) );
  INV_X1 U11535 ( .A(n9796), .ZN(n9815) );
  AND2_X2 U11536 ( .A1(n14577), .A2(n14578), .ZN(n14477) );
  NOR2_X2 U11537 ( .A1(n14490), .A2(n10209), .ZN(n14577) );
  INV_X1 U11538 ( .A(n13794), .ZN(n9816) );
  XNOR2_X2 U11539 ( .A(n11936), .B(n11935), .ZN(n12694) );
  NAND2_X2 U11540 ( .A1(n11818), .A2(n11817), .ZN(n11936) );
  OR3_X2 U11541 ( .A1(n11014), .A2(n21179), .A3(n18897), .ZN(n9842) );
  XNOR2_X2 U11542 ( .A(n11890), .B(n11889), .ZN(n11924) );
  NOR2_X4 U11543 ( .A1(n17481), .A2(n15789), .ZN(n16582) );
  NOR3_X2 U11544 ( .A1(n9909), .A2(n13836), .A3(n9908), .ZN(n17481) );
  OAI21_X2 U11545 ( .B1(n13817), .B2(n11757), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11844) );
  AND2_X2 U11546 ( .A1(n14354), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10678) );
  NAND2_X1 U11547 ( .A1(n11765), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11896) );
  NAND2_X1 U11548 ( .A1(n12475), .A2(n13824), .ZN(n12493) );
  AND2_X1 U11549 ( .A1(n20079), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13669) );
  OR2_X1 U11550 ( .A1(n11332), .A2(n10533), .ZN(n16398) );
  AND4_X1 U11551 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10766) );
  AND4_X1 U11552 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10765) );
  AND2_X1 U11553 ( .A1(n13498), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13499) );
  CLKBUF_X1 U11554 ( .A(n11729), .Z(n12261) );
  BUF_X1 U11555 ( .A(n11800), .Z(n12446) );
  AND2_X1 U11556 ( .A1(n13794), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12475) );
  OR2_X1 U11557 ( .A1(n11834), .A2(n11833), .ZN(n12686) );
  NAND2_X1 U11558 ( .A1(n10710), .A2(n10368), .ZN(n10076) );
  AND2_X1 U11559 ( .A1(n11367), .A2(n19970), .ZN(n11547) );
  AND2_X1 U11560 ( .A1(n18268), .A2(n17333), .ZN(n11250) );
  NAND2_X1 U11561 ( .A1(n13777), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12461) );
  NAND2_X1 U11562 ( .A1(n20168), .A2(n12697), .ZN(n12704) );
  OR2_X1 U11563 ( .A1(n12524), .A2(n20715), .ZN(n12434) );
  INV_X1 U11564 ( .A(n12076), .ZN(n12464) );
  INV_X1 U11565 ( .A(n13288), .ZN(n10059) );
  BUF_X1 U11566 ( .A(n11706), .Z(n13007) );
  NAND2_X1 U11567 ( .A1(n10204), .A2(n10202), .ZN(n11853) );
  NOR2_X1 U11568 ( .A1(n11838), .A2(n10203), .ZN(n10202) );
  INV_X1 U11569 ( .A(n11821), .ZN(n10203) );
  AOI21_X1 U11570 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19935), .A(
        n10527), .ZN(n10530) );
  INV_X1 U11571 ( .A(n15183), .ZN(n10090) );
  INV_X1 U11572 ( .A(n10147), .ZN(n10146) );
  OAI21_X1 U11573 ( .B1(n10148), .B2(n10150), .A(n13034), .ZN(n10147) );
  INV_X1 U11574 ( .A(n12995), .ZN(n10148) );
  INV_X1 U11575 ( .A(n13432), .ZN(n10135) );
  INV_X2 U11576 ( .A(n13570), .ZN(n10372) );
  INV_X1 U11577 ( .A(n16307), .ZN(n10095) );
  OAI21_X1 U11578 ( .B1(n13053), .B2(n13052), .A(n9865), .ZN(n10131) );
  INV_X1 U11579 ( .A(n16945), .ZN(n11014) );
  NAND2_X1 U11580 ( .A1(n11120), .A2(n11297), .ZN(n11121) );
  INV_X1 U11581 ( .A(n12529), .ZN(n12530) );
  OR2_X1 U11582 ( .A1(n12521), .A2(n12520), .ZN(n14388) );
  INV_X1 U11583 ( .A(n19992), .ZN(n14397) );
  INV_X1 U11584 ( .A(n12434), .ZN(n12635) );
  INV_X1 U11585 ( .A(n12659), .ZN(n14394) );
  XNOR2_X1 U11587 ( .A(n14023), .B(n13924), .ZN(n15056) );
  INV_X1 U11588 ( .A(n15698), .ZN(n13048) );
  NOR3_X1 U11589 ( .A1(n9899), .A2(n10157), .A3(n10156), .ZN(n10155) );
  INV_X1 U11590 ( .A(n11542), .ZN(n10157) );
  INV_X1 U11591 ( .A(n15246), .ZN(n10156) );
  NOR2_X1 U11592 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  NAND2_X1 U11593 ( .A1(n13995), .A2(n9896), .ZN(n14035) );
  NAND2_X1 U11594 ( .A1(n15310), .A2(n14051), .ZN(n14040) );
  NAND2_X1 U11595 ( .A1(n9997), .A2(n13961), .ZN(n13921) );
  NOR2_X1 U11596 ( .A1(n9991), .A2(n10940), .ZN(n9990) );
  INV_X1 U11597 ( .A(n10937), .ZN(n9991) );
  AND2_X1 U11598 ( .A1(n11358), .A2(n12969), .ZN(n11585) );
  AOI21_X1 U11599 ( .B1(n13712), .B2(n13141), .A(n12993), .ZN(n13046) );
  NOR2_X1 U11600 ( .A1(n13839), .A2(n15791), .ZN(n15886) );
  NOR3_X1 U11601 ( .A1(n13837), .A2(n17333), .A3(n13836), .ZN(n13839) );
  INV_X1 U11602 ( .A(n11256), .ZN(n9909) );
  INV_X1 U11603 ( .A(n11119), .ZN(n9932) );
  INV_X1 U11604 ( .A(n17852), .ZN(n9931) );
  INV_X1 U11605 ( .A(n18272), .ZN(n18933) );
  NAND2_X1 U11606 ( .A1(n17774), .A2(n17787), .ZN(n17761) );
  NOR2_X1 U11607 ( .A1(n18291), .A2(n15807), .ZN(n15806) );
  NOR2_X1 U11608 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16945) );
  OR2_X1 U11609 ( .A1(n20878), .A2(n12650), .ZN(n20079) );
  NAND2_X1 U11610 ( .A1(n19999), .A2(n12681), .ZN(n14805) );
  NAND2_X1 U11611 ( .A1(n11961), .A2(n11960), .ZN(n11971) );
  NAND2_X1 U11612 ( .A1(n9919), .A2(n11994), .ZN(n12016) );
  INV_X1 U11613 ( .A(n11993), .ZN(n9919) );
  AND2_X1 U11614 ( .A1(n12006), .A2(n12005), .ZN(n12017) );
  AND2_X1 U11615 ( .A1(n11759), .A2(n11753), .ZN(n11706) );
  AOI22_X1 U11616 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11897), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U11617 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11801), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11670) );
  OR2_X1 U11618 ( .A1(n11908), .A2(n11907), .ZN(n12724) );
  AND2_X1 U11619 ( .A1(n10009), .A2(n10008), .ZN(n10007) );
  NOR2_X1 U11620 ( .A1(n19970), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11372) );
  NAND2_X1 U11621 ( .A1(n11245), .A2(n17333), .ZN(n11251) );
  INV_X1 U11622 ( .A(n11778), .ZN(n11783) );
  INV_X1 U11623 ( .A(n11754), .ZN(n11761) );
  AND2_X1 U11624 ( .A1(n14422), .A2(n10225), .ZN(n10224) );
  AND2_X1 U11625 ( .A1(n12372), .A2(n10226), .ZN(n10225) );
  INV_X1 U11626 ( .A(n14439), .ZN(n10226) );
  NOR2_X1 U11627 ( .A1(n14568), .A2(n10218), .ZN(n10217) );
  INV_X1 U11628 ( .A(n14479), .ZN(n10218) );
  NAND2_X1 U11629 ( .A1(n12189), .A2(n10213), .ZN(n10212) );
  INV_X1 U11630 ( .A(n14595), .ZN(n10213) );
  NOR2_X1 U11631 ( .A1(n14820), .A2(n10072), .ZN(n9921) );
  INV_X1 U11632 ( .A(n12768), .ZN(n9922) );
  INV_X1 U11633 ( .A(n12765), .ZN(n10072) );
  NAND2_X1 U11634 ( .A1(n9894), .A2(n9834), .ZN(n10221) );
  XNOR2_X1 U11635 ( .A(n12757), .B(n12021), .ZN(n12750) );
  INV_X1 U11636 ( .A(n11929), .ZN(n10208) );
  AOI21_X1 U11637 ( .B1(n11929), .B2(n10207), .A(n10206), .ZN(n10205) );
  OAI21_X1 U11638 ( .B1(n12689), .B2(n20238), .A(n9846), .ZN(n12695) );
  AND2_X1 U11639 ( .A1(n12687), .A2(n11753), .ZN(n9914) );
  OR2_X1 U11640 ( .A1(n12688), .A2(n20874), .ZN(n9915) );
  AND2_X1 U11641 ( .A1(n12529), .A2(n12659), .ZN(n12603) );
  AND2_X1 U11642 ( .A1(n12655), .A2(n12659), .ZN(n12615) );
  NAND2_X1 U11643 ( .A1(n10176), .A2(n14526), .ZN(n10175) );
  INV_X1 U11644 ( .A(n10177), .ZN(n10176) );
  OR2_X1 U11645 ( .A1(n12659), .A2(n12568), .ZN(n12590) );
  INV_X1 U11646 ( .A(n12603), .ZN(n12623) );
  INV_X1 U11647 ( .A(n12746), .ZN(n12758) );
  INV_X1 U11648 ( .A(n12742), .ZN(n10067) );
  INV_X1 U11649 ( .A(n12740), .ZN(n10062) );
  INV_X1 U11650 ( .A(n16023), .ZN(n10063) );
  NAND2_X1 U11651 ( .A1(n11758), .A2(n11753), .ZN(n12754) );
  OR2_X1 U11652 ( .A1(n12755), .A2(n12758), .ZN(n11821) );
  INV_X1 U11653 ( .A(n12686), .ZN(n11851) );
  NAND2_X1 U11654 ( .A1(n20249), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12755) );
  OAI21_X1 U11655 ( .B1(n11930), .B2(n12689), .A(n11853), .ZN(n11925) );
  NAND2_X1 U11656 ( .A1(n11866), .A2(n11865), .ZN(n11892) );
  INV_X1 U11657 ( .A(n13228), .ZN(n15844) );
  NAND2_X1 U11658 ( .A1(n10877), .A2(n15213), .ZN(n10885) );
  INV_X1 U11659 ( .A(n13969), .ZN(n10014) );
  AND2_X1 U11660 ( .A1(n14064), .A2(n15210), .ZN(n10099) );
  INV_X1 U11661 ( .A(n13644), .ZN(n10144) );
  INV_X1 U11662 ( .A(n13036), .ZN(n14288) );
  NOR2_X1 U11663 ( .A1(n9925), .A2(n9924), .ZN(n9923) );
  INV_X1 U11664 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U11665 ( .A1(n10621), .A2(n10601), .ZN(n10603) );
  INV_X1 U11666 ( .A(n13920), .ZN(n9996) );
  INV_X1 U11667 ( .A(n15317), .ZN(n9988) );
  AND2_X1 U11668 ( .A1(n10154), .A2(n10153), .ZN(n10152) );
  INV_X1 U11669 ( .A(n15106), .ZN(n10153) );
  NAND2_X1 U11670 ( .A1(n10451), .A2(n10023), .ZN(n10022) );
  INV_X1 U11671 ( .A(n13389), .ZN(n10023) );
  INV_X1 U11672 ( .A(n10868), .ZN(n9985) );
  AND2_X1 U11673 ( .A1(n9848), .A2(n9987), .ZN(n9986) );
  INV_X1 U11674 ( .A(n15631), .ZN(n9987) );
  OR2_X1 U11675 ( .A1(n19078), .A2(n10959), .ZN(n10875) );
  INV_X1 U11676 ( .A(n13325), .ZN(n10451) );
  INV_X1 U11677 ( .A(n10094), .ZN(n10093) );
  NAND2_X1 U11678 ( .A1(n10989), .A2(n10931), .ZN(n10994) );
  INV_X1 U11679 ( .A(n10990), .ZN(n10989) );
  NAND2_X1 U11680 ( .A1(n9975), .A2(n10971), .ZN(n10973) );
  INV_X1 U11681 ( .A(n13438), .ZN(n9976) );
  BUF_X1 U11682 ( .A(n10400), .Z(n15728) );
  NAND2_X1 U11683 ( .A1(n10086), .A2(n13042), .ZN(n13043) );
  NAND2_X1 U11684 ( .A1(n13148), .A2(n13147), .ZN(n13150) );
  AND2_X1 U11685 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13149) );
  NAND2_X1 U11686 ( .A1(n13150), .A2(n13149), .ZN(n13186) );
  NAND2_X1 U11687 ( .A1(n10129), .A2(n10127), .ZN(n10345) );
  AND2_X1 U11688 ( .A1(n13712), .A2(n10073), .ZN(n10636) );
  NAND2_X1 U11689 ( .A1(n10620), .A2(n10619), .ZN(n9972) );
  NOR2_X1 U11690 ( .A1(n19976), .A2(n19204), .ZN(n16388) );
  AOI21_X1 U11691 ( .B1(n17231), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n11103), .ZN(n11104) );
  NOR2_X1 U11692 ( .A1(n17151), .A2(n18304), .ZN(n11103) );
  NAND2_X1 U11693 ( .A1(n17577), .A2(n9835), .ZN(n11270) );
  NOR2_X1 U11694 ( .A1(n17417), .A2(n11115), .ZN(n11120) );
  XNOR2_X1 U11695 ( .A(n17433), .B(n17430), .ZN(n11110) );
  NAND2_X1 U11696 ( .A1(n13284), .A2(n13283), .ZN(n13320) );
  AND2_X1 U11697 ( .A1(n13171), .A2(n13170), .ZN(n13284) );
  INV_X1 U11698 ( .A(n11773), .ZN(n14395) );
  AND2_X1 U11699 ( .A1(n20715), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12634) );
  NOR2_X2 U11700 ( .A1(n12465), .A2(n12466), .ZN(n12637) );
  AND2_X1 U11701 ( .A1(n14720), .A2(n12076), .ZN(n12436) );
  AND2_X1 U11702 ( .A1(n14560), .A2(n10215), .ZN(n10214) );
  AND2_X1 U11703 ( .A1(n12224), .A2(n12223), .ZN(n14588) );
  CLKBUF_X1 U11704 ( .A(n13448), .Z(n13449) );
  NOR2_X1 U11705 ( .A1(n12522), .A2(n12999), .ZN(n14385) );
  NAND2_X1 U11706 ( .A1(n10060), .A2(n10057), .ZN(n20154) );
  AND2_X1 U11707 ( .A1(n10058), .A2(n20155), .ZN(n10057) );
  NAND2_X1 U11708 ( .A1(n10056), .A2(n12714), .ZN(n10060) );
  NAND2_X1 U11709 ( .A1(n13791), .A2(n13790), .ZN(n13832) );
  OAI211_X1 U11710 ( .C1(n12493), .C2(n13417), .A(n11820), .B(n11819), .ZN(
        n11935) );
  AND2_X1 U11711 ( .A1(n9913), .A2(n9912), .ZN(n9910) );
  AND2_X1 U11712 ( .A1(n20481), .A2(n20367), .ZN(n20449) );
  OAI22_X2 U11713 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15014), .B1(n15864), 
        .B2(n20875), .ZN(n20269) );
  NOR2_X1 U11714 ( .A1(n20370), .A2(n20538), .ZN(n20681) );
  NAND2_X1 U11715 ( .A1(n9817), .A2(n13403), .ZN(n20448) );
  INV_X2 U11716 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20715) );
  INV_X1 U11717 ( .A(n14388), .ZN(n15862) );
  OAI22_X1 U11718 ( .A1(n19964), .A2(n10590), .B1(n11584), .B2(n19961), .ZN(
        n11354) );
  NAND2_X1 U11719 ( .A1(n10888), .A2(n10887), .ZN(n10905) );
  AND2_X1 U11720 ( .A1(n14050), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9928) );
  AND3_X1 U11721 ( .A1(n11473), .A2(n11472), .A3(n11471), .ZN(n15617) );
  AND2_X1 U11722 ( .A1(n13393), .A2(n13391), .ZN(n13466) );
  OR2_X1 U11723 ( .A1(n15128), .A2(n10102), .ZN(n10101) );
  NAND2_X1 U11724 ( .A1(n14290), .A2(n14291), .ZN(n14292) );
  AND2_X1 U11725 ( .A1(n9893), .A2(n10088), .ZN(n10087) );
  INV_X1 U11726 ( .A(n15175), .ZN(n10088) );
  AND2_X1 U11727 ( .A1(n11609), .A2(n11611), .ZN(n15501) );
  NOR2_X1 U11728 ( .A1(n13157), .A2(n16324), .ZN(n13275) );
  NAND2_X1 U11729 ( .A1(n10136), .A2(n9861), .ZN(n10134) );
  INV_X1 U11730 ( .A(n11391), .ZN(n10136) );
  INV_X1 U11731 ( .A(n18965), .ZN(n12969) );
  OR2_X1 U11732 ( .A1(n16398), .A2(n12858), .ZN(n13539) );
  NOR2_X1 U11733 ( .A1(n13981), .A2(n10596), .ZN(n15050) );
  NAND2_X1 U11734 ( .A1(n9929), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13981) );
  NOR2_X1 U11735 ( .A1(n15045), .A2(n15321), .ZN(n15046) );
  AOI21_X1 U11736 ( .B1(n10191), .B2(n10189), .A(n10188), .ZN(n10187) );
  INV_X1 U11737 ( .A(n10191), .ZN(n10190) );
  INV_X1 U11738 ( .A(n11591), .ZN(n10188) );
  NOR2_X1 U11739 ( .A1(n15027), .A2(n16298), .ZN(n15026) );
  NAND2_X1 U11740 ( .A1(n10441), .A2(n10440), .ZN(n13263) );
  INV_X1 U11741 ( .A(n13183), .ZN(n10440) );
  NOR2_X1 U11742 ( .A1(n9855), .A2(n14018), .ZN(n14019) );
  AND2_X1 U11743 ( .A1(n10952), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15319) );
  OR3_X1 U11744 ( .A1(n16227), .A2(n10959), .A3(n20965), .ZN(n10937) );
  XNOR2_X1 U11745 ( .A(n10936), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15484) );
  NAND2_X1 U11746 ( .A1(n13418), .A2(n10151), .ZN(n15289) );
  AND2_X1 U11747 ( .A1(n10152), .A2(n15290), .ZN(n10151) );
  NOR2_X1 U11748 ( .A1(n15217), .A2(n10029), .ZN(n15206) );
  NAND2_X1 U11749 ( .A1(n10030), .A2(n10472), .ZN(n10029) );
  INV_X1 U11750 ( .A(n10032), .ZN(n10030) );
  AND2_X1 U11751 ( .A1(n15366), .A2(n15367), .ZN(n15370) );
  NAND2_X1 U11752 ( .A1(n10200), .A2(n15425), .ZN(n15416) );
  NAND2_X1 U11753 ( .A1(n13458), .A2(n13464), .ZN(n15217) );
  AND2_X1 U11754 ( .A1(n10856), .A2(n10195), .ZN(n10194) );
  INV_X1 U11755 ( .A(n15646), .ZN(n10195) );
  AND2_X1 U11756 ( .A1(n11407), .A2(n11406), .ZN(n12995) );
  AND2_X1 U11757 ( .A1(n11568), .A2(n16358), .ZN(n19298) );
  AND2_X1 U11758 ( .A1(n12973), .A2(n12974), .ZN(n11381) );
  NAND2_X1 U11759 ( .A1(n10614), .A2(n10613), .ZN(n10074) );
  NOR2_X1 U11760 ( .A1(n11391), .A2(n10133), .ZN(n10132) );
  INV_X1 U11761 ( .A(n13349), .ZN(n10133) );
  NAND2_X1 U11762 ( .A1(n13050), .A2(n13049), .ZN(n13138) );
  INV_X1 U11764 ( .A(n10721), .ZN(n19546) );
  OR2_X1 U11765 ( .A1(n19565), .A2(n19598), .ZN(n19540) );
  NOR2_X2 U11766 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19924) );
  OR2_X1 U11767 ( .A1(n19354), .A2(n15124), .ZN(n19697) );
  OR2_X1 U11768 ( .A1(n19938), .A2(n19944), .ZN(n19696) );
  NAND2_X1 U11769 ( .A1(n10255), .A2(n16379), .ZN(n10262) );
  NAND2_X1 U11770 ( .A1(n10260), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10261) );
  OR2_X1 U11771 ( .A1(n19938), .A2(n13715), .ZN(n19719) );
  OR2_X1 U11772 ( .A1(n19354), .A2(n19955), .ZN(n19720) );
  INV_X1 U11773 ( .A(n19719), .ZN(n19781) );
  NAND2_X1 U11774 ( .A1(n11335), .A2(n11333), .ZN(n16402) );
  NOR2_X1 U11775 ( .A1(n9815), .A2(n11247), .ZN(n15789) );
  OAI21_X1 U11776 ( .B1(n11262), .B2(n11261), .A(n11260), .ZN(n18725) );
  NAND2_X1 U11777 ( .A1(n9959), .A2(n9958), .ZN(n9960) );
  AOI21_X1 U11778 ( .B1(n9952), .B2(n17566), .A(n16633), .ZN(n9958) );
  NAND2_X1 U11779 ( .A1(n16642), .A2(n9952), .ZN(n9959) );
  OR2_X1 U11780 ( .A1(n16642), .A2(n17566), .ZN(n9961) );
  NAND2_X1 U11781 ( .A1(n9955), .A2(n9954), .ZN(n9956) );
  AOI21_X1 U11782 ( .B1(n9952), .B2(n17602), .A(n17590), .ZN(n9954) );
  NAND2_X1 U11783 ( .A1(n16665), .A2(n9952), .ZN(n9955) );
  OR2_X1 U11784 ( .A1(n16665), .A2(n17602), .ZN(n9957) );
  OR2_X1 U11785 ( .A1(n9952), .A2(n17638), .ZN(n9951) );
  OR2_X1 U11786 ( .A1(n16695), .A2(n9886), .ZN(n9950) );
  OR2_X1 U11787 ( .A1(n16695), .A2(n16696), .ZN(n9953) );
  NAND2_X1 U11788 ( .A1(n11192), .A2(n10046), .ZN(n10045) );
  AOI21_X1 U11789 ( .B1(n17230), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n10047), .ZN(n10046) );
  NOR2_X1 U11790 ( .A1(n9811), .A2(n18618), .ZN(n10047) );
  NOR3_X1 U11791 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18916), .ZN(n11006) );
  OR2_X1 U11792 ( .A1(n10055), .A2(n11064), .ZN(n10054) );
  NOR2_X1 U11793 ( .A1(n10244), .A2(n20981), .ZN(n9934) );
  INV_X1 U11794 ( .A(n11062), .ZN(n9935) );
  NOR2_X1 U11795 ( .A1(n11270), .A2(n17910), .ZN(n16445) );
  NAND2_X1 U11796 ( .A1(n17705), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17673) );
  INV_X1 U11797 ( .A(n17748), .ZN(n9945) );
  NOR2_X1 U11798 ( .A1(n17777), .A2(n17847), .ZN(n17817) );
  NAND2_X1 U11799 ( .A1(n17862), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17777) );
  AND2_X1 U11800 ( .A1(n11125), .A2(n10051), .ZN(n10050) );
  NOR2_X1 U11801 ( .A1(n17820), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10051) );
  XNOR2_X1 U11802 ( .A(n11118), .B(n11116), .ZN(n17858) );
  NAND2_X1 U11803 ( .A1(n17858), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17857) );
  XNOR2_X1 U11804 ( .A(n17433), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17906) );
  AOI211_X2 U11805 ( .C1(n17195), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n11203), .B(n11202), .ZN(n18268) );
  NAND2_X1 U11806 ( .A1(n18113), .A2(n10038), .ZN(n10037) );
  INV_X1 U11807 ( .A(n18730), .ZN(n10038) );
  NAND2_X1 U11808 ( .A1(n18796), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18784) );
  NAND2_X1 U11809 ( .A1(n13669), .A2(n12662), .ZN(n20080) );
  INV_X1 U11810 ( .A(n20080), .ZN(n20084) );
  AND2_X1 U11811 ( .A1(n20079), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20087) );
  NAND2_X1 U11812 ( .A1(n13669), .A2(n12668), .ZN(n20043) );
  NAND2_X1 U11813 ( .A1(n13669), .A2(n12660), .ZN(n20098) );
  XNOR2_X1 U11814 ( .A(n12653), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13498) );
  NOR2_X1 U11815 ( .A1(n12652), .A2(n14401), .ZN(n12653) );
  INV_X1 U11816 ( .A(n14805), .ZN(n20165) );
  AND2_X1 U11817 ( .A1(n14805), .A2(n12683), .ZN(n20171) );
  XNOR2_X1 U11818 ( .A(n12658), .B(n12657), .ZN(n14546) );
  MUX2_X1 U11819 ( .A(n12656), .B(n12655), .S(n14410), .Z(n12658) );
  XNOR2_X1 U11820 ( .A(n12788), .B(n12787), .ZN(n13959) );
  CLKBUF_X1 U11822 ( .A(n13097), .Z(n20612) );
  INV_X1 U11823 ( .A(n19924), .ZN(n19722) );
  NAND2_X1 U11824 ( .A1(n10142), .A2(n10140), .ZN(n10139) );
  NOR2_X1 U11825 ( .A1(n15055), .A2(n10141), .ZN(n10140) );
  NAND2_X1 U11826 ( .A1(n15056), .A2(n19129), .ZN(n10142) );
  NOR2_X1 U11827 ( .A1(n19158), .A2(n15053), .ZN(n10141) );
  NAND2_X1 U11828 ( .A1(n16179), .A2(n19075), .ZN(n15051) );
  NAND2_X1 U11829 ( .A1(n15051), .A2(n15299), .ZN(n16174) );
  NAND2_X1 U11830 ( .A1(n16180), .A2(n16181), .ZN(n16179) );
  NAND2_X1 U11831 ( .A1(n13941), .A2(n14047), .ZN(n15054) );
  AND2_X1 U11832 ( .A1(n19288), .A2(n19942), .ZN(n19278) );
  INV_X1 U11833 ( .A(n16292), .ZN(n19276) );
  XNOR2_X1 U11834 ( .A(n14047), .B(n14046), .ZN(n19161) );
  NOR2_X1 U11835 ( .A1(n14055), .A2(n14054), .ZN(n14056) );
  XNOR2_X1 U11836 ( .A(n9978), .B(n14050), .ZN(n14058) );
  XNOR2_X1 U11837 ( .A(n14035), .B(n14034), .ZN(n16171) );
  NAND2_X1 U11838 ( .A1(n13921), .A2(n13920), .ZN(n14021) );
  NAND2_X1 U11839 ( .A1(n11579), .A2(n11578), .ZN(n11580) );
  INV_X1 U11840 ( .A(n11567), .ZN(n11579) );
  OR2_X1 U11841 ( .A1(n9880), .A2(n16337), .ZN(n10114) );
  NAND2_X1 U11842 ( .A1(n10122), .A2(n10111), .ZN(n10110) );
  NAND2_X1 U11843 ( .A1(n10118), .A2(n10120), .ZN(n10111) );
  INV_X1 U11844 ( .A(n10123), .ZN(n10122) );
  NAND2_X1 U11845 ( .A1(n15561), .A2(n10121), .ZN(n10120) );
  AOI21_X1 U11846 ( .B1(n15561), .B2(n10119), .A(n10125), .ZN(n10118) );
  NOR2_X1 U11847 ( .A1(n15563), .A2(n9889), .ZN(n10119) );
  OR2_X1 U11848 ( .A1(n15556), .A2(n9880), .ZN(n10115) );
  AOI21_X1 U11849 ( .B1(n15558), .B2(n9889), .A(n10117), .ZN(n10116) );
  INV_X1 U11850 ( .A(n15561), .ZN(n10117) );
  NAND2_X1 U11851 ( .A1(n10193), .A2(n15403), .ZN(n15394) );
  NAND2_X1 U11852 ( .A1(n11589), .A2(n15402), .ZN(n10193) );
  AND2_X1 U11853 ( .A1(n11585), .A2(n19962), .ZN(n16337) );
  INV_X1 U11854 ( .A(n19296), .ZN(n16339) );
  AND2_X1 U11855 ( .A1(n11585), .A2(n11363), .ZN(n19301) );
  AND2_X1 U11856 ( .A1(n11585), .A2(n19963), .ZN(n19303) );
  OR2_X1 U11857 ( .A1(n19289), .A2(n15559), .ZN(n16364) );
  INV_X1 U11858 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19935) );
  INV_X1 U11859 ( .A(n19676), .ZN(n19681) );
  INV_X1 U11860 ( .A(n16617), .ZN(n9966) );
  NOR2_X1 U11861 ( .A1(n16616), .A2(n9964), .ZN(n9963) );
  NAND2_X1 U11862 ( .A1(n16619), .A2(n9965), .ZN(n9964) );
  OR2_X1 U11863 ( .A1(n16628), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9965) );
  INV_X1 U11864 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17252) );
  INV_X1 U11865 ( .A(n17284), .ZN(n13841) );
  OR2_X1 U11866 ( .A1(n17372), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U11867 ( .A1(n17294), .A2(n17438), .ZN(n17292) );
  NAND2_X1 U11868 ( .A1(n17333), .A2(n17429), .ZN(n17438) );
  INV_X1 U11869 ( .A(n10040), .ZN(n10039) );
  AOI21_X1 U11870 ( .B1(n17667), .B2(n16913), .A(n16461), .ZN(n10041) );
  NAND2_X1 U11871 ( .A1(n11273), .A2(n11269), .ZN(n10043) );
  NAND2_X1 U11872 ( .A1(n17410), .A2(n11274), .ZN(n17753) );
  NAND2_X1 U11873 ( .A1(n17916), .A2(n17816), .ZN(n17911) );
  OAI22_X1 U11874 ( .A1(n11143), .A2(n11142), .B1(n11141), .B2(n11140), .ZN(
        n16469) );
  INV_X1 U11875 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10201) );
  CLKBUF_X1 U11876 ( .A(n14159), .Z(n14275) );
  XNOR2_X1 U11877 ( .A(n10372), .B(n10768), .ZN(n11346) );
  NAND2_X1 U11878 ( .A1(n11972), .A2(n11971), .ZN(n11993) );
  INV_X1 U11879 ( .A(n11948), .ZN(n10206) );
  OR2_X1 U11880 ( .A1(n11959), .A2(n11958), .ZN(n12725) );
  NAND2_X1 U11881 ( .A1(n13179), .A2(n12679), .ZN(n13006) );
  AND2_X2 U11882 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U11883 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11801), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11702) );
  XNOR2_X1 U11884 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10520) );
  AND2_X1 U11885 ( .A1(n10519), .A2(n10520), .ZN(n10527) );
  OAI211_X1 U11886 ( .C1(n9809), .C2(n10357), .A(n10356), .B(n10355), .ZN(
        n10385) );
  NAND4_X1 U11887 ( .A1(n19340), .A2(n13570), .A3(n10942), .A4(n10354), .ZN(
        n11545) );
  AND2_X1 U11888 ( .A1(n10543), .A2(n16379), .ZN(n10679) );
  AOI21_X1 U11889 ( .B1(n14031), .B2(P2_EBX_REG_0__SCAN_IN), .A(n9866), .ZN(
        n10389) );
  NAND2_X1 U11890 ( .A1(n11114), .A2(n11280), .ZN(n11115) );
  INV_X1 U11891 ( .A(n15802), .ZN(n11241) );
  NOR2_X1 U11892 ( .A1(n16582), .A2(n11255), .ZN(n15783) );
  NAND2_X1 U11893 ( .A1(n12755), .A2(n11896), .ZN(n12518) );
  NOR2_X1 U11894 ( .A1(n14466), .A2(n10216), .ZN(n10215) );
  INV_X1 U11895 ( .A(n10217), .ZN(n10216) );
  NOR2_X1 U11896 ( .A1(n12238), .A2(n15934), .ZN(n12239) );
  INV_X1 U11897 ( .A(n12461), .ZN(n12431) );
  NAND2_X1 U11898 ( .A1(n14610), .A2(n10220), .ZN(n10219) );
  INV_X1 U11899 ( .A(n10221), .ZN(n10220) );
  INV_X1 U11900 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12117) );
  INV_X1 U11901 ( .A(n13716), .ZN(n10222) );
  INV_X1 U11902 ( .A(n13127), .ZN(n11947) );
  AND2_X1 U11903 ( .A1(n9891), .A2(n10182), .ZN(n10181) );
  INV_X1 U11904 ( .A(n14447), .ZN(n10182) );
  NAND2_X1 U11905 ( .A1(n10168), .A2(n12602), .ZN(n10167) );
  NOR2_X1 U11906 ( .A1(n14589), .A2(n10169), .ZN(n10168) );
  INV_X1 U11907 ( .A(n14580), .ZN(n10169) );
  NAND2_X1 U11908 ( .A1(n10178), .A2(n14622), .ZN(n10177) );
  INV_X1 U11909 ( .A(n13773), .ZN(n10178) );
  OR2_X1 U11910 ( .A1(n12004), .A2(n12003), .ZN(n12744) );
  INV_X1 U11911 ( .A(n13320), .ZN(n10164) );
  NAND2_X1 U11913 ( .A1(n11764), .A2(n13786), .ZN(n9913) );
  XNOR2_X1 U11914 ( .A(n11845), .B(n11844), .ZN(n20334) );
  AND4_X2 U11915 ( .A1(n11643), .A2(n11642), .A3(n9845), .A4(n11641), .ZN(
        n11754) );
  INV_X1 U11916 ( .A(n12694), .ZN(n13403) );
  NAND2_X1 U11917 ( .A1(n10001), .A2(n10876), .ZN(n10899) );
  INV_X1 U11918 ( .A(n10893), .ZN(n10001) );
  NAND2_X1 U11919 ( .A1(n10007), .A2(n10449), .ZN(n10006) );
  INV_X1 U11920 ( .A(n10007), .ZN(n10005) );
  OR2_X1 U11921 ( .A1(n10829), .A2(n10828), .ZN(n10839) );
  INV_X1 U11922 ( .A(n10774), .ZN(n10783) );
  MUX2_X1 U11923 ( .A(n10771), .B(n10407), .S(n14024), .Z(n10787) );
  NAND2_X1 U11924 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19958), .ZN(
        n10531) );
  BUF_X1 U11925 ( .A(n10550), .Z(n14359) );
  NOR2_X1 U11926 ( .A1(n15128), .A2(n10105), .ZN(n10104) );
  INV_X1 U11927 ( .A(n10107), .ZN(n10105) );
  INV_X1 U11928 ( .A(n15132), .ZN(n10102) );
  NAND2_X1 U11929 ( .A1(n10098), .A2(n15156), .ZN(n10096) );
  OR2_X1 U11930 ( .A1(n14179), .A2(n14207), .ZN(n10097) );
  NOR2_X1 U11931 ( .A1(n10744), .A2(n10743), .ZN(n11403) );
  NOR2_X1 U11932 ( .A1(n15393), .A2(n10192), .ZN(n10191) );
  INV_X1 U11933 ( .A(n15403), .ZN(n10192) );
  INV_X1 U11934 ( .A(n15402), .ZN(n10189) );
  INV_X1 U11935 ( .A(n10979), .ZN(n10980) );
  NOR2_X1 U11936 ( .A1(n10013), .A2(n10015), .ZN(n10011) );
  AND4_X1 U11937 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10767) );
  NAND2_X1 U11938 ( .A1(n10949), .A2(n10948), .ZN(n13961) );
  AND2_X1 U11939 ( .A1(n11532), .A2(n11531), .ZN(n15254) );
  NAND2_X1 U11940 ( .A1(n11605), .A2(n9895), .ZN(n10028) );
  INV_X1 U11941 ( .A(n15165), .ZN(n10024) );
  NOR2_X1 U11942 ( .A1(n10026), .A2(n15170), .ZN(n10025) );
  INV_X1 U11943 ( .A(n11606), .ZN(n10026) );
  NAND2_X1 U11944 ( .A1(n10464), .A2(n10033), .ZN(n10032) );
  INV_X1 U11945 ( .A(n15100), .ZN(n10033) );
  AND2_X1 U11946 ( .A1(n11513), .A2(n11512), .ZN(n15106) );
  AND2_X1 U11947 ( .A1(n15585), .A2(n13503), .ZN(n10154) );
  NOR2_X1 U11948 ( .A1(n15636), .A2(n16278), .ZN(n10126) );
  NAND2_X1 U11949 ( .A1(n13309), .A2(n10018), .ZN(n10017) );
  INV_X1 U11950 ( .A(n14031), .ZN(n10507) );
  NAND2_X1 U11951 ( .A1(n10781), .A2(n10780), .ZN(n9977) );
  NAND2_X1 U11952 ( .A1(n10328), .A2(n10540), .ZN(n9971) );
  NAND2_X1 U11953 ( .A1(n11546), .A2(n10342), .ZN(n10350) );
  AND2_X1 U11954 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13044) );
  NAND2_X1 U11955 ( .A1(n13043), .A2(n13044), .ZN(n13137) );
  NAND2_X1 U11956 ( .A1(n10338), .A2(n16379), .ZN(n10339) );
  AND4_X1 U11957 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n10295) );
  NAND3_X1 U11958 ( .A1(n19924), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19777), 
        .ZN(n13514) );
  INV_X1 U11959 ( .A(n11330), .ZN(n11335) );
  AOI21_X1 U11960 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18261), .A(
        n11161), .ZN(n11260) );
  NOR3_X1 U11961 ( .A1(n18916), .A2(n9798), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11015) );
  OR2_X1 U11962 ( .A1(n11248), .A2(n18734), .ZN(n13837) );
  NOR2_X1 U11963 ( .A1(n11251), .A2(n9796), .ZN(n11256) );
  NOR2_X1 U11964 ( .A1(n17554), .A2(n9947), .ZN(n9946) );
  INV_X1 U11965 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9947) );
  OR2_X1 U11966 ( .A1(n11134), .A2(n11133), .ZN(n11135) );
  OAI21_X1 U11967 ( .B1(n17761), .B2(n9901), .A(n11132), .ZN(n11129) );
  NOR2_X1 U11968 ( .A1(n21098), .A2(n9862), .ZN(n15819) );
  AND2_X1 U11969 ( .A1(n17426), .A2(n11284), .ZN(n11114) );
  NOR2_X1 U11970 ( .A1(n11253), .A2(n11252), .ZN(n18733) );
  AND2_X1 U11971 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11234) );
  OR2_X1 U11972 ( .A1(n11014), .A2(n11010), .ZN(n9841) );
  AOI211_X1 U11973 ( .C1(n17216), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n11211), .B(n11210), .ZN(n11212) );
  INV_X1 U11974 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14532) );
  INV_X1 U11975 ( .A(n20031), .ZN(n20062) );
  NOR2_X1 U11976 ( .A1(n9874), .A2(n14467), .ZN(n14565) );
  AND2_X1 U11977 ( .A1(n12593), .A2(n12592), .ZN(n14597) );
  NAND2_X1 U11978 ( .A1(n10164), .A2(n10163), .ZN(n13400) );
  NOR2_X1 U11979 ( .A1(n13339), .A2(n13319), .ZN(n10163) );
  AND2_X1 U11980 ( .A1(n12245), .A2(n12244), .ZN(n14578) );
  OR2_X1 U11981 ( .A1(n15997), .A2(n12464), .ZN(n12244) );
  NAND2_X1 U11982 ( .A1(n14704), .A2(n12801), .ZN(n13425) );
  NOR2_X1 U11983 ( .A1(n12439), .A2(n14718), .ZN(n12651) );
  AND2_X1 U11984 ( .A1(n10224), .A2(n14412), .ZN(n10223) );
  NAND2_X1 U11985 ( .A1(n12367), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12368) );
  INV_X1 U11986 ( .A(n12366), .ZN(n12367) );
  OR2_X1 U11987 ( .A1(n12368), .A2(n14455), .ZN(n12411) );
  NAND2_X1 U11988 ( .A1(n12324), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12326) );
  NAND2_X1 U11989 ( .A1(n12276), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12277) );
  NOR2_X1 U11990 ( .A1(n12277), .A2(n15916), .ZN(n12324) );
  AND2_X1 U11991 ( .A1(n12260), .A2(n12259), .ZN(n14479) );
  AND2_X1 U11992 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n12239), .ZN(
        n12276) );
  OR2_X1 U11993 ( .A1(n10212), .A2(n10210), .ZN(n10209) );
  INV_X1 U11994 ( .A(n14588), .ZN(n10210) );
  NOR2_X1 U11995 ( .A1(n12205), .A2(n14502), .ZN(n12206) );
  NAND2_X1 U11996 ( .A1(n12206), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12238) );
  NAND2_X1 U11997 ( .A1(n10070), .A2(n10069), .ZN(n14815) );
  AND2_X1 U11998 ( .A1(n12169), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12170) );
  OR2_X1 U11999 ( .A1(n12122), .A2(n14532), .ZN(n12123) );
  INV_X1 U12000 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n21036) );
  OR2_X1 U12002 ( .A1(n12118), .A2(n12117), .ZN(n12122) );
  AND2_X1 U12003 ( .A1(n12074), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12075) );
  NAND2_X1 U12004 ( .A1(n12075), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12118) );
  OR2_X1 U12005 ( .A1(n10207), .A2(n12089), .ZN(n14520) );
  OR2_X1 U12006 ( .A1(n12042), .A2(n13736), .ZN(n12057) );
  AND2_X1 U12007 ( .A1(n12041), .A2(n12040), .ZN(n13488) );
  NAND2_X1 U12008 ( .A1(n12022), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12042) );
  AND2_X1 U12009 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n12007), .ZN(
        n12022) );
  INV_X1 U12010 ( .A(n12008), .ZN(n12007) );
  AOI21_X1 U12011 ( .B1(n12733), .B2(n12054), .A(n12013), .ZN(n13399) );
  INV_X1 U12012 ( .A(n11986), .ZN(n11987) );
  NAND2_X1 U12013 ( .A1(n11966), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11986) );
  NOR2_X1 U12014 ( .A1(n11916), .A2(n11915), .ZN(n11966) );
  INV_X1 U12015 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11915) );
  XNOR2_X1 U12016 ( .A(n12704), .B(n20204), .ZN(n13134) );
  NAND2_X1 U12017 ( .A1(n20166), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20168) );
  NAND2_X1 U12018 ( .A1(n14740), .A2(n14888), .ZN(n14721) );
  OR2_X1 U12019 ( .A1(n14421), .A2(n14408), .ZN(n14410) );
  NAND2_X1 U12020 ( .A1(n14436), .A2(n14419), .ZN(n14421) );
  AOI21_X1 U12021 ( .B1(n16013), .B2(n14750), .A(n14770), .ZN(n14729) );
  AND2_X1 U12022 ( .A1(n14565), .A2(n10179), .ZN(n14436) );
  AND2_X1 U12023 ( .A1(n10181), .A2(n10180), .ZN(n10179) );
  INV_X1 U12024 ( .A(n14435), .ZN(n10180) );
  NAND2_X1 U12025 ( .A1(n14565), .A2(n10181), .ZN(n14449) );
  OR2_X1 U12026 ( .A1(n14937), .A2(n13954), .ZN(n14909) );
  AND2_X1 U12027 ( .A1(n14565), .A2(n14564), .ZN(n14562) );
  NAND2_X1 U12028 ( .A1(n14565), .A2(n9891), .ZN(n14556) );
  NOR2_X1 U12029 ( .A1(n9873), .A2(n10166), .ZN(n14582) );
  INV_X1 U12030 ( .A(n10168), .ZN(n10166) );
  NOR2_X1 U12031 ( .A1(n9873), .A2(n14589), .ZN(n14590) );
  AND2_X1 U12033 ( .A1(n12584), .A2(n12583), .ZN(n14602) );
  NOR2_X1 U12034 ( .A1(n14603), .A2(n14602), .ZN(n14604) );
  NAND2_X1 U12035 ( .A1(n10174), .A2(n10173), .ZN(n14512) );
  NOR2_X1 U12036 ( .A1(n10175), .A2(n13827), .ZN(n10173) );
  INV_X1 U12037 ( .A(n13772), .ZN(n10174) );
  OR2_X1 U12038 ( .A1(n14512), .A2(n14511), .ZN(n14603) );
  AND2_X1 U12039 ( .A1(n12573), .A2(n12572), .ZN(n14526) );
  NOR2_X1 U12040 ( .A1(n13772), .A2(n10177), .ZN(n14625) );
  NOR2_X1 U12041 ( .A1(n13772), .A2(n13773), .ZN(n14623) );
  AND3_X1 U12042 ( .A1(n12564), .A2(n12590), .A3(n12563), .ZN(n13720) );
  OR2_X1 U12043 ( .A1(n13721), .A2(n13720), .ZN(n13772) );
  NOR2_X1 U12044 ( .A1(n13320), .A2(n10161), .ZN(n13695) );
  NAND2_X1 U12045 ( .A1(n10162), .A2(n9833), .ZN(n10161) );
  INV_X1 U12046 ( .A(n13339), .ZN(n10162) );
  NAND2_X1 U12047 ( .A1(n10064), .A2(n10065), .ZN(n13734) );
  NAND2_X1 U12048 ( .A1(n10067), .A2(n16023), .ZN(n10066) );
  NAND2_X1 U12049 ( .A1(n19990), .A2(n16155), .ZN(n12680) );
  NAND2_X1 U12050 ( .A1(n20154), .A2(n12722), .ZN(n16036) );
  NAND2_X1 U12051 ( .A1(n10164), .A2(n12546), .ZN(n13338) );
  OR2_X1 U12052 ( .A1(n20845), .A2(n12754), .ZN(n12712) );
  NAND2_X1 U12053 ( .A1(n11840), .A2(n11853), .ZN(n11930) );
  OR2_X1 U12054 ( .A1(n12755), .A2(n11851), .ZN(n11852) );
  INV_X1 U12055 ( .A(n13015), .ZN(n13777) );
  NAND2_X1 U12056 ( .A1(n9920), .A2(n20365), .ZN(n13229) );
  AND2_X1 U12057 ( .A1(n13029), .A2(n13028), .ZN(n15838) );
  OR2_X1 U12058 ( .A1(n9817), .A2(n13403), .ZN(n20607) );
  AND2_X1 U12059 ( .A1(n9817), .A2(n12694), .ZN(n20533) );
  INV_X1 U12060 ( .A(n20580), .ZN(n20584) );
  CLKBUF_X2 U12061 ( .A(n11754), .Z(n20258) );
  AOI21_X1 U12062 ( .B1(n20863), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20370), 
        .ZN(n20722) );
  NOR2_X2 U12063 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20846) );
  INV_X1 U12064 ( .A(n12524), .ZN(n20264) );
  INV_X1 U12065 ( .A(n20236), .ZN(n20267) );
  OR2_X1 U12066 ( .A1(n10538), .A2(n19969), .ZN(n11584) );
  AND2_X1 U12067 ( .A1(n15501), .A2(n15502), .ZN(n15504) );
  NOR2_X1 U12068 ( .A1(n10004), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U12069 ( .A1(n10888), .A2(n10003), .ZN(n10909) );
  NAND2_X1 U12070 ( .A1(n15032), .A2(n9926), .ZN(n15034) );
  NOR2_X1 U12071 ( .A1(n15409), .A2(n9927), .ZN(n9926) );
  INV_X1 U12072 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9927) );
  AND2_X1 U12073 ( .A1(n13995), .A2(n10011), .ZN(n13930) );
  NAND2_X1 U12074 ( .A1(n13995), .A2(n10503), .ZN(n13998) );
  AND2_X1 U12075 ( .A1(n14063), .A2(n14062), .ZN(n14064) );
  AND2_X1 U12076 ( .A1(n13467), .A2(n13466), .ZN(n13469) );
  AND2_X1 U12077 ( .A1(n10108), .A2(n15132), .ZN(n10107) );
  XNOR2_X1 U12078 ( .A(n14233), .B(n14235), .ZN(n15152) );
  NAND2_X1 U12079 ( .A1(n15504), .A2(n15268), .ZN(n15267) );
  OR2_X1 U12080 ( .A1(n14129), .A2(n14128), .ZN(n15179) );
  AND2_X1 U12081 ( .A1(n11523), .A2(n11522), .ZN(n15515) );
  AND2_X1 U12082 ( .A1(n11520), .A2(n11519), .ZN(n15279) );
  OR2_X1 U12083 ( .A1(n14085), .A2(n14084), .ZN(n15204) );
  CLKBUF_X1 U12084 ( .A(n15197), .Z(n15203) );
  AND2_X1 U12085 ( .A1(n9823), .A2(n13158), .ZN(n10143) );
  AND3_X1 U12086 ( .A1(n11420), .A2(n11419), .A3(n11418), .ZN(n13644) );
  AND2_X1 U12087 ( .A1(n10145), .A2(n9823), .ZN(n13643) );
  INV_X1 U12088 ( .A(n11331), .ZN(n19208) );
  NAND2_X1 U12089 ( .A1(n15043), .A2(n9836), .ZN(n15045) );
  NAND2_X1 U12090 ( .A1(n15043), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15044) );
  INV_X1 U12091 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15339) );
  AND2_X1 U12092 ( .A1(n15039), .A2(n10592), .ZN(n15042) );
  NAND2_X1 U12093 ( .A1(n15042), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15041) );
  NOR2_X1 U12094 ( .A1(n15034), .A2(n15398), .ZN(n15037) );
  AND2_X1 U12095 ( .A1(n15037), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15039) );
  NOR2_X1 U12096 ( .A1(n15031), .A2(n15429), .ZN(n15032) );
  NAND2_X1 U12097 ( .A1(n15032), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15036) );
  NOR2_X1 U12098 ( .A1(n15030), .A2(n19085), .ZN(n15029) );
  NAND2_X1 U12099 ( .A1(n15026), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15030) );
  NAND2_X1 U12100 ( .A1(n13639), .A2(n9885), .ZN(n15027) );
  AND2_X1 U12101 ( .A1(n13639), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13637) );
  NAND2_X1 U12102 ( .A1(n13622), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13621) );
  NOR2_X1 U12103 ( .A1(n19287), .A2(n13623), .ZN(n13622) );
  OAI21_X1 U12104 ( .B1(n10607), .B2(n10606), .A(n10605), .ZN(n10611) );
  AND2_X1 U12105 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13443) );
  INV_X1 U12106 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13553) );
  AND2_X1 U12107 ( .A1(n9995), .A2(n10948), .ZN(n9993) );
  NOR2_X1 U12108 ( .A1(n10959), .A2(n14039), .ZN(n10010) );
  OR2_X1 U12109 ( .A1(n13937), .A2(n11543), .ZN(n16177) );
  AOI21_X1 U12110 ( .B1(n10953), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15319), .ZN(n13963) );
  NAND2_X1 U12111 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10083) );
  INV_X1 U12112 ( .A(n13995), .ZN(n15144) );
  NAND2_X1 U12113 ( .A1(n9980), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9979) );
  INV_X1 U12114 ( .A(n10083), .ZN(n9980) );
  NOR2_X1 U12115 ( .A1(n15493), .A2(n15474), .ZN(n15332) );
  NAND2_X1 U12116 ( .A1(n11605), .A2(n10025), .ZN(n15172) );
  OR2_X1 U12117 ( .A1(n18992), .A2(n10959), .ZN(n10882) );
  NAND2_X1 U12118 ( .A1(n15366), .A2(n10197), .ZN(n15347) );
  NOR2_X1 U12119 ( .A1(n10199), .A2(n10198), .ZN(n10197) );
  INV_X1 U12120 ( .A(n15367), .ZN(n10198) );
  INV_X1 U12121 ( .A(n15359), .ZN(n10199) );
  AND2_X1 U12122 ( .A1(n11518), .A2(n11517), .ZN(n15088) );
  INV_X1 U12123 ( .A(n15087), .ZN(n15280) );
  NAND2_X1 U12124 ( .A1(n15206), .A2(n15084), .ZN(n15191) );
  INV_X1 U12125 ( .A(n15563), .ZN(n10121) );
  OAI21_X1 U12126 ( .B1(n15564), .B2(n16369), .A(n10124), .ZN(n10123) );
  AOI21_X1 U12127 ( .B1(n19033), .B2(n16339), .A(n15557), .ZN(n10124) );
  NAND2_X1 U12128 ( .A1(n13418), .A2(n10154), .ZN(n15107) );
  AND2_X1 U12129 ( .A1(n13418), .A2(n15585), .ZN(n15587) );
  NAND2_X1 U12130 ( .A1(n10031), .A2(n10464), .ZN(n15215) );
  INV_X1 U12131 ( .A(n15217), .ZN(n10031) );
  NAND2_X1 U12132 ( .A1(n10020), .A2(n13459), .ZN(n10019) );
  INV_X1 U12133 ( .A(n10022), .ZN(n10020) );
  AND2_X1 U12134 ( .A1(n9983), .A2(n15612), .ZN(n9982) );
  OR2_X1 U12135 ( .A1(n9986), .A2(n9984), .ZN(n9983) );
  OR2_X1 U12136 ( .A1(n15611), .A2(n9985), .ZN(n9984) );
  NAND2_X1 U12137 ( .A1(n10196), .A2(n9986), .ZN(n9981) );
  NAND2_X1 U12138 ( .A1(n10021), .A2(n10451), .ZN(n13324) );
  INV_X1 U12139 ( .A(n13326), .ZN(n10021) );
  NAND2_X1 U12140 ( .A1(n15440), .A2(n10079), .ZN(n10081) );
  NOR2_X1 U12141 ( .A1(n10095), .A2(n10080), .ZN(n10079) );
  INV_X1 U12142 ( .A(n15439), .ZN(n10080) );
  NAND2_X1 U12143 ( .A1(n10093), .A2(n10095), .ZN(n10091) );
  NAND2_X1 U12144 ( .A1(n15658), .A2(n10093), .ZN(n10092) );
  AND2_X1 U12145 ( .A1(n15674), .A2(n11571), .ZN(n16334) );
  NAND2_X1 U12146 ( .A1(n10973), .A2(n10974), .ZN(n13475) );
  AND3_X1 U12147 ( .A1(n11400), .A2(n11399), .A3(n11398), .ZN(n13432) );
  NAND2_X1 U12148 ( .A1(n9977), .A2(n10972), .ZN(n13439) );
  NAND2_X1 U12149 ( .A1(n11361), .A2(n10085), .ZN(n15744) );
  INV_X1 U12150 ( .A(n10363), .ZN(n10085) );
  NAND2_X1 U12151 ( .A1(n11371), .A2(n11370), .ZN(n12973) );
  NAND2_X1 U12152 ( .A1(n10351), .A2(n10400), .ZN(n11359) );
  NAND2_X1 U12153 ( .A1(n10380), .A2(n19970), .ZN(n10351) );
  AND2_X1 U12154 ( .A1(n11585), .A2(n11563), .ZN(n15559) );
  AND2_X1 U12155 ( .A1(n20977), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13141) );
  NAND2_X1 U12156 ( .A1(n12956), .A2(n19951), .ZN(n13146) );
  CLKBUF_X1 U12157 ( .A(n15710), .Z(n15724) );
  CLKBUF_X1 U12158 ( .A(n10380), .Z(n15748) );
  XNOR2_X1 U12159 ( .A(n15698), .B(n13047), .ZN(n13045) );
  OAI21_X1 U12160 ( .B1(n13139), .B2(n13138), .A(n13137), .ZN(n13153) );
  AND2_X1 U12161 ( .A1(n11334), .A2(n10345), .ZN(n10317) );
  BUF_X1 U12162 ( .A(n10718), .Z(n13519) );
  AND2_X1 U12163 ( .A1(n19938), .A2(n13715), .ZN(n19355) );
  NAND2_X1 U12164 ( .A1(n19354), .A2(n19955), .ZN(n19518) );
  INV_X1 U12165 ( .A(n19697), .ZN(n13572) );
  NOR2_X1 U12166 ( .A1(n14372), .A2(n13514), .ZN(n19344) );
  NOR2_X1 U12167 ( .A1(n14376), .A2(n13514), .ZN(n19343) );
  INV_X1 U12168 ( .A(n19344), .ZN(n19335) );
  INV_X1 U12169 ( .A(n19343), .ZN(n19337) );
  NAND2_X1 U12170 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19777), .ZN(n19339) );
  AND3_X1 U12171 ( .A1(n15706), .A2(n15705), .A3(n15704), .ZN(n16404) );
  NAND2_X1 U12172 ( .A1(n20977), .A2(n16419), .ZN(n19980) );
  INV_X1 U12173 ( .A(n10036), .ZN(n18724) );
  AND2_X1 U12174 ( .A1(n9960), .A2(n9952), .ZN(n16621) );
  NAND2_X1 U12175 ( .A1(n18951), .A2(n17444), .ZN(n12851) );
  NAND2_X1 U12176 ( .A1(n17112), .A2(n10233), .ZN(n17068) );
  INV_X1 U12177 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16769) );
  NAND2_X1 U12178 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17189), .ZN(n15770) );
  NOR2_X1 U12179 ( .A1(n17364), .A2(n9907), .ZN(n17329) );
  NAND2_X1 U12180 ( .A1(n9837), .A2(P3_EAX_REG_18__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U12181 ( .A1(n11012), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9941) );
  INV_X1 U12182 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17212) );
  AOI21_X1 U12183 ( .B1(n18747), .B2(n15781), .A(n15784), .ZN(n15888) );
  AND2_X1 U12184 ( .A1(n11109), .A2(n11108), .ZN(n11276) );
  NOR2_X1 U12185 ( .A1(n11246), .A2(n18287), .ZN(n18760) );
  INV_X1 U12186 ( .A(n18268), .ZN(n17444) );
  NOR2_X1 U12187 ( .A1(n17443), .A2(n17442), .ZN(n17461) );
  NOR2_X1 U12188 ( .A1(n18784), .A2(n18725), .ZN(n17480) );
  AND2_X1 U12189 ( .A1(n10042), .A2(n9870), .ZN(n16429) );
  NAND2_X1 U12190 ( .A1(n11272), .A2(n16614), .ZN(n10042) );
  NAND2_X1 U12191 ( .A1(n17577), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17553) );
  NOR2_X1 U12192 ( .A1(n17639), .A2(n17640), .ZN(n17618) );
  NOR2_X1 U12193 ( .A1(n17673), .A2(n17674), .ZN(n17662) );
  NAND2_X1 U12194 ( .A1(n9942), .A2(n17817), .ZN(n17712) );
  AND2_X1 U12195 ( .A1(n16786), .A2(n9850), .ZN(n9942) );
  INV_X1 U12196 ( .A(n16425), .ZN(n18112) );
  INV_X1 U12197 ( .A(n15819), .ZN(n18110) );
  INV_X1 U12198 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16849) );
  NOR2_X1 U12199 ( .A1(n11296), .A2(n17859), .ZN(n17843) );
  NOR2_X1 U12200 ( .A1(n17892), .A2(n17877), .ZN(n17862) );
  NOR2_X1 U12201 ( .A1(n18272), .A2(n16583), .ZN(n11274) );
  NAND2_X1 U12202 ( .A1(n9937), .A2(n9936), .ZN(n15800) );
  AND2_X1 U12203 ( .A1(n17928), .A2(n17551), .ZN(n9936) );
  OAI211_X1 U12204 ( .C1(n11076), .C2(n17252), .A(n11024), .B(n11023), .ZN(
        n16471) );
  INV_X1 U12205 ( .A(n11136), .ZN(n9937) );
  NAND2_X1 U12206 ( .A1(n17659), .A2(n17651), .ZN(n17688) );
  AOI21_X1 U12207 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n11128), .A(
        n9939), .ZN(n17698) );
  NAND2_X1 U12208 ( .A1(n11129), .A2(n9940), .ZN(n9939) );
  NAND2_X1 U12209 ( .A1(n17820), .A2(n18050), .ZN(n9940) );
  NAND2_X1 U12210 ( .A1(n17698), .A2(n18040), .ZN(n17697) );
  NOR2_X1 U12211 ( .A1(n11127), .A2(n17737), .ZN(n18057) );
  NOR2_X1 U12212 ( .A1(n18080), .A2(n18077), .ZN(n18055) );
  NAND2_X1 U12213 ( .A1(n18733), .A2(n10034), .ZN(n18759) );
  NAND2_X1 U12214 ( .A1(n12835), .A2(n10035), .ZN(n10034) );
  INV_X1 U12215 ( .A(n18734), .ZN(n10035) );
  NOR2_X1 U12216 ( .A1(n9849), .A2(n21098), .ZN(n17819) );
  INV_X1 U12217 ( .A(n11124), .ZN(n11122) );
  OR2_X1 U12218 ( .A1(n18735), .A2(n11265), .ZN(n13838) );
  NAND2_X1 U12219 ( .A1(n17915), .A2(n17906), .ZN(n17905) );
  NAND2_X1 U12220 ( .A1(n15806), .A2(n15788), .ZN(n15818) );
  NOR2_X1 U12221 ( .A1(n12834), .A2(n12833), .ZN(n18761) );
  NAND2_X1 U12222 ( .A1(n12835), .A2(n12834), .ZN(n18747) );
  NOR2_X1 U12223 ( .A1(n16578), .A2(n16580), .ZN(n18564) );
  INV_X1 U12224 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18626) );
  INV_X1 U12225 ( .A(n11238), .ZN(n18287) );
  NAND2_X1 U12226 ( .A1(n18936), .A2(n18266), .ZN(n18459) );
  NOR2_X1 U12227 ( .A1(n18948), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n17744) );
  NOR2_X1 U12228 ( .A1(n18933), .A2(n15782), .ZN(n18786) );
  INV_X1 U12229 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14502) );
  INV_X1 U12230 ( .A(n20022), .ZN(n20069) );
  XNOR2_X1 U12231 ( .A(n12533), .B(n13181), .ZN(n13666) );
  INV_X1 U12232 ( .A(n20098), .ZN(n20056) );
  INV_X1 U12233 ( .A(n20091), .ZN(n14545) );
  NAND2_X1 U12234 ( .A1(n12528), .A2(n14397), .ZN(n14612) );
  NAND2_X1 U12235 ( .A1(n13029), .A2(n12527), .ZN(n12528) );
  INV_X1 U12236 ( .A(n14612), .ZN(n14626) );
  NAND2_X1 U12237 ( .A1(n14704), .A2(n13424), .ZN(n15984) );
  NAND2_X1 U12238 ( .A1(n13789), .A2(n13020), .ZN(n12798) );
  AND2_X1 U12239 ( .A1(n15984), .A2(n13425), .ZN(n14706) );
  INV_X2 U12240 ( .A(n15988), .ZN(n14708) );
  AND2_X1 U12241 ( .A1(n13789), .A2(n13061), .ZN(n20104) );
  INV_X1 U12242 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15916) );
  INV_X1 U12243 ( .A(n14681), .ZN(n15994) );
  INV_X1 U12244 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15934) );
  INV_X1 U12246 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U12247 ( .A1(n13832), .A2(n14385), .ZN(n16116) );
  AND2_X1 U12248 ( .A1(n13947), .A2(n13948), .ZN(n14963) );
  INV_X1 U12249 ( .A(n9916), .ZN(n14835) );
  NOR2_X1 U12250 ( .A1(n20206), .A2(n16118), .ZN(n16135) );
  NAND2_X1 U12251 ( .A1(n10068), .A2(n12742), .ZN(n16025) );
  NAND2_X1 U12252 ( .A1(n16031), .A2(n12740), .ZN(n10068) );
  INV_X1 U12253 ( .A(n16116), .ZN(n20206) );
  AND2_X1 U12254 ( .A1(n13832), .A2(n13822), .ZN(n20228) );
  INV_X1 U12255 ( .A(n20846), .ZN(n20859) );
  INV_X1 U12256 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20539) );
  INV_X1 U12257 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20234) );
  NAND2_X1 U12258 ( .A1(n13241), .A2(n20370), .ZN(n20864) );
  INV_X1 U12259 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13079) );
  NOR2_X1 U12260 ( .A1(n20615), .A2(n15862), .ZN(n13240) );
  CLKBUF_X1 U12261 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15019) );
  INV_X1 U12262 ( .A(n13240), .ZN(n15014) );
  OAI22_X1 U12263 ( .A1(n20310), .A2(n20309), .B1(n20479), .B2(n20308), .ZN(
        n20328) );
  OAI21_X1 U12264 ( .B1(n20310), .B2(n20307), .A(n20306), .ZN(n20329) );
  OAI21_X1 U12265 ( .B1(n20389), .B2(n20371), .A(n20681), .ZN(n20391) );
  INV_X1 U12266 ( .A(n20387), .ZN(n20390) );
  NOR2_X1 U12267 ( .A1(n20863), .A2(n20453), .ZN(n20471) );
  OAI211_X1 U12268 ( .C1(n20502), .C2(n20615), .A(n20541), .B(n20486), .ZN(
        n20504) );
  INV_X1 U12269 ( .A(n20545), .ZN(n20569) );
  NOR2_X1 U12270 ( .A1(n20580), .A2(n20675), .ZN(n20587) );
  INV_X1 U12271 ( .A(n20275), .ZN(n20718) );
  INV_X1 U12272 ( .A(n20548), .ZN(n20717) );
  INV_X1 U12273 ( .A(n20551), .ZN(n20728) );
  INV_X1 U12274 ( .A(n20557), .ZN(n20740) );
  INV_X1 U12275 ( .A(n20560), .ZN(n20746) );
  INV_X1 U12276 ( .A(n20775), .ZN(n20761) );
  INV_X1 U12277 ( .A(n20566), .ZN(n20758) );
  NOR2_X1 U12278 ( .A1(n20863), .A2(n20716), .ZN(n20768) );
  OR2_X1 U12279 ( .A1(n20676), .A2(n20448), .ZN(n20775) );
  INV_X1 U12280 ( .A(n20764), .ZN(n20771) );
  OR2_X1 U12281 ( .A1(n20778), .A2(n16155), .ZN(n19992) );
  INV_X1 U12282 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16162) );
  INV_X1 U12283 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n16155) );
  NAND2_X1 U12284 ( .A1(n16162), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20778) );
  NAND2_X1 U12285 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20880) );
  NAND2_X1 U12286 ( .A1(n15062), .A2(n19075), .ZN(n16180) );
  NAND2_X1 U12287 ( .A1(n16192), .A2(n19075), .ZN(n15064) );
  NAND2_X1 U12288 ( .A1(n15064), .A2(n15063), .ZN(n15062) );
  NAND2_X1 U12289 ( .A1(n16193), .A2(n16194), .ZN(n16192) );
  NAND2_X1 U12290 ( .A1(n16215), .A2(n19075), .ZN(n16205) );
  NAND2_X1 U12291 ( .A1(n16205), .A2(n16206), .ZN(n16204) );
  NAND2_X1 U12292 ( .A1(n15080), .A2(n19075), .ZN(n16216) );
  NAND2_X1 U12293 ( .A1(n16216), .A2(n16217), .ZN(n16215) );
  NAND2_X1 U12294 ( .A1(n16229), .A2(n19075), .ZN(n15081) );
  NAND2_X1 U12295 ( .A1(n15081), .A2(n15334), .ZN(n15080) );
  NAND2_X1 U12296 ( .A1(n16230), .A2(n16231), .ZN(n16229) );
  NAND2_X1 U12297 ( .A1(n18995), .A2(n13635), .ZN(n15829) );
  NAND2_X1 U12298 ( .A1(n13635), .A2(n10232), .ZN(n19000) );
  NAND2_X1 U12299 ( .A1(n19000), .A2(n18996), .ZN(n18995) );
  AND2_X1 U12300 ( .A1(n10906), .A2(n10908), .ZN(n15095) );
  INV_X1 U12301 ( .A(n19158), .ZN(n19138) );
  NAND2_X1 U12302 ( .A1(n16166), .A2(n13542), .ZN(n19128) );
  NAND2_X1 U12303 ( .A1(n19133), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19158) );
  INV_X1 U12304 ( .A(n19150), .ZN(n19089) );
  INV_X1 U12305 ( .A(n10074), .ZN(n10616) );
  OR2_X1 U12306 ( .A1(n11469), .A2(n11468), .ZN(n13393) );
  OR2_X1 U12307 ( .A1(n11443), .A2(n11442), .ZN(n13208) );
  INV_X1 U12308 ( .A(n15219), .ZN(n15199) );
  INV_X1 U12309 ( .A(n15224), .ZN(n15205) );
  INV_X1 U12310 ( .A(n19944), .ZN(n13715) );
  NAND2_X1 U12311 ( .A1(n13048), .A2(n12961), .ZN(n15124) );
  NAND2_X1 U12312 ( .A1(n15701), .A2(n15727), .ZN(n12955) );
  NOR2_X1 U12313 ( .A1(n15126), .A2(n14345), .ZN(n14368) );
  NAND2_X1 U12314 ( .A1(n14315), .A2(n15132), .ZN(n10106) );
  NOR2_X1 U12315 ( .A1(n14179), .A2(n15162), .ZN(n15157) );
  INV_X1 U12316 ( .A(n15292), .ZN(n19167) );
  INV_X1 U12317 ( .A(n19160), .ZN(n19168) );
  OAI21_X1 U12318 ( .B1(n12996), .B2(n12995), .A(n10149), .ZN(n13035) );
  OR2_X1 U12319 ( .A1(n19190), .A2(n11367), .ZN(n19171) );
  NAND2_X1 U12320 ( .A1(n12970), .A2(n12969), .ZN(n19190) );
  OR2_X1 U12321 ( .A1(n15699), .A2(n12968), .ZN(n12970) );
  INV_X1 U12322 ( .A(n19170), .ZN(n16246) );
  INV_X1 U12323 ( .A(n19171), .ZN(n19194) );
  AND2_X1 U12324 ( .A1(n19205), .A2(n19972), .ZN(n19270) );
  CLKBUF_X1 U12325 ( .A(n13531), .Z(n13538) );
  OAI21_X1 U12326 ( .B1(n14294), .B2(n19983), .A(n18956), .ZN(n12905) );
  NOR2_X1 U12327 ( .A1(n13539), .A2(n14316), .ZN(n13531) );
  INV_X1 U12328 ( .A(n12989), .ZN(n12932) );
  INV_X1 U12329 ( .A(n13531), .ZN(n19201) );
  XNOR2_X1 U12330 ( .A(n13527), .B(n13526), .ZN(n14037) );
  NAND2_X1 U12331 ( .A1(n15050), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13527) );
  INV_X1 U12332 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15321) );
  INV_X1 U12333 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15409) );
  NAND2_X1 U12334 ( .A1(n16308), .A2(n16307), .ZN(n16306) );
  NAND2_X1 U12335 ( .A1(n15658), .A2(n10993), .ZN(n16308) );
  AND2_X1 U12336 ( .A1(n13263), .A2(n13184), .ZN(n16338) );
  INV_X1 U12337 ( .A(n19274), .ZN(n16314) );
  INV_X1 U12338 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16323) );
  OR2_X1 U12339 ( .A1(n18967), .A2(n19970), .ZN(n16292) );
  INV_X1 U12340 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13705) );
  NAND2_X1 U12341 ( .A1(n18967), .A2(n10591), .ZN(n19288) );
  AND2_X1 U12342 ( .A1(n19288), .A2(n12867), .ZN(n19274) );
  INV_X1 U12343 ( .A(n19278), .ZN(n16317) );
  INV_X1 U12344 ( .A(n19288), .ZN(n16299) );
  NAND2_X1 U12345 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U12346 ( .A1(n9989), .A2(n10939), .ZN(n15316) );
  NAND2_X1 U12347 ( .A1(n10938), .A2(n10937), .ZN(n15331) );
  AND2_X1 U12348 ( .A1(n10196), .A2(n10194), .ZN(n16280) );
  NAND2_X1 U12349 ( .A1(n10196), .A2(n10856), .ZN(n15648) );
  CLKBUF_X1 U12350 ( .A(n15669), .Z(n15670) );
  INV_X1 U12351 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19958) );
  INV_X1 U12352 ( .A(n15124), .ZN(n19955) );
  INV_X1 U12353 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19950) );
  NOR2_X1 U12354 ( .A1(n13251), .A2(n11391), .ZN(n13350) );
  INV_X1 U12355 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16419) );
  XNOR2_X1 U12356 ( .A(n13046), .B(n13045), .ZN(n19944) );
  XNOR2_X1 U12357 ( .A(n13139), .B(n13138), .ZN(n19938) );
  INV_X1 U12358 ( .A(n16394), .ZN(n15796) );
  INV_X1 U12359 ( .A(n19373), .ZN(n19378) );
  OAI21_X1 U12360 ( .B1(n13750), .B2(n19722), .A(n13749), .ZN(n19448) );
  INV_X1 U12361 ( .A(n19487), .ZN(n19506) );
  NOR2_X1 U12362 ( .A1(n19719), .A2(n19483), .ZN(n19535) );
  OAI21_X1 U12363 ( .B1(n19517), .B2(n19923), .A(n19516), .ZN(n19536) );
  OAI21_X1 U12364 ( .B1(n19564), .B2(n19543), .A(n19777), .ZN(n19567) );
  OAI21_X1 U12365 ( .B1(n19615), .B2(n19614), .A(n19777), .ZN(n19634) );
  NOR2_X1 U12366 ( .A1(n13569), .A2(n13568), .ZN(n19652) );
  INV_X1 U12367 ( .A(n19663), .ZN(n19682) );
  INV_X1 U12368 ( .A(n19763), .ZN(n19721) );
  NOR2_X2 U12369 ( .A1(n19697), .A2(n19696), .ZN(n19763) );
  INV_X1 U12370 ( .A(n19736), .ZN(n19775) );
  INV_X1 U12371 ( .A(n19744), .ZN(n19794) );
  AND2_X1 U12372 ( .A1(n10344), .A2(n19319), .ZN(n19799) );
  INV_X1 U12373 ( .A(n19752), .ZN(n19806) );
  INV_X1 U12374 ( .A(n19834), .ZN(n19814) );
  INV_X1 U12375 ( .A(n19370), .ZN(n19811) );
  AND2_X1 U12376 ( .A1(n13570), .A2(n19319), .ZN(n19819) );
  INV_X1 U12377 ( .A(n19760), .ZN(n19820) );
  AOI22_X1 U12378 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19344), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19343), .ZN(n19835) );
  NAND2_X1 U12379 ( .A1(n19837), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n18965) );
  AND2_X1 U12380 ( .A1(n16419), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19837) );
  NOR2_X1 U12381 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19977) );
  NAND2_X1 U12382 ( .A1(n19849), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19986) );
  INV_X2 U12383 ( .A(n19986), .ZN(n19988) );
  INV_X1 U12384 ( .A(n17480), .ZN(n17443) );
  NAND2_X1 U12385 ( .A1(n11255), .A2(n11254), .ZN(n18950) );
  AOI21_X1 U12386 ( .B1(n18724), .B2(n18747), .A(n17443), .ZN(n18951) );
  AND2_X1 U12387 ( .A1(n9961), .A2(n9952), .ZN(n16632) );
  AND2_X1 U12388 ( .A1(n9956), .A2(n9952), .ZN(n12849) );
  AND2_X1 U12389 ( .A1(n9957), .A2(n9952), .ZN(n16652) );
  NOR2_X1 U12390 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16678), .ZN(n16663) );
  INV_X1 U12391 ( .A(n16935), .ZN(n16943) );
  NAND2_X1 U12392 ( .A1(n9950), .A2(n9951), .ZN(n16686) );
  AND2_X1 U12393 ( .A1(n9953), .A2(n9952), .ZN(n16687) );
  NOR2_X1 U12394 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16719), .ZN(n16705) );
  NOR2_X1 U12395 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16815), .ZN(n16800) );
  INV_X1 U12396 ( .A(n16939), .ZN(n16938) );
  INV_X1 U12397 ( .A(n16954), .ZN(n16947) );
  NOR2_X2 U12398 ( .A1(n18626), .A2(n16950), .ZN(n16939) );
  NOR2_X1 U12399 ( .A1(n16658), .A2(n17014), .ZN(n17017) );
  NOR2_X1 U12400 ( .A1(n17023), .A2(n16679), .ZN(n17027) );
  AND2_X1 U12401 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17066), .ZN(n17052) );
  NOR2_X1 U12402 ( .A1(n16721), .A2(n17068), .ZN(n17083) );
  NAND2_X1 U12403 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17157), .ZN(n17136) );
  NOR2_X1 U12404 ( .A1(n16795), .A2(n15770), .ZN(n17157) );
  INV_X1 U12405 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17208) );
  NAND2_X1 U12406 ( .A1(n17258), .A2(n13842), .ZN(n17248) );
  INV_X1 U12407 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17249) );
  NOR2_X1 U12408 ( .A1(n17248), .A2(n17249), .ZN(n17247) );
  NOR2_X1 U12409 ( .A1(n11193), .A2(n10045), .ZN(n10044) );
  OR3_X1 U12410 ( .A1(n18272), .A2(n18268), .A3(n18784), .ZN(n13840) );
  INV_X1 U12411 ( .A(P3_EAX_REG_31__SCAN_IN), .ZN(n9905) );
  NOR2_X1 U12412 ( .A1(n17503), .A2(n17308), .ZN(n17304) );
  NAND2_X1 U12413 ( .A1(n17312), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17308) );
  NOR2_X1 U12414 ( .A1(n17318), .A2(n17499), .ZN(n17312) );
  NAND2_X1 U12415 ( .A1(n17323), .A2(n18297), .ZN(n17317) );
  OR2_X1 U12416 ( .A1(n17497), .A2(n17317), .ZN(n17318) );
  NOR2_X1 U12417 ( .A1(n17324), .A2(n17495), .ZN(n17323) );
  NAND2_X1 U12418 ( .A1(n17329), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17324) );
  NOR2_X1 U12419 ( .A1(n17486), .A2(n17357), .ZN(n17351) );
  INV_X1 U12420 ( .A(n17367), .ZN(n17356) );
  NAND2_X1 U12421 ( .A1(n17368), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17364) );
  INV_X1 U12422 ( .A(n17438), .ZN(n17394) );
  INV_X1 U12423 ( .A(n17333), .ZN(n18297) );
  NOR2_X1 U12424 ( .A1(n17374), .A2(n17428), .ZN(n17412) );
  INV_X1 U12425 ( .A(n17435), .ZN(n17425) );
  OR2_X1 U12426 ( .A1(n17373), .A2(n17372), .ZN(n17428) );
  NOR2_X1 U12427 ( .A1(n10054), .A2(n10053), .ZN(n10052) );
  OAI21_X1 U12428 ( .B1(n15888), .B2(n15887), .A(n18939), .ZN(n17436) );
  NOR3_X1 U12429 ( .A1(n15886), .A2(n17444), .A3(n18933), .ZN(n15887) );
  NAND2_X1 U12430 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11057) );
  INV_X1 U12431 ( .A(n17436), .ZN(n17429) );
  NOR2_X1 U12432 ( .A1(n15889), .A2(n17436), .ZN(n17434) );
  OAI211_X1 U12433 ( .C1(n18272), .C2(n18809), .A(n17481), .B(n17480), .ZN(
        n17539) );
  NOR2_X1 U12435 ( .A1(n16428), .A2(n17630), .ZN(n17573) );
  NOR2_X1 U12436 ( .A1(n17591), .A2(n17592), .ZN(n17577) );
  INV_X1 U12437 ( .A(n17720), .ZN(n17702) );
  AND2_X1 U12438 ( .A1(n9821), .A2(n17817), .ZN(n17705) );
  INV_X1 U12439 ( .A(n17713), .ZN(n9943) );
  NAND2_X1 U12440 ( .A1(n17786), .A2(n16426), .ZN(n17720) );
  AND2_X1 U12441 ( .A1(n9944), .A2(n17817), .ZN(n17731) );
  AND2_X1 U12442 ( .A1(n16786), .A2(n9945), .ZN(n9944) );
  OAI22_X1 U12443 ( .A1(n17753), .A2(n18110), .B1(n17920), .B2(n18112), .ZN(
        n17786) );
  INV_X1 U12444 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17834) );
  INV_X1 U12445 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17847) );
  NAND2_X1 U12446 ( .A1(n17857), .A2(n11119), .ZN(n17851) );
  INV_X1 U12447 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17877) );
  NAND2_X1 U12448 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17892) );
  INV_X1 U12449 ( .A(n18666), .ZN(n18392) );
  INV_X1 U12450 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17910) );
  NAND2_X1 U12451 ( .A1(n16583), .A2(n9900), .ZN(n17916) );
  INV_X1 U12452 ( .A(n17909), .ZN(n17920) );
  NAND2_X1 U12453 ( .A1(n9937), .A2(n17928), .ZN(n17568) );
  INV_X1 U12454 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18948) );
  INV_X1 U12455 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18040) );
  NOR2_X1 U12456 ( .A1(n17761), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17754) );
  NOR3_X2 U12457 ( .A1(n15818), .A2(n18245), .A3(n17410), .ZN(n18139) );
  INV_X1 U12458 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18181) );
  INV_X1 U12459 ( .A(n18113), .ZN(n18723) );
  AOI21_X2 U12460 ( .B1(n15812), .B2(n15811), .A(n18784), .ZN(n18224) );
  AOI211_X1 U12461 ( .C1(n15806), .C2(n15805), .A(n15804), .B(n15803), .ZN(
        n15812) );
  NAND2_X1 U12462 ( .A1(n16718), .A2(n18245), .ZN(n18230) );
  INV_X1 U12463 ( .A(n18224), .ZN(n18245) );
  INV_X1 U12464 ( .A(n18761), .ZN(n18739) );
  INV_X1 U12465 ( .A(n18175), .ZN(n18244) );
  INV_X1 U12466 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18767) );
  INV_X1 U12467 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18772) );
  INV_X1 U12468 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18261) );
  AOI211_X1 U12469 ( .C1(n18939), .C2(n18758), .A(n18267), .B(n15792), .ZN(
        n18917) );
  INV_X1 U12470 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18506) );
  INV_X1 U12471 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n21093) );
  NOR2_X1 U12472 ( .A1(n18936), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18796) );
  INV_X1 U12473 ( .A(n17744), .ZN(n18803) );
  NOR3_X1 U12474 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18829), .A3(n18806), 
        .ZN(n18932) );
  NAND2_X1 U12475 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18820), .ZN(n18946) );
  AND2_X2 U12476 ( .A1(n12811), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14628)
         );
  CLKBUF_X1 U12477 ( .A(n16569), .Z(n16566) );
  OAI21_X1 U12478 ( .B1(n14546), .B2(n20098), .A(n12675), .ZN(n12676) );
  AND4_X1 U12479 ( .A1(n20095), .A2(n20094), .A3(n20093), .A4(n20092), .ZN(
        n20096) );
  OAI21_X1 U12480 ( .B1(n13959), .B2(n19999), .A(n12789), .ZN(P1_U2968) );
  OAI21_X1 U12481 ( .B1(n13959), .B2(n16049), .A(n10170), .ZN(P1_U3000) );
  INV_X1 U12482 ( .A(n10171), .ZN(n10170) );
  OAI21_X1 U12483 ( .B1(n14546), .B2(n20224), .A(n10172), .ZN(n10171) );
  NOR3_X1 U12484 ( .A1(n13958), .A2(n13957), .A3(n13956), .ZN(n10172) );
  OR2_X1 U12485 ( .A1(n15054), .A2(n19150), .ZN(n10137) );
  AOI21_X1 U12486 ( .B1(n15301), .B2(n19109), .A(n10139), .ZN(n10138) );
  NOR2_X1 U12487 ( .A1(n10600), .A2(n10599), .ZN(n11005) );
  AOI21_X1 U12488 ( .B1(n16171), .B2(n16339), .A(n14057), .ZN(n14060) );
  OAI21_X1 U12489 ( .B1(n19161), .B2(n16360), .A(n14056), .ZN(n14057) );
  AOI211_X1 U12490 ( .C1(n15301), .C2(n16339), .A(n13943), .B(n13942), .ZN(
        n13945) );
  NOR2_X1 U12491 ( .A1(n11581), .A2(n11580), .ZN(n11587) );
  NAND2_X1 U12492 ( .A1(n10115), .A2(n10113), .ZN(n10112) );
  AND2_X1 U12493 ( .A1(n10114), .A2(n9903), .ZN(n10113) );
  INV_X1 U12494 ( .A(n10116), .ZN(n15570) );
  AND2_X1 U12495 ( .A1(n9966), .A2(n9963), .ZN(n9962) );
  INV_X1 U12496 ( .A(n16613), .ZN(n9968) );
  AOI21_X1 U12497 ( .B1(n17287), .B2(P3_EAX_REG_30__SCAN_IN), .A(n9904), .ZN(
        n17288) );
  AOI21_X1 U12498 ( .B1(n17292), .B2(n9906), .A(n9905), .ZN(n9904) );
  AND2_X1 U12499 ( .A1(n11308), .A2(n11307), .ZN(n11309) );
  AND2_X1 U12500 ( .A1(n10043), .A2(n10039), .ZN(n11308) );
  BUF_X1 U12501 ( .A(n12291), .Z(n12209) );
  INV_X1 U12502 ( .A(n12291), .ZN(n11734) );
  INV_X2 U12503 ( .A(n9841), .ZN(n17105) );
  AND2_X2 U12504 ( .A1(n14354), .A2(n16379), .ZN(n11447) );
  AND2_X1 U12505 ( .A1(n13140), .A2(n10642), .ZN(n9818) );
  NAND2_X1 U12506 ( .A1(n10089), .A2(n9893), .ZN(n15173) );
  AND2_X1 U12507 ( .A1(n12373), .A2(n10224), .ZN(n14411) );
  OR2_X1 U12508 ( .A1(n15191), .A2(n15190), .ZN(n9819) );
  AND2_X1 U12509 ( .A1(n9989), .A2(n9892), .ZN(n15306) );
  AND2_X1 U12510 ( .A1(n14477), .A2(n10215), .ZN(n14465) );
  NAND2_X1 U12511 ( .A1(n14477), .A2(n14479), .ZN(n14478) );
  NAND2_X1 U12512 ( .A1(n10222), .A2(n12078), .ZN(n13769) );
  AND2_X1 U12513 ( .A1(n13140), .A2(n10644), .ZN(n9820) );
  INV_X1 U12514 ( .A(n13037), .ZN(n10655) );
  NOR2_X1 U12515 ( .A1(n13991), .A2(n9899), .ZN(n11541) );
  OR2_X1 U12516 ( .A1(n13763), .A2(n9867), .ZN(n14855) );
  AND2_X1 U12517 ( .A1(n16786), .A2(n9864), .ZN(n9821) );
  AND2_X1 U12518 ( .A1(n15308), .A2(n9892), .ZN(n9822) );
  AND2_X1 U12519 ( .A1(n10146), .A2(n10144), .ZN(n9823) );
  AND2_X1 U12520 ( .A1(n10277), .A2(n10275), .ZN(n9824) );
  AND2_X1 U12521 ( .A1(n10281), .A2(n10279), .ZN(n9825) );
  AND2_X1 U12522 ( .A1(n10077), .A2(n9884), .ZN(n9826) );
  AND2_X1 U12523 ( .A1(n11774), .A2(n20238), .ZN(n9827) );
  OR2_X1 U12524 ( .A1(n10036), .A2(n9869), .ZN(n12833) );
  AND2_X1 U12525 ( .A1(n10845), .A2(n9887), .ZN(n9828) );
  NAND2_X1 U12526 ( .A1(n14035), .A2(n13931), .ZN(n15058) );
  INV_X1 U12527 ( .A(n15058), .ZN(n15301) );
  NAND4_X1 U12528 ( .A1(n13811), .A2(n14819), .A3(n12776), .A4(n14822), .ZN(
        n9829) );
  AND2_X1 U12529 ( .A1(n15372), .A2(n9902), .ZN(n15386) );
  AND2_X1 U12530 ( .A1(n9951), .A2(n9952), .ZN(n9830) );
  NOR2_X1 U12531 ( .A1(n10017), .A2(n13342), .ZN(n9831) );
  AND2_X1 U12532 ( .A1(n13452), .A2(n13453), .ZN(n9832) );
  AND2_X1 U12533 ( .A1(n12546), .A2(n9832), .ZN(n9833) );
  OR2_X1 U12534 ( .A1(n12090), .A2(n12078), .ZN(n9834) );
  AND2_X1 U12535 ( .A1(n9946), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9835) );
  AND2_X1 U12536 ( .A1(n9923), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9836) );
  AND4_X1 U12537 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(P3_EAX_REG_21__SCAN_IN), .ZN(n9837)
         );
  AND2_X1 U12538 ( .A1(n10126), .A2(n15373), .ZN(n9838) );
  AND2_X2 U12539 ( .A1(n14353), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10560) );
  NAND2_X1 U12540 ( .A1(n9941), .A2(n18897), .ZN(n11055) );
  OR2_X1 U12541 ( .A1(n12972), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9839) );
  INV_X1 U12542 ( .A(n10073), .ZN(n15695) );
  INV_X1 U12543 ( .A(n11076), .ZN(n13906) );
  AND2_X2 U12544 ( .A1(n14353), .A2(n16379), .ZN(n10759) );
  AND2_X1 U12545 ( .A1(n10837), .A2(n10988), .ZN(n10979) );
  AND2_X2 U12546 ( .A1(n14357), .A2(n16379), .ZN(n10669) );
  NAND2_X1 U12547 ( .A1(n14855), .A2(n12765), .ZN(n13810) );
  INV_X1 U12549 ( .A(n13794), .ZN(n11765) );
  INV_X1 U12550 ( .A(n11246), .ZN(n18291) );
  NAND2_X1 U12551 ( .A1(n15247), .A2(n15246), .ZN(n13991) );
  NAND2_X1 U12552 ( .A1(n10093), .A2(n10081), .ZN(n15371) );
  AND2_X2 U12553 ( .A1(n14359), .A2(n16379), .ZN(n10686) );
  NAND2_X1 U12554 ( .A1(n10846), .A2(n10845), .ZN(n15435) );
  AND2_X1 U12555 ( .A1(n15372), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9843) );
  AND3_X1 U12556 ( .A1(n13798), .A2(n11782), .A3(n11781), .ZN(n9844) );
  AND4_X1 U12557 ( .A1(n11633), .A2(n11632), .A3(n11631), .A4(n11630), .ZN(
        n9845) );
  OAI21_X1 U12558 ( .B1(n9802), .B2(n10101), .A(n10100), .ZN(n15126) );
  AND2_X1 U12559 ( .A1(n9915), .A2(n9914), .ZN(n9846) );
  AND2_X1 U12560 ( .A1(n14477), .A2(n10214), .ZN(n14552) );
  NAND2_X1 U12561 ( .A1(n10211), .A2(n12189), .ZN(n14492) );
  NOR2_X1 U12562 ( .A1(n14490), .A2(n10212), .ZN(n14586) );
  NAND2_X1 U12563 ( .A1(n14477), .A2(n10217), .ZN(n9847) );
  AND2_X1 U12564 ( .A1(n10194), .A2(n16282), .ZN(n9848) );
  AND2_X1 U12565 ( .A1(n17831), .A2(n11125), .ZN(n9849) );
  NAND2_X1 U12566 ( .A1(n9981), .A2(n10868), .ZN(n15610) );
  OAI21_X1 U12567 ( .B1(n15423), .B2(n10924), .A(n10923), .ZN(n15497) );
  AND2_X1 U12568 ( .A1(n9945), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9850) );
  OR2_X1 U12569 ( .A1(n10893), .A2(n9999), .ZN(n9851) );
  NAND2_X1 U12570 ( .A1(n9818), .A2(n10654), .ZN(n10701) );
  AND2_X1 U12571 ( .A1(n13995), .A2(n10012), .ZN(n9852) );
  NAND2_X1 U12572 ( .A1(n10078), .A2(n10656), .ZN(n10726) );
  AND2_X1 U12573 ( .A1(n19970), .A2(n19951), .ZN(n11375) );
  OR2_X1 U12574 ( .A1(n13930), .A2(n10513), .ZN(n15125) );
  AND2_X1 U12575 ( .A1(n10888), .A2(n10002), .ZN(n9853) );
  NOR2_X1 U12576 ( .A1(n10617), .A2(n10629), .ZN(n10644) );
  OR2_X1 U12577 ( .A1(n10075), .A2(n19282), .ZN(n9854) );
  AND2_X1 U12578 ( .A1(n15056), .A2(n10010), .ZN(n9855) );
  AND2_X1 U12579 ( .A1(n9950), .A2(n9830), .ZN(n9856) );
  OR2_X1 U12580 ( .A1(n13991), .A2(n13992), .ZN(n9857) );
  NAND2_X1 U12581 ( .A1(n10196), .A2(n9848), .ZN(n15627) );
  AND2_X1 U12582 ( .A1(n10106), .A2(n10103), .ZN(n15127) );
  AND3_X1 U12583 ( .A1(n10276), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10278), .ZN(n9858) );
  AND3_X1 U12584 ( .A1(n10280), .A2(n16379), .A3(n10282), .ZN(n9859) );
  AND2_X1 U12585 ( .A1(n11125), .A2(n11132), .ZN(n9860) );
  AND2_X1 U12586 ( .A1(n10135), .A2(n13349), .ZN(n9861) );
  INV_X1 U12587 ( .A(n14490), .ZN(n10211) );
  AND2_X1 U12588 ( .A1(n17831), .A2(n9860), .ZN(n9862) );
  OR2_X1 U12589 ( .A1(n10858), .A2(n10005), .ZN(n9863) );
  AND2_X1 U12590 ( .A1(n9850), .A2(n9943), .ZN(n9864) );
  INV_X1 U12591 ( .A(n10150), .ZN(n10149) );
  OR2_X1 U12592 ( .A1(n11381), .A2(n11382), .ZN(n9865) );
  AND2_X1 U12593 ( .A1(n15247), .A2(n10155), .ZN(n13937) );
  NAND2_X1 U12594 ( .A1(n10089), .A2(n10087), .ZN(n14178) );
  NAND2_X1 U12595 ( .A1(n19980), .A2(n10388), .ZN(n9866) );
  NAND2_X1 U12596 ( .A1(n15372), .A2(n9838), .ZN(n15417) );
  NOR2_X1 U12597 ( .A1(n16013), .A2(n13764), .ZN(n9867) );
  NOR2_X1 U12598 ( .A1(n15145), .A2(n14260), .ZN(n14290) );
  AND3_X1 U12599 ( .A1(n14292), .A2(n9802), .A3(n10108), .ZN(n9868) );
  AND3_X1 U12600 ( .A1(n11250), .A2(n18272), .A3(n11249), .ZN(n9869) );
  NOR2_X1 U12601 ( .A1(n16446), .A2(n16452), .ZN(n9870) );
  NAND2_X1 U12602 ( .A1(n11547), .A2(n11545), .ZN(n10391) );
  NOR2_X1 U12603 ( .A1(n11061), .A2(n9934), .ZN(n9871) );
  NOR2_X1 U12604 ( .A1(n14020), .A2(n9996), .ZN(n9995) );
  AND2_X1 U12605 ( .A1(n10099), .A2(n15204), .ZN(n9872) );
  INV_X1 U12606 ( .A(n10084), .ZN(n14374) );
  AND2_X1 U12607 ( .A1(n10343), .A2(n12972), .ZN(n10084) );
  AND2_X2 U12608 ( .A1(n11635), .A2(n13070), .ZN(n11876) );
  OR2_X1 U12609 ( .A1(n14598), .A2(n14597), .ZN(n9873) );
  OR3_X1 U12610 ( .A1(n9873), .A2(n10167), .A3(n14570), .ZN(n9874) );
  NOR2_X1 U12611 ( .A1(n15167), .A2(n15166), .ZN(n9875) );
  NAND2_X1 U12612 ( .A1(n12766), .A2(n14990), .ZN(n9916) );
  INV_X2 U12613 ( .A(n10368), .ZN(n19970) );
  NAND2_X1 U12614 ( .A1(n12996), .A2(n10149), .ZN(n10145) );
  NAND2_X1 U12615 ( .A1(n10145), .A2(n10143), .ZN(n13157) );
  OAI21_X1 U12616 ( .B1(n13044), .B2(n13043), .A(n13137), .ZN(n13139) );
  NOR2_X1 U12617 ( .A1(n13326), .A2(n10022), .ZN(n13388) );
  NOR2_X1 U12618 ( .A1(n15516), .A2(n15515), .ZN(n11609) );
  NOR2_X1 U12619 ( .A1(n15182), .A2(n15183), .ZN(n15178) );
  NAND2_X1 U12620 ( .A1(n10145), .A2(n10146), .ZN(n13033) );
  NOR2_X1 U12621 ( .A1(n10786), .A2(n10783), .ZN(n10782) );
  NOR2_X1 U12622 ( .A1(n10028), .A2(n10027), .ZN(n15070) );
  NAND2_X1 U12623 ( .A1(n16394), .A2(n16397), .ZN(n11340) );
  OR2_X1 U12624 ( .A1(n13716), .A2(n10221), .ZN(n9876) );
  AND2_X1 U12625 ( .A1(n15043), .A2(n9923), .ZN(n9877) );
  OR2_X1 U12626 ( .A1(n15217), .A2(n10032), .ZN(n9878) );
  NOR2_X1 U12627 ( .A1(n9819), .A2(n15185), .ZN(n11605) );
  BUF_X1 U12628 ( .A(n10352), .Z(n11337) );
  NOR2_X1 U12629 ( .A1(n10799), .A2(n10775), .ZN(n10840) );
  OR2_X1 U12630 ( .A1(n10559), .A2(n10558), .ZN(n11397) );
  AND2_X1 U12631 ( .A1(n14065), .A2(n10099), .ZN(n15202) );
  AND2_X1 U12632 ( .A1(n13418), .A2(n10152), .ZN(n9879) );
  AND2_X1 U12634 ( .A1(n15575), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9880) );
  XNOR2_X1 U12635 ( .A(n10844), .B(n15675), .ZN(n15668) );
  NAND2_X1 U12636 ( .A1(n12764), .A2(n12763), .ZN(n13763) );
  NOR2_X1 U12637 ( .A1(n13326), .A2(n10019), .ZN(n13458) );
  AND2_X1 U12639 ( .A1(n15616), .A2(n13420), .ZN(n13418) );
  AND2_X1 U12640 ( .A1(n14065), .A2(n14064), .ZN(n9881) );
  OR2_X1 U12641 ( .A1(n15818), .A2(n18728), .ZN(n9882) );
  NOR2_X1 U12642 ( .A1(n15157), .A2(n15156), .ZN(n9883) );
  AND2_X1 U12643 ( .A1(n10694), .A2(n11397), .ZN(n9884) );
  INV_X1 U12644 ( .A(n10892), .ZN(n10876) );
  INV_X1 U12645 ( .A(n15182), .ZN(n10089) );
  AND2_X1 U12646 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9885) );
  INV_X1 U12647 ( .A(n10165), .ZN(n14571) );
  NOR2_X1 U12648 ( .A1(n9873), .A2(n10167), .ZN(n10165) );
  INV_X1 U12649 ( .A(n10004), .ZN(n10003) );
  NAND2_X1 U12650 ( .A1(n10887), .A2(n9898), .ZN(n10004) );
  INV_X1 U12651 ( .A(n10000), .ZN(n9999) );
  NOR2_X1 U12652 ( .A1(n10892), .A2(n10897), .ZN(n10000) );
  NOR2_X1 U12653 ( .A1(n15289), .A2(n15088), .ZN(n15087) );
  OR2_X1 U12654 ( .A1(n17638), .A2(n16696), .ZN(n9886) );
  NAND2_X1 U12655 ( .A1(n11605), .A2(n11606), .ZN(n11604) );
  INV_X1 U12656 ( .A(n13319), .ZN(n12546) );
  NOR2_X1 U12657 ( .A1(n11779), .A2(n11728), .ZN(n12645) );
  AND2_X1 U12658 ( .A1(n16302), .A2(n16300), .ZN(n9887) );
  AND2_X1 U12659 ( .A1(n10000), .A2(n10890), .ZN(n9888) );
  OR2_X1 U12660 ( .A1(n14075), .A2(n14074), .ZN(n15210) );
  INV_X1 U12661 ( .A(n10541), .ZN(n14272) );
  INV_X1 U12662 ( .A(n16913), .ZN(n16884) );
  NAND2_X1 U12663 ( .A1(n9971), .A2(n11340), .ZN(n11360) );
  AND2_X1 U12664 ( .A1(n20258), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12054) );
  INV_X1 U12665 ( .A(n12054), .ZN(n10207) );
  NAND2_X1 U12666 ( .A1(n13252), .A2(n10132), .ZN(n13351) );
  INV_X1 U12667 ( .A(n19109), .ZN(n19151) );
  OR2_X1 U12668 ( .A1(n16337), .A2(n19289), .ZN(n9889) );
  OR2_X1 U12669 ( .A1(n13269), .A2(n10017), .ZN(n13308) );
  NOR2_X1 U12670 ( .A1(n13099), .A2(n14395), .ZN(n9890) );
  AND2_X1 U12671 ( .A1(n14564), .A2(n14554), .ZN(n9891) );
  AND2_X1 U12672 ( .A1(n9988), .A2(n10939), .ZN(n9892) );
  AND2_X1 U12673 ( .A1(n10090), .A2(n15179), .ZN(n9893) );
  INV_X1 U12674 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21098) );
  AND2_X1 U12675 ( .A1(n13789), .A2(n15847), .ZN(n20169) );
  INV_X1 U12676 ( .A(n20169), .ZN(n19999) );
  AND2_X1 U12677 ( .A1(n14618), .A2(n14523), .ZN(n9894) );
  AND2_X1 U12678 ( .A1(n10025), .A2(n10024), .ZN(n9895) );
  AND2_X1 U12679 ( .A1(n10011), .A2(n13929), .ZN(n9896) );
  OR2_X1 U12680 ( .A1(n13772), .A2(n10175), .ZN(n9897) );
  NAND2_X1 U12681 ( .A1(n11970), .A2(n11913), .ZN(n20845) );
  NAND2_X1 U12682 ( .A1(n11895), .A2(n11894), .ZN(n20365) );
  INV_X1 U12683 ( .A(n9929), .ZN(n14008) );
  NOR2_X1 U12684 ( .A1(n15048), .A2(n16186), .ZN(n9929) );
  INV_X1 U12685 ( .A(n10013), .ZN(n10012) );
  NAND2_X1 U12686 ( .A1(n10503), .A2(n10014), .ZN(n10013) );
  INV_X1 U12687 ( .A(n14207), .ZN(n10098) );
  NAND2_X1 U12688 ( .A1(n10942), .A2(n10880), .ZN(n9898) );
  OR2_X1 U12689 ( .A1(n13992), .A2(n13970), .ZN(n9899) );
  INV_X1 U12690 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10008) );
  OR2_X1 U12691 ( .A1(n18938), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U12692 ( .A1(n16393), .A2(n10341), .ZN(n12966) );
  NAND2_X1 U12693 ( .A1(n10236), .A2(n21108), .ZN(n9901) );
  NAND2_X1 U12694 ( .A1(n17577), .A2(n9946), .ZN(n9949) );
  INV_X1 U12695 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9925) );
  AND2_X1 U12696 ( .A1(n9838), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9902) );
  INV_X1 U12697 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9948) );
  INV_X1 U12698 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10009) );
  AND4_X1 U12699 ( .A1(n18948), .A2(n18936), .A3(n16580), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n16941) );
  INV_X1 U12700 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15474) );
  INV_X1 U12701 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10125) );
  AND2_X1 U12702 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n10125), .ZN(
        n9903) );
  NOR2_X1 U12703 ( .A1(n18666), .A2(n19316), .ZN(n18680) );
  NAND2_X1 U12704 ( .A1(n18625), .A2(n18564), .ZN(n18666) );
  AOI22_X2 U12705 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20267), .B1(DATAI_28_), 
        .B2(n20266), .ZN(n20751) );
  NOR2_X4 U12706 ( .A1(n20884), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20830) );
  AOI22_X2 U12707 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20267), .B1(DATAI_24_), 
        .B2(n20266), .ZN(n20727) );
  INV_X1 U12708 ( .A(n20235), .ZN(n20266) );
  INV_X1 U12709 ( .A(n14043), .ZN(n11528) );
  AND2_X2 U12710 ( .A1(n11375), .A2(n10084), .ZN(n14043) );
  NAND3_X1 U12711 ( .A1(n17444), .A2(n18287), .A3(n18291), .ZN(n9908) );
  INV_X2 U12712 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18916) );
  NAND3_X1 U12713 ( .A1(n21179), .A2(n16945), .A3(n18897), .ZN(n17151) );
  NAND2_X1 U12714 ( .A1(n17304), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n17300) );
  NAND2_X1 U12715 ( .A1(n11675), .A2(n11674), .ZN(n9912) );
  INV_X1 U12716 ( .A(n11728), .ZN(n9911) );
  NAND3_X1 U12717 ( .A1(n9912), .A2(n9913), .A3(n11774), .ZN(n11779) );
  NAND2_X1 U12718 ( .A1(n12525), .A2(n11753), .ZN(n11663) );
  AOI21_X1 U12719 ( .B1(n14986), .B2(n9916), .A(n14985), .ZN(n14989) );
  XNOR2_X2 U12720 ( .A(n9917), .B(n14877), .ZN(n14876) );
  MUX2_X1 U12721 ( .A(n16013), .B(n14722), .S(n14721), .Z(n9917) );
  NAND2_X1 U12722 ( .A1(n14753), .A2(n14739), .ZN(n14740) );
  INV_X1 U12723 ( .A(n11892), .ZN(n9920) );
  AND2_X2 U12725 ( .A1(n9922), .A2(n9921), .ZN(n10071) );
  AOI21_X2 U12726 ( .B1(n14037), .B2(n20977), .A(n9928), .ZN(n13635) );
  OR2_X2 U12727 ( .A1(n9933), .A2(n11060), .ZN(n17433) );
  NAND3_X1 U12728 ( .A1(n9935), .A2(n11063), .A3(n9871), .ZN(n9933) );
  NAND2_X1 U12729 ( .A1(n10049), .A2(n17871), .ZN(n9938) );
  NAND2_X1 U12730 ( .A1(n17817), .A2(n16786), .ZN(n17746) );
  INV_X1 U12731 ( .A(n9949), .ZN(n16444) );
  INV_X1 U12732 ( .A(n9953), .ZN(n16694) );
  INV_X1 U12733 ( .A(n16884), .ZN(n9952) );
  INV_X1 U12734 ( .A(n9957), .ZN(n16664) );
  INV_X1 U12735 ( .A(n9956), .ZN(n16651) );
  INV_X1 U12736 ( .A(n9961), .ZN(n16641) );
  INV_X1 U12737 ( .A(n9960), .ZN(n16631) );
  OAI21_X1 U12738 ( .B1(n9967), .B2(n18800), .A(n9962), .ZN(P3_U2641) );
  XNOR2_X1 U12739 ( .A(n9969), .B(n9968), .ZN(n9967) );
  NOR2_X1 U12740 ( .A1(n16620), .A2(n16884), .ZN(n9969) );
  NAND3_X1 U12741 ( .A1(n9971), .A2(n11340), .A3(n9970), .ZN(n10380) );
  NAND3_X1 U12742 ( .A1(n16393), .A2(n10341), .A3(n10084), .ZN(n9970) );
  NOR2_X2 U12743 ( .A1(n9972), .A2(n10654), .ZN(n19659) );
  NAND2_X2 U12744 ( .A1(n9974), .A2(n9973), .ZN(n10364) );
  NAND2_X1 U12745 ( .A1(n9858), .A2(n9824), .ZN(n9973) );
  NAND2_X1 U12746 ( .A1(n9859), .A2(n9825), .ZN(n9974) );
  NAND3_X1 U12747 ( .A1(n9977), .A2(n10972), .A3(n9976), .ZN(n9975) );
  NAND2_X2 U12748 ( .A1(n10778), .A2(n10779), .ZN(n10972) );
  NOR2_X2 U12749 ( .A1(n14040), .A2(n14039), .ZN(n9978) );
  NOR2_X2 U12750 ( .A1(n15493), .A2(n9979), .ZN(n15310) );
  AND2_X2 U12751 ( .A1(n10077), .A2(n10694), .ZN(n10778) );
  NAND2_X2 U12752 ( .A1(n10076), .A2(n10711), .ZN(n10779) );
  INV_X1 U12753 ( .A(n10956), .ZN(n9997) );
  NAND2_X1 U12754 ( .A1(n10956), .A2(n9995), .ZN(n9992) );
  NAND3_X1 U12755 ( .A1(n9992), .A2(n9994), .A3(n14019), .ZN(n14029) );
  NAND2_X1 U12756 ( .A1(n10949), .A2(n9993), .ZN(n9994) );
  AND2_X2 U12757 ( .A1(n14358), .A2(n16379), .ZN(n10677) );
  AND3_X4 U12758 ( .A1(n15725), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n9998), .ZN(n14358) );
  NAND2_X1 U12759 ( .A1(n10001), .A2(n9888), .ZN(n10883) );
  NAND2_X1 U12760 ( .A1(n9853), .A2(n15180), .ZN(n10928) );
  OR2_X1 U12761 ( .A1(n10858), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10861) );
  INV_X1 U12762 ( .A(n10512), .ZN(n10015) );
  INV_X1 U12763 ( .A(n13269), .ZN(n10016) );
  NAND2_X1 U12764 ( .A1(n10016), .A2(n9831), .ZN(n13182) );
  NOR2_X1 U12765 ( .A1(n13269), .A2(n13268), .ZN(n13270) );
  INV_X1 U12766 ( .A(n13268), .ZN(n10018) );
  INV_X1 U12767 ( .A(n10028), .ZN(n15166) );
  INV_X1 U12768 ( .A(n15072), .ZN(n10027) );
  NAND2_X2 U12769 ( .A1(n10617), .A2(n10405), .ZN(n10417) );
  OR2_X2 U12770 ( .A1(n15783), .A2(n17481), .ZN(n10036) );
  NAND2_X1 U12771 ( .A1(n17871), .A2(n17870), .ZN(n17869) );
  NAND2_X1 U12772 ( .A1(n17870), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10048) );
  INV_X1 U12773 ( .A(n16485), .ZN(n17569) );
  AND2_X2 U12774 ( .A1(n11136), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16485) );
  NOR2_X1 U12775 ( .A1(n17579), .A2(n11135), .ZN(n11136) );
  NAND2_X2 U12776 ( .A1(n17831), .A2(n10050), .ZN(n17802) );
  NAND3_X1 U12777 ( .A1(n10052), .A2(n11070), .A3(n11072), .ZN(n17430) );
  NAND3_X1 U12778 ( .A1(n11073), .A2(n11068), .A3(n11067), .ZN(n10053) );
  NAND3_X1 U12779 ( .A1(n11071), .A2(n11069), .A3(n10235), .ZN(n10055) );
  INV_X2 U12780 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18897) );
  NOR2_X4 U12781 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13069) );
  INV_X1 U12782 ( .A(n13289), .ZN(n10056) );
  NAND2_X1 U12783 ( .A1(n12714), .A2(n10059), .ZN(n10058) );
  NAND2_X1 U12784 ( .A1(n13287), .A2(n12714), .ZN(n20156) );
  NAND2_X1 U12785 ( .A1(n13289), .A2(n13288), .ZN(n13287) );
  NAND2_X1 U12786 ( .A1(n16031), .A2(n10061), .ZN(n10064) );
  NOR2_X1 U12787 ( .A1(n10063), .A2(n10062), .ZN(n10061) );
  NAND2_X1 U12788 ( .A1(n13763), .A2(n10071), .ZN(n10070) );
  NAND2_X1 U12789 ( .A1(n10628), .A2(n10074), .ZN(n10073) );
  OR2_X1 U12790 ( .A1(n10075), .A2(n19295), .ZN(n10247) );
  NAND2_X1 U12791 ( .A1(n11003), .A2(n14040), .ZN(n10075) );
  NAND4_X1 U12792 ( .A1(n10662), .A2(n10663), .A3(n10660), .A4(n10661), .ZN(
        n10077) );
  NAND3_X1 U12793 ( .A1(n10078), .A2(n10656), .A3(
        P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10657) );
  XNOR2_X2 U12794 ( .A(n10992), .B(n15664), .ZN(n15440) );
  OR3_X1 U12796 ( .A1(n15493), .A2(n15325), .A3(n15474), .ZN(n15309) );
  NAND3_X1 U12797 ( .A1(n10360), .A2(n10084), .A3(n10372), .ZN(n10352) );
  NAND2_X1 U12799 ( .A1(n13037), .A2(n13141), .ZN(n10086) );
  NAND3_X1 U12800 ( .A1(n10092), .A2(n10091), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15644) );
  OAI21_X2 U12801 ( .B1(n10097), .B2(n15162), .A(n10096), .ZN(n14233) );
  NAND2_X1 U12802 ( .A1(n14065), .A2(n9872), .ZN(n15197) );
  NAND3_X1 U12803 ( .A1(n14292), .A2(n10104), .A3(n9802), .ZN(n10100) );
  NAND3_X1 U12804 ( .A1(n14292), .A2(n9802), .A3(n10107), .ZN(n10103) );
  NAND2_X1 U12805 ( .A1(n14292), .A2(n9802), .ZN(n15138) );
  INV_X1 U12806 ( .A(n15137), .ZN(n10108) );
  AOI21_X1 U12807 ( .B1(n15556), .B2(n16337), .A(n9880), .ZN(n15566) );
  NAND2_X1 U12808 ( .A1(n10112), .A2(n10109), .ZN(P2_U3029) );
  AND2_X1 U12809 ( .A1(n15372), .A2(n10126), .ZN(n15625) );
  NAND2_X1 U12810 ( .A1(n10128), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10127) );
  NAND4_X1 U12811 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10286), .ZN(
        n10128) );
  NAND2_X1 U12812 ( .A1(n10130), .A2(n16379), .ZN(n10129) );
  NAND4_X1 U12813 ( .A1(n10289), .A2(n10288), .A3(n10290), .A4(n10287), .ZN(
        n10130) );
  XNOR2_X1 U12814 ( .A(n11381), .B(n11382), .ZN(n13053) );
  NOR2_X1 U12815 ( .A1(n13250), .A2(n13249), .ZN(n13251) );
  NAND3_X1 U12816 ( .A1(n15057), .A2(n10138), .A3(n10137), .ZN(P2_U2825) );
  NOR2_X1 U12817 ( .A1(n10959), .A2(n11511), .ZN(n10150) );
  NAND2_X1 U12818 ( .A1(n10158), .A2(n10159), .ZN(n12533) );
  NAND3_X1 U12819 ( .A1(n10160), .A2(n12655), .A3(n12531), .ZN(n10158) );
  NAND2_X1 U12820 ( .A1(n12659), .A2(n13094), .ZN(n10160) );
  NAND3_X1 U12821 ( .A1(n12529), .A2(n13094), .A3(n12659), .ZN(n10159) );
  NAND2_X1 U12822 ( .A1(n9820), .A2(n10654), .ZN(n10700) );
  NAND4_X1 U12823 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10704) );
  NAND3_X1 U12824 ( .A1(n9820), .A2(n10654), .A3(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10183) );
  NAND3_X1 U12825 ( .A1(n9818), .A2(n10654), .A3(
        P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10184) );
  NAND3_X1 U12826 ( .A1(n9818), .A2(n10645), .A3(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10185) );
  NAND3_X1 U12827 ( .A1(n9820), .A2(n10645), .A3(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10186) );
  INV_X1 U12828 ( .A(n15384), .ZN(n11594) );
  NAND2_X1 U12829 ( .A1(n11596), .A2(n11595), .ZN(n15366) );
  NAND2_X1 U12830 ( .A1(n15347), .A2(n11597), .ZN(n11598) );
  NAND2_X1 U12831 ( .A1(n15423), .A2(n15424), .ZN(n10200) );
  INV_X1 U12832 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U12833 ( .A1(n11936), .A2(n11935), .ZN(n10204) );
  NAND2_X1 U12834 ( .A1(n10204), .A2(n11821), .ZN(n11839) );
  OAI21_X1 U12835 ( .B1(n12698), .B2(n10208), .A(n10205), .ZN(n13127) );
  NOR2_X2 U12836 ( .A1(n13716), .A2(n10219), .ZN(n14506) );
  NAND2_X1 U12837 ( .A1(n12373), .A2(n10223), .ZN(n12465) );
  AND2_X1 U12838 ( .A1(n12373), .A2(n10225), .ZN(n14423) );
  NAND2_X1 U12839 ( .A1(n12373), .A2(n12372), .ZN(n14438) );
  INV_X1 U12840 ( .A(n15501), .ZN(n11610) );
  AND2_X4 U12841 ( .A1(n11634), .A2(n11636), .ZN(n11800) );
  NAND2_X1 U12842 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11718) );
  AND2_X1 U12843 ( .A1(n13037), .A2(n13712), .ZN(n10641) );
  NAND2_X1 U12844 ( .A1(n14058), .A2(n16337), .ZN(n14059) );
  NOR2_X2 U12845 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15733) );
  AND2_X2 U12846 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15710) );
  NAND2_X1 U12847 ( .A1(n11053), .A2(n11052), .ZN(n11061) );
  CLKBUF_X1 U12848 ( .A(n13140), .Z(n15755) );
  AOI22_X1 U12849 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U12850 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U12851 ( .A1(n15224), .A2(n12972), .ZN(n15219) );
  OR2_X1 U12852 ( .A1(n19190), .A2(n12972), .ZN(n19170) );
  NAND2_X1 U12853 ( .A1(n13570), .A2(n12972), .ZN(n10358) );
  NOR2_X1 U12855 ( .A1(n10650), .A2(n10649), .ZN(n10718) );
  NOR2_X2 U12856 ( .A1(n10650), .A2(n10637), .ZN(n13617) );
  AND4_X2 U12857 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n10250) );
  NAND2_X1 U12858 ( .A1(n13152), .A2(n13153), .ZN(n13188) );
  OAI21_X1 U12859 ( .B1(n13153), .B2(n13152), .A(n13188), .ZN(n19354) );
  NOR2_X2 U12860 ( .A1(n15164), .A2(n15163), .ZN(n15162) );
  XNOR2_X1 U12861 ( .A(n11930), .B(n12689), .ZN(n13242) );
  NAND2_X1 U12862 ( .A1(n13129), .A2(n11948), .ZN(n13281) );
  NAND2_X1 U12863 ( .A1(n20845), .A2(n20848), .ZN(n20333) );
  NOR3_X1 U12864 ( .A1(n9853), .A2(n15180), .A3(n13515), .ZN(n10881) );
  NAND2_X1 U12865 ( .A1(n12800), .A2(n20050), .ZN(n12678) );
  INV_X1 U12866 ( .A(n14704), .ZN(n15985) );
  NAND2_X2 U12867 ( .A1(n12798), .A2(n12797), .ZN(n14704) );
  BUF_X1 U12868 ( .A(n11828), .Z(n12441) );
  INV_X1 U12869 ( .A(n10685), .ZN(n10738) );
  INV_X1 U12870 ( .A(n17661), .ZN(n17620) );
  OR2_X2 U12871 ( .A1(n11013), .A2(n11012), .ZN(n10227) );
  OR2_X1 U12872 ( .A1(n16013), .A2(n14890), .ZN(n10228) );
  AND2_X1 U12873 ( .A1(n15359), .A2(n15358), .ZN(n10229) );
  AND4_X1 U12874 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n10230) );
  AND2_X1 U12875 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10231) );
  OR2_X1 U12876 ( .A1(n19001), .A2(n19004), .ZN(n10232) );
  AND3_X1 U12877 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .A3(P3_EBX_REG_17__SCAN_IN), .ZN(n10233) );
  NOR2_X2 U12878 ( .A1(n17410), .A2(n11121), .ZN(n17820) );
  INV_X1 U12879 ( .A(n17820), .ZN(n11132) );
  INV_X1 U12880 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12784) );
  AND2_X1 U12881 ( .A1(n15369), .A2(n15358), .ZN(n10234) );
  OR2_X1 U12882 ( .A1(n17186), .A2(n11066), .ZN(n10235) );
  AND3_X1 U12883 ( .A1(n18080), .A2(n17756), .A3(n11127), .ZN(n10236) );
  INV_X1 U12884 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13038) );
  OR2_X1 U12885 ( .A1(n15560), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10237) );
  OR2_X1 U12886 ( .A1(n17433), .A2(n20976), .ZN(n10238) );
  AND2_X1 U12887 ( .A1(n10297), .A2(n10296), .ZN(n10239) );
  INV_X1 U12888 ( .A(n14627), .ZN(n14584) );
  OR2_X1 U12889 ( .A1(n21022), .A2(n18803), .ZN(n18940) );
  AND4_X1 U12890 ( .A1(n11600), .A2(n11590), .A3(n10903), .A4(n15349), .ZN(
        n10240) );
  AND2_X1 U12891 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .ZN(n10241) );
  AND2_X1 U12892 ( .A1(n10390), .A2(n10389), .ZN(n10242) );
  INV_X1 U12893 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11127) );
  INV_X1 U12894 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15885) );
  OR2_X1 U12895 ( .A1(n19270), .A2(n19269), .ZN(n19272) );
  INV_X1 U12896 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12787) );
  INV_X1 U12897 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20024) );
  INV_X2 U12898 ( .A(n12766), .ZN(n14858) );
  AND2_X1 U12899 ( .A1(n14258), .A2(n14288), .ZN(n10243) );
  AND2_X1 U12900 ( .A1(n11600), .A2(n11599), .ZN(n10245) );
  OR2_X1 U12901 ( .A1(n17852), .A2(n18181), .ZN(n10246) );
  INV_X1 U12902 ( .A(n14316), .ZN(n14294) );
  AND2_X1 U12903 ( .A1(n13960), .A2(n13963), .ZN(n10248) );
  AND2_X1 U12904 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10249) );
  INV_X1 U12905 ( .A(n10423), .ZN(n13199) );
  INV_X1 U12906 ( .A(n11372), .ZN(n11524) );
  AOI21_X1 U12907 ( .B1(n12487), .B2(n12486), .A(n12485), .ZN(n12499) );
  INV_X1 U12908 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11620) );
  OR2_X1 U12909 ( .A1(n11982), .A2(n11981), .ZN(n12735) );
  AOI22_X1 U12910 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11876), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U12911 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10286) );
  AND2_X1 U12912 ( .A1(n11549), .A2(n13570), .ZN(n10341) );
  NAND2_X1 U12913 ( .A1(n11545), .A2(n10346), .ZN(n10374) );
  INV_X1 U12914 ( .A(n10344), .ZN(n10346) );
  AOI22_X1 U12915 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10282) );
  OR2_X1 U12916 ( .A1(n12361), .A2(n12360), .ZN(n12374) );
  INV_X1 U12917 ( .A(n14520), .ZN(n12090) );
  INV_X1 U12918 ( .A(n11760), .ZN(n11781) );
  OR2_X1 U12919 ( .A1(n11799), .A2(n11798), .ZN(n12691) );
  NAND2_X1 U12920 ( .A1(n10375), .A2(n10374), .ZN(n10392) );
  AND2_X1 U12921 ( .A1(n10371), .A2(n12972), .ZN(n10342) );
  AND2_X1 U12922 ( .A1(n12503), .A2(n12504), .ZN(n12502) );
  OR2_X1 U12923 ( .A1(n12320), .A2(n12319), .ZN(n12331) );
  INV_X1 U12924 ( .A(n14453), .ZN(n12372) );
  INV_X1 U12925 ( .A(n14494), .ZN(n12189) );
  INV_X1 U12926 ( .A(n14606), .ZN(n12173) );
  INV_X1 U12927 ( .A(n13399), .ZN(n12014) );
  INV_X1 U12928 ( .A(n12687), .ZN(n12679) );
  INV_X1 U12929 ( .A(n12017), .ZN(n12018) );
  INV_X1 U12930 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11619) );
  AND2_X1 U12931 ( .A1(n14259), .A2(n10243), .ZN(n14260) );
  INV_X1 U12932 ( .A(n14234), .ZN(n14235) );
  INV_X1 U12933 ( .A(n15194), .ZN(n14108) );
  AOI22_X1 U12934 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10334) );
  NAND2_X1 U12935 ( .A1(n10240), .A2(n10234), .ZN(n10924) );
  NOR2_X1 U12936 ( .A1(n10581), .A2(n10580), .ZN(n10582) );
  INV_X1 U12937 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11329) );
  OAI21_X1 U12938 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21179), .A(
        n11156), .ZN(n11157) );
  AOI21_X1 U12939 ( .B1(n15019), .B2(n20574), .A(n12502), .ZN(n12501) );
  NOR2_X1 U12940 ( .A1(n12493), .A2(n12754), .ZN(n12519) );
  INV_X1 U12941 ( .A(n11846), .ZN(n11784) );
  AND2_X1 U12942 ( .A1(n12577), .A2(n12576), .ZN(n13827) );
  INV_X1 U12943 ( .A(n12615), .ZN(n12621) );
  INV_X1 U12944 ( .A(n12493), .ZN(n12514) );
  NAND2_X1 U12945 ( .A1(n14236), .A2(n14235), .ZN(n14237) );
  INV_X1 U12946 ( .A(n15198), .ZN(n14096) );
  AND4_X1 U12947 ( .A1(n10763), .A2(n10762), .A3(n10761), .A4(n10760), .ZN(
        n10764) );
  AOI22_X1 U12948 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10271) );
  NAND2_X1 U12949 ( .A1(n10307), .A2(n16379), .ZN(n10315) );
  INV_X1 U12950 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17143) );
  INV_X1 U12951 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17201) );
  INV_X1 U12952 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13851) );
  INV_X1 U12953 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17213) );
  INV_X1 U12954 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17071) );
  INV_X1 U12955 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n21086) );
  AOI221_X1 U12956 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12501), 
        .C1(n11963), .C2(n12501), .A(n12468), .ZN(n12642) );
  AOI21_X1 U12957 ( .B1(n12518), .B2(n12642), .A(n12517), .ZN(n12521) );
  AND2_X1 U12958 ( .A1(n12618), .A2(n12617), .ZN(n14554) );
  AND4_X1 U12959 ( .A1(n11718), .A2(n11717), .A3(n11716), .A4(n11715), .ZN(
        n11719) );
  INV_X1 U12960 ( .A(n13126), .ZN(n11946) );
  AND2_X1 U12961 ( .A1(n16013), .A2(n12760), .ZN(n13732) );
  AND2_X1 U12962 ( .A1(n11841), .A2(n11861), .ZN(n20536) );
  INV_X1 U12963 ( .A(n15218), .ZN(n10464) );
  OR2_X1 U12964 ( .A1(n14285), .A2(n14284), .ZN(n14287) );
  NOR2_X1 U12965 ( .A1(n14178), .A2(n14206), .ZN(n14179) );
  INV_X1 U12966 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13526) );
  OR2_X1 U12967 ( .A1(n16187), .A2(n10959), .ZN(n13962) );
  OR3_X1 U12968 ( .A1(n15824), .A2(n10959), .A3(n10999), .ZN(n15498) );
  OR2_X1 U12969 ( .A1(n10912), .A2(n15534), .ZN(n15359) );
  INV_X1 U12970 ( .A(n15634), .ZN(n15652) );
  XNOR2_X1 U12971 ( .A(n10994), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16307) );
  INV_X1 U12972 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15693) );
  INV_X1 U12973 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17234) );
  NAND2_X1 U12974 ( .A1(n17481), .A2(n18933), .ZN(n15781) );
  AND2_X1 U12975 ( .A1(n18900), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11137) );
  INV_X1 U12976 ( .A(n18092), .ZN(n18111) );
  NOR2_X1 U12977 ( .A1(n11107), .A2(n11106), .ZN(n11108) );
  INV_X1 U12978 ( .A(n18744), .ZN(n11009) );
  OR2_X1 U12979 ( .A1(n11234), .A2(n11233), .ZN(n11235) );
  INV_X1 U12980 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12325) );
  AND2_X1 U12981 ( .A1(n12607), .A2(n12606), .ZN(n14570) );
  NOR2_X1 U12982 ( .A1(n13498), .A2(n16162), .ZN(n12654) );
  INV_X1 U12983 ( .A(n20087), .ZN(n20025) );
  AND2_X1 U12984 ( .A1(n12620), .A2(n12619), .ZN(n14447) );
  AND2_X1 U12985 ( .A1(n15895), .A2(n12076), .ZN(n12346) );
  AND4_X1 U12986 ( .A1(n11725), .A2(n11724), .A3(n11723), .A4(n11722), .ZN(
        n11726) );
  OR2_X1 U12987 ( .A1(n12413), .A2(n14426), .ZN(n12439) );
  OR2_X1 U12988 ( .A1(n12371), .A2(n12370), .ZN(n14453) );
  NOR2_X1 U12989 ( .A1(n21036), .A2(n12123), .ZN(n12169) );
  NOR2_X1 U12990 ( .A1(n12057), .A2(n20024), .ZN(n12074) );
  NAND2_X1 U12991 ( .A1(n11923), .A2(n11922), .ZN(n13282) );
  AND2_X1 U12992 ( .A1(n13022), .A2(n13007), .ZN(n15847) );
  AND2_X1 U12993 ( .A1(n13946), .A2(n16116), .ZN(n20215) );
  INV_X1 U12994 ( .A(n20613), .ZN(n20678) );
  OR2_X1 U12995 ( .A1(n20845), .A2(n20481), .ZN(n20580) );
  NAND2_X1 U12996 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20269), .ZN(n20265) );
  INV_X1 U12997 ( .A(n13637), .ZN(n13638) );
  INV_X1 U12998 ( .A(n19129), .ZN(n19142) );
  AOI221_X1 U12999 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10530), 
        .C1(n11329), .C2(n10530), .A(n10529), .ZN(n11332) );
  OR2_X1 U13000 ( .A1(n16402), .A2(n15744), .ZN(n15701) );
  AND2_X1 U13001 ( .A1(n13470), .A2(n13469), .ZN(n14062) );
  XNOR2_X1 U13002 ( .A(n14178), .B(n14206), .ZN(n15164) );
  OR2_X1 U13003 ( .A1(n19190), .A2(n14377), .ZN(n15292) );
  INV_X1 U13004 ( .A(n11511), .ZN(n11470) );
  OAI21_X1 U13005 ( .B1(n12830), .B2(n12829), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12831) );
  INV_X1 U13006 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16186) );
  INV_X1 U13007 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15398) );
  INV_X1 U13008 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15429) );
  OR2_X1 U13009 ( .A1(n16227), .A2(n10959), .ZN(n10936) );
  INV_X1 U13010 ( .A(n16364), .ZN(n15562) );
  AND2_X1 U13011 ( .A1(n15579), .A2(n10237), .ZN(n15561) );
  AND2_X1 U13012 ( .A1(n16334), .A2(n11573), .ZN(n15649) );
  INV_X1 U13013 ( .A(n15471), .ZN(n15446) );
  INV_X1 U13014 ( .A(n19301), .ZN(n16360) );
  NAND2_X1 U13015 ( .A1(n15695), .A2(n13141), .ZN(n12958) );
  AND2_X1 U13016 ( .A1(n11561), .A2(n11560), .ZN(n15715) );
  INV_X1 U13017 ( .A(n19925), .ZN(n13742) );
  INV_X1 U13018 ( .A(n13610), .ZN(n19483) );
  INV_X1 U13019 ( .A(n19355), .ZN(n19577) );
  AND2_X1 U13020 ( .A1(n10700), .A2(n13562), .ZN(n13569) );
  INV_X1 U13021 ( .A(n19339), .ZN(n19319) );
  NOR2_X1 U13022 ( .A1(n17444), .A2(n18272), .ZN(n11267) );
  INV_X1 U13023 ( .A(n12833), .ZN(n12835) );
  NOR2_X1 U13024 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16746), .ZN(n16733) );
  NOR2_X1 U13025 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16794), .ZN(n16776) );
  NOR2_X1 U13026 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16830), .ZN(n16829) );
  INV_X1 U13027 ( .A(n16956), .ZN(n16902) );
  INV_X1 U13028 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17194) );
  INV_X1 U13029 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17170) );
  OAI21_X1 U13030 ( .B1(n15783), .B2(n18786), .A(n18932), .ZN(n17442) );
  NAND2_X1 U13031 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17618), .ZN(
        n17591) );
  NAND2_X1 U13032 ( .A1(n11305), .A2(n17821), .ZN(n16425) );
  AND2_X1 U13033 ( .A1(n17433), .A2(n17430), .ZN(n11284) );
  NOR2_X1 U13034 ( .A1(n18110), .A2(n18031), .ZN(n18058) );
  INV_X1 U13035 ( .A(n18220), .ZN(n18752) );
  NAND2_X1 U13036 ( .A1(n18722), .A2(n18802), .ZN(n18266) );
  INV_X1 U13037 ( .A(n18459), .ZN(n18625) );
  NOR2_X1 U13038 ( .A1(n18626), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18660) );
  AND2_X1 U13039 ( .A1(n14388), .A2(n14397), .ZN(n13789) );
  NAND2_X1 U13040 ( .A1(n13114), .A2(n12870), .ZN(n20878) );
  OR2_X1 U13041 ( .A1(n12326), .A2(n12325), .ZN(n12366) );
  NOR2_X1 U13042 ( .A1(n13727), .A2(n20037), .ZN(n20027) );
  AND2_X1 U13043 ( .A1(n20079), .A2(n12654), .ZN(n20050) );
  OAI22_X1 U13044 ( .A1(n14867), .A2(n14608), .B1(n14400), .B2(n14626), .ZN(
        n12631) );
  INV_X1 U13045 ( .A(n14608), .ZN(n14614) );
  INV_X1 U13046 ( .A(n15992), .ZN(n14689) );
  AND2_X1 U13047 ( .A1(n14704), .A2(n13422), .ZN(n15988) );
  INV_X1 U13048 ( .A(n13177), .ZN(n20136) );
  AND2_X1 U13049 ( .A1(n20874), .A2(n20781), .ZN(n13113) );
  AND2_X1 U13050 ( .A1(n9847), .A2(n14569), .ZN(n15922) );
  NAND2_X1 U13051 ( .A1(n12170), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12205) );
  AND2_X1 U13052 ( .A1(n14617), .A2(n14618), .ZN(n14619) );
  NAND2_X1 U13053 ( .A1(n11987), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12008) );
  AND2_X1 U13054 ( .A1(n13129), .A2(n13128), .ZN(n20090) );
  AND2_X1 U13055 ( .A1(n16156), .A2(n20846), .ZN(n20159) );
  INV_X1 U13056 ( .A(n16070), .ZN(n16056) );
  INV_X1 U13057 ( .A(n20215), .ZN(n16095) );
  INV_X1 U13058 ( .A(n20224), .ZN(n20186) );
  INV_X1 U13059 ( .A(n13946), .ZN(n16114) );
  INV_X1 U13060 ( .A(n20269), .ZN(n20370) );
  NOR2_X1 U13061 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19990) );
  OAI22_X1 U13062 ( .A1(n13410), .A2(n13409), .B1(n20366), .B2(n20479), .ZN(
        n20271) );
  OR2_X1 U13063 ( .A1(n9817), .A2(n12694), .ZN(n20512) );
  INV_X1 U13064 ( .A(n20325), .ZN(n20326) );
  INV_X1 U13065 ( .A(n20356), .ZN(n20359) );
  AND2_X1 U13066 ( .A1(n20449), .A2(n20640), .ZN(n20442) );
  AND2_X1 U13067 ( .A1(n20449), .A2(n20533), .ZN(n20472) );
  INV_X1 U13068 ( .A(n20532), .ZN(n20503) );
  INV_X1 U13069 ( .A(n20607), .ZN(n20482) );
  NOR2_X2 U13070 ( .A1(n20580), .A2(n20512), .ZN(n20568) );
  INV_X1 U13071 ( .A(n20639), .ZN(n20602) );
  OAI22_X1 U13072 ( .A1(n20619), .A2(n20618), .B1(n20673), .B2(n20617), .ZN(
        n20635) );
  INV_X1 U13073 ( .A(n20608), .ZN(n20668) );
  OAI211_X1 U13074 ( .C1(n20706), .C2(n20682), .A(n20681), .B(n20680), .ZN(
        n20708) );
  INV_X1 U13075 ( .A(n20512), .ZN(n20640) );
  INV_X1 U13076 ( .A(n20554), .ZN(n20734) );
  INV_X1 U13077 ( .A(n20563), .ZN(n20752) );
  INV_X1 U13078 ( .A(n20572), .ZN(n20767) );
  INV_X1 U13079 ( .A(n20880), .ZN(n20781) );
  INV_X1 U13080 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21063) );
  NOR2_X1 U13081 ( .A1(n16397), .A2(n18965), .ZN(n12857) );
  OR2_X1 U13082 ( .A1(n13930), .A2(n13929), .ZN(n13931) );
  AND2_X1 U13083 ( .A1(n13536), .A2(n13535), .ZN(n19129) );
  INV_X1 U13084 ( .A(n13635), .ZN(n19147) );
  OR2_X1 U13085 ( .A1(n19981), .A2(n13534), .ZN(n19133) );
  AND2_X1 U13086 ( .A1(n13536), .A2(n13532), .ZN(n19109) );
  OR2_X1 U13087 ( .A1(n11483), .A2(n11482), .ZN(n13467) );
  OR2_X1 U13088 ( .A1(n11430), .A2(n11429), .ZN(n13261) );
  INV_X1 U13089 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n15119) );
  INV_X1 U13090 ( .A(n13505), .ZN(n19192) );
  NOR2_X4 U13091 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19206), .ZN(n19269) );
  INV_X1 U13092 ( .A(n12831), .ZN(n14372) );
  NAND2_X1 U13093 ( .A1(n15029), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15031) );
  NOR2_X1 U13094 ( .A1(n13990), .A2(n14002), .ZN(n13989) );
  NOR2_X1 U13095 ( .A1(n15675), .A2(n15676), .ZN(n16342) );
  AND2_X1 U13096 ( .A1(n11585), .A2(n15743), .ZN(n19289) );
  AND2_X1 U13097 ( .A1(n18957), .A2(n20977), .ZN(n19088) );
  AND2_X1 U13098 ( .A1(n16402), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16413) );
  OAI21_X1 U13099 ( .B1(n13522), .B2(n13521), .A(n13520), .ZN(n19345) );
  AND2_X1 U13100 ( .A1(n19354), .A2(n15124), .ZN(n13610) );
  NOR2_X2 U13101 ( .A1(n19577), .A2(n19518), .ZN(n19401) );
  NOR2_X2 U13102 ( .A1(n19483), .A2(n13742), .ZN(n19430) );
  NOR2_X2 U13103 ( .A1(n19518), .A2(n13742), .ZN(n19449) );
  NOR2_X2 U13104 ( .A1(n19483), .A2(n19696), .ZN(n19475) );
  INV_X1 U13105 ( .A(n19500), .ZN(n19505) );
  INV_X1 U13106 ( .A(n19561), .ZN(n19565) );
  NOR2_X2 U13107 ( .A1(n19720), .A2(n19577), .ZN(n19598) );
  INV_X1 U13108 ( .A(n19650), .ZN(n19653) );
  AND2_X1 U13109 ( .A1(n19938), .A2(n19944), .ZN(n19925) );
  NOR2_X1 U13110 ( .A1(n19720), .A2(n19696), .ZN(n19715) );
  INV_X1 U13111 ( .A(n9793), .ZN(n19777) );
  INV_X1 U13112 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20977) );
  INV_X1 U13113 ( .A(n19983), .ZN(n19976) );
  INV_X1 U13114 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19861) );
  NOR2_X1 U13115 ( .A1(n21158), .A2(n16599), .ZN(n16640) );
  NOR2_X1 U13116 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16700), .ZN(n16685) );
  NOR2_X1 U13117 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16767), .ZN(n16755) );
  INV_X1 U13118 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16795) );
  NOR2_X1 U13119 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16862), .ZN(n16839) );
  NOR2_X1 U13120 ( .A1(n12850), .A2(n12851), .ZN(n16935) );
  NAND2_X1 U13121 ( .A1(n17052), .A2(n10241), .ZN(n17023) );
  INV_X1 U13122 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17263) );
  INV_X1 U13123 ( .A(n17300), .ZN(n17295) );
  AND3_X1 U13124 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n17351), .ZN(n17338) );
  NOR2_X1 U13125 ( .A1(n17531), .A2(n17399), .ZN(n17393) );
  OAI211_X1 U13126 ( .C1(n10244), .C2(n18506), .A(n11094), .B(n11093), .ZN(
        n11297) );
  NOR2_X1 U13127 ( .A1(n17438), .A2(n18760), .ZN(n17435) );
  INV_X1 U13128 ( .A(n17769), .ZN(n17667) );
  NOR2_X2 U13129 ( .A1(n17919), .A2(n17410), .ZN(n17812) );
  NAND2_X1 U13130 ( .A1(n16479), .A2(n16478), .ZN(n16480) );
  INV_X1 U13131 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21108) );
  INV_X1 U13132 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17787) );
  XNOR2_X1 U13133 ( .A(n11123), .B(n11122), .ZN(n17832) );
  NOR2_X2 U13134 ( .A1(n18950), .A2(n13838), .ZN(n18220) );
  INV_X1 U13135 ( .A(n18230), .ZN(n18225) );
  NOR2_X1 U13136 ( .A1(n15818), .A2(n18245), .ZN(n18242) );
  NOR2_X1 U13137 ( .A1(n18626), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n18911) );
  INV_X1 U13138 ( .A(n18343), .ZN(n18342) );
  INV_X1 U13139 ( .A(n18354), .ZN(n18361) );
  INV_X1 U13140 ( .A(n18382), .ZN(n18384) );
  INV_X1 U13141 ( .A(n18435), .ZN(n18420) );
  INV_X1 U13142 ( .A(n18483), .ZN(n18508) );
  NOR2_X1 U13143 ( .A1(n18765), .A2(n18484), .ZN(n18534) );
  INV_X1 U13144 ( .A(n18587), .ZN(n18576) );
  INV_X1 U13145 ( .A(n18671), .ZN(n18620) );
  INV_X1 U13146 ( .A(n18784), .ZN(n18939) );
  INV_X1 U13147 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18936) );
  AND2_X1 U13148 ( .A1(n18945), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18829) );
  INV_X1 U13149 ( .A(U212), .ZN(n20886) );
  NAND2_X1 U13150 ( .A1(n13789), .A2(n14391), .ZN(n13114) );
  INV_X1 U13151 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20847) );
  OR2_X1 U13152 ( .A1(n14612), .A2(n12524), .ZN(n14608) );
  OR2_X1 U13153 ( .A1(n13425), .A2(n13411), .ZN(n15992) );
  INV_X1 U13154 ( .A(n13292), .ZN(n13690) );
  INV_X1 U13155 ( .A(n20104), .ZN(n20123) );
  NOR2_X1 U13156 ( .A1(n13114), .A2(n13113), .ZN(n13176) );
  OAI21_X1 U13157 ( .B1(n14619), .B2(n14523), .A(n9876), .ZN(n14854) );
  INV_X1 U13158 ( .A(n20228), .ZN(n16049) );
  AND2_X1 U13159 ( .A1(n20218), .A2(n13808), .ZN(n16082) );
  NAND2_X1 U13160 ( .A1(n13832), .A2(n13826), .ZN(n20224) );
  NOR2_X1 U13161 ( .A1(n20220), .A2(n20227), .ZN(n20218) );
  INV_X1 U13162 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20863) );
  OR2_X1 U13163 ( .A1(n20333), .A2(n20607), .ZN(n20292) );
  OR2_X1 U13164 ( .A1(n20333), .A2(n20512), .ZN(n20325) );
  NAND2_X1 U13165 ( .A1(n20303), .A2(n20533), .ZN(n20356) );
  OR2_X1 U13166 ( .A1(n20333), .A2(n20448), .ZN(n20387) );
  NAND2_X1 U13167 ( .A1(n20449), .A2(n20482), .ZN(n20417) );
  AOI22_X1 U13168 ( .A1(n20426), .A2(n20423), .B1(n20422), .B2(n20421), .ZN(
        n20447) );
  NAND2_X1 U13169 ( .A1(n20449), .A2(n20583), .ZN(n20507) );
  NAND2_X1 U13170 ( .A1(n20584), .A2(n20482), .ZN(n20532) );
  AOI22_X1 U13171 ( .A1(n20544), .A2(n20540), .B1(n20538), .B2(n20537), .ZN(
        n20573) );
  INV_X1 U13172 ( .A(n20587), .ZN(n20606) );
  NAND2_X1 U13173 ( .A1(n20584), .A2(n20583), .ZN(n20639) );
  NAND2_X1 U13174 ( .A1(n20854), .A2(n20640), .ZN(n20711) );
  OR2_X1 U13175 ( .A1(n20676), .A2(n20675), .ZN(n20764) );
  INV_X1 U13176 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20615) );
  INV_X1 U13177 ( .A(n20844), .ZN(n20780) );
  AND2_X1 U13178 ( .A1(n21063), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20873) );
  INV_X1 U13179 ( .A(n20834), .ZN(n20832) );
  NAND2_X1 U13180 ( .A1(n13539), .A2(n18958), .ZN(n19981) );
  NAND2_X1 U13181 ( .A1(n11354), .A2(n12857), .ZN(n18967) );
  NAND2_X1 U13182 ( .A1(n13531), .A2(n13530), .ZN(n19150) );
  OR2_X1 U13183 ( .A1(n16398), .A2(n19202), .ZN(n18958) );
  NAND2_X1 U13184 ( .A1(n12955), .A2(n12969), .ZN(n15212) );
  INV_X1 U13185 ( .A(n15212), .ZN(n15224) );
  INV_X1 U13186 ( .A(n19190), .ZN(n15286) );
  NOR2_X1 U13187 ( .A1(n19194), .A2(n16246), .ZN(n19200) );
  OR2_X1 U13188 ( .A1(n19190), .A2(n12971), .ZN(n13505) );
  NAND2_X1 U13189 ( .A1(n19270), .A2(n19208), .ZN(n19237) );
  INV_X1 U13190 ( .A(n19270), .ZN(n19267) );
  INV_X1 U13191 ( .A(n12905), .ZN(n12989) );
  INV_X1 U13192 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19085) );
  INV_X1 U13193 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16298) );
  INV_X1 U13194 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19287) );
  INV_X1 U13195 ( .A(n16337), .ZN(n19295) );
  INV_X1 U13196 ( .A(n19303), .ZN(n16369) );
  AOI21_X1 U13197 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15883), .A(n15707), .ZN(
        n15795) );
  INV_X1 U13198 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19313) );
  AND2_X1 U13199 ( .A1(n13513), .A2(n13512), .ZN(n19349) );
  NAND2_X1 U13200 ( .A1(n19355), .A2(n13610), .ZN(n19373) );
  AOI211_X2 U13201 ( .C1(n13615), .C2(n19924), .A(n9793), .B(n13614), .ZN(
        n19405) );
  AOI21_X1 U13202 ( .B1(n19412), .B2(n19410), .A(n19409), .ZN(n19434) );
  AOI211_X2 U13203 ( .C1(n13747), .C2(n13750), .A(n9793), .B(n13746), .ZN(
        n19452) );
  AOI21_X1 U13204 ( .B1(n19459), .B2(n19454), .A(n19453), .ZN(n19479) );
  OR2_X1 U13205 ( .A1(n19518), .A2(n19696), .ZN(n19500) );
  INV_X1 U13206 ( .A(n19535), .ZN(n19531) );
  OR2_X1 U13207 ( .A1(n19518), .A2(n19719), .ZN(n19561) );
  AND2_X1 U13208 ( .A1(n19576), .A2(n19575), .ZN(n19599) );
  INV_X1 U13209 ( .A(n19633), .ZN(n19628) );
  NAND2_X1 U13210 ( .A1(n13571), .A2(n19925), .ZN(n19650) );
  NAND2_X1 U13211 ( .A1(n13572), .A2(n19925), .ZN(n19676) );
  INV_X1 U13212 ( .A(n19715), .ZN(n19710) );
  AOI21_X1 U13213 ( .B1(n19729), .B2(n19726), .A(n19725), .ZN(n19768) );
  INV_X1 U13214 ( .A(n19830), .ZN(n19817) );
  NAND2_X1 U13215 ( .A1(n13572), .A2(n19781), .ZN(n19834) );
  INV_X1 U13216 ( .A(n19922), .ZN(n19843) );
  INV_X1 U13217 ( .A(n16946), .ZN(n18953) );
  INV_X1 U13218 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16580) );
  INV_X1 U13219 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16823) );
  INV_X1 U13220 ( .A(n16955), .ZN(n16942) );
  NOR2_X1 U13221 ( .A1(n16967), .A2(n16966), .ZN(n16994) );
  NAND2_X1 U13222 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17247), .ZN(n17227) );
  INV_X1 U13223 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17264) );
  AND2_X1 U13224 ( .A1(n17284), .A2(n17333), .ZN(n17281) );
  INV_X1 U13225 ( .A(n16471), .ZN(n17410) );
  INV_X1 U13226 ( .A(n17434), .ZN(n17422) );
  NAND2_X1 U13227 ( .A1(n17461), .A2(n17444), .ZN(n17460) );
  INV_X1 U13228 ( .A(n17461), .ZN(n17479) );
  INV_X1 U13229 ( .A(n17635), .ZN(n17719) );
  INV_X1 U13230 ( .A(n17812), .ZN(n17823) );
  INV_X1 U13231 ( .A(n11274), .ZN(n17919) );
  NAND2_X1 U13232 ( .A1(n16480), .A2(n16718), .ZN(n16490) );
  INV_X1 U13233 ( .A(n16718), .ZN(n18140) );
  INV_X1 U13234 ( .A(n18139), .ZN(n18161) );
  INV_X1 U13235 ( .A(n18242), .ZN(n18238) );
  INV_X1 U13236 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18765) );
  INV_X1 U13237 ( .A(n18409), .ZN(n18407) );
  INV_X1 U13238 ( .A(n18450), .ZN(n18457) );
  INV_X1 U13239 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18463) );
  INV_X1 U13240 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n20981) );
  INV_X1 U13241 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18500) );
  INV_X1 U13242 ( .A(n18534), .ZN(n18527) );
  INV_X1 U13243 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18542) );
  INV_X1 U13244 ( .A(n18558), .ZN(n18553) );
  INV_X1 U13245 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n21111) );
  INV_X1 U13246 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18618) );
  INV_X1 U13247 ( .A(n18700), .ZN(n18648) );
  INV_X1 U13248 ( .A(n18631), .ZN(n18677) );
  INV_X1 U13249 ( .A(n18691), .ZN(n18720) );
  INV_X1 U13250 ( .A(n16941), .ZN(n18800) );
  INV_X1 U13251 ( .A(n18888), .ZN(n18805) );
  INV_X1 U13252 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18820) );
  INV_X1 U13253 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18837) );
  NOR2_X1 U13254 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12832), .ZN(n16569)
         );
  INV_X1 U13255 ( .A(n20887), .ZN(n16536) );
  INV_X1 U13256 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n21024) );
  OAI21_X1 U13257 ( .B1(n12633), .B2(n14627), .A(n12632), .ZN(P1_U2842) );
  OR4_X1 U13258 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n12853), .ZN(
        P3_U2645) );
  NOR2_X4 U13259 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15709) );
  AND2_X4 U13260 ( .A1(n15709), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10541) );
  AND3_X4 U13261 ( .A1(n10379), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U13262 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10254) );
  INV_X2 U13263 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16370) );
  AND2_X4 U13264 ( .A1(n15710), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10544) );
  AOI22_X1 U13265 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10253) );
  AND2_X4 U13266 ( .A1(n15709), .A2(n16370), .ZN(n10545) );
  AND2_X2 U13267 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15722) );
  AND2_X4 U13268 ( .A1(n15722), .A2(n15693), .ZN(n10542) );
  AOI22_X1 U13269 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10252) );
  AND2_X4 U13270 ( .A1(n15733), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10550) );
  AOI22_X1 U13271 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10251) );
  NAND4_X1 U13272 ( .A1(n10254), .A2(n10253), .A3(n10252), .A4(n10251), .ZN(
        n10255) );
  AOI22_X1 U13273 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U13274 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13275 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13276 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10256) );
  NAND4_X1 U13277 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10260) );
  AOI22_X1 U13278 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13279 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U13280 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U13281 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10263) );
  NAND4_X1 U13282 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(n10263), .ZN(
        n10267) );
  NAND2_X1 U13283 ( .A1(n10267), .A2(n16379), .ZN(n10274) );
  AOI22_X1 U13284 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U13285 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U13286 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10268) );
  NAND4_X1 U13287 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n10272) );
  NAND2_X1 U13288 ( .A1(n10272), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10273) );
  NAND2_X4 U13289 ( .A1(n10274), .A2(n10273), .ZN(n12972) );
  INV_X1 U13290 ( .A(n10358), .ZN(n14371) );
  AOI22_X1 U13291 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13292 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13293 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13294 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13295 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13296 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13297 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U13298 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U13299 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13300 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13301 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13302 ( .A1(n10542), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13303 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13304 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13305 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13306 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13307 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U13308 ( .A1(n10295), .A2(n16379), .ZN(n10302) );
  AOI22_X1 U13309 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13310 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13311 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U13312 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10298) );
  INV_X1 U13313 ( .A(n10354), .ZN(n10371) );
  AOI22_X1 U13314 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13315 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13316 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13317 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10303) );
  NAND4_X1 U13318 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10307) );
  AOI22_X1 U13319 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13320 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13321 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13322 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10309) );
  NAND4_X1 U13323 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n10309), .ZN(
        n10313) );
  NAND2_X1 U13324 ( .A1(n10313), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10314) );
  NOR2_X1 U13325 ( .A1(n10371), .A2(n10344), .ZN(n10316) );
  AOI22_X1 U13326 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13327 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13328 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13329 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10318) );
  NAND4_X1 U13330 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10327) );
  AOI22_X1 U13331 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13332 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13333 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10322) );
  NAND4_X1 U13334 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10326) );
  MUX2_X2 U13335 ( .A(n10327), .B(n10326), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19971) );
  INV_X4 U13336 ( .A(n19971), .ZN(n16397) );
  INV_X1 U13337 ( .A(n16397), .ZN(n10540) );
  AOI22_X1 U13338 ( .A1(n10308), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13339 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13340 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13341 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10329) );
  NAND4_X1 U13342 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10333) );
  NAND2_X1 U13343 ( .A1(n10333), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10340) );
  AOI22_X1 U13344 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13345 ( .A1(n10541), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13346 ( .A1(n10550), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10335) );
  NAND4_X1 U13347 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n10338) );
  INV_X2 U13348 ( .A(n10343), .ZN(n10768) );
  NAND2_X2 U13349 ( .A1(n10372), .A2(n10768), .ZN(n11367) );
  NAND2_X1 U13350 ( .A1(n11367), .A2(n10344), .ZN(n10365) );
  INV_X2 U13351 ( .A(n10345), .ZN(n10942) );
  NAND3_X1 U13352 ( .A1(n10942), .A2(n10372), .A3(n16397), .ZN(n10347) );
  NAND2_X1 U13353 ( .A1(n10347), .A2(n10346), .ZN(n10348) );
  NAND2_X1 U13354 ( .A1(n10365), .A2(n10348), .ZN(n10349) );
  NOR2_X4 U13355 ( .A1(n10350), .A2(n10349), .ZN(n11361) );
  NAND2_X1 U13356 ( .A1(n11361), .A2(n11549), .ZN(n10400) );
  INV_X1 U13357 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10357) );
  NOR2_X1 U13358 ( .A1(n13570), .A2(n20977), .ZN(n12959) );
  CLKBUF_X3 U13359 ( .A(n10368), .Z(n14316) );
  NAND2_X1 U13360 ( .A1(n12959), .A2(n14316), .ZN(n13036) );
  AND2_X4 U13362 ( .A1(n10328), .A2(n10353), .ZN(n14030) );
  AOI22_X1 U13363 ( .A1(n14030), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10356) );
  INV_X1 U13364 ( .A(n11582), .ZN(n10376) );
  NAND2_X1 U13365 ( .A1(n11549), .A2(n10376), .ZN(n10396) );
  NOR2_X2 U13366 ( .A1(n10396), .A2(n11545), .ZN(n11562) );
  AND2_X4 U13367 ( .A1(n11562), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14031) );
  NAND2_X1 U13368 ( .A1(n14031), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10355) );
  INV_X1 U13369 ( .A(n10385), .ZN(n10384) );
  NOR2_X1 U13370 ( .A1(n10358), .A2(n10942), .ZN(n10359) );
  NAND2_X1 U13371 ( .A1(n10360), .A2(n10359), .ZN(n10538) );
  NOR2_X1 U13372 ( .A1(n19970), .A2(n11334), .ZN(n10361) );
  NAND2_X1 U13373 ( .A1(n10538), .A2(n10361), .ZN(n10362) );
  NAND2_X1 U13374 ( .A1(n10363), .A2(n10540), .ZN(n10370) );
  NAND3_X1 U13375 ( .A1(n10365), .A2(n10364), .A3(n12972), .ZN(n10367) );
  MUX2_X1 U13376 ( .A(n10354), .B(n10768), .S(n13570), .Z(n10366) );
  NAND2_X1 U13377 ( .A1(n10391), .A2(n11555), .ZN(n10369) );
  NAND3_X1 U13378 ( .A1(n10370), .A2(n11553), .A3(n10369), .ZN(n10393) );
  INV_X1 U13379 ( .A(n10393), .ZN(n10378) );
  NAND2_X1 U13380 ( .A1(n11367), .A2(n10371), .ZN(n11341) );
  AND2_X1 U13381 ( .A1(n11341), .A2(n12972), .ZN(n10373) );
  NAND2_X1 U13382 ( .A1(n11346), .A2(n10354), .ZN(n11347) );
  NAND2_X1 U13383 ( .A1(n11557), .A2(n10344), .ZN(n10375) );
  NAND2_X1 U13384 ( .A1(n10392), .A2(n10376), .ZN(n10377) );
  NAND2_X1 U13385 ( .A1(n10378), .A2(n10377), .ZN(n10399) );
  NAND2_X1 U13386 ( .A1(n10399), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10413) );
  NOR2_X1 U13387 ( .A1(n19980), .A2(n19950), .ZN(n10381) );
  OAI21_X2 U13388 ( .B1(n10413), .B2(n15711), .A(n10382), .ZN(n10386) );
  INV_X1 U13389 ( .A(n10386), .ZN(n10383) );
  NAND2_X2 U13390 ( .A1(n10384), .A2(n10383), .ZN(n10405) );
  NAND2_X1 U13391 ( .A1(n10386), .A2(n10385), .ZN(n10387) );
  NAND2_X1 U13392 ( .A1(n14030), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10390) );
  NAND2_X1 U13393 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10388) );
  INV_X1 U13394 ( .A(n10391), .ZN(n12967) );
  AND2_X1 U13395 ( .A1(n10392), .A2(n10391), .ZN(n10394) );
  OAI21_X1 U13396 ( .B1(n10394), .B2(n10393), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10395) );
  INV_X1 U13397 ( .A(n10396), .ZN(n10398) );
  AND2_X1 U13398 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10397) );
  OAI22_X1 U13399 ( .A1(n10399), .A2(n10398), .B1(n14031), .B2(n10397), .ZN(
        n10404) );
  INV_X1 U13400 ( .A(n15728), .ZN(n10402) );
  NOR2_X1 U13401 ( .A1(n19980), .A2(n19958), .ZN(n10401) );
  AOI21_X1 U13402 ( .B1(n10402), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10401), 
        .ZN(n10403) );
  NAND2_X1 U13403 ( .A1(n10404), .A2(n10403), .ZN(n10613) );
  INV_X4 U13404 ( .A(n10406), .ZN(n10509) );
  NAND2_X1 U13405 ( .A1(n14030), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10409) );
  INV_X1 U13406 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10407) );
  AOI21_X1 U13407 ( .B1(n14031), .B2(P2_EBX_REG_2__SCAN_IN), .A(n10249), .ZN(
        n10408) );
  NAND2_X1 U13408 ( .A1(n10409), .A2(n10408), .ZN(n10410) );
  AOI21_X2 U13409 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10410), .ZN(n10621) );
  INV_X1 U13410 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16356) );
  AOI22_X1 U13411 ( .A1(n14030), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10412) );
  NAND2_X1 U13412 ( .A1(n14031), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10411) );
  INV_X1 U13413 ( .A(n10606), .ZN(n10609) );
  OAI21_X1 U13414 ( .B1(n10417), .B2(n10621), .A(n10609), .ZN(n10422) );
  INV_X1 U13415 ( .A(n10413), .ZN(n10414) );
  NAND2_X1 U13416 ( .A1(n10414), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10416) );
  AOI21_X1 U13417 ( .B1(n20977), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10415) );
  INV_X1 U13418 ( .A(n10622), .ZN(n10601) );
  AOI21_X1 U13419 ( .B1(n10417), .B2(n10621), .A(n10601), .ZN(n10421) );
  OR2_X1 U13420 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  OAI21_X1 U13421 ( .B1(n10422), .B2(n10421), .A(n10420), .ZN(n10423) );
  INV_X1 U13422 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13482) );
  AOI22_X1 U13423 ( .A1(n14030), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10426) );
  NAND2_X1 U13424 ( .A1(n14031), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10425) );
  OAI211_X1 U13425 ( .C1(n10406), .C2(n13482), .A(n10426), .B(n10425), .ZN(
        n13200) );
  NAND2_X1 U13426 ( .A1(n13199), .A2(n13200), .ZN(n13269) );
  INV_X1 U13427 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10429) );
  NAND2_X1 U13428 ( .A1(n14030), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10428) );
  NAND2_X1 U13429 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10427) );
  OAI211_X1 U13430 ( .C1(n10507), .C2(n10429), .A(n10428), .B(n10427), .ZN(
        n10430) );
  AOI21_X1 U13431 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10430), .ZN(n13268) );
  INV_X1 U13432 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15675) );
  AOI22_X1 U13433 ( .A1(n14030), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10432) );
  NAND2_X1 U13434 ( .A1(n14031), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10431) );
  OAI211_X1 U13435 ( .C1(n10406), .C2(n15675), .A(n10432), .B(n10431), .ZN(
        n13309) );
  INV_X1 U13436 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U13437 ( .A1(n14030), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10434) );
  NAND2_X1 U13438 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10433) );
  OAI211_X1 U13439 ( .C1(n10507), .C2(n10847), .A(n10434), .B(n10433), .ZN(
        n10435) );
  AOI21_X1 U13440 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10435), .ZN(n13342) );
  INV_X1 U13441 ( .A(n13182), .ZN(n10441) );
  INV_X1 U13442 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U13443 ( .A1(n14030), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10437) );
  NAND2_X1 U13444 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10436) );
  OAI211_X1 U13445 ( .C1(n10507), .C2(n10438), .A(n10437), .B(n10436), .ZN(
        n10439) );
  AOI21_X1 U13446 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10439), .ZN(n13183) );
  NAND2_X1 U13447 ( .A1(n14030), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10443) );
  NAND2_X1 U13448 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10442) );
  OAI211_X1 U13449 ( .C1(n10507), .C2(n10008), .A(n10443), .B(n10442), .ZN(
        n10444) );
  AOI21_X1 U13450 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10444), .ZN(n13262) );
  INV_X1 U13451 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16278) );
  AOI22_X1 U13452 ( .A1(n14030), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10446) );
  NAND2_X1 U13453 ( .A1(n14031), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10445) );
  OAI211_X1 U13454 ( .C1(n10424), .C2(n16278), .A(n10446), .B(n10445), .ZN(
        n13210) );
  NAND2_X1 U13455 ( .A1(n13264), .A2(n13210), .ZN(n13326) );
  INV_X1 U13456 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10449) );
  NAND2_X1 U13457 ( .A1(n14030), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10448) );
  NAND2_X1 U13458 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10447) );
  OAI211_X1 U13459 ( .C1(n10507), .C2(n10449), .A(n10448), .B(n10447), .ZN(
        n10450) );
  AOI21_X1 U13460 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10450), .ZN(n13325) );
  INV_X1 U13461 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10454) );
  NAND2_X1 U13462 ( .A1(n14030), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10453) );
  NAND2_X1 U13463 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10452) );
  OAI211_X1 U13464 ( .C1(n10507), .C2(n10454), .A(n10453), .B(n10452), .ZN(
        n10455) );
  AOI21_X1 U13465 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10455), .ZN(n13389) );
  INV_X1 U13466 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13467 ( .A1(n14030), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10457) );
  NAND2_X1 U13468 ( .A1(n14031), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10456) );
  OAI211_X1 U13469 ( .C1(n10424), .C2(n10895), .A(n10457), .B(n10456), .ZN(
        n13459) );
  INV_X1 U13470 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15588) );
  AOI22_X1 U13471 ( .A1(n14030), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10459) );
  NAND2_X1 U13472 ( .A1(n14031), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10458) );
  OAI211_X1 U13473 ( .C1(n10424), .C2(n15588), .A(n10459), .B(n10458), .ZN(
        n13464) );
  INV_X1 U13474 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U13475 ( .A1(n14030), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U13476 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10460) );
  OAI211_X1 U13477 ( .C1(n10507), .C2(n10462), .A(n10461), .B(n10460), .ZN(
        n10463) );
  AOI21_X1 U13478 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10463), .ZN(n15218) );
  INV_X1 U13479 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n15213) );
  NAND2_X1 U13480 ( .A1(n14030), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10466) );
  NAND2_X1 U13481 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10465) );
  OAI211_X1 U13482 ( .C1(n10507), .C2(n15213), .A(n10466), .B(n10465), .ZN(
        n10467) );
  AOI21_X1 U13483 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10467), .ZN(n15100) );
  INV_X1 U13484 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U13485 ( .A1(n14030), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U13486 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10468) );
  OAI211_X1 U13487 ( .C1(n10507), .C2(n10470), .A(n10469), .B(n10468), .ZN(
        n10471) );
  AOI21_X1 U13488 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10471), .ZN(n15207) );
  INV_X1 U13489 ( .A(n15207), .ZN(n10472) );
  INV_X1 U13490 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15377) );
  AOI22_X1 U13491 ( .A1(n14030), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10474) );
  NAND2_X1 U13492 ( .A1(n14031), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10473) );
  OAI211_X1 U13493 ( .C1(n10424), .C2(n15377), .A(n10474), .B(n10473), .ZN(
        n15084) );
  INV_X1 U13494 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10879) );
  NAND2_X1 U13495 ( .A1(n14030), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10476) );
  NAND2_X1 U13496 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10475) );
  OAI211_X1 U13497 ( .C1(n10507), .C2(n10879), .A(n10476), .B(n10475), .ZN(
        n10477) );
  AOI21_X1 U13498 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10477), .ZN(n15190) );
  INV_X1 U13499 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15189) );
  NAND2_X1 U13500 ( .A1(n14030), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10479) );
  NAND2_X1 U13501 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10478) );
  OAI211_X1 U13502 ( .C1(n10507), .C2(n15189), .A(n10479), .B(n10478), .ZN(
        n10480) );
  AOI21_X1 U13503 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10480), .ZN(n15185) );
  INV_X1 U13504 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U13505 ( .A1(n14030), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10482) );
  NAND2_X1 U13506 ( .A1(n14031), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10481) );
  OAI211_X1 U13507 ( .C1(n10424), .C2(n11612), .A(n10482), .B(n10481), .ZN(
        n11606) );
  INV_X1 U13508 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n10485) );
  NAND2_X1 U13509 ( .A1(n14030), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10484) );
  NAND2_X1 U13510 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10483) );
  OAI211_X1 U13511 ( .C1(n10507), .C2(n10485), .A(n10484), .B(n10483), .ZN(
        n10486) );
  AOI21_X1 U13512 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10486), .ZN(n15170) );
  INV_X1 U13513 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U13514 ( .A1(n14030), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U13515 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10487) );
  OAI211_X1 U13516 ( .C1(n10507), .C2(n10489), .A(n10488), .B(n10487), .ZN(
        n10490) );
  AOI21_X1 U13517 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10490), .ZN(n15165) );
  AOI22_X1 U13518 ( .A1(n14030), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10492) );
  NAND2_X1 U13519 ( .A1(n14031), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10491) );
  OAI211_X1 U13520 ( .C1(n10424), .C2(n15474), .A(n10492), .B(n10491), .ZN(
        n15072) );
  INV_X1 U13521 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15325) );
  AOI22_X1 U13522 ( .A1(n14030), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10494) );
  NAND2_X1 U13523 ( .A1(n14031), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10493) );
  OAI211_X1 U13524 ( .C1(n10424), .C2(n15325), .A(n10494), .B(n10493), .ZN(
        n15153) );
  NAND2_X1 U13525 ( .A1(n15070), .A2(n15153), .ZN(n15141) );
  INV_X1 U13526 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10497) );
  NAND2_X1 U13527 ( .A1(n14030), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10496) );
  NAND2_X1 U13528 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10495) );
  OAI211_X1 U13529 ( .C1(n10507), .C2(n10497), .A(n10496), .B(n10495), .ZN(
        n10498) );
  AOI21_X1 U13530 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10498), .ZN(n15142) );
  INV_X1 U13531 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n10501) );
  NAND2_X1 U13532 ( .A1(n14030), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10500) );
  NAND2_X1 U13533 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10499) );
  OAI211_X1 U13534 ( .C1(n10507), .C2(n10501), .A(n10500), .B(n10499), .ZN(
        n10502) );
  AOI21_X1 U13535 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10502), .ZN(n13996) );
  INV_X1 U13536 ( .A(n13996), .ZN(n10503) );
  INV_X1 U13537 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U13538 ( .A1(n14030), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10505) );
  NAND2_X1 U13539 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10504) );
  OAI211_X1 U13540 ( .C1(n10507), .C2(n10506), .A(n10505), .B(n10504), .ZN(
        n10508) );
  AOI21_X1 U13541 ( .B1(n10509), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10508), .ZN(n13969) );
  INV_X1 U13542 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U13543 ( .A1(n14030), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10511) );
  NAND2_X1 U13544 ( .A1(n14031), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10510) );
  OAI211_X1 U13545 ( .C1(n10424), .C2(n11000), .A(n10511), .B(n10510), .ZN(
        n10512) );
  NOR2_X1 U13546 ( .A1(n9852), .A2(n10512), .ZN(n10513) );
  OAI21_X1 U13547 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19958), .A(
        n10531), .ZN(n11314) );
  XNOR2_X1 U13548 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10586) );
  INV_X1 U13549 ( .A(n10531), .ZN(n10514) );
  NAND2_X1 U13550 ( .A1(n10586), .A2(n10514), .ZN(n10516) );
  NAND2_X1 U13551 ( .A1(n19950), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10515) );
  NAND2_X1 U13552 ( .A1(n10516), .A2(n10515), .ZN(n10526) );
  MUX2_X1 U13553 ( .A(n13038), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10525) );
  NAND2_X1 U13554 ( .A1(n10526), .A2(n10525), .ZN(n10518) );
  NAND2_X1 U13555 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13038), .ZN(
        n10517) );
  NAND2_X1 U13556 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  INV_X1 U13557 ( .A(n10527), .ZN(n10524) );
  INV_X1 U13558 ( .A(n10519), .ZN(n10522) );
  INV_X1 U13559 ( .A(n10520), .ZN(n10521) );
  NAND2_X1 U13560 ( .A1(n10522), .A2(n10521), .ZN(n10523) );
  NAND2_X1 U13561 ( .A1(n10524), .A2(n10523), .ZN(n11321) );
  XNOR2_X1 U13562 ( .A(n10526), .B(n10525), .ZN(n11319) );
  NAND3_X1 U13563 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10530), .A3(
        n11329), .ZN(n11310) );
  INV_X1 U13564 ( .A(n11310), .ZN(n10528) );
  NOR3_X1 U13565 ( .A1(n11321), .A2(n11319), .A3(n10528), .ZN(n10532) );
  INV_X1 U13566 ( .A(n10532), .ZN(n10535) );
  NOR2_X1 U13567 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15885), .ZN(
        n10529) );
  XNOR2_X1 U13568 ( .A(n10586), .B(n10531), .ZN(n11315) );
  AND2_X1 U13569 ( .A1(n11315), .A2(n10532), .ZN(n10533) );
  INV_X1 U13570 ( .A(n16398), .ZN(n10534) );
  OAI21_X1 U13571 ( .B1(n11314), .B2(n10535), .A(n10534), .ZN(n10537) );
  AND2_X2 U13572 ( .A1(n14357), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10573) );
  INV_X1 U13573 ( .A(n10573), .ZN(n10536) );
  NAND3_X1 U13574 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10552) );
  AND2_X1 U13575 ( .A1(n11329), .A2(n10552), .ZN(n16391) );
  AOI21_X1 U13576 ( .B1(n10536), .B2(n16391), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n16417) );
  MUX2_X1 U13577 ( .A(n10537), .B(n16417), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19964) );
  INV_X1 U13578 ( .A(n10538), .ZN(n10539) );
  NAND2_X1 U13579 ( .A1(n10539), .A2(n14316), .ZN(n10590) );
  NAND2_X1 U13580 ( .A1(n10540), .A2(n14294), .ZN(n19969) );
  AOI22_X1 U13581 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10549) );
  INV_X1 U13582 ( .A(n14272), .ZN(n10543) );
  AND2_X2 U13583 ( .A1(n9807), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14130) );
  AND2_X2 U13584 ( .A1(n14352), .A2(n16379), .ZN(n14142) );
  AOI22_X1 U13585 ( .A1(n14130), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14142), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10548) );
  AND2_X1 U13586 ( .A1(n14351), .A2(n16379), .ZN(n10676) );
  AND2_X2 U13587 ( .A1(n14352), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10684) );
  AOI22_X1 U13588 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14143), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13589 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10546) );
  NAND4_X1 U13590 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10559) );
  INV_X1 U13591 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14261) );
  AND2_X2 U13592 ( .A1(n14359), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10685) );
  INV_X1 U13593 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14269) );
  OAI22_X1 U13594 ( .A1(n14261), .A2(n10668), .B1(n10738), .B2(n14269), .ZN(
        n10551) );
  INV_X1 U13595 ( .A(n10551), .ZN(n10557) );
  INV_X1 U13596 ( .A(n10552), .ZN(n10553) );
  AOI22_X1 U13597 ( .A1(n10677), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n14151), .ZN(n10556) );
  AOI22_X1 U13598 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10555) );
  AND2_X1 U13599 ( .A1(n14358), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10565) );
  AOI22_X1 U13600 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10669), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10554) );
  NAND4_X1 U13601 ( .A1(n10557), .A2(n10556), .A3(n10555), .A4(n10554), .ZN(
        n10558) );
  MUX2_X1 U13602 ( .A(n11397), .B(n11310), .S(n11582), .Z(n10770) );
  AOI22_X1 U13603 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13604 ( .A1(n10679), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13605 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13606 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14142), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10561) );
  NAND4_X1 U13607 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n10571) );
  AOI22_X1 U13608 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n14151), .ZN(n10569) );
  INV_X1 U13609 ( .A(n10686), .ZN(n10668) );
  AOI22_X1 U13610 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13611 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13612 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10566) );
  NAND4_X1 U13613 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10570) );
  INV_X1 U13614 ( .A(n11321), .ZN(n10572) );
  MUX2_X1 U13615 ( .A(n11392), .B(n10572), .S(n11582), .Z(n10773) );
  NAND2_X1 U13616 ( .A1(n10770), .A2(n10773), .ZN(n11325) );
  INV_X1 U13617 ( .A(n11319), .ZN(n10585) );
  AOI22_X1 U13618 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14142), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13619 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n14151), .ZN(n10577) );
  AOI22_X1 U13620 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13621 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U13622 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10669), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13623 ( .A1(n14130), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U13624 ( .A1(n10679), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10578) );
  INV_X1 U13625 ( .A(n10578), .ZN(n10581) );
  AOI22_X1 U13626 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10676), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10579) );
  INV_X1 U13627 ( .A(n10579), .ZN(n10580) );
  NAND4_X1 U13628 ( .A1(n10584), .A2(n10230), .A3(n10583), .A4(n10582), .ZN(
        n11383) );
  MUX2_X1 U13629 ( .A(n10585), .B(n11383), .S(n10376), .Z(n10771) );
  INV_X1 U13630 ( .A(n10586), .ZN(n11313) );
  NOR2_X1 U13631 ( .A1(n11313), .A2(n11314), .ZN(n10587) );
  NOR2_X1 U13632 ( .A1(n10771), .A2(n10587), .ZN(n10588) );
  NOR2_X1 U13633 ( .A1(n11325), .A2(n10588), .ZN(n10589) );
  OR2_X1 U13634 ( .A1(n10589), .A2(n11332), .ZN(n19961) );
  NOR2_X1 U13635 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15719) );
  OR2_X1 U13636 ( .A1(n19924), .A2(n15719), .ZN(n19954) );
  NAND2_X1 U13637 ( .A1(n19954), .A2(n20977), .ZN(n10591) );
  AND2_X1 U13638 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19942) );
  NOR2_X1 U13639 ( .A1(n15125), .A2(n16317), .ZN(n10600) );
  INV_X1 U13640 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10596) );
  NAND2_X1 U13641 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13443), .ZN(
        n13623) );
  AND2_X1 U13642 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U13643 ( .A1(n15046), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15048) );
  INV_X1 U13644 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13979) );
  AOI21_X1 U13645 ( .B1(n10596), .B2(n13981), .A(n15050), .ZN(n15020) );
  INV_X1 U13646 ( .A(n13141), .ZN(n10595) );
  INV_X1 U13647 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n10593) );
  NAND2_X1 U13648 ( .A1(n10593), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10594) );
  NAND2_X1 U13649 ( .A1(n10595), .A2(n10594), .ZN(n12867) );
  INV_X1 U13650 ( .A(n19977), .ZN(n13510) );
  NOR2_X1 U13651 ( .A1(n13510), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18957) );
  NAND2_X1 U13652 ( .A1(n19088), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11566) );
  OAI21_X1 U13653 ( .B1(n19288), .B2(n10596), .A(n11566), .ZN(n10597) );
  AOI21_X1 U13654 ( .B1(n15020), .B2(n19274), .A(n10597), .ZN(n10598) );
  INV_X1 U13655 ( .A(n10598), .ZN(n10599) );
  INV_X1 U13656 ( .A(n10417), .ZN(n10602) );
  NAND3_X1 U13657 ( .A1(n10602), .A2(n10606), .A3(n10603), .ZN(n10612) );
  INV_X1 U13658 ( .A(n10603), .ZN(n10607) );
  INV_X1 U13659 ( .A(n10621), .ZN(n10604) );
  NAND2_X1 U13660 ( .A1(n10622), .A2(n10604), .ZN(n10608) );
  NAND2_X1 U13661 ( .A1(n10608), .A2(n10606), .ZN(n10605) );
  NAND3_X1 U13662 ( .A1(n10417), .A2(n10609), .A3(n10608), .ZN(n10610) );
  NAND3_X2 U13663 ( .A1(n10612), .A2(n10611), .A3(n10610), .ZN(n13140) );
  NAND2_X1 U13664 ( .A1(n13140), .A2(n10073), .ZN(n10640) );
  INV_X1 U13665 ( .A(n10640), .ZN(n10620) );
  INV_X1 U13666 ( .A(n10615), .ZN(n10624) );
  NAND2_X1 U13667 ( .A1(n10624), .A2(n10616), .ZN(n10618) );
  INV_X1 U13668 ( .A(n13712), .ZN(n10619) );
  XNOR2_X1 U13669 ( .A(n10622), .B(n10621), .ZN(n10623) );
  XNOR2_X2 U13670 ( .A(n10417), .B(n10623), .ZN(n13037) );
  INV_X1 U13671 ( .A(n10705), .ZN(n10721) );
  INV_X1 U13672 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10625) );
  AND2_X2 U13673 ( .A1(n13154), .A2(n13037), .ZN(n10635) );
  INV_X1 U13674 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14183) );
  OAI22_X1 U13675 ( .A1(n10721), .A2(n10625), .B1(n19456), .B2(n14183), .ZN(
        n10633) );
  NOR2_X1 U13676 ( .A1(n13712), .A2(n15695), .ZN(n10648) );
  INV_X1 U13677 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14181) );
  INV_X1 U13678 ( .A(n13037), .ZN(n10626) );
  NAND2_X2 U13679 ( .A1(n10627), .A2(n10626), .ZN(n10650) );
  INV_X1 U13680 ( .A(n10650), .ZN(n10630) );
  INV_X1 U13681 ( .A(n10628), .ZN(n10629) );
  NAND2_X2 U13682 ( .A1(n10630), .A2(n10644), .ZN(n10713) );
  INV_X1 U13683 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10631) );
  OAI22_X1 U13684 ( .A1(n13745), .A2(n14181), .B1(n10713), .B2(n10631), .ZN(
        n10632) );
  NOR2_X1 U13685 ( .A1(n10633), .A2(n10632), .ZN(n10663) );
  INV_X1 U13686 ( .A(n10712), .ZN(n19481) );
  INV_X1 U13687 ( .A(n10642), .ZN(n10634) );
  NOR2_X2 U13688 ( .A1(n10650), .A2(n10634), .ZN(n19351) );
  AOI22_X1 U13689 ( .A1(n19481), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n19351), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10639) );
  AND2_X2 U13690 ( .A1(n10635), .A2(n10644), .ZN(n10717) );
  INV_X1 U13691 ( .A(n10636), .ZN(n10637) );
  AOI22_X1 U13692 ( .A1(n10717), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13617), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10638) );
  AND2_X1 U13693 ( .A1(n10639), .A2(n10638), .ZN(n10662) );
  INV_X1 U13694 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14189) );
  INV_X1 U13695 ( .A(n10640), .ZN(n10656) );
  INV_X1 U13696 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14191) );
  OAI22_X1 U13697 ( .A1(n14189), .A2(n19731), .B1(n10701), .B2(n14191), .ZN(
        n10643) );
  AOI21_X1 U13698 ( .B1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n19659), .A(
        n10643), .ZN(n10661) );
  INV_X1 U13700 ( .A(n19770), .ZN(n10646) );
  NAND2_X1 U13701 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10653) );
  INV_X1 U13702 ( .A(n19686), .ZN(n10647) );
  NAND2_X1 U13703 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10652) );
  INV_X1 U13704 ( .A(n10648), .ZN(n10649) );
  NAND2_X1 U13705 ( .A1(n10718), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10651) );
  NAND3_X1 U13706 ( .A1(n10653), .A2(n10652), .A3(n10651), .ZN(n10659) );
  INV_X1 U13707 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13582) );
  INV_X1 U13708 ( .A(n13037), .ZN(n10654) );
  OAI211_X1 U13709 ( .C1(n13582), .C2(n10700), .A(n10657), .B(n14316), .ZN(
        n10658) );
  NOR2_X1 U13710 ( .A1(n10659), .A2(n10658), .ZN(n10660) );
  AOI22_X1 U13711 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10684), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13712 ( .A1(n14130), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13713 ( .A1(n10573), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n14151), .ZN(n10665) );
  AOI22_X1 U13714 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10664) );
  NAND4_X1 U13715 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10675) );
  AOI22_X1 U13716 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14142), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13717 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13718 ( .A1(n10679), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13719 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10670) );
  NAND4_X1 U13720 ( .A1(n10673), .A2(n10672), .A3(n10671), .A4(n10670), .ZN(
        n10674) );
  NOR2_X1 U13721 ( .A1(n10675), .A2(n10674), .ZN(n10963) );
  OR2_X1 U13722 ( .A1(n10963), .A2(n14316), .ZN(n10693) );
  AOI22_X1 U13723 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13724 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13725 ( .A1(n10573), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13726 ( .A1(n10679), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10680) );
  NAND4_X1 U13727 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(
        n10692) );
  AOI22_X1 U13728 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14142), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13729 ( .A1(n14130), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13730 ( .A1(n10684), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13731 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10685), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10687) );
  NAND4_X1 U13732 ( .A1(n10690), .A2(n10689), .A3(n10688), .A4(n10687), .ZN(
        n10691) );
  NOR2_X1 U13733 ( .A1(n10692), .A2(n10691), .ZN(n12863) );
  NOR2_X1 U13734 ( .A1(n10693), .A2(n12863), .ZN(n10967) );
  OR2_X1 U13735 ( .A1(n10967), .A2(n11383), .ZN(n10694) );
  AOI22_X1 U13736 ( .A1(n10717), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n10718), .ZN(n10696) );
  AOI22_X1 U13737 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13617), .B1(
        n19351), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10695) );
  AND2_X1 U13738 ( .A1(n10696), .A2(n10695), .ZN(n10709) );
  INV_X1 U13739 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14241) );
  INV_X1 U13740 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14239) );
  OAI22_X1 U13741 ( .A1(n14241), .A2(n19456), .B1(n13745), .B2(n14239), .ZN(
        n10699) );
  INV_X1 U13742 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14238) );
  INV_X1 U13743 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10697) );
  OAI22_X1 U13744 ( .A1(n10712), .A2(n14238), .B1(n10713), .B2(n10697), .ZN(
        n10698) );
  NOR2_X1 U13745 ( .A1(n10699), .A2(n10698), .ZN(n10708) );
  INV_X1 U13746 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14249) );
  INV_X1 U13747 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14250) );
  INV_X1 U13748 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10702) );
  INV_X1 U13749 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14247) );
  OAI22_X1 U13750 ( .A1(n10702), .A2(n10726), .B1(n19731), .B2(n14247), .ZN(
        n10703) );
  NOR2_X1 U13751 ( .A1(n10704), .A2(n10703), .ZN(n10707) );
  AOI22_X1 U13752 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10705), .B1(
        n19659), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10706) );
  NAND4_X1 U13753 ( .A1(n10709), .A2(n10708), .A3(n10707), .A4(n10706), .ZN(
        n10710) );
  NAND2_X1 U13754 ( .A1(n11392), .A2(n14294), .ZN(n10711) );
  INV_X1 U13755 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14298) );
  INV_X1 U13756 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14296) );
  OAI22_X1 U13757 ( .A1(n14298), .A2(n19456), .B1(n13745), .B2(n14296), .ZN(
        n10716) );
  INV_X1 U13758 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14295) );
  INV_X1 U13759 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10714) );
  OAI22_X1 U13760 ( .A1(n10712), .A2(n14295), .B1(n10713), .B2(n10714), .ZN(
        n10715) );
  NOR2_X1 U13761 ( .A1(n10716), .A2(n10715), .ZN(n10733) );
  AOI22_X1 U13762 ( .A1(n10717), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13519), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13763 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n13617), .B1(
        n19351), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10719) );
  AND2_X1 U13764 ( .A1(n10720), .A2(n10719), .ZN(n10732) );
  AOI22_X1 U13765 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19546), .B1(
        n19659), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10731) );
  INV_X1 U13766 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10723) );
  INV_X1 U13767 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10722) );
  OAI22_X1 U13768 ( .A1(n10723), .A2(n10700), .B1(n19770), .B2(n10722), .ZN(
        n10725) );
  INV_X1 U13769 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14307) );
  INV_X1 U13770 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14306) );
  OAI22_X1 U13771 ( .A1(n14307), .A2(n19686), .B1(n10701), .B2(n14306), .ZN(
        n10724) );
  OR2_X1 U13772 ( .A1(n10725), .A2(n10724), .ZN(n10729) );
  INV_X1 U13773 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10727) );
  INV_X1 U13774 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14304) );
  OAI22_X1 U13775 ( .A1(n10727), .A2(n10726), .B1(n19731), .B2(n14304), .ZN(
        n10728) );
  NOR2_X1 U13776 ( .A1(n10729), .A2(n10728), .ZN(n10730) );
  NAND4_X1 U13777 ( .A1(n10733), .A2(n10732), .A3(n10731), .A4(n10730), .ZN(
        n10746) );
  AOI22_X1 U13778 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13779 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13780 ( .A1(n10684), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13781 ( .A1(n14142), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10734) );
  NAND4_X1 U13782 ( .A1(n10737), .A2(n10736), .A3(n10735), .A4(n10734), .ZN(
        n10744) );
  AOI22_X1 U13783 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13784 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13785 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13786 ( .A1(n10573), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10739) );
  NAND4_X1 U13787 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n10743) );
  NAND2_X1 U13788 ( .A1(n11403), .A2(n14294), .ZN(n10745) );
  NAND2_X1 U13789 ( .A1(n14130), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10750) );
  NAND2_X1 U13790 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10749) );
  NAND2_X1 U13791 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10748) );
  NAND2_X1 U13792 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10747) );
  NAND2_X1 U13793 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10754) );
  NAND2_X1 U13794 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10753) );
  INV_X1 U13795 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19348) );
  NAND2_X1 U13796 ( .A1(n14151), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10752) );
  NAND2_X1 U13797 ( .A1(n10573), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10751) );
  NAND2_X1 U13798 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10758) );
  NAND2_X1 U13799 ( .A1(n14143), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10757) );
  NAND2_X1 U13800 ( .A1(n10684), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10756) );
  NAND2_X1 U13801 ( .A1(n14142), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10755) );
  NAND2_X1 U13802 ( .A1(n10677), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10763) );
  NAND2_X1 U13803 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10762) );
  NAND2_X1 U13804 ( .A1(n10669), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10761) );
  NAND2_X1 U13805 ( .A1(n10565), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10760) );
  NAND4_X2 U13806 ( .A1(n10767), .A2(n10766), .A3(n10765), .A4(n10764), .ZN(
        n10931) );
  NAND2_X1 U13807 ( .A1(n10978), .A2(n10959), .ZN(n10777) );
  INV_X1 U13808 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10769) );
  MUX2_X1 U13809 ( .A(n10770), .B(n10769), .S(n14024), .Z(n10800) );
  AND2_X1 U13810 ( .A1(n10942), .A2(n15119), .ZN(n10789) );
  INV_X1 U13811 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13706) );
  NAND2_X1 U13812 ( .A1(n10789), .A2(n13706), .ZN(n10772) );
  NAND2_X1 U13813 ( .A1(n11380), .A2(n10772), .ZN(n10793) );
  NAND2_X1 U13814 ( .A1(n10787), .A2(n10793), .ZN(n10786) );
  INV_X1 U13815 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13543) );
  MUX2_X1 U13816 ( .A(n10773), .B(n13543), .S(n14024), .Z(n10774) );
  NAND2_X1 U13817 ( .A1(n10800), .A2(n10782), .ZN(n10799) );
  MUX2_X1 U13818 ( .A(n11403), .B(P2_EBX_REG_5__SCAN_IN), .S(n14024), .Z(
        n10775) );
  AND2_X1 U13819 ( .A1(n10799), .A2(n10775), .ZN(n10776) );
  OR2_X1 U13820 ( .A1(n10776), .A2(n10840), .ZN(n19141) );
  XNOR2_X1 U13821 ( .A(n10802), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13583) );
  INV_X1 U13822 ( .A(n10778), .ZN(n10781) );
  INV_X1 U13823 ( .A(n10779), .ZN(n10780) );
  INV_X1 U13824 ( .A(n10782), .ZN(n10785) );
  NAND2_X1 U13825 ( .A1(n10786), .A2(n10783), .ZN(n10784) );
  NAND2_X1 U13826 ( .A1(n10785), .A2(n10784), .ZN(n13537) );
  OAI21_X2 U13827 ( .B1(n13439), .B2(n10931), .A(n13537), .ZN(n13442) );
  OAI21_X1 U13828 ( .B1(n10787), .B2(n10793), .A(n10786), .ZN(n13552) );
  INV_X1 U13829 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19297) );
  MUX2_X1 U13830 ( .A(n11314), .B(n12863), .S(n10376), .Z(n10788) );
  NAND2_X1 U13831 ( .A1(n10788), .A2(n13515), .ZN(n10791) );
  INV_X1 U13832 ( .A(n10789), .ZN(n10790) );
  NAND2_X1 U13833 ( .A1(n10791), .A2(n10790), .ZN(n15118) );
  INV_X1 U13834 ( .A(n15118), .ZN(n10792) );
  NAND2_X1 U13835 ( .A1(n10792), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12936) );
  INV_X1 U13836 ( .A(n10793), .ZN(n10795) );
  NAND3_X1 U13837 ( .A1(n10942), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10794) );
  NAND2_X1 U13838 ( .A1(n10795), .A2(n10794), .ZN(n13710) );
  NOR2_X1 U13839 ( .A1(n12936), .A2(n13710), .ZN(n10796) );
  NAND2_X1 U13840 ( .A1(n12936), .A2(n13710), .ZN(n12935) );
  OAI21_X1 U13841 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10796), .A(
        n12935), .ZN(n12946) );
  XNOR2_X1 U13842 ( .A(n13552), .B(n19297), .ZN(n12945) );
  OR2_X1 U13843 ( .A1(n12946), .A2(n12945), .ZN(n12943) );
  OAI21_X1 U13844 ( .B1(n13552), .B2(n19297), .A(n12943), .ZN(n13440) );
  OAI21_X1 U13845 ( .B1(n13442), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13440), .ZN(n10798) );
  NAND2_X1 U13846 ( .A1(n13442), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10797) );
  NAND2_X1 U13847 ( .A1(n10798), .A2(n10797), .ZN(n13480) );
  OAI21_X1 U13848 ( .B1(n10782), .B2(n10800), .A(n10799), .ZN(n13661) );
  XNOR2_X1 U13849 ( .A(n13661), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13478) );
  NOR2_X1 U13850 ( .A1(n13661), .A2(n13482), .ZN(n10801) );
  NAND2_X1 U13851 ( .A1(n10802), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10803) );
  OAI21_X1 U13852 ( .B1(n13583), .B2(n13584), .A(n10803), .ZN(n15669) );
  NAND2_X1 U13853 ( .A1(n10836), .A2(n10834), .ZN(n10832) );
  INV_X1 U13854 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14321) );
  INV_X1 U13855 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14319) );
  OAI22_X1 U13856 ( .A1(n14321), .A2(n19456), .B1(n13745), .B2(n14319), .ZN(
        n10807) );
  INV_X1 U13857 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14318) );
  INV_X1 U13858 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10805) );
  OAI22_X1 U13859 ( .A1(n10712), .A2(n14318), .B1(n10713), .B2(n10805), .ZN(
        n10806) );
  NOR2_X1 U13860 ( .A1(n10807), .A2(n10806), .ZN(n10819) );
  AOI22_X1 U13861 ( .A1(n10717), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13617), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13862 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13519), .B1(
        n19351), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10808) );
  AND2_X1 U13863 ( .A1(n10809), .A2(n10808), .ZN(n10818) );
  AOI22_X1 U13864 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19546), .B1(
        n19659), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10817) );
  INV_X1 U13865 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10810) );
  INV_X1 U13866 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14333) );
  OAI22_X1 U13867 ( .A1(n10810), .A2(n19770), .B1(n19686), .B2(n14333), .ZN(
        n10812) );
  INV_X1 U13868 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13577) );
  INV_X1 U13869 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14327) );
  OAI22_X1 U13870 ( .A1(n13577), .A2(n10700), .B1(n10701), .B2(n14327), .ZN(
        n10811) );
  OR2_X1 U13871 ( .A1(n10812), .A2(n10811), .ZN(n10815) );
  INV_X1 U13872 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10813) );
  INV_X1 U13873 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14331) );
  OAI22_X1 U13874 ( .A1(n10813), .A2(n10726), .B1(n19731), .B2(n14331), .ZN(
        n10814) );
  NOR2_X1 U13875 ( .A1(n10815), .A2(n10814), .ZN(n10816) );
  NAND4_X1 U13876 ( .A1(n10819), .A2(n10818), .A3(n10817), .A4(n10816), .ZN(
        n10831) );
  AOI22_X1 U13877 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13878 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13879 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13880 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14142), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10820) );
  NAND4_X1 U13881 ( .A1(n10823), .A2(n10822), .A3(n10821), .A4(n10820), .ZN(
        n10829) );
  AOI22_X1 U13882 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n14151), .ZN(n10827) );
  AOI22_X1 U13883 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13884 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13885 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10824) );
  NAND4_X1 U13886 ( .A1(n10827), .A2(n10826), .A3(n10825), .A4(n10824), .ZN(
        n10828) );
  INV_X1 U13887 ( .A(n10839), .ZN(n11404) );
  NAND2_X1 U13888 ( .A1(n11404), .A2(n14294), .ZN(n10830) );
  NAND2_X1 U13889 ( .A1(n10831), .A2(n10830), .ZN(n10981) );
  NAND2_X1 U13890 ( .A1(n10832), .A2(n10981), .ZN(n10837) );
  INV_X1 U13891 ( .A(n10981), .ZN(n10833) );
  NAND2_X1 U13892 ( .A1(n10836), .A2(n10835), .ZN(n10988) );
  NAND2_X1 U13893 ( .A1(n10979), .A2(n10959), .ZN(n10843) );
  INV_X1 U13894 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10838) );
  MUX2_X1 U13895 ( .A(n10839), .B(n10838), .S(n14024), .Z(n10841) );
  NOR2_X1 U13896 ( .A1(n10840), .A2(n10841), .ZN(n10842) );
  OR2_X1 U13897 ( .A1(n10853), .A2(n10842), .ZN(n13630) );
  NAND2_X1 U13898 ( .A1(n15669), .A2(n15668), .ZN(n10846) );
  NAND2_X1 U13899 ( .A1(n10844), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10845) );
  MUX2_X1 U13900 ( .A(n10931), .B(n10847), .S(n14024), .Z(n10851) );
  AND2_X2 U13901 ( .A1(n10853), .A2(n10851), .ZN(n10859) );
  NAND2_X1 U13902 ( .A1(n14024), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10848) );
  OR2_X1 U13903 ( .A1(n10859), .A2(n10848), .ZN(n10849) );
  AND2_X1 U13904 ( .A1(n10849), .A2(n10858), .ZN(n13642) );
  AND2_X1 U13905 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10850) );
  NAND2_X1 U13906 ( .A1(n13642), .A2(n10850), .ZN(n16302) );
  INV_X1 U13907 ( .A(n10851), .ZN(n10852) );
  XNOR2_X1 U13908 ( .A(n10853), .B(n10852), .ZN(n19130) );
  NAND2_X1 U13909 ( .A1(n19130), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16300) );
  INV_X1 U13910 ( .A(n13642), .ZN(n10854) );
  INV_X1 U13911 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16333) );
  OAI21_X1 U13912 ( .B1(n10854), .B2(n10959), .A(n16333), .ZN(n16303) );
  INV_X1 U13913 ( .A(n19130), .ZN(n10855) );
  INV_X1 U13914 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15664) );
  NAND2_X1 U13915 ( .A1(n10855), .A2(n15664), .ZN(n15436) );
  AND2_X1 U13916 ( .A1(n16303), .A2(n15436), .ZN(n10856) );
  NAND2_X1 U13917 ( .A1(n14024), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10857) );
  XNOR2_X1 U13918 ( .A(n10858), .B(n10857), .ZN(n19117) );
  NAND2_X1 U13919 ( .A1(n19117), .A2(n10931), .ZN(n10866) );
  INV_X1 U13920 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21028) );
  AND2_X1 U13921 ( .A1(n10866), .A2(n21028), .ZN(n15646) );
  NAND3_X1 U13922 ( .A1(n10861), .A2(P2_EBX_REG_10__SCAN_IN), .A3(n10942), 
        .ZN(n10860) );
  OAI211_X1 U13923 ( .C1(n10861), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10860), .B(
        n10941), .ZN(n19103) );
  OAI21_X1 U13924 ( .B1(n19103), .B2(n10959), .A(n16278), .ZN(n16282) );
  INV_X1 U13925 ( .A(n10869), .ZN(n10863) );
  NAND3_X1 U13926 ( .A1(n10942), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n9863), .ZN(
        n10862) );
  AND2_X1 U13927 ( .A1(n10863), .A2(n10862), .ZN(n19086) );
  AOI21_X1 U13928 ( .B1(n19086), .B2(n10931), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15631) );
  INV_X1 U13929 ( .A(n19103), .ZN(n10865) );
  AND2_X1 U13930 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10864) );
  NAND2_X1 U13931 ( .A1(n10865), .A2(n10864), .ZN(n16281) );
  OR2_X1 U13932 ( .A1(n10866), .A2(n21028), .ZN(n15645) );
  AND2_X1 U13933 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10867) );
  NAND2_X1 U13934 ( .A1(n19086), .A2(n10867), .ZN(n15629) );
  AND3_X1 U13935 ( .A1(n16281), .A2(n15645), .A3(n15629), .ZN(n10868) );
  NAND2_X1 U13936 ( .A1(n14024), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10870) );
  NAND2_X1 U13937 ( .A1(n10869), .A2(n10870), .ZN(n10893) );
  INV_X1 U13938 ( .A(n10870), .ZN(n10872) );
  NAND2_X1 U13939 ( .A1(n10872), .A2(n10871), .ZN(n10873) );
  NAND2_X1 U13940 ( .A1(n10893), .A2(n10873), .ZN(n19078) );
  INV_X1 U13941 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10874) );
  NOR2_X1 U13942 ( .A1(n10875), .A2(n10874), .ZN(n15611) );
  NAND2_X1 U13943 ( .A1(n10875), .A2(n10874), .ZN(n15612) );
  AND2_X1 U13944 ( .A1(n10942), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10892) );
  AND2_X1 U13945 ( .A1(n10942), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10897) );
  NAND2_X1 U13946 ( .A1(n14024), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10890) );
  INV_X1 U13947 ( .A(n10883), .ZN(n10877) );
  NAND2_X1 U13948 ( .A1(n14024), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10887) );
  INV_X1 U13949 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10878) );
  NAND2_X1 U13950 ( .A1(n10879), .A2(n10878), .ZN(n10880) );
  INV_X1 U13951 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15180) );
  NAND2_X1 U13952 ( .A1(n10928), .A2(n10941), .ZN(n10925) );
  OR2_X1 U13953 ( .A1(n10925), .A2(n10881), .ZN(n18992) );
  NAND2_X1 U13954 ( .A1(n10882), .A2(n11612), .ZN(n11600) );
  NAND3_X1 U13955 ( .A1(n10883), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n14024), 
        .ZN(n10884) );
  NAND3_X1 U13956 ( .A1(n10885), .A2(n10941), .A3(n10884), .ZN(n15110) );
  OR2_X1 U13957 ( .A1(n15110), .A2(n10959), .ZN(n10886) );
  XNOR2_X1 U13958 ( .A(n10886), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11590) );
  OR2_X1 U13959 ( .A1(n10888), .A2(n10887), .ZN(n10889) );
  NAND2_X1 U13960 ( .A1(n10905), .A2(n10889), .ZN(n19031) );
  OAI21_X1 U13961 ( .B1(n19031), .B2(n10959), .A(n10125), .ZN(n11595) );
  XNOR2_X1 U13962 ( .A(n9851), .B(n10890), .ZN(n19043) );
  NAND2_X1 U13963 ( .A1(n19043), .A2(n10931), .ZN(n10891) );
  INV_X1 U13964 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15578) );
  NAND2_X1 U13965 ( .A1(n10891), .A2(n15578), .ZN(n15403) );
  NAND2_X1 U13966 ( .A1(n10893), .A2(n10892), .ZN(n10894) );
  NAND2_X1 U13967 ( .A1(n10899), .A2(n10894), .ZN(n19066) );
  OR2_X1 U13968 ( .A1(n19066), .A2(n10959), .ZN(n10896) );
  NAND2_X1 U13969 ( .A1(n10896), .A2(n10895), .ZN(n15425) );
  INV_X1 U13970 ( .A(n10897), .ZN(n10898) );
  XNOR2_X1 U13971 ( .A(n10899), .B(n10898), .ZN(n19054) );
  NAND2_X1 U13972 ( .A1(n19054), .A2(n10931), .ZN(n10900) );
  NAND2_X1 U13973 ( .A1(n10900), .A2(n15588), .ZN(n15414) );
  AND4_X1 U13974 ( .A1(n11595), .A2(n15403), .A3(n15425), .A4(n15414), .ZN(
        n10903) );
  NAND2_X1 U13975 ( .A1(n14024), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10901) );
  XNOR2_X1 U13976 ( .A(n10909), .B(n10901), .ZN(n19002) );
  NAND2_X1 U13977 ( .A1(n19002), .A2(n10931), .ZN(n10902) );
  INV_X1 U13978 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15527) );
  NAND2_X1 U13979 ( .A1(n10902), .A2(n15527), .ZN(n15349) );
  NAND2_X1 U13980 ( .A1(n10905), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10904) );
  MUX2_X1 U13981 ( .A(n10905), .B(n10904), .S(n14024), .Z(n10906) );
  OR2_X1 U13982 ( .A1(n10905), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10908) );
  NAND2_X1 U13983 ( .A1(n15095), .A2(n10931), .ZN(n10907) );
  NAND2_X1 U13984 ( .A1(n10907), .A2(n15377), .ZN(n15369) );
  NAND3_X1 U13985 ( .A1(n10908), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n10942), 
        .ZN(n10910) );
  AND2_X1 U13986 ( .A1(n10910), .A2(n10909), .ZN(n19014) );
  NAND2_X1 U13987 ( .A1(n19014), .A2(n10931), .ZN(n10912) );
  INV_X1 U13988 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15534) );
  NAND2_X1 U13989 ( .A1(n10912), .A2(n15534), .ZN(n15358) );
  NAND2_X1 U13990 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10911) );
  OR2_X1 U13991 ( .A1(n18992), .A2(n10911), .ZN(n11599) );
  NAND2_X1 U13992 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10913) );
  OR2_X1 U13993 ( .A1(n15110), .A2(n10913), .ZN(n11591) );
  AND2_X1 U13994 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10914) );
  NAND2_X1 U13995 ( .A1(n19043), .A2(n10914), .ZN(n15402) );
  NAND2_X1 U13996 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10915) );
  OR2_X1 U13997 ( .A1(n19066), .A2(n10915), .ZN(n15424) );
  AND2_X1 U13998 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10916) );
  NAND2_X1 U13999 ( .A1(n19054), .A2(n10916), .ZN(n15413) );
  AND4_X1 U14000 ( .A1(n11591), .A2(n15402), .A3(n15424), .A4(n15413), .ZN(
        n10919) );
  INV_X1 U14001 ( .A(n19031), .ZN(n10918) );
  AND2_X1 U14002 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10917) );
  NAND2_X1 U14003 ( .A1(n10918), .A2(n10917), .ZN(n11592) );
  AND3_X1 U14004 ( .A1(n15359), .A2(n10919), .A3(n11592), .ZN(n10922) );
  AND2_X1 U14005 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10920) );
  NAND2_X1 U14006 ( .A1(n19002), .A2(n10920), .ZN(n15348) );
  AND2_X1 U14007 ( .A1(n10931), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10921) );
  NAND2_X1 U14008 ( .A1(n15095), .A2(n10921), .ZN(n15367) );
  AND4_X1 U14009 ( .A1(n11599), .A2(n10922), .A3(n15348), .A4(n15367), .ZN(
        n10923) );
  NAND2_X1 U14010 ( .A1(n14024), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10926) );
  NAND2_X1 U14011 ( .A1(n10925), .A2(n10926), .ZN(n10934) );
  INV_X1 U14012 ( .A(n10926), .ZN(n10927) );
  NAND2_X1 U14013 ( .A1(n10928), .A2(n10927), .ZN(n10929) );
  NAND2_X1 U14014 ( .A1(n10934), .A2(n10929), .ZN(n15824) );
  OR2_X1 U14015 ( .A1(n15824), .A2(n10959), .ZN(n10930) );
  INV_X1 U14016 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10999) );
  NAND2_X1 U14017 ( .A1(n10930), .A2(n10999), .ZN(n15499) );
  NAND2_X1 U14018 ( .A1(n15497), .A2(n15499), .ZN(n10932) );
  NAND2_X1 U14019 ( .A1(n10932), .A2(n15498), .ZN(n15483) );
  AND2_X1 U14020 ( .A1(n10942), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10933) );
  OR2_X2 U14021 ( .A1(n10934), .A2(n10933), .ZN(n15076) );
  NAND2_X1 U14022 ( .A1(n10934), .A2(n10933), .ZN(n10935) );
  NAND2_X1 U14023 ( .A1(n15076), .A2(n10935), .ZN(n16227) );
  NAND2_X1 U14024 ( .A1(n15483), .A2(n15484), .ZN(n10938) );
  INV_X1 U14025 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20965) );
  NAND2_X1 U14026 ( .A1(n10941), .A2(n10931), .ZN(n15329) );
  NOR2_X1 U14027 ( .A1(n15329), .A2(n15474), .ZN(n10940) );
  NAND2_X1 U14028 ( .A1(n15329), .A2(n15474), .ZN(n10939) );
  AND2_X1 U14029 ( .A1(n15329), .A2(n15325), .ZN(n15317) );
  NOR2_X2 U14030 ( .A1(n15076), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16220) );
  INV_X1 U14031 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16219) );
  NAND2_X1 U14032 ( .A1(n16220), .A2(n16219), .ZN(n16218) );
  OR2_X2 U14033 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n16218), .ZN(n10945) );
  AND3_X1 U14034 ( .A1(n10942), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n16218), .ZN(
        n10943) );
  NOR2_X1 U14035 ( .A1(n14022), .A2(n10943), .ZN(n16199) );
  NAND2_X1 U14036 ( .A1(n16199), .A2(n10931), .ZN(n10951) );
  XNOR2_X1 U14037 ( .A(n10951), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15308) );
  INV_X1 U14038 ( .A(n13964), .ZN(n10949) );
  NAND2_X1 U14039 ( .A1(n14024), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10944) );
  INV_X1 U14040 ( .A(n10944), .ZN(n10946) );
  NAND2_X1 U14041 ( .A1(n10946), .A2(n10945), .ZN(n10947) );
  NAND2_X1 U14042 ( .A1(n10958), .A2(n10947), .ZN(n16187) );
  INV_X1 U14043 ( .A(n13962), .ZN(n10948) );
  NAND2_X1 U14044 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11002) );
  NOR2_X1 U14045 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13973) );
  NAND2_X1 U14046 ( .A1(n14024), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10950) );
  XNOR2_X1 U14047 ( .A(n10958), .B(n10950), .ZN(n15065) );
  NAND2_X1 U14048 ( .A1(n15065), .A2(n10931), .ZN(n13966) );
  INV_X1 U14049 ( .A(n10951), .ZN(n10953) );
  INV_X1 U14050 ( .A(n15329), .ZN(n10952) );
  OAI21_X1 U14051 ( .B1(n13973), .B2(n13966), .A(n13963), .ZN(n10954) );
  INV_X1 U14052 ( .A(n10954), .ZN(n10955) );
  AND2_X1 U14053 ( .A1(n14024), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10957) );
  NAND2_X1 U14054 ( .A1(n14024), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13922) );
  XNOR2_X1 U14055 ( .A(n13923), .B(n13922), .ZN(n10960) );
  INV_X1 U14056 ( .A(n10960), .ZN(n16176) );
  NAND3_X1 U14057 ( .A1(n16176), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10931), .ZN(n14017) );
  OAI21_X1 U14058 ( .B1(n10960), .B2(n10959), .A(n11000), .ZN(n13920) );
  NAND2_X1 U14059 ( .A1(n14017), .A2(n13920), .ZN(n10961) );
  XNOR2_X1 U14060 ( .A(n13921), .B(n10961), .ZN(n11583) );
  NAND2_X1 U14061 ( .A1(n11583), .A2(n19276), .ZN(n11004) );
  OR2_X1 U14062 ( .A1(n12863), .A2(n14316), .ZN(n10962) );
  NAND2_X1 U14063 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12862) );
  INV_X1 U14064 ( .A(n12862), .ZN(n10964) );
  XOR2_X1 U14065 ( .A(n12863), .B(n10963), .Z(n10965) );
  NAND2_X1 U14066 ( .A1(n10964), .A2(n10965), .ZN(n10966) );
  XOR2_X1 U14067 ( .A(n10965), .B(n10964), .Z(n12939) );
  NAND2_X1 U14068 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12939), .ZN(
        n12938) );
  NAND2_X1 U14069 ( .A1(n10966), .A2(n12938), .ZN(n10968) );
  XNOR2_X1 U14070 ( .A(n19297), .B(n10968), .ZN(n12949) );
  XNOR2_X1 U14071 ( .A(n11383), .B(n10967), .ZN(n12948) );
  NAND2_X1 U14072 ( .A1(n12949), .A2(n12948), .ZN(n12947) );
  NAND2_X1 U14073 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10968), .ZN(
        n10969) );
  NAND2_X1 U14074 ( .A1(n12947), .A2(n10969), .ZN(n10970) );
  XNOR2_X1 U14075 ( .A(n10970), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13438) );
  NAND2_X1 U14076 ( .A1(n10970), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10971) );
  NAND2_X1 U14077 ( .A1(n13475), .A2(n13482), .ZN(n10977) );
  INV_X1 U14078 ( .A(n10973), .ZN(n10976) );
  INV_X1 U14079 ( .A(n10974), .ZN(n10975) );
  NAND2_X1 U14080 ( .A1(n10976), .A2(n10975), .ZN(n13476) );
  NAND2_X1 U14081 ( .A1(n10977), .A2(n13476), .ZN(n13597) );
  NAND2_X1 U14082 ( .A1(n10979), .A2(n13595), .ZN(n10984) );
  NAND2_X1 U14083 ( .A1(n13596), .A2(n10980), .ZN(n10983) );
  INV_X1 U14084 ( .A(n13595), .ZN(n13599) );
  NAND2_X1 U14085 ( .A1(n13599), .A2(n10981), .ZN(n10982) );
  OAI211_X1 U14086 ( .C1(n13596), .C2(n10984), .A(n10983), .B(n10982), .ZN(
        n15672) );
  NAND2_X1 U14087 ( .A1(n15672), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15671) );
  INV_X1 U14088 ( .A(n13596), .ZN(n10985) );
  NAND2_X1 U14089 ( .A1(n10985), .A2(n13595), .ZN(n10986) );
  NAND2_X1 U14090 ( .A1(n10986), .A2(n10979), .ZN(n10987) );
  NAND2_X2 U14091 ( .A1(n15671), .A2(n10987), .ZN(n10992) );
  NAND2_X1 U14092 ( .A1(n10990), .A2(n10959), .ZN(n10991) );
  AND2_X1 U14093 ( .A1(n10994), .A2(n10991), .ZN(n15439) );
  NAND2_X1 U14094 ( .A1(n10992), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10993) );
  INV_X1 U14095 ( .A(n10994), .ZN(n10995) );
  NAND2_X1 U14096 ( .A1(n10995), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10996) );
  AND2_X1 U14097 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15635) );
  AND2_X1 U14098 ( .A1(n15635), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15522) );
  NAND3_X1 U14099 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15525) );
  NOR2_X1 U14100 ( .A1(n15525), .A2(n15377), .ZN(n10997) );
  NAND2_X1 U14101 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15590) );
  NOR2_X1 U14102 ( .A1(n15590), .A2(n15588), .ZN(n15523) );
  AND3_X1 U14103 ( .A1(n15522), .A2(n10997), .A3(n15523), .ZN(n15526) );
  AND3_X1 U14104 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10998) );
  NAND2_X1 U14105 ( .A1(n15526), .A2(n10998), .ZN(n11575) );
  INV_X1 U14106 ( .A(n11575), .ZN(n11608) );
  OR3_X4 U14107 ( .A1(n15511), .A2(n20965), .A3(n10999), .ZN(n15493) );
  INV_X1 U14108 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15311) );
  INV_X1 U14109 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11001) );
  OAI21_X1 U14110 ( .B1(n9840), .B2(n11001), .A(n11000), .ZN(n11003) );
  INV_X1 U14111 ( .A(n11002), .ZN(n13971) );
  AND2_X1 U14112 ( .A1(n13971), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14051) );
  NOR2_X1 U14113 ( .A1(n18967), .A2(n14316), .ZN(n16287) );
  INV_X1 U14114 ( .A(n16287), .ZN(n19282) );
  NAND3_X1 U14115 ( .A1(n11005), .A2(n11004), .A3(n9854), .ZN(P2_U2985) );
  INV_X1 U14116 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18900) );
  NAND3_X1 U14117 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15793) );
  INV_X2 U14118 ( .A(n11056), .ZN(n17216) );
  NAND2_X2 U14119 ( .A1(n18897), .A2(n11015), .ZN(n11037) );
  INV_X2 U14120 ( .A(n11037), .ZN(n11065) );
  AOI22_X1 U14121 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11065), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11024) );
  NAND4_X2 U14122 ( .A1(n18910), .A2(n21179), .A3(n18897), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17163) );
  INV_X1 U14123 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U14124 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U14125 ( .A1(n21179), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11013) );
  INV_X2 U14126 ( .A(n17072), .ZN(n11051) );
  AOI22_X1 U14127 ( .A1(n9801), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11007) );
  OAI211_X1 U14128 ( .C1(n17246), .C2(n17126), .A(n11008), .B(n11007), .ZN(
        n11022) );
  INV_X2 U14129 ( .A(n17186), .ZN(n17230) );
  AOI22_X1 U14130 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n9806), .ZN(n11020) );
  NOR2_X2 U14131 ( .A1(n11010), .A2(n11012), .ZN(n11011) );
  INV_X1 U14132 ( .A(n17177), .ZN(n17229) );
  AOI22_X1 U14133 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11019) );
  INV_X2 U14134 ( .A(n9842), .ZN(n17236) );
  AOI22_X1 U14135 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11018) );
  INV_X1 U14136 ( .A(n11015), .ZN(n11016) );
  NAND2_X1 U14137 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11017) );
  NAND4_X1 U14138 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11021) );
  AOI211_X1 U14139 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11022), .B(n11021), .ZN(n11023) );
  INV_X1 U14140 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15760) );
  AOI22_X1 U14141 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11011), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11025) );
  OAI21_X1 U14142 ( .B1(n17151), .B2(n15760), .A(n11025), .ZN(n11035) );
  INV_X1 U14143 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U14144 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11032) );
  INV_X1 U14145 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n21130) );
  OAI22_X1 U14146 ( .A1(n17163), .A2(n21130), .B1(n11038), .B2(n21086), .ZN(
        n11030) );
  AOI22_X1 U14147 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11028) );
  INV_X1 U14148 ( .A(n11076), .ZN(n17235) );
  INV_X2 U14149 ( .A(n9841), .ZN(n17192) );
  AOI22_X1 U14150 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14151 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11026) );
  NAND3_X1 U14152 ( .A1(n11028), .A2(n11027), .A3(n11026), .ZN(n11029) );
  AOI211_X1 U14153 ( .C1(n11065), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n11030), .B(n11029), .ZN(n11031) );
  OAI211_X1 U14154 ( .C1(n11054), .C2(n11033), .A(n11032), .B(n11031), .ZN(
        n11034) );
  INV_X1 U14155 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U14156 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11036) );
  OAI21_X1 U14157 ( .B1(n11076), .B2(n17268), .A(n11036), .ZN(n11047) );
  AOI22_X1 U14158 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11045) );
  INV_X1 U14159 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U14160 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11039) );
  OAI21_X1 U14161 ( .B1(n9811), .B2(n17178), .A(n11039), .ZN(n11043) );
  INV_X1 U14162 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U14163 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U14164 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11040) );
  OAI211_X1 U14165 ( .C1(n17163), .C2(n17070), .A(n11041), .B(n11040), .ZN(
        n11042) );
  AOI211_X1 U14166 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n11043), .B(n11042), .ZN(n11044) );
  OAI211_X1 U14167 ( .C1(n11037), .C2(n17071), .A(n11045), .B(n11044), .ZN(
        n11046) );
  AOI211_X2 U14168 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n11047), .B(n11046), .ZN(n11282) );
  INV_X1 U14169 ( .A(n11282), .ZN(n17426) );
  AOI22_X1 U14170 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11065), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11063) );
  INV_X1 U14171 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U14172 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U14173 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11048) );
  OAI211_X1 U14174 ( .C1(n17163), .C2(n11050), .A(n11049), .B(n11048), .ZN(
        n11062) );
  AOI22_X1 U14175 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14176 ( .A1(n9801), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11052) );
  AOI22_X1 U14177 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11059) );
  NAND2_X1 U14178 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11058) );
  NAND3_X1 U14179 ( .A1(n11059), .A2(n11058), .A3(n11057), .ZN(n11060) );
  AOI22_X1 U14180 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U14181 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14182 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11071) );
  OAI22_X1 U14183 ( .A1(n9811), .A2(n17194), .B1(n10227), .B2(n21093), .ZN(
        n11064) );
  AOI22_X1 U14184 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11011), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14185 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11067) );
  INV_X1 U14186 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14187 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11070) );
  NAND2_X1 U14188 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11069) );
  AOI22_X1 U14189 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11065), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14190 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11075) );
  AOI22_X1 U14191 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11074) );
  OAI211_X1 U14192 ( .C1(n17246), .C2(n13851), .A(n11075), .B(n11074), .ZN(
        n11082) );
  AOI22_X1 U14193 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U14194 ( .A1(n9799), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U14195 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U14196 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11077) );
  NAND4_X1 U14197 ( .A1(n11080), .A2(n11079), .A3(n11078), .A4(n11077), .ZN(
        n11081) );
  AOI211_X1 U14198 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n11082), .B(n11081), .ZN(n11083) );
  OAI211_X1 U14199 ( .C1(n10244), .C2(n18500), .A(n11084), .B(n11083), .ZN(
        n11280) );
  AOI22_X1 U14200 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11094) );
  INV_X1 U14201 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U14202 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14203 ( .A1(n9799), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11085) );
  OAI211_X1 U14204 ( .C1(n17163), .C2(n17150), .A(n11086), .B(n11085), .ZN(
        n11092) );
  AOI22_X1 U14205 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14206 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14207 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11088) );
  NAND2_X1 U14208 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11087) );
  NAND4_X1 U14209 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n11091) );
  AOI211_X1 U14210 ( .C1(n17216), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n11092), .B(n11091), .ZN(n11093) );
  XOR2_X1 U14211 ( .A(n18900), .B(n11132), .Z(n11143) );
  INV_X1 U14212 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17950) );
  NOR2_X1 U14213 ( .A1(n17820), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17686) );
  INV_X1 U14214 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17681) );
  NAND2_X1 U14215 ( .A1(n17686), .A2(n17681), .ZN(n11095) );
  NOR2_X1 U14216 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11095), .ZN(
        n17653) );
  INV_X1 U14217 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17655) );
  NAND2_X1 U14218 ( .A1(n17653), .A2(n17655), .ZN(n17631) );
  NOR3_X1 U14219 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17631), .ZN(n11130) );
  INV_X1 U14220 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18050) );
  NOR2_X1 U14221 ( .A1(n18050), .A2(n18040), .ZN(n18025) );
  NAND2_X1 U14222 ( .A1(n18025), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17632) );
  INV_X1 U14223 ( .A(n17632), .ZN(n17996) );
  AND2_X1 U14224 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18000) );
  NAND2_X1 U14225 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18000), .ZN(
        n17983) );
  INV_X1 U14226 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17990) );
  NOR2_X1 U14227 ( .A1(n17983), .A2(n17990), .ZN(n16482) );
  NAND2_X1 U14228 ( .A1(n17996), .A2(n16482), .ZN(n16427) );
  INV_X1 U14229 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17973) );
  NOR2_X1 U14230 ( .A1(n16427), .A2(n17973), .ZN(n17606) );
  INV_X1 U14231 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18216) );
  XOR2_X1 U14232 ( .A(n18216), .B(n11110), .Z(n17897) );
  INV_X1 U14233 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n21045) );
  OAI22_X1 U14234 ( .A1(n17186), .A2(n18463), .B1(n17072), .B2(n21045), .ZN(
        n11101) );
  AOI22_X1 U14235 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14236 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17235), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14237 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11097) );
  NAND3_X1 U14238 ( .A1(n11099), .A2(n11098), .A3(n11097), .ZN(n11100) );
  AOI211_X1 U14239 ( .C1(n17237), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n11101), .B(n11100), .ZN(n11109) );
  INV_X1 U14240 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18593) );
  AOI22_X1 U14241 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11102) );
  OAI21_X1 U14242 ( .B1(n9842), .B2(n18593), .A(n11102), .ZN(n11107) );
  AOI22_X1 U14243 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11105) );
  INV_X1 U14244 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18304) );
  NAND2_X1 U14245 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  INV_X1 U14246 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18913) );
  NOR2_X1 U14247 ( .A1(n11276), .A2(n18913), .ZN(n17915) );
  INV_X1 U14248 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20976) );
  NAND2_X1 U14249 ( .A1(n17905), .A2(n10238), .ZN(n17896) );
  NAND2_X1 U14250 ( .A1(n17897), .A2(n17896), .ZN(n17895) );
  OR2_X1 U14251 ( .A1(n18216), .A2(n11110), .ZN(n11111) );
  NAND2_X1 U14252 ( .A1(n17895), .A2(n11111), .ZN(n11112) );
  INV_X1 U14253 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18195) );
  XNOR2_X1 U14254 ( .A(n11112), .B(n18195), .ZN(n17884) );
  XOR2_X1 U14255 ( .A(n11284), .B(n17426), .Z(n17883) );
  NAND2_X1 U14256 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11112), .ZN(
        n11113) );
  XOR2_X1 U14257 ( .A(n11114), .B(n11280), .Z(n17870) );
  INV_X1 U14258 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18194) );
  XOR2_X1 U14259 ( .A(n11115), .B(n17417), .Z(n11117) );
  INV_X1 U14260 ( .A(n11117), .ZN(n11116) );
  NAND2_X1 U14261 ( .A1(n11118), .A2(n11117), .ZN(n11119) );
  XNOR2_X1 U14262 ( .A(n18181), .B(n11297), .ZN(n17845) );
  XOR2_X1 U14263 ( .A(n11120), .B(n17845), .Z(n17852) );
  AOI21_X1 U14264 ( .B1(n17410), .B2(n11121), .A(n17820), .ZN(n11124) );
  NAND2_X1 U14265 ( .A1(n11124), .A2(n11123), .ZN(n11125) );
  NOR2_X1 U14266 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17801) );
  INV_X1 U14267 ( .A(n17801), .ZN(n11126) );
  NOR2_X2 U14268 ( .A1(n17802), .A2(n11126), .ZN(n17774) );
  INV_X1 U14269 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18080) );
  INV_X1 U14270 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17756) );
  NAND2_X1 U14271 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18117) );
  NOR2_X1 U14272 ( .A1(n18117), .A2(n17787), .ZN(n18090) );
  INV_X1 U14273 ( .A(n18090), .ZN(n17762) );
  NOR2_X1 U14274 ( .A1(n21108), .A2(n17762), .ZN(n18100) );
  NAND2_X1 U14275 ( .A1(n18100), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18077) );
  NAND2_X1 U14276 ( .A1(n18055), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18031) );
  INV_X1 U14277 ( .A(n18031), .ZN(n16426) );
  NAND2_X1 U14278 ( .A1(n16426), .A2(n17819), .ZN(n11128) );
  NAND2_X1 U14279 ( .A1(n11129), .A2(n11128), .ZN(n17709) );
  OAI221_X1 U14280 ( .B1(n11130), .B2(n17606), .C1(n11130), .C2(n17709), .A(
        n17659), .ZN(n17608) );
  NOR2_X2 U14281 ( .A1(n17608), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17607) );
  NAND2_X1 U14282 ( .A1(n18025), .A2(n17709), .ZN(n17651) );
  NAND3_X1 U14283 ( .A1(n16482), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17688), .ZN(n17615) );
  OR2_X1 U14284 ( .A1(n17820), .A2(n17607), .ZN(n17596) );
  OAI221_X1 U14285 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n11132), 
        .C1(n17950), .C2(n17597), .A(n17596), .ZN(n17580) );
  NOR2_X1 U14286 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17580), .ZN(
        n17579) );
  NOR2_X1 U14287 ( .A1(n17597), .A2(n11132), .ZN(n11134) );
  NAND2_X1 U14288 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17922) );
  INV_X1 U14289 ( .A(n17922), .ZN(n11131) );
  NOR2_X1 U14290 ( .A1(n11132), .A2(n11131), .ZN(n11133) );
  INV_X1 U14291 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17551) );
  NOR2_X1 U14292 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15800), .ZN(
        n15872) );
  NOR2_X1 U14293 ( .A1(n17820), .A2(n15872), .ZN(n11141) );
  NAND2_X1 U14294 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16453) );
  INV_X1 U14295 ( .A(n16453), .ZN(n15821) );
  NAND2_X1 U14296 ( .A1(n15821), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16458) );
  NOR2_X2 U14297 ( .A1(n16470), .A2(n16458), .ZN(n15871) );
  OR2_X1 U14298 ( .A1(n15871), .A2(n11137), .ZN(n11138) );
  OAI22_X1 U14299 ( .A1(n11141), .A2(n11138), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18900), .ZN(n11142) );
  OAI21_X1 U14300 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n15871), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U14301 ( .A1(n11143), .A2(n11139), .ZN(n11140) );
  AOI22_X1 U14302 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11144) );
  OAI21_X1 U14303 ( .B1(n9842), .B2(n17212), .A(n11144), .ZN(n11154) );
  AOI22_X1 U14304 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11152) );
  AOI22_X1 U14305 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11146) );
  OAI21_X1 U14306 ( .B1(n11054), .B2(n21111), .A(n11146), .ZN(n11150) );
  AOI22_X1 U14307 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14308 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11147) );
  OAI211_X1 U14309 ( .C1(n17246), .C2(n20981), .A(n11148), .B(n11147), .ZN(
        n11149) );
  AOI211_X1 U14310 ( .C1(n17216), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n11150), .B(n11149), .ZN(n11151) );
  OAI211_X1 U14311 ( .C1(n11076), .C2(n17213), .A(n11152), .B(n11151), .ZN(
        n11153) );
  AOI211_X4 U14312 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n11154), .B(n11153), .ZN(n18272) );
  AOI22_X1 U14313 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18767), .B2(n18910), .ZN(
        n11258) );
  AOI22_X1 U14314 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18772), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n9798), .ZN(n11162) );
  NAND2_X1 U14315 ( .A1(n18765), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11259) );
  OR2_X1 U14316 ( .A1(n11258), .A2(n11259), .ZN(n11155) );
  OAI21_X1 U14317 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18910), .A(
        n11155), .ZN(n11163) );
  NAND2_X1 U14318 ( .A1(n11162), .A2(n11163), .ZN(n11156) );
  OAI22_X1 U14319 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18261), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11157), .ZN(n11159) );
  NOR2_X1 U14320 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18261), .ZN(
        n11158) );
  NAND2_X1 U14321 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11157), .ZN(
        n11160) );
  AOI22_X1 U14322 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11159), .B1(
        n11158), .B2(n11160), .ZN(n11164) );
  OAI211_X1 U14323 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18765), .A(
        n11164), .B(n11259), .ZN(n11263) );
  AOI21_X1 U14324 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11160), .A(
        n11159), .ZN(n11161) );
  XOR2_X1 U14325 ( .A(n11163), .B(n11162), .Z(n11257) );
  NAND2_X1 U14326 ( .A1(n11164), .A2(n11257), .ZN(n11261) );
  OAI211_X1 U14327 ( .C1(n11258), .C2(n11263), .A(n11260), .B(n11261), .ZN(
        n18730) );
  AOI22_X1 U14328 ( .A1(n9801), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11165) );
  OAI21_X1 U14329 ( .B1(n17151), .B2(n17264), .A(n11165), .ZN(n11174) );
  AOI22_X1 U14330 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11172) );
  OAI22_X1 U14331 ( .A1(n10227), .A2(n13851), .B1(n17246), .B2(n18500), .ZN(
        n11170) );
  AOI22_X1 U14332 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U14333 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14334 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11166) );
  NAND3_X1 U14335 ( .A1(n11168), .A2(n11167), .A3(n11166), .ZN(n11169) );
  AOI211_X1 U14336 ( .C1(n17237), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n11170), .B(n11169), .ZN(n11171) );
  OAI211_X1 U14337 ( .C1(n17186), .C2(n17170), .A(n11172), .B(n11171), .ZN(
        n11173) );
  AOI211_X4 U14338 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n11174), .B(n11173), .ZN(n18282) );
  AOI22_X1 U14339 ( .A1(n17105), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11175) );
  OAI21_X1 U14340 ( .B1(n17177), .B2(n17071), .A(n11175), .ZN(n11184) );
  AOI22_X1 U14341 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11182) );
  INV_X1 U14342 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U14343 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11176) );
  OAI21_X1 U14344 ( .B1(n10244), .B2(n17176), .A(n11176), .ZN(n11180) );
  INV_X1 U14345 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18497) );
  AOI22_X1 U14346 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11178) );
  AOI22_X1 U14347 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11177) );
  OAI211_X1 U14348 ( .C1(n17246), .C2(n18497), .A(n11178), .B(n11177), .ZN(
        n11179) );
  AOI211_X1 U14349 ( .C1(n17216), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n11180), .B(n11179), .ZN(n11181) );
  OAI211_X1 U14350 ( .C1(n11055), .C2(n17070), .A(n11182), .B(n11181), .ZN(
        n11183) );
  AOI211_X2 U14351 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n11184), .B(n11183), .ZN(n18278) );
  AOI22_X1 U14352 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n11051), .ZN(n11185) );
  OAI21_X1 U14353 ( .B1(n17151), .B2(n17252), .A(n11185), .ZN(n11193) );
  AOI22_X1 U14354 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13905), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11192) );
  INV_X1 U14355 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U14356 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17216), .B1(
        n11065), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11186) );
  OAI21_X1 U14357 ( .B1(n17177), .B2(n16988), .A(n11186), .ZN(n11190) );
  INV_X1 U14358 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U14359 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n9801), .ZN(n11188) );
  AOI22_X1 U14360 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n9799), .ZN(n11187) );
  OAI211_X1 U14361 ( .C1(n16981), .C2(n17163), .A(n11188), .B(n11187), .ZN(
        n11189) );
  AOI211_X1 U14362 ( .C1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .C2(n17215), .A(
        n11190), .B(n11189), .ZN(n11191) );
  AOI22_X1 U14363 ( .A1(n17236), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11194) );
  OAI21_X1 U14364 ( .B1(n10244), .B2(n18463), .A(n11194), .ZN(n11203) );
  AOI22_X1 U14365 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11201) );
  INV_X1 U14366 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18489) );
  OAI22_X1 U14367 ( .A1(n17246), .A2(n18489), .B1(n11038), .B2(n18542), .ZN(
        n11199) );
  AOI22_X1 U14368 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14369 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17235), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14370 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11195) );
  NAND3_X1 U14371 ( .A1(n11197), .A2(n11196), .A3(n11195), .ZN(n11198) );
  AOI211_X1 U14372 ( .C1(n17237), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n11199), .B(n11198), .ZN(n11200) );
  OAI211_X1 U14373 ( .C1(n17151), .C2(n17234), .A(n11201), .B(n11200), .ZN(
        n11202) );
  AOI22_X1 U14374 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14375 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14376 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11204) );
  OAI211_X1 U14377 ( .C1(n17163), .C2(n17143), .A(n11205), .B(n11204), .ZN(
        n11211) );
  AOI22_X1 U14378 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14379 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14380 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11207) );
  NAND2_X1 U14381 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11206) );
  NAND4_X1 U14382 ( .A1(n11209), .A2(n11208), .A3(n11207), .A4(n11206), .ZN(
        n11210) );
  OAI211_X1 U14383 ( .C1(n17246), .C2(n18506), .A(n11213), .B(n11212), .ZN(
        n11246) );
  AOI22_X1 U14384 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14385 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14386 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11221) );
  INV_X1 U14387 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17041) );
  OAI22_X1 U14388 ( .A1(n17177), .A2(n17041), .B1(n9842), .B2(n21086), .ZN(
        n11219) );
  AOI22_X1 U14389 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14390 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14391 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U14392 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11214) );
  NAND4_X1 U14393 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(
        n11218) );
  AOI211_X1 U14394 ( .C1(n11065), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n11219), .B(n11218), .ZN(n11220) );
  NAND4_X1 U14395 ( .A1(n11223), .A2(n11222), .A3(n11221), .A4(n11220), .ZN(
        n11238) );
  NAND2_X1 U14396 ( .A1(n11246), .A2(n11238), .ZN(n15802) );
  NAND4_X1 U14397 ( .A1(n18282), .A2(n18278), .A3(n11250), .A4(n11241), .ZN(
        n11247) );
  INV_X1 U14398 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U14399 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11065), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11232) );
  AOI22_X1 U14400 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14401 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U14402 ( .A1(n11225), .A2(n11224), .ZN(n11230) );
  INV_X1 U14403 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18494) );
  AOI22_X1 U14404 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14405 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11227) );
  OAI211_X1 U14406 ( .C1(n17246), .C2(n18494), .A(n11228), .B(n11227), .ZN(
        n11229) );
  AOI211_X1 U14407 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n11230), .B(n11229), .ZN(n11231) );
  OAI211_X1 U14408 ( .C1(n17186), .C2(n17193), .A(n11232), .B(n11231), .ZN(
        n11236) );
  OAI22_X1 U14409 ( .A1(n9841), .A2(n17201), .B1(n11038), .B2(n21093), .ZN(
        n11233) );
  NAND2_X1 U14410 ( .A1(n13836), .A2(n18291), .ZN(n18735) );
  NOR2_X1 U14411 ( .A1(n11238), .A2(n18291), .ZN(n11266) );
  INV_X1 U14412 ( .A(n11266), .ZN(n11248) );
  NAND3_X1 U14413 ( .A1(n9815), .A2(n18735), .A3(n11248), .ZN(n11237) );
  NAND2_X1 U14414 ( .A1(n9815), .A2(n11238), .ZN(n15809) );
  INV_X1 U14415 ( .A(n18760), .ZN(n15889) );
  NAND2_X1 U14416 ( .A1(n18272), .A2(n17444), .ZN(n11254) );
  AOI21_X1 U14417 ( .B1(n17333), .B2(n15889), .A(n11254), .ZN(n15785) );
  AOI21_X1 U14418 ( .B1(n11237), .B2(n15809), .A(n15785), .ZN(n11244) );
  INV_X1 U14419 ( .A(n18278), .ZN(n11245) );
  OAI22_X1 U14420 ( .A1(n11250), .A2(n11245), .B1(n17444), .B2(n11237), .ZN(
        n11243) );
  AOI211_X1 U14421 ( .C1(n18282), .C2(n11238), .A(n11267), .B(n9796), .ZN(
        n11240) );
  OAI21_X1 U14422 ( .B1(n11241), .B2(n18297), .A(n13836), .ZN(n11239) );
  OAI21_X1 U14423 ( .B1(n11241), .B2(n11240), .A(n11239), .ZN(n11242) );
  NOR2_X1 U14424 ( .A1(n11243), .A2(n11242), .ZN(n15787) );
  OAI21_X1 U14425 ( .B1(n18278), .B2(n11244), .A(n15787), .ZN(n11252) );
  INV_X1 U14426 ( .A(n11267), .ZN(n11255) );
  NAND2_X1 U14427 ( .A1(n9815), .A2(n18278), .ZN(n18734) );
  INV_X1 U14428 ( .A(n13837), .ZN(n11249) );
  AND3_X1 U14429 ( .A1(n18933), .A2(n18724), .A3(n11251), .ZN(n11253) );
  OAI21_X1 U14430 ( .B1(n18282), .B2(n18760), .A(n11256), .ZN(n11265) );
  INV_X1 U14431 ( .A(n11257), .ZN(n11264) );
  XNOR2_X1 U14432 ( .A(n11259), .B(n11258), .ZN(n11262) );
  INV_X1 U14433 ( .A(n18725), .ZN(n15810) );
  OAI21_X1 U14434 ( .B1(n11264), .B2(n11263), .A(n15810), .ZN(n18728) );
  NAND2_X1 U14435 ( .A1(n9815), .A2(n18933), .ZN(n15807) );
  NOR3_X1 U14436 ( .A1(n11267), .A2(n11266), .A3(n11265), .ZN(n15788) );
  INV_X1 U14437 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n21022) );
  NAND2_X1 U14438 ( .A1(n21022), .A2(n18626), .ZN(n18892) );
  INV_X1 U14439 ( .A(n18892), .ZN(n18949) );
  NAND2_X1 U14440 ( .A1(n18948), .A2(n18626), .ZN(n16578) );
  INV_X1 U14441 ( .A(n16578), .ZN(n11268) );
  NOR2_X1 U14442 ( .A1(n18949), .A2(n11268), .ZN(n18938) );
  NAND2_X1 U14443 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17816) );
  INV_X1 U14444 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11269) );
  NOR2_X1 U14445 ( .A1(n17834), .A2(n16849), .ZN(n17778) );
  INV_X1 U14446 ( .A(n17778), .ZN(n17826) );
  NAND3_X1 U14447 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17780) );
  NOR2_X1 U14448 ( .A1(n17826), .A2(n17780), .ZN(n16786) );
  NAND2_X1 U14449 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17748) );
  NAND2_X1 U14450 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17713) );
  NAND2_X1 U14451 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17674) );
  NAND2_X1 U14452 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17662), .ZN(
        n17639) );
  NAND2_X1 U14453 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17640) );
  NAND2_X1 U14454 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17592) );
  NAND2_X1 U14455 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17554) );
  NAND2_X1 U14456 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16445), .ZN(
        n16431) );
  XOR2_X2 U14457 ( .A(n11269), .B(n16431), .Z(n16913) );
  INV_X1 U14458 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18878) );
  NOR2_X1 U14459 ( .A1(n18878), .A2(n16718), .ZN(n16461) );
  INV_X1 U14460 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16614) );
  INV_X1 U14461 ( .A(n18911), .ZN(n18722) );
  AOI22_X1 U14462 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18948), .B1(
        P3_STATE2_REG_2__SCAN_IN), .B2(n21022), .ZN(n18802) );
  INV_X1 U14463 ( .A(n11272), .ZN(n16430) );
  NOR2_X1 U14464 ( .A1(n16614), .A2(n16430), .ZN(n11273) );
  NOR2_X1 U14465 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17661), .ZN(
        n16446) );
  NAND2_X1 U14466 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16444), .ZN(
        n16605) );
  INV_X1 U14467 ( .A(n16605), .ZN(n11271) );
  NAND2_X1 U14468 ( .A1(n18392), .A2(n11270), .ZN(n16449) );
  OAI211_X1 U14469 ( .C1(n11271), .C2(n18803), .A(n17916), .B(n16449), .ZN(
        n16452) );
  NAND2_X1 U14470 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17942) );
  INV_X1 U14471 ( .A(n17942), .ZN(n17945) );
  NAND3_X1 U14472 ( .A1(n17945), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16428) );
  NOR2_X1 U14473 ( .A1(n16427), .A2(n16428), .ZN(n16464) );
  NAND2_X1 U14474 ( .A1(n18058), .A2(n16464), .ZN(n17923) );
  NOR2_X1 U14475 ( .A1(n17923), .A2(n16458), .ZN(n16437) );
  NAND2_X1 U14476 ( .A1(n16437), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11275) );
  XOR2_X1 U14477 ( .A(n18900), .B(n11275), .Z(n16466) );
  NOR2_X4 U14478 ( .A1(n18933), .A2(n16583), .ZN(n17909) );
  INV_X1 U14479 ( .A(n11276), .ZN(n15890) );
  NAND2_X1 U14480 ( .A1(n17433), .A2(n15890), .ZN(n11285) );
  INV_X1 U14481 ( .A(n11285), .ZN(n11277) );
  NOR2_X1 U14482 ( .A1(n11277), .A2(n17430), .ZN(n11283) );
  NOR2_X1 U14483 ( .A1(n11282), .A2(n11283), .ZN(n11281) );
  NAND2_X1 U14484 ( .A1(n11281), .A2(n11280), .ZN(n11279) );
  NOR2_X1 U14485 ( .A1(n17417), .A2(n11279), .ZN(n17844) );
  NAND2_X1 U14486 ( .A1(n17844), .A2(n11297), .ZN(n11278) );
  NOR2_X1 U14487 ( .A1(n17410), .A2(n11278), .ZN(n11304) );
  XOR2_X1 U14488 ( .A(n17410), .B(n11278), .Z(n11300) );
  XOR2_X1 U14489 ( .A(n17417), .B(n11279), .Z(n11294) );
  AND2_X1 U14490 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11294), .ZN(
        n11296) );
  INV_X1 U14491 ( .A(n11280), .ZN(n17421) );
  XNOR2_X1 U14492 ( .A(n17421), .B(n11281), .ZN(n11292) );
  AND2_X1 U14493 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11292), .ZN(
        n11293) );
  XOR2_X1 U14494 ( .A(n11283), .B(n11282), .Z(n11290) );
  AND2_X1 U14495 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11290), .ZN(
        n11291) );
  AOI21_X1 U14496 ( .B1(n11284), .B2(n15890), .A(n11283), .ZN(n11287) );
  NOR2_X1 U14497 ( .A1(n11287), .A2(n18216), .ZN(n11289) );
  OR2_X1 U14498 ( .A1(n17433), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11286) );
  INV_X1 U14499 ( .A(n17906), .ZN(n17908) );
  NOR2_X1 U14500 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15890), .ZN(
        n17914) );
  NAND2_X1 U14501 ( .A1(n17908), .A2(n17914), .ZN(n17907) );
  NAND3_X1 U14502 ( .A1(n11286), .A2(n11285), .A3(n17907), .ZN(n17899) );
  XNOR2_X1 U14503 ( .A(n18216), .B(n11287), .ZN(n17898) );
  NOR2_X1 U14504 ( .A1(n17899), .A2(n17898), .ZN(n11288) );
  NOR2_X1 U14505 ( .A1(n11289), .A2(n11288), .ZN(n17887) );
  XOR2_X1 U14506 ( .A(n18195), .B(n11290), .Z(n17886) );
  NOR2_X1 U14507 ( .A1(n17887), .A2(n17886), .ZN(n17885) );
  NOR2_X1 U14508 ( .A1(n11291), .A2(n17885), .ZN(n17876) );
  XOR2_X1 U14509 ( .A(n18194), .B(n11292), .Z(n17875) );
  NOR2_X1 U14510 ( .A1(n17876), .A2(n17875), .ZN(n17874) );
  NOR2_X1 U14511 ( .A1(n11293), .A2(n17874), .ZN(n17861) );
  INV_X1 U14512 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11295) );
  XOR2_X1 U14513 ( .A(n11295), .B(n11294), .Z(n17860) );
  NOR2_X1 U14514 ( .A1(n17861), .A2(n17860), .ZN(n17859) );
  INV_X1 U14515 ( .A(n11297), .ZN(n17414) );
  INV_X1 U14516 ( .A(n17844), .ZN(n17842) );
  XNOR2_X1 U14517 ( .A(n17414), .B(n17842), .ZN(n11298) );
  AOI222_X1 U14518 ( .A1(n17843), .A2(n18181), .B1(n17843), .B2(n11298), .C1(
        n18181), .C2(n11298), .ZN(n11301) );
  NOR2_X1 U14519 ( .A1(n11300), .A2(n11301), .ZN(n17836) );
  INV_X1 U14520 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21142) );
  NOR2_X1 U14521 ( .A1(n17836), .A2(n21142), .ZN(n11299) );
  NAND2_X1 U14522 ( .A1(n11304), .A2(n11299), .ZN(n11305) );
  INV_X1 U14523 ( .A(n11299), .ZN(n11303) );
  AND2_X1 U14524 ( .A1(n11301), .A2(n11300), .ZN(n17837) );
  AOI21_X1 U14525 ( .B1(n11304), .B2(n11303), .A(n17837), .ZN(n11302) );
  OAI21_X1 U14526 ( .B1(n11304), .B2(n11303), .A(n11302), .ZN(n17822) );
  NAND2_X1 U14527 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17822), .ZN(
        n17821) );
  NAND2_X1 U14528 ( .A1(n18055), .A2(n16425), .ZN(n17737) );
  NAND2_X1 U14529 ( .A1(n16464), .A2(n18057), .ZN(n17924) );
  NOR2_X1 U14530 ( .A1(n16458), .A2(n17924), .ZN(n16436) );
  NAND2_X1 U14531 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16436), .ZN(
        n11306) );
  XOR2_X1 U14532 ( .A(n18900), .B(n11306), .Z(n16465) );
  AOI22_X1 U14533 ( .A1(n17825), .A2(n16466), .B1(n17909), .B2(n16465), .ZN(
        n11307) );
  OAI21_X1 U14534 ( .B1(n16469), .B2(n17823), .A(n11309), .ZN(P3_U2799) );
  NOR2_X1 U14535 ( .A1(n11310), .A2(n11582), .ZN(n11311) );
  OR2_X1 U14536 ( .A1(n11332), .A2(n11311), .ZN(n11327) );
  OAI21_X1 U14537 ( .B1(n11313), .B2(n11314), .A(n10376), .ZN(n11318) );
  INV_X1 U14538 ( .A(n11314), .ZN(n11316) );
  OAI211_X1 U14539 ( .C1(n14316), .C2(n11316), .A(n11555), .B(n11315), .ZN(
        n11317) );
  OAI211_X1 U14540 ( .C1(n11312), .C2(n11319), .A(n11318), .B(n11317), .ZN(
        n11323) );
  NAND2_X1 U14541 ( .A1(n10540), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U14542 ( .A1(n11331), .A2(n14316), .ZN(n11320) );
  MUX2_X1 U14543 ( .A(n11582), .B(n11320), .S(n11319), .Z(n11322) );
  AOI21_X1 U14544 ( .B1(n11323), .B2(n11322), .A(n11321), .ZN(n11324) );
  AOI21_X1 U14545 ( .B1(n11325), .B2(n11582), .A(n11324), .ZN(n11326) );
  NOR2_X1 U14546 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  MUX2_X1 U14547 ( .A(n11329), .B(n11328), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n11330) );
  NAND2_X1 U14548 ( .A1(n11332), .A2(n19208), .ZN(n11333) );
  NAND2_X1 U14549 ( .A1(n16402), .A2(n14316), .ZN(n19203) );
  NAND2_X1 U14550 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19983) );
  INV_X1 U14551 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19849) );
  NAND2_X2 U14552 ( .A1(n19988), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19911) );
  NOR2_X1 U14553 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19845) );
  INV_X1 U14554 ( .A(n19845), .ZN(n19855) );
  NAND3_X1 U14555 ( .A1(n19849), .A2(n19911), .A3(n19855), .ZN(n19204) );
  NAND2_X1 U14556 ( .A1(n11334), .A2(n16388), .ZN(n11357) );
  AOI21_X1 U14557 ( .B1(n11335), .B2(n11555), .A(n10354), .ZN(n11336) );
  NAND2_X1 U14558 ( .A1(n19203), .A2(n11336), .ZN(n11356) );
  MUX2_X1 U14559 ( .A(n11337), .B(n10364), .S(n14294), .Z(n11338) );
  OR2_X1 U14560 ( .A1(n11338), .A2(n19976), .ZN(n11352) );
  NAND2_X1 U14561 ( .A1(n10328), .A2(n16388), .ZN(n11339) );
  OR2_X1 U14562 ( .A1(n16398), .A2(n11339), .ZN(n11351) );
  NAND2_X1 U14563 ( .A1(n11341), .A2(n10364), .ZN(n11342) );
  NAND2_X1 U14564 ( .A1(n11340), .A2(n11342), .ZN(n11349) );
  OAI21_X1 U14565 ( .B1(n14316), .B2(n10354), .A(n11555), .ZN(n11343) );
  NAND2_X1 U14566 ( .A1(n11343), .A2(n12972), .ZN(n11344) );
  AOI21_X1 U14567 ( .B1(n11344), .B2(n10364), .A(n11549), .ZN(n11348) );
  INV_X1 U14568 ( .A(n19969), .ZN(n11345) );
  OAI21_X1 U14569 ( .B1(n11346), .B2(n19340), .A(n11345), .ZN(n11558) );
  AND4_X1 U14570 ( .A1(n11349), .A2(n11348), .A3(n11558), .A4(n11347), .ZN(
        n11350) );
  AND2_X1 U14571 ( .A1(n11351), .A2(n11350), .ZN(n15700) );
  OAI21_X1 U14572 ( .B1(n16398), .B2(n11352), .A(n15700), .ZN(n11353) );
  NOR2_X1 U14573 ( .A1(n11354), .A2(n11353), .ZN(n11355) );
  OAI211_X1 U14574 ( .C1(n19203), .C2(n11357), .A(n11356), .B(n11355), .ZN(
        n11358) );
  NAND2_X1 U14575 ( .A1(n11585), .A2(n11359), .ZN(n19296) );
  NOR2_X1 U14576 ( .A1(n15125), .A2(n19296), .ZN(n11581) );
  NAND2_X1 U14577 ( .A1(n11360), .A2(n14316), .ZN(n11362) );
  NAND2_X1 U14578 ( .A1(n11362), .A2(n15744), .ZN(n11363) );
  NAND2_X1 U14579 ( .A1(n14043), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11366) );
  NAND2_X1 U14580 ( .A1(n12972), .A2(n19951), .ZN(n11376) );
  INV_X1 U14581 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12987) );
  NAND2_X1 U14582 ( .A1(n19951), .A2(n12987), .ZN(n11364) );
  AOI22_X1 U14583 ( .A1(n14316), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n11376), .B2(n11364), .ZN(n11365) );
  NAND2_X1 U14584 ( .A1(n11366), .A2(n11365), .ZN(n12974) );
  INV_X1 U14585 ( .A(n11367), .ZN(n11368) );
  NAND2_X1 U14586 ( .A1(n11372), .A2(n11368), .ZN(n11384) );
  OAI21_X1 U14587 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19951), .A(
        n11376), .ZN(n11369) );
  AND2_X1 U14588 ( .A1(n11384), .A2(n11369), .ZN(n11371) );
  OR2_X1 U14589 ( .A1(n12863), .A2(n11511), .ZN(n11370) );
  INV_X2 U14590 ( .A(n9839), .ZN(n13934) );
  AOI22_X1 U14591 ( .A1(n11372), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n11374) );
  INV_X1 U14592 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19862) );
  NAND2_X1 U14593 ( .A1(n14043), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U14594 ( .A1(n11374), .A2(n11373), .ZN(n11382) );
  INV_X1 U14595 ( .A(n11375), .ZN(n11379) );
  INV_X1 U14596 ( .A(n11376), .ZN(n11377) );
  AOI22_X1 U14597 ( .A1(n11367), .A2(n11377), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11378) );
  OAI21_X1 U14598 ( .B1(n11380), .B2(n11379), .A(n11378), .ZN(n13052) );
  INV_X1 U14599 ( .A(n11383), .ZN(n11386) );
  NAND2_X1 U14600 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11385) );
  OAI211_X1 U14601 ( .C1(n11511), .C2(n11386), .A(n11385), .B(n11384), .ZN(
        n11389) );
  XNOR2_X1 U14602 ( .A(n11390), .B(n11389), .ZN(n13250) );
  AOI22_X1 U14603 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n11388) );
  NAND2_X1 U14604 ( .A1(n14043), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11387) );
  NAND2_X1 U14605 ( .A1(n11388), .A2(n11387), .ZN(n13249) );
  NOR2_X1 U14606 ( .A1(n11390), .A2(n11389), .ZN(n11391) );
  NAND2_X1 U14607 ( .A1(n11470), .A2(n11392), .ZN(n11396) );
  NAND2_X1 U14608 ( .A1(n14043), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14609 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11394) );
  NAND2_X1 U14610 ( .A1(n13934), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11393) );
  NAND4_X1 U14611 ( .A1(n11396), .A2(n11395), .A3(n11394), .A4(n11393), .ZN(
        n13349) );
  NAND2_X1 U14612 ( .A1(n11470), .A2(n11397), .ZN(n11400) );
  NAND2_X1 U14613 ( .A1(n14043), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14614 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14615 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11402) );
  NAND2_X1 U14616 ( .A1(n14043), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11401) );
  OAI211_X1 U14617 ( .C1(n11403), .C2(n11511), .A(n11402), .B(n11401), .ZN(
        n13588) );
  NOR2_X1 U14618 ( .A1(n11511), .A2(n11404), .ZN(n11405) );
  AOI21_X1 U14619 ( .B1(n13587), .B2(n13588), .A(n11405), .ZN(n12996) );
  NAND2_X1 U14620 ( .A1(n14043), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11407) );
  INV_X2 U14621 ( .A(n11524), .ZN(n11516) );
  AOI22_X1 U14622 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n11406) );
  INV_X1 U14623 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19254) );
  INV_X1 U14624 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19872) );
  OAI222_X1 U14625 ( .A1(n11524), .A2(n15664), .B1(n9839), .B2(n19254), .C1(
        n11528), .C2(n19872), .ZN(n13034) );
  AOI22_X1 U14626 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14627 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14628 ( .A1(n14142), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14629 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11408) );
  NAND4_X1 U14630 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(
        n11417) );
  AOI22_X1 U14631 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14632 ( .A1(n10573), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14633 ( .A1(n14130), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14634 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11412) );
  NAND4_X1 U14635 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(
        n11416) );
  OR2_X1 U14636 ( .A1(n11417), .A2(n11416), .ZN(n13192) );
  NAND2_X1 U14637 ( .A1(n11470), .A2(n13192), .ZN(n11420) );
  NAND2_X1 U14638 ( .A1(n14043), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14639 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14640 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14641 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14642 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14643 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14142), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11421) );
  NAND4_X1 U14644 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .ZN(
        n11430) );
  AOI22_X1 U14645 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n14151), .ZN(n11428) );
  AOI22_X1 U14646 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14647 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14648 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11425) );
  NAND4_X1 U14649 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(
        n11429) );
  AOI22_X1 U14650 ( .A1(n11470), .A2(n13261), .B1(n14043), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14651 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11431) );
  NAND2_X1 U14652 ( .A1(n11432), .A2(n11431), .ZN(n13158) );
  AOI22_X1 U14653 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14141), .B1(
        n10678), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14654 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14655 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10684), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14656 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14142), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U14657 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n11443) );
  INV_X1 U14658 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14212) );
  INV_X1 U14659 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14221) );
  OAI22_X1 U14660 ( .A1(n14212), .A2(n10668), .B1(n10738), .B2(n14221), .ZN(
        n11437) );
  INV_X1 U14661 ( .A(n11437), .ZN(n11441) );
  AOI22_X1 U14662 ( .A1(n10573), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n14151), .ZN(n11440) );
  AOI22_X1 U14663 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14664 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11438) );
  NAND4_X1 U14665 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n11442) );
  INV_X1 U14666 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14667 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n11444) );
  OAI21_X1 U14668 ( .B1(n11528), .B2(n11445), .A(n11444), .ZN(n11446) );
  AOI21_X1 U14669 ( .B1(n11470), .B2(n13208), .A(n11446), .ZN(n16324) );
  AOI22_X1 U14670 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14671 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14672 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14673 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14142), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11448) );
  NAND4_X1 U14674 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11457) );
  AOI22_X1 U14675 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14151), .ZN(n11455) );
  AOI22_X1 U14676 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14677 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14678 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11452) );
  NAND4_X1 U14679 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11456) );
  NOR2_X1 U14680 ( .A1(n11457), .A2(n11456), .ZN(n13331) );
  AOI22_X1 U14681 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11459) );
  NAND2_X1 U14682 ( .A1(n14043), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11458) );
  OAI211_X1 U14683 ( .C1(n13331), .C2(n11511), .A(n11459), .B(n11458), .ZN(
        n13276) );
  NAND2_X1 U14684 ( .A1(n13275), .A2(n13276), .ZN(n13274) );
  AOI22_X1 U14685 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14686 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14142), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14687 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10684), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14688 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11460) );
  NAND4_X1 U14689 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(
        n11469) );
  AOI22_X1 U14690 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n14151), .ZN(n11467) );
  AOI22_X1 U14691 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10669), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U14692 ( .A1(n14130), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14693 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11464) );
  NAND4_X1 U14694 ( .A1(n11467), .A2(n11466), .A3(n11465), .A4(n11464), .ZN(
        n11468) );
  NAND2_X1 U14695 ( .A1(n11470), .A2(n13393), .ZN(n11473) );
  NAND2_X1 U14696 ( .A1(n14043), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14697 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n11471) );
  NOR2_X2 U14698 ( .A1(n13274), .A2(n15617), .ZN(n15616) );
  AOI22_X1 U14699 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14700 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14701 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14702 ( .A1(n14142), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11474) );
  NAND4_X1 U14703 ( .A1(n11477), .A2(n11476), .A3(n11475), .A4(n11474), .ZN(
        n11483) );
  AOI22_X1 U14704 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14705 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14706 ( .A1(n10669), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14707 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11478) );
  NAND4_X1 U14708 ( .A1(n11481), .A2(n11480), .A3(n11479), .A4(n11478), .ZN(
        n11482) );
  INV_X1 U14709 ( .A(n13467), .ZN(n11486) );
  AOI22_X1 U14710 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11485) );
  NAND2_X1 U14711 ( .A1(n14043), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11484) );
  OAI211_X1 U14712 ( .C1(n11486), .C2(n11511), .A(n11485), .B(n11484), .ZN(
        n13420) );
  AOI22_X1 U14713 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14141), .B1(
        n10678), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14714 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14715 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10684), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14716 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n14142), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11487) );
  NAND4_X1 U14717 ( .A1(n11490), .A2(n11489), .A3(n11488), .A4(n11487), .ZN(
        n11496) );
  AOI22_X1 U14718 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n14151), .ZN(n11494) );
  AOI22_X1 U14719 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14720 ( .A1(n14130), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U14721 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11491) );
  NAND4_X1 U14722 ( .A1(n11494), .A2(n11493), .A3(n11492), .A4(n11491), .ZN(
        n11495) );
  NOR2_X1 U14723 ( .A1(n11496), .A2(n11495), .ZN(n13468) );
  AOI22_X1 U14724 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11498) );
  NAND2_X1 U14725 ( .A1(n14043), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11497) );
  OAI211_X1 U14726 ( .C1(n13468), .C2(n11511), .A(n11498), .B(n11497), .ZN(
        n15585) );
  AOI22_X1 U14727 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14728 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14729 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14730 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14142), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11499) );
  NAND4_X1 U14731 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n11508) );
  AOI22_X1 U14732 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n14151), .ZN(n11506) );
  AOI22_X1 U14733 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14734 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14735 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11503) );
  NAND4_X1 U14736 ( .A1(n11506), .A2(n11505), .A3(n11504), .A4(n11503), .ZN(
        n11507) );
  NOR2_X1 U14737 ( .A1(n11508), .A2(n11507), .ZN(n15221) );
  AOI22_X1 U14738 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U14739 ( .A1(n14043), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11509) );
  OAI211_X1 U14740 ( .C1(n15221), .C2(n11511), .A(n11510), .B(n11509), .ZN(
        n13503) );
  NAND2_X1 U14741 ( .A1(n14043), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14742 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14743 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U14744 ( .A1(n14043), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11514) );
  NAND2_X1 U14745 ( .A1(n11515), .A2(n11514), .ZN(n15290) );
  NAND2_X1 U14746 ( .A1(n14043), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14747 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n11517) );
  NAND2_X1 U14748 ( .A1(n14043), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14749 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n11519) );
  INV_X1 U14750 ( .A(n15279), .ZN(n11521) );
  NAND2_X1 U14751 ( .A1(n15087), .A2(n11521), .ZN(n15516) );
  NAND2_X1 U14752 ( .A1(n14043), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14753 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n11522) );
  INV_X1 U14754 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19893) );
  INV_X1 U14755 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19228) );
  OAI222_X1 U14756 ( .A1(n11528), .A2(n19893), .B1(n9839), .B2(n19228), .C1(
        n11612), .C2(n11524), .ZN(n11611) );
  AOI22_X1 U14757 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11526) );
  NAND2_X1 U14758 ( .A1(n14043), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U14759 ( .A1(n11526), .A2(n11525), .ZN(n15502) );
  INV_X1 U14760 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U14761 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11527) );
  OAI21_X1 U14762 ( .B1(n19897), .B2(n11528), .A(n11527), .ZN(n15268) );
  NAND2_X1 U14763 ( .A1(n14043), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14764 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n11529) );
  AND2_X1 U14765 ( .A1(n11530), .A2(n11529), .ZN(n15073) );
  OR2_X2 U14766 ( .A1(n15267), .A2(n15073), .ZN(n15253) );
  NAND2_X1 U14767 ( .A1(n14043), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14768 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n11531) );
  NOR2_X2 U14769 ( .A1(n15253), .A2(n15254), .ZN(n15247) );
  AOI22_X1 U14770 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11534) );
  NAND2_X1 U14771 ( .A1(n14043), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U14772 ( .A1(n11534), .A2(n11533), .ZN(n15246) );
  NAND2_X1 U14773 ( .A1(n14043), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14774 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11535) );
  AND2_X1 U14775 ( .A1(n11536), .A2(n11535), .ZN(n13992) );
  NAND2_X1 U14776 ( .A1(n14043), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14777 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n11537) );
  AND2_X1 U14778 ( .A1(n11538), .A2(n11537), .ZN(n13970) );
  AOI22_X1 U14779 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n11540) );
  NAND2_X1 U14780 ( .A1(n14043), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11539) );
  NAND2_X1 U14781 ( .A1(n11540), .A2(n11539), .ZN(n11542) );
  NOR2_X1 U14782 ( .A1(n11541), .A2(n11542), .ZN(n11543) );
  INV_X1 U14783 ( .A(n14051), .ZN(n13932) );
  NAND2_X1 U14784 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15448) );
  NOR2_X1 U14785 ( .A1(n15474), .A2(n15448), .ZN(n11577) );
  NOR2_X1 U14786 ( .A1(n20965), .A2(n10999), .ZN(n15486) );
  INV_X1 U14787 ( .A(n15486), .ZN(n11574) );
  NOR2_X1 U14788 ( .A1(n16333), .A2(n15664), .ZN(n11572) );
  NAND2_X1 U14789 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13585) );
  INV_X1 U14790 ( .A(n13585), .ZN(n11564) );
  AND3_X1 U14791 ( .A1(n13515), .A2(n10364), .A3(n14294), .ZN(n11544) );
  AND2_X1 U14792 ( .A1(n11361), .A2(n11544), .ZN(n15743) );
  NAND2_X1 U14793 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19306) );
  NOR2_X1 U14794 ( .A1(n19297), .A2(n19306), .ZN(n19291) );
  NAND2_X1 U14795 ( .A1(n19297), .A2(n19306), .ZN(n11569) );
  INV_X1 U14796 ( .A(n11545), .ZN(n11548) );
  OAI21_X1 U14797 ( .B1(n11548), .B2(n11547), .A(n11546), .ZN(n11552) );
  INV_X1 U14798 ( .A(n11549), .ZN(n11550) );
  OAI21_X1 U14799 ( .B1(n11546), .B2(n10354), .A(n11550), .ZN(n11551) );
  NAND2_X1 U14800 ( .A1(n11552), .A2(n11551), .ZN(n11554) );
  OAI211_X1 U14801 ( .C1(n10364), .C2(n11555), .A(n11554), .B(n11553), .ZN(
        n11556) );
  INV_X1 U14802 ( .A(n11556), .ZN(n11561) );
  NAND2_X1 U14803 ( .A1(n11557), .A2(n14316), .ZN(n15691) );
  NAND2_X1 U14804 ( .A1(n15691), .A2(n11558), .ZN(n11559) );
  NAND2_X1 U14805 ( .A1(n11559), .A2(n10344), .ZN(n11560) );
  INV_X1 U14806 ( .A(n11562), .ZN(n15727) );
  NAND2_X1 U14807 ( .A1(n15715), .A2(n15727), .ZN(n11563) );
  OAI211_X1 U14808 ( .C1(n19289), .C2(n19291), .A(n11569), .B(n16364), .ZN(
        n16355) );
  NOR2_X1 U14809 ( .A1(n16356), .A2(n16355), .ZN(n13586) );
  NAND2_X1 U14810 ( .A1(n11564), .A2(n13586), .ZN(n15676) );
  NAND2_X1 U14811 ( .A1(n11572), .A2(n16342), .ZN(n15634) );
  NOR3_X1 U14812 ( .A1(n11575), .A2(n11574), .A3(n15634), .ZN(n15469) );
  NAND2_X1 U14813 ( .A1(n11577), .A2(n15469), .ZN(n13972) );
  INV_X1 U14814 ( .A(n13972), .ZN(n14049) );
  OAI211_X1 U14815 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n13971), .A(
        n13932), .B(n14049), .ZN(n11565) );
  OAI211_X1 U14816 ( .C1(n16360), .C2(n16177), .A(n11566), .B(n11565), .ZN(
        n11567) );
  NAND2_X1 U14817 ( .A1(n15559), .A2(n19306), .ZN(n11568) );
  OR2_X1 U14818 ( .A1(n11585), .A2(n19088), .ZN(n16358) );
  NAND2_X1 U14819 ( .A1(n15562), .A2(n19298), .ZN(n15471) );
  INV_X1 U14820 ( .A(n11569), .ZN(n19290) );
  NAND2_X1 U14821 ( .A1(n15559), .A2(n19297), .ZN(n19307) );
  NAND3_X1 U14822 ( .A1(n19298), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n19307), .ZN(n11570) );
  AOI21_X1 U14823 ( .B1(n19289), .B2(n19290), .A(n11570), .ZN(n16357) );
  NOR2_X1 U14824 ( .A1(n15446), .A2(n16357), .ZN(n13594) );
  AOI21_X1 U14825 ( .B1(n15471), .B2(n13585), .A(n13594), .ZN(n15674) );
  NAND2_X1 U14826 ( .A1(n16364), .A2(n15675), .ZN(n11571) );
  INV_X1 U14827 ( .A(n11572), .ZN(n16341) );
  NAND2_X1 U14828 ( .A1(n16364), .A2(n16341), .ZN(n11573) );
  NOR2_X1 U14829 ( .A1(n11575), .A2(n11574), .ZN(n11576) );
  NAND2_X1 U14830 ( .A1(n15649), .A2(n11576), .ZN(n15470) );
  INV_X1 U14831 ( .A(n15470), .ZN(n15447) );
  AOI21_X1 U14832 ( .B1(n15447), .B2(n11577), .A(n15446), .ZN(n14001) );
  NAND2_X1 U14833 ( .A1(n14001), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11578) );
  NOR2_X1 U14834 ( .A1(n10538), .A2(n11582), .ZN(n19963) );
  NAND2_X1 U14835 ( .A1(n11583), .A2(n19303), .ZN(n11586) );
  INV_X1 U14836 ( .A(n11584), .ZN(n19962) );
  NAND3_X1 U14837 ( .A1(n11587), .A2(n11586), .A3(n10247), .ZN(P2_U3017) );
  INV_X1 U14838 ( .A(n15414), .ZN(n11588) );
  INV_X1 U14839 ( .A(n15404), .ZN(n11589) );
  INV_X1 U14840 ( .A(n11590), .ZN(n15393) );
  NAND2_X1 U14841 ( .A1(n11595), .A2(n11592), .ZN(n15385) );
  INV_X1 U14842 ( .A(n15385), .ZN(n11593) );
  NAND2_X1 U14843 ( .A1(n11594), .A2(n11593), .ZN(n11596) );
  AND2_X1 U14844 ( .A1(n10234), .A2(n15349), .ZN(n11597) );
  NAND2_X1 U14845 ( .A1(n11598), .A2(n15348), .ZN(n11601) );
  XNOR2_X1 U14846 ( .A(n11601), .B(n10245), .ZN(n15346) );
  NAND2_X1 U14847 ( .A1(n15371), .A2(n15526), .ZN(n15375) );
  AOI21_X1 U14848 ( .B1(n15361), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11603) );
  INV_X1 U14849 ( .A(n15511), .ZN(n11602) );
  NOR2_X1 U14850 ( .A1(n11603), .A2(n11602), .ZN(n15344) );
  OR2_X1 U14851 ( .A1(n11605), .A2(n11606), .ZN(n11607) );
  NAND2_X1 U14852 ( .A1(n11604), .A2(n11607), .ZN(n18989) );
  OAI21_X1 U14853 ( .B1(n11608), .B2(n15562), .A(n15649), .ZN(n15510) );
  OAI21_X1 U14854 ( .B1(n11609), .B2(n11611), .A(n11610), .ZN(n18999) );
  NAND3_X1 U14855 ( .A1(n15652), .A2(n15526), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15520) );
  NOR2_X1 U14856 ( .A1(n15520), .A2(n15527), .ZN(n15485) );
  NAND2_X1 U14857 ( .A1(n15485), .A2(n11612), .ZN(n11613) );
  NAND2_X1 U14858 ( .A1(n19088), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15338) );
  OAI211_X1 U14859 ( .C1(n16360), .C2(n18999), .A(n11613), .B(n15338), .ZN(
        n11614) );
  AOI21_X1 U14860 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15510), .A(
        n11614), .ZN(n11615) );
  OAI21_X1 U14861 ( .B1(n18989), .B2(n19296), .A(n11615), .ZN(n11616) );
  AOI21_X1 U14862 ( .B1(n15344), .B2(n16337), .A(n11616), .ZN(n11617) );
  OAI21_X1 U14863 ( .B1(n15346), .B2(n16369), .A(n11617), .ZN(P2_U3025) );
  AND2_X4 U14864 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13070) );
  AND2_X4 U14865 ( .A1(n13215), .A2(n13070), .ZN(n11897) );
  NAND2_X1 U14866 ( .A1(n11897), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11624) );
  AND2_X4 U14867 ( .A1(n11619), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13218) );
  AND2_X4 U14868 ( .A1(n13218), .A2(n13070), .ZN(n11875) );
  NAND2_X1 U14869 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11623) );
  AND2_X4 U14870 ( .A1(n11629), .A2(n13218), .ZN(n12291) );
  NAND2_X1 U14871 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11622) );
  NAND2_X1 U14872 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11621) );
  AND2_X4 U14873 ( .A1(n13218), .A2(n13069), .ZN(n11801) );
  NAND2_X1 U14874 ( .A1(n11801), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11628) );
  AND2_X4 U14875 ( .A1(n11634), .A2(n13218), .ZN(n11827) );
  NAND2_X1 U14876 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11627) );
  AND2_X4 U14877 ( .A1(n13215), .A2(n11629), .ZN(n11902) );
  NAND2_X1 U14878 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11626) );
  AND2_X2 U14879 ( .A1(n13069), .A2(n11636), .ZN(n11807) );
  NAND2_X1 U14880 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11625) );
  NAND2_X1 U14881 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11633) );
  AND2_X4 U14882 ( .A1(n11629), .A2(n11636), .ZN(n11828) );
  NAND2_X1 U14883 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11632) );
  AND2_X2 U14884 ( .A1(n11629), .A2(n11635), .ZN(n11802) );
  NAND2_X1 U14885 ( .A1(n11802), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11631) );
  NAND2_X1 U14886 ( .A1(n11729), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11630) );
  AND2_X2 U14887 ( .A1(n13215), .A2(n13069), .ZN(n11785) );
  NAND2_X1 U14888 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11640) );
  NAND2_X1 U14889 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11639) );
  NAND2_X1 U14890 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11638) );
  AND2_X4 U14891 ( .A1(n11636), .A2(n13070), .ZN(n11822) );
  NAND2_X1 U14892 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11637) );
  INV_X1 U14893 ( .A(n11754), .ZN(n12525) );
  AOI22_X1 U14894 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14895 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14896 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11828), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14897 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11897), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11644) );
  AND4_X2 U14898 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11653) );
  AOI22_X1 U14899 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11802), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14900 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11807), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14901 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14902 ( .A1(n11801), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11876), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11648) );
  NAND2_X2 U14904 ( .A1(n11653), .A2(n11652), .ZN(n11753) );
  AOI22_X1 U14905 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11897), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14906 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14907 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14908 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14909 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11828), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14910 ( .A1(n11802), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11807), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14911 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11801), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11658) );
  NAND3_X2 U14912 ( .A1(n10250), .A2(n11662), .A3(n11661), .ZN(n13779) );
  NAND2_X1 U14913 ( .A1(n11663), .A2(n13784), .ZN(n11675) );
  AOI22_X1 U14914 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14915 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14916 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11876), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14917 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11828), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14918 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14919 ( .A1(n11802), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11807), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11668) );
  NAND2_X1 U14920 ( .A1(n13779), .A2(n11706), .ZN(n11674) );
  NAND2_X1 U14921 ( .A1(n11801), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11679) );
  NAND2_X1 U14922 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11678) );
  NAND2_X1 U14923 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11677) );
  NAND2_X1 U14924 ( .A1(n11729), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11676) );
  NAND2_X1 U14925 ( .A1(n11897), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11683) );
  NAND2_X1 U14926 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11682) );
  NAND2_X1 U14927 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11681) );
  NAND2_X1 U14928 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11680) );
  NAND2_X1 U14929 ( .A1(n11802), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11687) );
  NAND2_X1 U14930 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11686) );
  NAND2_X1 U14931 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11685) );
  NAND2_X1 U14932 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11684) );
  NAND2_X1 U14933 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11691) );
  NAND2_X1 U14934 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11690) );
  NAND2_X1 U14935 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11689) );
  NAND2_X1 U14936 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11688) );
  NAND2_X2 U14937 ( .A1(n12524), .A2(n11761), .ZN(n13786) );
  NAND2_X1 U14938 ( .A1(n13824), .A2(n12524), .ZN(n11764) );
  NAND2_X1 U14939 ( .A1(n11754), .A2(n11753), .ZN(n12523) );
  AOI22_X1 U14940 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14941 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11807), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14942 ( .A1(n11802), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11828), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14943 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11897), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14944 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14945 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U14946 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11700) );
  NAND2_X1 U14947 ( .A1(n12523), .A2(n12690), .ZN(n11774) );
  NAND2_X1 U14948 ( .A1(n11801), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11710) );
  NAND2_X1 U14949 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11709) );
  NAND2_X1 U14950 ( .A1(n11802), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11708) );
  NAND2_X1 U14951 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11707) );
  NAND2_X1 U14952 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11714) );
  NAND2_X1 U14953 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11713) );
  NAND2_X1 U14954 ( .A1(n11897), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11712) );
  NAND2_X1 U14955 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11711) );
  NAND2_X1 U14956 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11717) );
  NAND2_X1 U14957 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11716) );
  NAND2_X1 U14958 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11715) );
  NAND2_X1 U14959 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11725) );
  NAND2_X1 U14960 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11724) );
  NAND2_X1 U14961 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11723) );
  NAND2_X1 U14962 ( .A1(n11729), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11722) );
  NAND2_X4 U14963 ( .A1(n11727), .A2(n11726), .ZN(n13794) );
  NAND2_X1 U14964 ( .A1(n13007), .A2(n9816), .ZN(n11728) );
  NAND2_X1 U14965 ( .A1(n11729), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11732) );
  NAND2_X1 U14966 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U14967 ( .A1(n11802), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11730) );
  NAND3_X1 U14968 ( .A1(n11732), .A2(n11731), .A3(n11730), .ZN(n11736) );
  INV_X1 U14969 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11733) );
  NAND2_X1 U14970 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11740) );
  NAND2_X1 U14971 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U14972 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11738) );
  NAND2_X1 U14973 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11737) );
  NAND2_X1 U14974 ( .A1(n11801), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11744) );
  NAND2_X1 U14975 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11743) );
  NAND2_X1 U14976 ( .A1(n11897), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U14977 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11741) );
  NAND2_X1 U14978 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U14979 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11747) );
  NAND2_X1 U14980 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11746) );
  NAND2_X1 U14981 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11745) );
  NAND4_X4 U14982 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n11758) );
  INV_X2 U14983 ( .A(n11753), .ZN(n20254) );
  NAND2_X1 U14984 ( .A1(n20254), .A2(n11759), .ZN(n12474) );
  NAND2_X1 U14985 ( .A1(n20258), .A2(n12524), .ZN(n11755) );
  NOR2_X1 U14986 ( .A1(n12474), .A2(n11755), .ZN(n11756) );
  AND2_X2 U14987 ( .A1(n11756), .A2(n12687), .ZN(n15858) );
  AND2_X4 U14988 ( .A1(n11758), .A2(n13794), .ZN(n12659) );
  NAND2_X1 U14989 ( .A1(n15858), .A2(n12659), .ZN(n12790) );
  NAND2_X1 U14990 ( .A1(n12793), .A2(n12790), .ZN(n13817) );
  NAND2_X2 U14991 ( .A1(n15858), .A2(n13794), .ZN(n12638) );
  NAND2_X1 U14992 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20793) );
  OAI21_X1 U14993 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20793), .ZN(n12661) );
  NOR2_X2 U14994 ( .A1(n9797), .A2(n9805), .ZN(n11773) );
  NOR2_X2 U14995 ( .A1(n12690), .A2(n13779), .ZN(n12998) );
  NAND3_X1 U14996 ( .A1(n11773), .A2(n20254), .A3(n12998), .ZN(n13010) );
  INV_X1 U14998 ( .A(n12690), .ZN(n20245) );
  NAND2_X1 U14999 ( .A1(n20245), .A2(n13794), .ZN(n12551) );
  NAND2_X2 U15000 ( .A1(n12551), .A2(n12530), .ZN(n13179) );
  NAND2_X2 U15001 ( .A1(n20238), .A2(n13794), .ZN(n20874) );
  NAND2_X1 U15002 ( .A1(n13007), .A2(n12529), .ZN(n13795) );
  NAND2_X1 U15003 ( .A1(n13779), .A2(n13794), .ZN(n13792) );
  OAI211_X1 U15004 ( .C1(n20249), .C2(n20874), .A(n13795), .B(n13792), .ZN(
        n11760) );
  NAND2_X1 U15005 ( .A1(n20254), .A2(n11761), .ZN(n11762) );
  AND2_X1 U15006 ( .A1(n11762), .A2(n12524), .ZN(n11777) );
  OR2_X1 U15007 ( .A1(n12523), .A2(n13824), .ZN(n11763) );
  NAND2_X1 U15008 ( .A1(n13001), .A2(n13015), .ZN(n11768) );
  INV_X1 U15009 ( .A(n12998), .ZN(n13099) );
  NAND2_X1 U15010 ( .A1(n13099), .A2(n20238), .ZN(n11766) );
  OAI21_X1 U15011 ( .B1(n11779), .B2(n11766), .A(n11765), .ZN(n11767) );
  NAND4_X1 U15012 ( .A1(n13006), .A2(n11781), .A3(n11768), .A4(n11767), .ZN(
        n12522) );
  NAND2_X1 U15013 ( .A1(n12522), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U15014 ( .A1(n11858), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11772) );
  INV_X1 U15015 ( .A(n20778), .ZN(n11770) );
  MUX2_X1 U15016 ( .A(n11770), .B(n12680), .S(n20863), .Z(n11771) );
  NAND2_X1 U15017 ( .A1(n12985), .A2(n11774), .ZN(n11776) );
  NAND2_X1 U15018 ( .A1(n11765), .A2(n11758), .ZN(n13667) );
  AND3_X1 U15019 ( .A1(n13667), .A2(n19990), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11775) );
  OAI211_X1 U15020 ( .C1(n11777), .C2(n20874), .A(n11776), .B(n11775), .ZN(
        n11778) );
  NAND2_X1 U15021 ( .A1(n11779), .A2(n11773), .ZN(n13013) );
  NAND2_X1 U15022 ( .A1(n12998), .A2(n20258), .ZN(n11780) );
  NAND3_X1 U15023 ( .A1(n13001), .A2(n11758), .A3(n13015), .ZN(n11782) );
  NAND2_X1 U15024 ( .A1(n11938), .A2(n16155), .ZN(n11818) );
  INV_X1 U15025 ( .A(n12755), .ZN(n11816) );
  AOI22_X1 U15026 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U15027 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U15029 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U15030 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11786) );
  NAND4_X1 U15031 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11799) );
  BUF_X1 U15032 ( .A(n11897), .Z(n11790) );
  AOI22_X1 U15033 ( .A1(n11790), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11801), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U15035 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U15036 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11795) );
  BUF_X1 U15038 ( .A(n11822), .Z(n11792) );
  AOI22_X1 U15039 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11794) );
  NAND4_X1 U15040 ( .A1(n11797), .A2(n11796), .A3(n11795), .A4(n11794), .ZN(
        n11798) );
  INV_X1 U15041 ( .A(n12691), .ZN(n11814) );
  AOI22_X1 U15042 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U15043 ( .A1(n12448), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U15044 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U15045 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11803) );
  NAND4_X1 U15046 ( .A1(n11806), .A2(n11805), .A3(n11804), .A4(n11803), .ZN(
        n11813) );
  AOI22_X1 U15047 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U15048 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U15049 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U15050 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11808) );
  NAND4_X1 U15051 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11812) );
  XNOR2_X1 U15052 ( .A(n11814), .B(n12746), .ZN(n11815) );
  NAND2_X1 U15053 ( .A1(n11816), .A2(n11815), .ZN(n11817) );
  INV_X1 U15054 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13417) );
  AOI21_X1 U15055 ( .B1(n20249), .B2(n12746), .A(n16155), .ZN(n11820) );
  NAND2_X1 U15056 ( .A1(n11765), .A2(n12691), .ZN(n11819) );
  INV_X1 U15057 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11837) );
  OR2_X1 U15058 ( .A1(n12755), .A2(n12746), .ZN(n11836) );
  AOI22_X1 U15059 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U15060 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U15061 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12209), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U15062 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11823) );
  NAND4_X1 U15063 ( .A1(n11826), .A2(n11825), .A3(n11824), .A4(n11823), .ZN(
        n11834) );
  AOI22_X1 U15064 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11793), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U15065 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U15066 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U15067 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11829) );
  NAND4_X1 U15068 ( .A1(n11832), .A2(n11831), .A3(n11830), .A4(n11829), .ZN(
        n11833) );
  OR2_X1 U15069 ( .A1(n11896), .A2(n11851), .ZN(n11835) );
  OAI211_X1 U15070 ( .C1(n12493), .C2(n11837), .A(n11836), .B(n11835), .ZN(
        n11838) );
  NAND2_X1 U15071 ( .A1(n11839), .A2(n11838), .ZN(n11840) );
  NAND2_X1 U15072 ( .A1(n11858), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11843) );
  INV_X1 U15073 ( .A(n12680), .ZN(n11893) );
  NAND2_X1 U15074 ( .A1(n20539), .A2(n20863), .ZN(n11841) );
  NAND2_X1 U15075 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11861) );
  AND2_X1 U15076 ( .A1(n20778), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11854) );
  AOI21_X1 U15077 ( .B1(n11893), .B2(n20536), .A(n11854), .ZN(n11842) );
  NAND2_X1 U15078 ( .A1(n11843), .A2(n11842), .ZN(n11845) );
  INV_X1 U15079 ( .A(n20334), .ZN(n11849) );
  INV_X1 U15080 ( .A(n11850), .ZN(n11848) );
  NAND2_X2 U15081 ( .A1(n20334), .A2(n11850), .ZN(n11872) );
  NAND2_X1 U15082 ( .A1(n20276), .A2(n11872), .ZN(n13068) );
  OAI21_X2 U15083 ( .B1(n13068), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11852), 
        .ZN(n12689) );
  INV_X1 U15084 ( .A(n11925), .ZN(n11891) );
  INV_X1 U15085 ( .A(n11844), .ZN(n11857) );
  INV_X1 U15086 ( .A(n11854), .ZN(n11855) );
  NAND2_X1 U15087 ( .A1(n11855), .A2(n13079), .ZN(n11856) );
  NAND2_X1 U15088 ( .A1(n11857), .A2(n11856), .ZN(n11870) );
  NAND2_X1 U15089 ( .A1(n11872), .A2(n11870), .ZN(n11866) );
  NAND2_X1 U15090 ( .A1(n11858), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11864) );
  INV_X1 U15091 ( .A(n11861), .ZN(n11860) );
  INV_X1 U15092 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11859) );
  NAND2_X1 U15093 ( .A1(n11860), .A2(n11859), .ZN(n20575) );
  NAND2_X1 U15094 ( .A1(n11861), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11862) );
  NAND2_X1 U15095 ( .A1(n20575), .A2(n11862), .ZN(n13408) );
  NAND2_X1 U15096 ( .A1(n11893), .A2(n13408), .ZN(n11863) );
  NAND2_X1 U15097 ( .A1(n11864), .A2(n11863), .ZN(n11867) );
  AND2_X1 U15098 ( .A1(n20778), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11868) );
  INV_X1 U15099 ( .A(n11867), .ZN(n11871) );
  INV_X1 U15100 ( .A(n11868), .ZN(n11869) );
  NAND4_X1 U15101 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11873) );
  NAND2_X1 U15102 ( .A1(n11892), .A2(n11873), .ZN(n13097) );
  AOI22_X1 U15103 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U15104 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U15105 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U15106 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11877) );
  NAND4_X1 U15107 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n11886) );
  AOI22_X1 U15108 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U15109 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U15110 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U15111 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11881) );
  NAND4_X1 U15112 ( .A1(n11884), .A2(n11883), .A3(n11882), .A4(n11881), .ZN(
        n11885) );
  NOR2_X1 U15113 ( .A1(n11886), .A2(n11885), .ZN(n12707) );
  OAI22_X2 U15114 ( .A1(n13097), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12707), 
        .B2(n12755), .ZN(n11890) );
  INV_X1 U15115 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11887) );
  OAI22_X1 U15116 ( .A1(n12493), .A2(n11887), .B1(n11896), .B2(n12707), .ZN(
        n11888) );
  INV_X1 U15117 ( .A(n11888), .ZN(n11889) );
  NAND2_X1 U15118 ( .A1(n11858), .A2(n15019), .ZN(n11895) );
  INV_X1 U15119 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20574) );
  NAND3_X1 U15120 ( .A1(n20574), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20453) );
  INV_X1 U15121 ( .A(n20471), .ZN(n20450) );
  NOR3_X1 U15122 ( .A1(n20574), .A2(n11859), .A3(n20539), .ZN(n20723) );
  INV_X1 U15123 ( .A(n20723), .ZN(n20716) );
  AOI21_X1 U15124 ( .B1(n20574), .B2(n20450), .A(n20768), .ZN(n20477) );
  AOI22_X1 U15125 ( .A1(n11893), .A2(n20477), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20778), .ZN(n11894) );
  NAND2_X1 U15126 ( .A1(n20476), .A2(n16155), .ZN(n11910) );
  INV_X1 U15127 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n21076) );
  AOI22_X1 U15128 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U15129 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U15130 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U15131 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11898) );
  NAND4_X1 U15132 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11908) );
  AOI22_X1 U15133 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U15134 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15135 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U15136 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11903) );
  NAND4_X1 U15137 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11907) );
  AOI22_X1 U15138 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12514), .B1(
        n12518), .B2(n12724), .ZN(n11909) );
  INV_X1 U15139 ( .A(n11911), .ZN(n11912) );
  INV_X1 U15140 ( .A(n13402), .ZN(n20367) );
  NAND2_X1 U15141 ( .A1(n11912), .A2(n20367), .ZN(n11913) );
  INV_X1 U15142 ( .A(n20845), .ZN(n11914) );
  NAND2_X1 U15143 ( .A1(n11914), .A2(n12054), .ZN(n11923) );
  NOR2_X1 U15144 ( .A1(n13786), .A2(n20715), .ZN(n11940) );
  INV_X1 U15145 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11920) );
  NOR2_X2 U15146 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12076) );
  NAND2_X1 U15147 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11916) );
  INV_X1 U15148 ( .A(n11916), .ZN(n11918) );
  INV_X1 U15149 ( .A(n11966), .ZN(n11917) );
  OAI21_X1 U15150 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11918), .A(
        n11917), .ZN(n13679) );
  AOI22_X1 U15151 ( .A1(n12076), .A2(n13679), .B1(n12634), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11919) );
  OAI21_X1 U15152 ( .B1(n12434), .B2(n11920), .A(n11919), .ZN(n11921) );
  AOI21_X1 U15153 ( .B1(n11940), .B2(n15019), .A(n11921), .ZN(n11922) );
  XNOR2_X1 U15154 ( .A(n11925), .B(n11924), .ZN(n12698) );
  INV_X1 U15155 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n11927) );
  XNOR2_X1 U15156 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13130) );
  AOI21_X1 U15157 ( .B1(n12076), .B2(n13130), .A(n12634), .ZN(n11926) );
  OAI21_X1 U15158 ( .B1(n12434), .B2(n11927), .A(n11926), .ZN(n11928) );
  AOI21_X1 U15159 ( .B1(n11940), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11928), .ZN(n11929) );
  NAND2_X1 U15160 ( .A1(n12634), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11948) );
  NAND2_X1 U15161 ( .A1(n13242), .A2(n12054), .ZN(n11934) );
  INV_X1 U15162 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11931) );
  INV_X1 U15163 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20170) );
  OAI22_X1 U15164 ( .A1(n12434), .A2(n11931), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20170), .ZN(n11932) );
  AOI21_X1 U15165 ( .B1(n11940), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11932), .ZN(n11933) );
  NAND2_X1 U15166 ( .A1(n11934), .A2(n11933), .ZN(n13092) );
  NAND2_X1 U15167 ( .A1(n12694), .A2(n20258), .ZN(n11937) );
  NAND2_X1 U15168 ( .A1(n11937), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13081) );
  INV_X1 U15170 ( .A(n11940), .ZN(n11964) );
  NAND2_X1 U15171 ( .A1(n20715), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11942) );
  NAND2_X1 U15172 ( .A1(n12635), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11941) );
  OAI211_X1 U15173 ( .C1(n11964), .C2(n13030), .A(n11942), .B(n11941), .ZN(
        n11943) );
  AOI21_X1 U15174 ( .B1(n11939), .B2(n12054), .A(n11943), .ZN(n13080) );
  OR2_X1 U15175 ( .A1(n13081), .A2(n13080), .ZN(n13083) );
  INV_X1 U15176 ( .A(n13080), .ZN(n11944) );
  OR2_X1 U15177 ( .A1(n11944), .A2(n12464), .ZN(n11945) );
  NAND2_X1 U15178 ( .A1(n13083), .A2(n11945), .ZN(n13091) );
  NAND2_X1 U15179 ( .A1(n13092), .A2(n13091), .ZN(n13126) );
  NAND2_X1 U15180 ( .A1(n11947), .A2(n11946), .ZN(n13129) );
  NAND2_X1 U15181 ( .A1(n13282), .A2(n13281), .ZN(n13317) );
  AOI22_X1 U15182 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U15183 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U15184 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12376), .B1(
        n12209), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U15185 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11950) );
  NAND4_X1 U15186 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n11959) );
  AOI22_X1 U15187 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12448), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15188 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U15189 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12441), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15190 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n9803), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11954) );
  NAND4_X1 U15191 ( .A1(n11957), .A2(n11956), .A3(n11955), .A4(n11954), .ZN(
        n11958) );
  NAND2_X1 U15192 ( .A1(n12518), .A2(n12725), .ZN(n11961) );
  INV_X1 U15193 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20253) );
  OR2_X1 U15194 ( .A1(n12493), .A2(n20253), .ZN(n11960) );
  XNOR2_X1 U15195 ( .A(n11970), .B(n11971), .ZN(n12715) );
  INV_X1 U15196 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15197 ( .A1(n12635), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20715), .ZN(n11962) );
  OAI21_X1 U15198 ( .B1(n11964), .B2(n11963), .A(n11962), .ZN(n11965) );
  NAND2_X1 U15199 ( .A1(n11965), .A2(n12464), .ZN(n11968) );
  OAI21_X1 U15200 ( .B1(n11966), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11986), .ZN(n20162) );
  NAND2_X1 U15201 ( .A1(n12076), .A2(n20162), .ZN(n11967) );
  NAND2_X1 U15202 ( .A1(n11968), .A2(n11967), .ZN(n11969) );
  AOI21_X1 U15203 ( .B1(n12715), .B2(n12054), .A(n11969), .ZN(n13318) );
  INV_X1 U15204 ( .A(n11970), .ZN(n11972) );
  AOI22_X1 U15205 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15206 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15207 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15208 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11973) );
  NAND4_X1 U15209 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11982) );
  AOI22_X1 U15210 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11980) );
  INV_X1 U15211 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n21062) );
  AOI22_X1 U15212 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15213 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15214 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11977) );
  NAND4_X1 U15215 ( .A1(n11980), .A2(n11979), .A3(n11978), .A4(n11977), .ZN(
        n11981) );
  NAND2_X1 U15216 ( .A1(n12518), .A2(n12735), .ZN(n11985) );
  INV_X1 U15217 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11983) );
  OR2_X1 U15218 ( .A1(n12493), .A2(n11983), .ZN(n11984) );
  NAND2_X1 U15219 ( .A1(n11985), .A2(n11984), .ZN(n11994) );
  XNOR2_X1 U15220 ( .A(n11993), .B(n11994), .ZN(n12723) );
  NAND2_X1 U15221 ( .A1(n12723), .A2(n12054), .ZN(n11992) );
  INV_X1 U15222 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11989) );
  OAI21_X1 U15223 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11987), .A(
        n12008), .ZN(n20066) );
  AOI22_X1 U15224 ( .A1(n12076), .A2(n20066), .B1(n12634), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11988) );
  OAI21_X1 U15225 ( .B1(n12434), .B2(n11989), .A(n11988), .ZN(n11990) );
  INV_X1 U15226 ( .A(n11990), .ZN(n11991) );
  NAND2_X1 U15227 ( .A1(n11992), .A2(n11991), .ZN(n13336) );
  NAND2_X1 U15228 ( .A1(n13316), .A2(n13336), .ZN(n13335) );
  INV_X1 U15229 ( .A(n13335), .ZN(n12015) );
  AOI22_X1 U15230 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15231 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15232 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15233 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11995) );
  NAND4_X1 U15234 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        n12004) );
  AOI22_X1 U15235 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15236 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15237 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15238 ( .A1(n11790), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11999) );
  NAND4_X1 U15239 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n12003) );
  NAND2_X1 U15240 ( .A1(n12518), .A2(n12744), .ZN(n12006) );
  INV_X1 U15241 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20262) );
  OR2_X1 U15242 ( .A1(n12493), .A2(n20262), .ZN(n12005) );
  NAND2_X1 U15243 ( .A1(n12016), .A2(n12017), .ZN(n12733) );
  INV_X1 U15244 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20114) );
  INV_X1 U15245 ( .A(n12022), .ZN(n12011) );
  INV_X1 U15246 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12009) );
  NAND2_X1 U15247 ( .A1(n12009), .A2(n12008), .ZN(n12010) );
  NAND2_X1 U15248 ( .A1(n12011), .A2(n12010), .ZN(n20053) );
  AOI22_X1 U15249 ( .A1(n20053), .A2(n12076), .B1(n12634), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12012) );
  OAI21_X1 U15250 ( .B1(n12434), .B2(n20114), .A(n12012), .ZN(n12013) );
  NAND2_X1 U15251 ( .A1(n12015), .A2(n12014), .ZN(n13398) );
  INV_X1 U15252 ( .A(n13398), .ZN(n12027) );
  INV_X1 U15253 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12020) );
  NAND2_X1 U15254 ( .A1(n12518), .A2(n12746), .ZN(n12019) );
  OAI21_X1 U15255 ( .B1(n12020), .B2(n12493), .A(n12019), .ZN(n12021) );
  INV_X1 U15256 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12024) );
  OAI21_X1 U15257 ( .B1(n12022), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n12042), .ZN(n20041) );
  AOI22_X1 U15258 ( .A1(n20041), .A2(n12076), .B1(n12634), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12023) );
  OAI21_X1 U15259 ( .B1(n12434), .B2(n12024), .A(n12023), .ZN(n12025) );
  AOI21_X1 U15260 ( .B1(n12750), .B2(n12054), .A(n12025), .ZN(n13451) );
  INV_X1 U15261 ( .A(n13451), .ZN(n12026) );
  NAND2_X1 U15262 ( .A1(n12027), .A2(n12026), .ZN(n13448) );
  XNOR2_X1 U15263 ( .A(n12042), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13738) );
  INV_X1 U15264 ( .A(n12634), .ZN(n12102) );
  OAI22_X1 U15265 ( .A1(n13738), .A2(n12464), .B1(n12102), .B2(n13736), .ZN(
        n12028) );
  AOI21_X1 U15266 ( .B1(n12635), .B2(P1_EAX_REG_8__SCAN_IN), .A(n12028), .ZN(
        n12041) );
  AOI22_X1 U15267 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15268 ( .A1(n11790), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15269 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15270 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12029) );
  NAND4_X1 U15271 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n12038) );
  AOI22_X1 U15272 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15273 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U15274 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15275 ( .A1(n12446), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12033) );
  NAND4_X1 U15276 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n12037) );
  NOR2_X1 U15277 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  OR2_X1 U15278 ( .A1(n10207), .A2(n12039), .ZN(n12040) );
  XOR2_X1 U15279 ( .A(n20024), .B(n12057), .Z(n20018) );
  AOI22_X1 U15280 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15281 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15282 ( .A1(n12446), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15283 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12043) );
  NAND4_X1 U15284 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12052) );
  AOI22_X1 U15285 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15286 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15287 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15288 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15289 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12051) );
  OR2_X1 U15290 ( .A1(n12052), .A2(n12051), .ZN(n12053) );
  AOI22_X1 U15291 ( .A1(n12054), .A2(n12053), .B1(n12634), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U15292 ( .A1(n12635), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12055) );
  OAI211_X1 U15293 ( .C1(n20018), .C2(n12464), .A(n12056), .B(n12055), .ZN(
        n13692) );
  XNOR2_X1 U15294 ( .A(n12074), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13719) );
  NAND2_X1 U15295 ( .A1(n13719), .A2(n12076), .ZN(n12073) );
  AOI22_X1 U15296 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15297 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12209), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15298 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15299 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12058) );
  NAND4_X1 U15300 ( .A1(n12061), .A2(n12060), .A3(n12059), .A4(n12058), .ZN(
        n12067) );
  AOI22_X1 U15301 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15302 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15303 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15304 ( .A1(n12448), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12062) );
  NAND4_X1 U15305 ( .A1(n12065), .A2(n12064), .A3(n12063), .A4(n12062), .ZN(
        n12066) );
  NOR2_X1 U15306 ( .A1(n12067), .A2(n12066), .ZN(n12070) );
  NAND2_X1 U15307 ( .A1(n12635), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12069) );
  NAND2_X1 U15308 ( .A1(n12634), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12068) );
  OAI211_X1 U15309 ( .C1(n10207), .C2(n12070), .A(n12069), .B(n12068), .ZN(
        n12071) );
  INV_X1 U15310 ( .A(n12071), .ZN(n12072) );
  NAND2_X1 U15311 ( .A1(n12073), .A2(n12072), .ZN(n13717) );
  INV_X1 U15312 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13775) );
  OAI21_X1 U15313 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12075), .A(
        n12118), .ZN(n16021) );
  AOI22_X1 U15314 ( .A1(n12076), .A2(n16021), .B1(n12634), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12077) );
  OAI21_X1 U15315 ( .B1(n12434), .B2(n13775), .A(n12077), .ZN(n12078) );
  INV_X1 U15316 ( .A(n12078), .ZN(n13770) );
  AOI22_X1 U15317 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15318 ( .A1(n11790), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15319 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15320 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12079) );
  NAND4_X1 U15321 ( .A1(n12082), .A2(n12081), .A3(n12080), .A4(n12079), .ZN(
        n12088) );
  AOI22_X1 U15322 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15323 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15324 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15325 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12083) );
  NAND4_X1 U15326 ( .A1(n12086), .A2(n12085), .A3(n12084), .A4(n12083), .ZN(
        n12087) );
  NOR2_X1 U15327 ( .A1(n12088), .A2(n12087), .ZN(n12089) );
  INV_X1 U15328 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14705) );
  AOI22_X1 U15329 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15330 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11790), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15331 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9803), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15332 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12209), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12091) );
  NAND4_X1 U15333 ( .A1(n12094), .A2(n12093), .A3(n12092), .A4(n12091), .ZN(
        n12100) );
  AOI22_X1 U15334 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12351), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15335 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12376), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15336 ( .A1(n12446), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15337 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15338 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12099) );
  NOR2_X1 U15339 ( .A1(n12100), .A2(n12099), .ZN(n12101) );
  OR2_X1 U15340 ( .A1(n10207), .A2(n12101), .ZN(n12105) );
  XNOR2_X1 U15341 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12118), .ZN(
        n16009) );
  OAI22_X1 U15342 ( .A1(n16009), .A2(n12464), .B1(n12102), .B2(n12117), .ZN(
        n12103) );
  INV_X1 U15343 ( .A(n12103), .ZN(n12104) );
  OAI211_X1 U15344 ( .C1(n14705), .C2(n12434), .A(n12105), .B(n12104), .ZN(
        n14618) );
  INV_X1 U15345 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14702) );
  AOI22_X1 U15346 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11793), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15347 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15348 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15349 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12106) );
  NAND4_X1 U15350 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12115) );
  AOI22_X1 U15351 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15352 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15353 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U15354 ( .A1(n12448), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12110) );
  NAND4_X1 U15355 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12114) );
  NOR2_X1 U15356 ( .A1(n12115), .A2(n12114), .ZN(n12116) );
  OR2_X1 U15357 ( .A1(n10207), .A2(n12116), .ZN(n12121) );
  INV_X1 U15358 ( .A(n12122), .ZN(n12119) );
  XNOR2_X1 U15359 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12119), .ZN(
        n14850) );
  AOI22_X1 U15360 ( .A1(n12076), .A2(n14850), .B1(n12634), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12120) );
  OAI211_X1 U15361 ( .C1(n12434), .C2(n14702), .A(n12121), .B(n12120), .ZN(
        n14523) );
  AOI21_X1 U15362 ( .B1(n21036), .B2(n12123), .A(n12169), .ZN(n16003) );
  OR2_X1 U15363 ( .A1(n16003), .A2(n12464), .ZN(n12139) );
  AOI22_X1 U15364 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15365 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15366 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15367 ( .A1(n12448), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12124) );
  NAND4_X1 U15368 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(
        n12133) );
  AOI22_X1 U15369 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15370 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15371 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15372 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12128) );
  NAND4_X1 U15373 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12132) );
  NOR2_X1 U15374 ( .A1(n12133), .A2(n12132), .ZN(n12136) );
  NAND2_X1 U15375 ( .A1(n12635), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12135) );
  NAND2_X1 U15376 ( .A1(n12634), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12134) );
  OAI211_X1 U15377 ( .C1(n10207), .C2(n12136), .A(n12135), .B(n12134), .ZN(
        n12137) );
  INV_X1 U15378 ( .A(n12137), .ZN(n12138) );
  NAND2_X1 U15379 ( .A1(n12139), .A2(n12138), .ZN(n14610) );
  XNOR2_X1 U15380 ( .A(n12169), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14838) );
  NAND2_X1 U15381 ( .A1(n14838), .A2(n12076), .ZN(n12155) );
  AOI22_X1 U15382 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15383 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15384 ( .A1(n11790), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15385 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12140) );
  NAND4_X1 U15386 ( .A1(n12143), .A2(n12142), .A3(n12141), .A4(n12140), .ZN(
        n12149) );
  AOI22_X1 U15387 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15388 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12209), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15389 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15390 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12144) );
  NAND4_X1 U15391 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12148) );
  NOR2_X1 U15392 ( .A1(n12149), .A2(n12148), .ZN(n12152) );
  NAND2_X1 U15393 ( .A1(n12635), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U15394 ( .A1(n12634), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12150) );
  OAI211_X1 U15395 ( .C1(n10207), .C2(n12152), .A(n12151), .B(n12150), .ZN(
        n12153) );
  INV_X1 U15396 ( .A(n12153), .ZN(n12154) );
  NAND2_X1 U15397 ( .A1(n12155), .A2(n12154), .ZN(n14509) );
  NAND2_X1 U15398 ( .A1(n14506), .A2(n14509), .ZN(n14508) );
  INV_X1 U15399 ( .A(n14508), .ZN(n12174) );
  AOI22_X1 U15400 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11897), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15401 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15402 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15403 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12156) );
  NAND4_X1 U15404 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12165) );
  AOI22_X1 U15405 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15406 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15407 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15408 ( .A1(n12420), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12160) );
  NAND4_X1 U15409 ( .A1(n12163), .A2(n12162), .A3(n12161), .A4(n12160), .ZN(
        n12164) );
  NOR2_X1 U15410 ( .A1(n12165), .A2(n12164), .ZN(n12168) );
  OAI21_X1 U15411 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20847), .A(
        n20715), .ZN(n12167) );
  NAND2_X1 U15412 ( .A1(n12635), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n12166) );
  OAI211_X1 U15413 ( .C1(n12461), .C2(n12168), .A(n12167), .B(n12166), .ZN(
        n12172) );
  OAI21_X1 U15414 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12170), .A(
        n12205), .ZN(n16002) );
  OR2_X1 U15415 ( .A1(n12464), .A2(n16002), .ZN(n12171) );
  NAND2_X1 U15416 ( .A1(n12172), .A2(n12171), .ZN(n14606) );
  NAND2_X1 U15417 ( .A1(n12174), .A2(n12173), .ZN(n14490) );
  AOI22_X1 U15418 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15419 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15420 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15421 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12175) );
  NAND4_X1 U15422 ( .A1(n12178), .A2(n12177), .A3(n12176), .A4(n12175), .ZN(
        n12184) );
  AOI22_X1 U15423 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15424 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15425 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15426 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12179) );
  NAND4_X1 U15427 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12183) );
  OR2_X1 U15428 ( .A1(n12184), .A2(n12183), .ZN(n12188) );
  INV_X1 U15429 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14686) );
  INV_X1 U15430 ( .A(n12205), .ZN(n12185) );
  XNOR2_X1 U15431 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12185), .ZN(
        n14827) );
  AOI22_X1 U15432 ( .A1(n12076), .A2(n14827), .B1(n12634), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12186) );
  OAI21_X1 U15433 ( .B1(n12434), .B2(n14686), .A(n12186), .ZN(n12187) );
  AOI21_X1 U15434 ( .B1(n12431), .B2(n12188), .A(n12187), .ZN(n14494) );
  AOI22_X1 U15435 ( .A1(n12446), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12351), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15436 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15437 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15438 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12190) );
  NAND4_X1 U15439 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n12199) );
  AOI22_X1 U15440 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15441 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15442 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15443 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12194) );
  NAND4_X1 U15444 ( .A1(n12197), .A2(n12196), .A3(n12195), .A4(n12194), .ZN(
        n12198) );
  NOR2_X1 U15445 ( .A1(n12199), .A2(n12198), .ZN(n12204) );
  INV_X1 U15446 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12201) );
  NAND2_X1 U15447 ( .A1(n20715), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12200) );
  OAI211_X1 U15448 ( .C1(n12434), .C2(n12201), .A(n12464), .B(n12200), .ZN(
        n12202) );
  INV_X1 U15449 ( .A(n12202), .ZN(n12203) );
  OAI21_X1 U15450 ( .B1(n12461), .B2(n12204), .A(n12203), .ZN(n12208) );
  OAI21_X1 U15451 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12206), .A(
        n12238), .ZN(n15943) );
  OR2_X1 U15452 ( .A1(n12464), .A2(n15943), .ZN(n12207) );
  NAND2_X1 U15453 ( .A1(n12208), .A2(n12207), .ZN(n14595) );
  AOI22_X1 U15454 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15455 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12209), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15456 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15457 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12210) );
  NAND4_X1 U15458 ( .A1(n12213), .A2(n12212), .A3(n12211), .A4(n12210), .ZN(
        n12219) );
  AOI22_X1 U15459 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15460 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15461 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15462 ( .A1(n12448), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12214) );
  NAND4_X1 U15463 ( .A1(n12217), .A2(n12216), .A3(n12215), .A4(n12214), .ZN(
        n12218) );
  NOR2_X1 U15464 ( .A1(n12219), .A2(n12218), .ZN(n12222) );
  OAI21_X1 U15465 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15934), .A(n12464), 
        .ZN(n12220) );
  AOI21_X1 U15466 ( .B1(n12635), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12220), .ZN(
        n12221) );
  OAI21_X1 U15467 ( .B1(n12461), .B2(n12222), .A(n12221), .ZN(n12224) );
  XNOR2_X1 U15468 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12238), .ZN(
        n15938) );
  NAND2_X1 U15469 ( .A1(n15938), .A2(n12076), .ZN(n12223) );
  AOI22_X1 U15470 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11827), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15471 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15472 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11828), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15473 ( .A1(n11897), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12225) );
  NAND4_X1 U15474 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12234) );
  AOI22_X1 U15475 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15476 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15477 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12376), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15478 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11791), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12229) );
  NAND4_X1 U15479 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12233) );
  NOR2_X1 U15480 ( .A1(n12234), .A2(n12233), .ZN(n12237) );
  OAI21_X1 U15481 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20847), .A(
        n20715), .ZN(n12236) );
  NAND2_X1 U15482 ( .A1(n12635), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n12235) );
  OAI211_X1 U15483 ( .C1(n12461), .C2(n12237), .A(n12236), .B(n12235), .ZN(
        n12245) );
  INV_X1 U15484 ( .A(n12276), .ZN(n12243) );
  INV_X1 U15485 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12241) );
  INV_X1 U15486 ( .A(n12239), .ZN(n12240) );
  NAND2_X1 U15487 ( .A1(n12241), .A2(n12240), .ZN(n12242) );
  NAND2_X1 U15488 ( .A1(n12243), .A2(n12242), .ZN(n15997) );
  AOI22_X1 U15489 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15490 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11793), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15491 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15492 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12209), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12246) );
  NAND4_X1 U15493 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12255) );
  AOI22_X1 U15494 ( .A1(n11897), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15495 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15496 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15497 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12250) );
  NAND4_X1 U15498 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12254) );
  NOR2_X1 U15499 ( .A1(n12255), .A2(n12254), .ZN(n12258) );
  INV_X1 U15500 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14793) );
  AOI21_X1 U15501 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14793), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12256) );
  AOI21_X1 U15502 ( .B1(n12635), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12256), .ZN(
        n12257) );
  OAI21_X1 U15503 ( .B1(n12461), .B2(n12258), .A(n12257), .ZN(n12260) );
  XNOR2_X1 U15504 ( .A(n12276), .B(n14793), .ZN(n14795) );
  NAND2_X1 U15505 ( .A1(n14795), .A2(n12076), .ZN(n12259) );
  AOI22_X1 U15506 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15507 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15508 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15509 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12262) );
  NAND4_X1 U15510 ( .A1(n12265), .A2(n12264), .A3(n12263), .A4(n12262), .ZN(
        n12271) );
  AOI22_X1 U15511 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15512 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11828), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15513 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15514 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12266) );
  NAND4_X1 U15515 ( .A1(n12269), .A2(n12268), .A3(n12267), .A4(n12266), .ZN(
        n12270) );
  NOR2_X1 U15516 ( .A1(n12271), .A2(n12270), .ZN(n12275) );
  INV_X1 U15517 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14666) );
  OAI21_X1 U15518 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20847), .A(
        n20715), .ZN(n12272) );
  OAI21_X1 U15519 ( .B1(n12434), .B2(n14666), .A(n12272), .ZN(n12273) );
  INV_X1 U15520 ( .A(n12273), .ZN(n12274) );
  OAI21_X1 U15521 ( .B1(n12461), .B2(n12275), .A(n12274), .ZN(n12280) );
  AND2_X1 U15522 ( .A1(n12277), .A2(n15916), .ZN(n12278) );
  NOR2_X1 U15523 ( .A1(n12324), .A2(n12278), .ZN(n15918) );
  NAND2_X1 U15524 ( .A1(n15918), .A2(n12076), .ZN(n12279) );
  NAND2_X1 U15525 ( .A1(n12280), .A2(n12279), .ZN(n14568) );
  AOI22_X1 U15526 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15527 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11897), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15528 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15529 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12281) );
  NAND4_X1 U15530 ( .A1(n12284), .A2(n12283), .A3(n12282), .A4(n12281), .ZN(
        n12290) );
  AOI22_X1 U15531 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15532 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15533 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15534 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12285) );
  NAND4_X1 U15535 ( .A1(n12288), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(
        n12289) );
  NOR2_X1 U15536 ( .A1(n12290), .A2(n12289), .ZN(n12310) );
  AOI22_X1 U15537 ( .A1(n11790), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15538 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15539 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15540 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12292) );
  NAND4_X1 U15541 ( .A1(n12295), .A2(n12294), .A3(n12293), .A4(n12292), .ZN(
        n12301) );
  AOI22_X1 U15542 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15543 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15544 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15545 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U15546 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12300) );
  NOR2_X1 U15547 ( .A1(n12301), .A2(n12300), .ZN(n12309) );
  XOR2_X1 U15548 ( .A(n12310), .B(n12309), .Z(n12302) );
  NAND2_X1 U15549 ( .A1(n12302), .A2(n12431), .ZN(n12306) );
  INV_X1 U15550 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14660) );
  NAND2_X1 U15551 ( .A1(n20715), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12303) );
  OAI211_X1 U15552 ( .C1(n12434), .C2(n14660), .A(n12464), .B(n12303), .ZN(
        n12304) );
  INV_X1 U15553 ( .A(n12304), .ZN(n12305) );
  NAND2_X1 U15554 ( .A1(n12306), .A2(n12305), .ZN(n12308) );
  INV_X1 U15555 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14781) );
  XNOR2_X1 U15556 ( .A(n12324), .B(n14781), .ZN(n14779) );
  NAND2_X1 U15557 ( .A1(n14779), .A2(n12076), .ZN(n12307) );
  NAND2_X1 U15558 ( .A1(n12308), .A2(n12307), .ZN(n14466) );
  NOR2_X1 U15559 ( .A1(n12310), .A2(n12309), .ZN(n12332) );
  AOI22_X1 U15560 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15561 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11897), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15562 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15563 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12311) );
  NAND4_X1 U15564 ( .A1(n12314), .A2(n12313), .A3(n12312), .A4(n12311), .ZN(
        n12320) );
  AOI22_X1 U15565 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15566 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11828), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15567 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15568 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12315) );
  NAND4_X1 U15569 ( .A1(n12318), .A2(n12317), .A3(n12316), .A4(n12315), .ZN(
        n12319) );
  INV_X1 U15570 ( .A(n12331), .ZN(n12321) );
  XNOR2_X1 U15571 ( .A(n12332), .B(n12321), .ZN(n12322) );
  NAND2_X1 U15572 ( .A1(n12322), .A2(n12431), .ZN(n12330) );
  OAI21_X1 U15573 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n12325), .A(n12464), 
        .ZN(n12323) );
  AOI21_X1 U15574 ( .B1(n12635), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12323), .ZN(
        n12329) );
  NAND2_X1 U15575 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  NAND2_X1 U15576 ( .A1(n12366), .A2(n12327), .ZN(n15911) );
  NOR2_X1 U15577 ( .A1(n15911), .A2(n12464), .ZN(n12328) );
  AOI21_X1 U15578 ( .B1(n12330), .B2(n12329), .A(n12328), .ZN(n14560) );
  NAND2_X1 U15579 ( .A1(n12332), .A2(n12331), .ZN(n12349) );
  AOI22_X1 U15580 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15581 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12209), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15582 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15583 ( .A1(n11790), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12333) );
  NAND4_X1 U15584 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12342) );
  AOI22_X1 U15585 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12351), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15586 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15587 ( .A1(n11828), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15588 ( .A1(n12448), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12337) );
  NAND4_X1 U15589 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(
        n12341) );
  NOR2_X1 U15590 ( .A1(n12342), .A2(n12341), .ZN(n12350) );
  XOR2_X1 U15591 ( .A(n12349), .B(n12350), .Z(n12343) );
  NAND2_X1 U15592 ( .A1(n12343), .A2(n12431), .ZN(n12348) );
  INV_X1 U15593 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14653) );
  NAND2_X1 U15594 ( .A1(n20715), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12344) );
  OAI211_X1 U15595 ( .C1(n12434), .C2(n14653), .A(n12464), .B(n12344), .ZN(
        n12345) );
  INV_X1 U15596 ( .A(n12345), .ZN(n12347) );
  XNOR2_X1 U15597 ( .A(n12366), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15895) );
  AOI21_X1 U15598 ( .B1(n12348), .B2(n12347), .A(n12346), .ZN(n14553) );
  NAND2_X1 U15599 ( .A1(n14552), .A2(n14553), .ZN(n14450) );
  INV_X1 U15600 ( .A(n14450), .ZN(n12373) );
  NOR2_X1 U15601 ( .A1(n12350), .A2(n12349), .ZN(n12375) );
  AOI22_X1 U15602 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15603 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11897), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15604 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15605 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12352) );
  NAND4_X1 U15606 ( .A1(n12355), .A2(n12354), .A3(n12353), .A4(n12352), .ZN(
        n12361) );
  AOI22_X1 U15607 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15608 ( .A1(n12209), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15609 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12261), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15610 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12356) );
  NAND4_X1 U15611 ( .A1(n12359), .A2(n12358), .A3(n12357), .A4(n12356), .ZN(
        n12360) );
  INV_X1 U15612 ( .A(n12374), .ZN(n12362) );
  XNOR2_X1 U15613 ( .A(n12375), .B(n12362), .ZN(n12365) );
  INV_X1 U15614 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14648) );
  NAND2_X1 U15615 ( .A1(n20715), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12363) );
  OAI211_X1 U15616 ( .C1(n12434), .C2(n14648), .A(n12464), .B(n12363), .ZN(
        n12364) );
  AOI21_X1 U15617 ( .B1(n12365), .B2(n12431), .A(n12364), .ZN(n12371) );
  INV_X1 U15618 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14455) );
  NAND2_X1 U15619 ( .A1(n12368), .A2(n14455), .ZN(n12369) );
  NAND2_X1 U15620 ( .A1(n12411), .A2(n12369), .ZN(n14757) );
  NOR2_X1 U15621 ( .A1(n14757), .A2(n12464), .ZN(n12370) );
  NAND2_X1 U15622 ( .A1(n12375), .A2(n12374), .ZN(n12394) );
  AOI22_X1 U15623 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15624 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12376), .B1(
        n12209), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U15625 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12351), .B1(
        n9803), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15626 ( .A1(n11790), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12377) );
  NAND4_X1 U15627 ( .A1(n12380), .A2(n12379), .A3(n12378), .A4(n12377), .ZN(
        n12386) );
  AOI22_X1 U15628 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12448), .B1(
        n11875), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15629 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15630 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11828), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15631 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12381) );
  NAND4_X1 U15632 ( .A1(n12384), .A2(n12383), .A3(n12382), .A4(n12381), .ZN(
        n12385) );
  NOR2_X1 U15633 ( .A1(n12386), .A2(n12385), .ZN(n12395) );
  XOR2_X1 U15634 ( .A(n12394), .B(n12395), .Z(n12387) );
  NAND2_X1 U15635 ( .A1(n12387), .A2(n12431), .ZN(n12391) );
  INV_X1 U15636 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14642) );
  NAND2_X1 U15637 ( .A1(n20715), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12388) );
  OAI211_X1 U15638 ( .C1(n12434), .C2(n14642), .A(n12464), .B(n12388), .ZN(
        n12389) );
  INV_X1 U15639 ( .A(n12389), .ZN(n12390) );
  NAND2_X1 U15640 ( .A1(n12391), .A2(n12390), .ZN(n12393) );
  XNOR2_X1 U15641 ( .A(n12411), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14747) );
  NAND2_X1 U15642 ( .A1(n14747), .A2(n12076), .ZN(n12392) );
  NAND2_X1 U15643 ( .A1(n12393), .A2(n12392), .ZN(n14439) );
  NOR2_X1 U15644 ( .A1(n12395), .A2(n12394), .ZN(n12419) );
  AOI22_X1 U15645 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15646 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11897), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15647 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15648 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12397) );
  NAND4_X1 U15649 ( .A1(n12400), .A2(n12399), .A3(n12398), .A4(n12397), .ZN(
        n12406) );
  AOI22_X1 U15650 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15651 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11828), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15652 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15653 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12401) );
  NAND4_X1 U15654 ( .A1(n12404), .A2(n12403), .A3(n12402), .A4(n12401), .ZN(
        n12405) );
  OR2_X1 U15655 ( .A1(n12406), .A2(n12405), .ZN(n12418) );
  INV_X1 U15656 ( .A(n12418), .ZN(n12407) );
  XNOR2_X1 U15657 ( .A(n12419), .B(n12407), .ZN(n12408) );
  NAND2_X1 U15658 ( .A1(n12408), .A2(n12431), .ZN(n12417) );
  INV_X1 U15659 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14638) );
  NAND2_X1 U15660 ( .A1(n20715), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12409) );
  OAI211_X1 U15661 ( .C1(n12434), .C2(n14638), .A(n12464), .B(n12409), .ZN(
        n12410) );
  INV_X1 U15662 ( .A(n12410), .ZN(n12416) );
  INV_X1 U15663 ( .A(n12411), .ZN(n12412) );
  NAND2_X1 U15664 ( .A1(n12412), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12413) );
  INV_X1 U15665 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14426) );
  NAND2_X1 U15666 ( .A1(n12413), .A2(n14426), .ZN(n12414) );
  NAND2_X1 U15667 ( .A1(n12439), .A2(n12414), .ZN(n14735) );
  NOR2_X1 U15668 ( .A1(n14735), .A2(n12464), .ZN(n12415) );
  AOI21_X1 U15669 ( .B1(n12417), .B2(n12416), .A(n12415), .ZN(n14422) );
  NAND2_X1 U15670 ( .A1(n12419), .A2(n12418), .ZN(n12455) );
  AOI22_X1 U15671 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U15672 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U15673 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15674 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11792), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12421) );
  NAND4_X1 U15675 ( .A1(n12424), .A2(n12423), .A3(n12422), .A4(n12421), .ZN(
        n12430) );
  AOI22_X1 U15676 ( .A1(n11793), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15677 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15678 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11828), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15679 ( .A1(n11827), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12425) );
  NAND4_X1 U15680 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        n12429) );
  NOR2_X1 U15681 ( .A1(n12430), .A2(n12429), .ZN(n12456) );
  XOR2_X1 U15682 ( .A(n12455), .B(n12456), .Z(n12432) );
  NAND2_X1 U15683 ( .A1(n12432), .A2(n12431), .ZN(n12438) );
  INV_X1 U15684 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14634) );
  NAND2_X1 U15685 ( .A1(n20715), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12433) );
  OAI211_X1 U15686 ( .C1(n12434), .C2(n14634), .A(n12464), .B(n12433), .ZN(
        n12435) );
  INV_X1 U15687 ( .A(n12435), .ZN(n12437) );
  XNOR2_X1 U15688 ( .A(n12439), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14720) );
  AOI21_X1 U15689 ( .B1(n12438), .B2(n12437), .A(n12436), .ZN(n14412) );
  INV_X1 U15690 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14718) );
  XNOR2_X1 U15691 ( .A(n12651), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14714) );
  AOI22_X1 U15692 ( .A1(n11897), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15693 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9804), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15694 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U15695 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12442) );
  NAND4_X1 U15696 ( .A1(n12445), .A2(n12444), .A3(n12443), .A4(n12442), .ZN(
        n12454) );
  AOI22_X1 U15697 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12446), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15698 ( .A1(n12351), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12448), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15699 ( .A1(n12376), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12291), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15700 ( .A1(n9803), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12420), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12449) );
  NAND4_X1 U15701 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        n12453) );
  NOR2_X1 U15702 ( .A1(n12454), .A2(n12453), .ZN(n12458) );
  NOR2_X1 U15703 ( .A1(n12456), .A2(n12455), .ZN(n12457) );
  XOR2_X1 U15704 ( .A(n12458), .B(n12457), .Z(n12462) );
  AOI21_X1 U15705 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20715), .A(
        n12076), .ZN(n12460) );
  NAND2_X1 U15706 ( .A1(n12635), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12459) );
  OAI211_X1 U15707 ( .C1(n12462), .C2(n12461), .A(n12460), .B(n12459), .ZN(
        n12463) );
  OAI21_X1 U15708 ( .B1(n12464), .B2(n14714), .A(n12463), .ZN(n12466) );
  INV_X1 U15709 ( .A(n14716), .ZN(n12633) );
  XNOR2_X1 U15710 ( .A(n13079), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12469) );
  NAND2_X1 U15711 ( .A1(n20863), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12473) );
  OAI22_X1 U15712 ( .A1(n12469), .A2(n12473), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n13079), .ZN(n12488) );
  MUX2_X1 U15713 ( .A(n11859), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12489) );
  NAND2_X1 U15714 ( .A1(n12488), .A2(n12489), .ZN(n12490) );
  NAND2_X1 U15715 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11859), .ZN(
        n12467) );
  NAND2_X1 U15716 ( .A1(n12490), .A2(n12467), .ZN(n12503) );
  MUX2_X1 U15717 ( .A(n20574), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n15019), .Z(n12504) );
  NOR2_X1 U15718 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20234), .ZN(
        n12468) );
  INV_X1 U15719 ( .A(n12518), .ZN(n12494) );
  NAND2_X1 U15720 ( .A1(n20254), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12480) );
  XNOR2_X1 U15721 ( .A(n12469), .B(n12473), .ZN(n12640) );
  NAND2_X1 U15722 ( .A1(n12514), .A2(n12640), .ZN(n12470) );
  OAI211_X1 U15723 ( .C1(n12494), .C2(n20238), .A(n12480), .B(n12470), .ZN(
        n12483) );
  INV_X1 U15724 ( .A(n12483), .ZN(n12487) );
  NAND2_X1 U15725 ( .A1(n20254), .A2(n13794), .ZN(n12471) );
  NAND2_X1 U15726 ( .A1(n12471), .A2(n20238), .ZN(n12495) );
  NAND2_X1 U15727 ( .A1(n13030), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12472) );
  AND2_X1 U15728 ( .A1(n12473), .A2(n12472), .ZN(n12477) );
  INV_X1 U15729 ( .A(n12477), .ZN(n12476) );
  OAI211_X1 U15730 ( .C1(n20249), .C2(n12476), .A(n12474), .B(n12475), .ZN(
        n12479) );
  AOI21_X1 U15731 ( .B1(n12477), .B2(n12518), .A(n12519), .ZN(n12478) );
  AOI21_X1 U15732 ( .B1(n12495), .B2(n12479), .A(n12478), .ZN(n12484) );
  INV_X1 U15733 ( .A(n12484), .ZN(n12486) );
  NAND2_X1 U15734 ( .A1(n12480), .A2(n11758), .ZN(n12481) );
  NOR2_X1 U15735 ( .A1(n12518), .A2(n12481), .ZN(n12510) );
  INV_X1 U15736 ( .A(n12640), .ZN(n12482) );
  AOI211_X1 U15737 ( .C1(n12484), .C2(n12483), .A(n12510), .B(n12482), .ZN(
        n12485) );
  OR2_X1 U15738 ( .A1(n12489), .A2(n12488), .ZN(n12491) );
  NAND2_X1 U15739 ( .A1(n12491), .A2(n12490), .ZN(n12641) );
  INV_X1 U15740 ( .A(n12641), .ZN(n12492) );
  OAI21_X1 U15741 ( .B1(n12493), .B2(n12492), .A(n12495), .ZN(n12498) );
  INV_X1 U15742 ( .A(n12499), .ZN(n12496) );
  AOI211_X1 U15743 ( .C1(n12496), .C2(n12495), .A(n12494), .B(n12641), .ZN(
        n12497) );
  AOI21_X1 U15744 ( .B1(n12499), .B2(n12498), .A(n12497), .ZN(n12512) );
  INV_X1 U15745 ( .A(n12512), .ZN(n12500) );
  AOI22_X1 U15746 ( .A1(n12500), .A2(n12514), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n16155), .ZN(n12516) );
  NAND3_X1 U15747 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12501), .A3(
        n11963), .ZN(n12643) );
  INV_X1 U15748 ( .A(n12502), .ZN(n12508) );
  INV_X1 U15749 ( .A(n12503), .ZN(n12506) );
  INV_X1 U15750 ( .A(n12504), .ZN(n12505) );
  NAND2_X1 U15751 ( .A1(n12506), .A2(n12505), .ZN(n12507) );
  NAND2_X1 U15752 ( .A1(n12508), .A2(n12507), .ZN(n12639) );
  INV_X1 U15753 ( .A(n12643), .ZN(n12509) );
  AOI22_X1 U15754 ( .A1(n12510), .A2(n12509), .B1(n12519), .B2(n12639), .ZN(
        n12511) );
  OAI21_X1 U15755 ( .B1(n12512), .B2(n12639), .A(n12511), .ZN(n12513) );
  OAI21_X1 U15756 ( .B1(n12514), .B2(n12643), .A(n12513), .ZN(n12515) );
  NAND2_X1 U15757 ( .A1(n12516), .A2(n12515), .ZN(n12517) );
  AND2_X1 U15758 ( .A1(n12642), .A2(n12519), .ZN(n12520) );
  OR2_X1 U15759 ( .A1(n12523), .A2(n20238), .ZN(n12999) );
  NAND2_X1 U15760 ( .A1(n15862), .A2(n14385), .ZN(n13029) );
  INV_X1 U15761 ( .A(n12474), .ZN(n12526) );
  NAND4_X1 U15762 ( .A1(n12526), .A2(n20264), .A3(n12998), .A4(n12525), .ZN(
        n12795) );
  OR2_X1 U15763 ( .A1(n12795), .A2(n14394), .ZN(n12527) );
  OR2_X2 U15764 ( .A1(n14612), .A2(n20264), .ZN(n14627) );
  AOI22_X1 U15765 ( .A1(n13179), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14394), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12656) );
  INV_X1 U15766 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13094) );
  BUF_X1 U15767 ( .A(n12551), .Z(n12568) );
  INV_X1 U15768 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20219) );
  NAND2_X1 U15769 ( .A1(n12568), .A2(n20219), .ZN(n12531) );
  NAND2_X1 U15770 ( .A1(n12568), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12532) );
  OAI21_X1 U15771 ( .B1(n12529), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12532), .ZN(
        n13181) );
  INV_X1 U15772 ( .A(n12533), .ZN(n12534) );
  AOI21_X1 U15773 ( .B1(n13666), .B2(n12659), .A(n12534), .ZN(n13171) );
  MUX2_X1 U15774 ( .A(n12623), .B(n12568), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12537) );
  NAND2_X1 U15775 ( .A1(n14394), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12535) );
  AND2_X1 U15776 ( .A1(n12535), .A2(n12590), .ZN(n12536) );
  NAND2_X1 U15777 ( .A1(n12537), .A2(n12536), .ZN(n13170) );
  INV_X1 U15778 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13684) );
  NAND2_X1 U15779 ( .A1(n12615), .A2(n13684), .ZN(n12540) );
  INV_X1 U15780 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12706) );
  NAND2_X1 U15781 ( .A1(n12659), .A2(n13684), .ZN(n12538) );
  OAI211_X1 U15782 ( .C1(n12529), .C2(n12706), .A(n12538), .B(n12568), .ZN(
        n12539) );
  AND2_X1 U15783 ( .A1(n12540), .A2(n12539), .ZN(n13283) );
  INV_X1 U15784 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n12541) );
  NAND2_X1 U15785 ( .A1(n12603), .A2(n12541), .ZN(n12545) );
  INV_X1 U15786 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12720) );
  NAND2_X1 U15787 ( .A1(n12568), .A2(n12720), .ZN(n12543) );
  NAND2_X1 U15788 ( .A1(n12659), .A2(n12541), .ZN(n12542) );
  NAND3_X1 U15789 ( .A1(n12543), .A2(n12655), .A3(n12542), .ZN(n12544) );
  AND2_X1 U15790 ( .A1(n12545), .A2(n12544), .ZN(n13319) );
  MUX2_X1 U15791 ( .A(n12621), .B(n12655), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12547) );
  OAI21_X1 U15792 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n13179), .A(
        n12547), .ZN(n13339) );
  INV_X1 U15793 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20033) );
  NAND2_X1 U15794 ( .A1(n12615), .A2(n20033), .ZN(n12550) );
  INV_X1 U15795 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U15796 ( .A1(n12659), .A2(n20033), .ZN(n12548) );
  OAI211_X1 U15797 ( .C1(n12529), .C2(n12751), .A(n12548), .B(n12568), .ZN(
        n12549) );
  AND2_X1 U15798 ( .A1(n12550), .A2(n12549), .ZN(n13452) );
  INV_X1 U15799 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20042) );
  NAND2_X1 U15800 ( .A1(n12603), .A2(n20042), .ZN(n12555) );
  INV_X1 U15801 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16028) );
  NAND2_X1 U15802 ( .A1(n12568), .A2(n16028), .ZN(n12553) );
  NAND2_X1 U15803 ( .A1(n12659), .A2(n20042), .ZN(n12552) );
  NAND3_X1 U15804 ( .A1(n12553), .A2(n12655), .A3(n12552), .ZN(n12554) );
  NAND2_X1 U15805 ( .A1(n12555), .A2(n12554), .ZN(n13453) );
  MUX2_X1 U15806 ( .A(n12623), .B(n12568), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12558) );
  NAND2_X1 U15807 ( .A1(n14394), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12556) );
  AND2_X1 U15808 ( .A1(n12590), .A2(n12556), .ZN(n12557) );
  NAND2_X1 U15809 ( .A1(n12558), .A2(n12557), .ZN(n13694) );
  INV_X1 U15810 ( .A(n13694), .ZN(n12561) );
  MUX2_X1 U15811 ( .A(n12621), .B(n12655), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12560) );
  OR2_X1 U15812 ( .A1(n13179), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12559) );
  NAND2_X1 U15813 ( .A1(n12560), .A2(n12559), .ZN(n13696) );
  NOR2_X1 U15814 ( .A1(n12561), .A2(n13696), .ZN(n12562) );
  NAND2_X1 U15815 ( .A1(n13695), .A2(n12562), .ZN(n13721) );
  MUX2_X1 U15816 ( .A(n12623), .B(n12568), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12564) );
  NAND2_X1 U15817 ( .A1(n14394), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12563) );
  OR2_X1 U15818 ( .A1(n12621), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n12567) );
  INV_X1 U15819 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16089) );
  INV_X1 U15820 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21107) );
  NAND2_X1 U15821 ( .A1(n12659), .A2(n21107), .ZN(n12565) );
  OAI211_X1 U15822 ( .C1(n12529), .C2(n16089), .A(n12565), .B(n12568), .ZN(
        n12566) );
  NAND2_X1 U15823 ( .A1(n12567), .A2(n12566), .ZN(n13773) );
  MUX2_X1 U15824 ( .A(n12623), .B(n12568), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12571) );
  NAND2_X1 U15825 ( .A1(n14394), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12569) );
  AND2_X1 U15826 ( .A1(n12590), .A2(n12569), .ZN(n12570) );
  NAND2_X1 U15827 ( .A1(n12571), .A2(n12570), .ZN(n14622) );
  MUX2_X1 U15828 ( .A(n12621), .B(n12655), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12573) );
  OR2_X1 U15829 ( .A1(n13179), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12572) );
  INV_X1 U15830 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15960) );
  NAND2_X1 U15831 ( .A1(n12603), .A2(n15960), .ZN(n12577) );
  INV_X1 U15832 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21132) );
  NAND2_X1 U15833 ( .A1(n12568), .A2(n21132), .ZN(n12575) );
  NAND2_X1 U15834 ( .A1(n12659), .A2(n15960), .ZN(n12574) );
  NAND3_X1 U15835 ( .A1(n12575), .A2(n12655), .A3(n12574), .ZN(n12576) );
  OR2_X1 U15836 ( .A1(n12621), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n12581) );
  INV_X1 U15837 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14990) );
  INV_X1 U15838 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n12578) );
  NAND2_X1 U15839 ( .A1(n12659), .A2(n12578), .ZN(n12579) );
  OAI211_X1 U15840 ( .C1(n12529), .C2(n14990), .A(n12579), .B(n12568), .ZN(
        n12580) );
  NAND2_X1 U15841 ( .A1(n12581), .A2(n12580), .ZN(n14511) );
  MUX2_X1 U15842 ( .A(n12623), .B(n12568), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12584) );
  NAND2_X1 U15843 ( .A1(n14394), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12582) );
  AND2_X1 U15844 ( .A1(n12590), .A2(n12582), .ZN(n12583) );
  INV_X1 U15845 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U15846 ( .A1(n12615), .A2(n12585), .ZN(n12589) );
  INV_X1 U15847 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12587) );
  NAND2_X1 U15848 ( .A1(n12659), .A2(n12585), .ZN(n12586) );
  OAI211_X1 U15849 ( .C1(n12529), .C2(n12587), .A(n12586), .B(n12568), .ZN(
        n12588) );
  AND2_X1 U15850 ( .A1(n12589), .A2(n12588), .ZN(n14498) );
  NAND2_X1 U15851 ( .A1(n14604), .A2(n14498), .ZN(n14598) );
  MUX2_X1 U15852 ( .A(n12623), .B(n12568), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12593) );
  INV_X1 U15853 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16055) );
  OAI21_X1 U15854 ( .B1(n12659), .B2(n16055), .A(n12590), .ZN(n12591) );
  INV_X1 U15855 ( .A(n12591), .ZN(n12592) );
  OR2_X1 U15856 ( .A1(n12621), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n12596) );
  INV_X1 U15857 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16045) );
  INV_X1 U15858 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14592) );
  NAND2_X1 U15859 ( .A1(n12659), .A2(n14592), .ZN(n12594) );
  OAI211_X1 U15860 ( .C1(n12529), .C2(n16045), .A(n12594), .B(n12568), .ZN(
        n12595) );
  NAND2_X1 U15861 ( .A1(n12596), .A2(n12595), .ZN(n14589) );
  INV_X1 U15862 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14970) );
  NAND2_X1 U15863 ( .A1(n12568), .A2(n14970), .ZN(n12598) );
  INV_X1 U15864 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15925) );
  NAND2_X1 U15865 ( .A1(n12659), .A2(n15925), .ZN(n12597) );
  NAND3_X1 U15866 ( .A1(n12598), .A2(n12655), .A3(n12597), .ZN(n12599) );
  OAI21_X1 U15867 ( .B1(n12623), .B2(P1_EBX_REG_20__SCAN_IN), .A(n12599), .ZN(
        n14580) );
  MUX2_X1 U15868 ( .A(n12621), .B(n12655), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12601) );
  OR2_X1 U15869 ( .A1(n13179), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12600) );
  NAND2_X1 U15870 ( .A1(n12601), .A2(n12600), .ZN(n14487) );
  INV_X1 U15871 ( .A(n14487), .ZN(n12602) );
  INV_X1 U15872 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14573) );
  NAND2_X1 U15873 ( .A1(n12603), .A2(n14573), .ZN(n12607) );
  INV_X1 U15874 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14952) );
  NAND2_X1 U15875 ( .A1(n12568), .A2(n14952), .ZN(n12605) );
  NAND2_X1 U15876 ( .A1(n12659), .A2(n14573), .ZN(n12604) );
  NAND3_X1 U15877 ( .A1(n12605), .A2(n12655), .A3(n12604), .ZN(n12606) );
  OR2_X1 U15878 ( .A1(n12621), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n12610) );
  INV_X1 U15879 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14931) );
  INV_X1 U15880 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21069) );
  NAND2_X1 U15881 ( .A1(n12659), .A2(n21069), .ZN(n12608) );
  OAI211_X1 U15882 ( .C1(n12529), .C2(n14931), .A(n12608), .B(n12568), .ZN(
        n12609) );
  NAND2_X1 U15883 ( .A1(n12610), .A2(n12609), .ZN(n14467) );
  INV_X1 U15884 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14930) );
  NAND2_X1 U15885 ( .A1(n12568), .A2(n14930), .ZN(n12613) );
  INV_X1 U15886 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n12611) );
  NAND2_X1 U15887 ( .A1(n12659), .A2(n12611), .ZN(n12612) );
  NAND3_X1 U15888 ( .A1(n12613), .A2(n12655), .A3(n12612), .ZN(n12614) );
  OAI21_X1 U15889 ( .B1(n12623), .B2(P1_EBX_REG_24__SCAN_IN), .A(n12614), .ZN(
        n14564) );
  INV_X1 U15890 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14557) );
  NAND2_X1 U15891 ( .A1(n12615), .A2(n14557), .ZN(n12618) );
  INV_X1 U15892 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14727) );
  NAND2_X1 U15893 ( .A1(n12659), .A2(n14557), .ZN(n12616) );
  OAI211_X1 U15894 ( .C1(n12529), .C2(n14727), .A(n12616), .B(n12568), .ZN(
        n12617) );
  MUX2_X1 U15895 ( .A(n12623), .B(n12568), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12620) );
  NAND2_X1 U15896 ( .A1(n14394), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12619) );
  MUX2_X1 U15897 ( .A(n12621), .B(n12655), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12622) );
  OAI21_X1 U15898 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13179), .A(
        n12622), .ZN(n14435) );
  MUX2_X1 U15899 ( .A(n12623), .B(n12568), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12625) );
  NAND2_X1 U15900 ( .A1(n14394), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12624) );
  NAND2_X1 U15901 ( .A1(n12625), .A2(n12624), .ZN(n14419) );
  OR2_X1 U15902 ( .A1(n13179), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12626) );
  INV_X1 U15903 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14547) );
  NAND2_X1 U15904 ( .A1(n12659), .A2(n14547), .ZN(n12627) );
  NAND2_X1 U15905 ( .A1(n12626), .A2(n12627), .ZN(n12628) );
  MUX2_X1 U15906 ( .A(n12628), .B(n12627), .S(n12529), .Z(n14408) );
  INV_X1 U15907 ( .A(n14410), .ZN(n12629) );
  OAI22_X1 U15908 ( .A1(n12629), .A2(n12655), .B1(n14421), .B2(n12628), .ZN(
        n12630) );
  XOR2_X1 U15909 ( .A(n12656), .B(n12630), .Z(n14867) );
  INV_X1 U15910 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14400) );
  INV_X1 U15911 ( .A(n12631), .ZN(n12632) );
  AOI22_X1 U15912 ( .A1(n12635), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12634), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12636) );
  INV_X1 U15913 ( .A(n12638), .ZN(n14391) );
  NOR3_X1 U15914 ( .A1(n12641), .A2(n12640), .A3(n12639), .ZN(n12644) );
  AOI21_X1 U15915 ( .B1(n12644), .B2(n12643), .A(n12642), .ZN(n14392) );
  AND2_X1 U15916 ( .A1(n12645), .A2(n14397), .ZN(n12646) );
  NAND2_X1 U15917 ( .A1(n14392), .A2(n12646), .ZN(n12870) );
  OR2_X2 U15918 ( .A1(n12680), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20208) );
  AND2_X1 U15919 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n16155), .ZN(n12648) );
  NAND3_X1 U15920 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20715), .A3(n16162), 
        .ZN(n15861) );
  INV_X1 U15921 ( .A(n15861), .ZN(n12647) );
  AOI22_X1 U15922 ( .A1(n12076), .A2(n12648), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n12647), .ZN(n12649) );
  NAND2_X1 U15923 ( .A1(n20208), .A2(n12649), .ZN(n12650) );
  INV_X1 U15924 ( .A(n12651), .ZN(n12652) );
  INV_X1 U15925 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14401) );
  AOI22_X1 U15926 ( .A1(n13179), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14394), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12657) );
  NAND2_X1 U15927 ( .A1(n12659), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12667) );
  AND2_X1 U15928 ( .A1(n20880), .A2(n20847), .ZN(n15855) );
  NOR2_X1 U15929 ( .A1(n12667), .A2(n15855), .ZN(n12660) );
  OR2_X1 U15930 ( .A1(n12661), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15880) );
  INV_X1 U15931 ( .A(n15880), .ZN(n15856) );
  OR2_X1 U15932 ( .A1(n11758), .A2(n15856), .ZN(n13785) );
  NAND2_X1 U15933 ( .A1(n13785), .A2(n15855), .ZN(n12666) );
  NOR2_X1 U15934 ( .A1(n12666), .A2(n11765), .ZN(n12662) );
  NAND2_X1 U15935 ( .A1(n20080), .A2(n20079), .ZN(n20031) );
  NAND2_X1 U15936 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n12672) );
  INV_X1 U15937 ( .A(n12672), .ZN(n12665) );
  INV_X1 U15938 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20822) );
  NAND4_X1 U15939 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .A3(P1_REIP_REG_19__SCAN_IN), .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n15913) );
  NAND4_X1 U15940 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(P1_REIP_REG_8__SCAN_IN), .A4(P1_REIP_REG_7__SCAN_IN), .ZN(n13493)
         );
  NAND3_X1 U15941 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14481) );
  INV_X1 U15942 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n13809) );
  NAND2_X1 U15943 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14525) );
  NAND3_X1 U15944 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n15958) );
  NOR3_X1 U15945 ( .A1(n13809), .A2(n14525), .A3(n15958), .ZN(n14495) );
  AND4_X1 U15946 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20054)
         );
  NAND3_X1 U15947 ( .A1(n14495), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n20054), 
        .ZN(n12663) );
  NOR4_X1 U15948 ( .A1(n15913), .A2(n13493), .A3(n14481), .A4(n12663), .ZN(
        n14470) );
  NAND2_X1 U15949 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14470), .ZN(n14464) );
  NOR2_X1 U15950 ( .A1(n20822), .A2(n14464), .ZN(n15897) );
  AND2_X1 U15951 ( .A1(n15897), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14454) );
  AND2_X1 U15952 ( .A1(n14454), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14427) );
  AND2_X1 U15953 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n12671) );
  NAND3_X1 U15954 ( .A1(n20079), .A2(n14427), .A3(n12671), .ZN(n12664) );
  NAND2_X1 U15955 ( .A1(n20031), .A2(n12664), .ZN(n14428) );
  OAI21_X1 U15956 ( .B1(n20062), .B2(n12665), .A(n14428), .ZN(n14404) );
  INV_X1 U15957 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n12670) );
  AND3_X1 U15958 ( .A1(n12667), .A2(n12666), .A3(n13794), .ZN(n12668) );
  INV_X1 U15959 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12669) );
  OAI22_X1 U15960 ( .A1(n12670), .A2(n20043), .B1(n20025), .B2(n12669), .ZN(
        n12674) );
  INV_X1 U15961 ( .A(n14427), .ZN(n14440) );
  NOR2_X1 U15962 ( .A1(n20080), .A2(n14440), .ZN(n14441) );
  NAND2_X1 U15963 ( .A1(n14441), .A2(n12671), .ZN(n14415) );
  NOR3_X1 U15964 ( .A1(n14415), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n12672), 
        .ZN(n12673) );
  AOI211_X1 U15965 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14404), .A(n12674), 
        .B(n12673), .ZN(n12675) );
  INV_X1 U15966 ( .A(n12676), .ZN(n12677) );
  NAND2_X1 U15967 ( .A1(n12678), .A2(n12677), .ZN(P1_U2809) );
  AND3_X1 U15968 ( .A1(n16155), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16156) );
  AOI21_X1 U15969 ( .B1(n13015), .B2(n11765), .A(n12679), .ZN(n12791) );
  AND2_X1 U15970 ( .A1(n12791), .A2(n13002), .ZN(n13022) );
  NAND2_X1 U15971 ( .A1(n20859), .A2(n12680), .ZN(n20879) );
  NAND2_X1 U15972 ( .A1(n20879), .A2(n16155), .ZN(n12681) );
  NAND2_X1 U15973 ( .A1(n16155), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20777) );
  NAND2_X1 U15974 ( .A1(n20847), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12682) );
  AND2_X1 U15975 ( .A1(n20777), .A2(n12682), .ZN(n13084) );
  INV_X1 U15976 ( .A(n13084), .ZN(n12683) );
  INV_X1 U15977 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20837) );
  NOR2_X1 U15978 ( .A1(n20208), .A2(n20837), .ZN(n13957) );
  AOI21_X1 U15979 ( .B1(n20165), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13957), .ZN(n12684) );
  OAI21_X1 U15980 ( .B1(n20163), .B2(n13498), .A(n12684), .ZN(n12685) );
  AOI21_X1 U15981 ( .B1(n12800), .B2(n20159), .A(n12685), .ZN(n12789) );
  NAND2_X1 U15982 ( .A1(n12686), .A2(n12691), .ZN(n12708) );
  OAI21_X1 U15983 ( .B1(n12691), .B2(n12686), .A(n12708), .ZN(n12688) );
  NAND2_X1 U15984 ( .A1(n11765), .A2(n12690), .ZN(n12699) );
  OAI21_X1 U15985 ( .B1(n20874), .B2(n12691), .A(n12699), .ZN(n12692) );
  INV_X1 U15986 ( .A(n12692), .ZN(n12693) );
  NAND2_X2 U15987 ( .A1(n13086), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13085) );
  INV_X1 U15988 ( .A(n12695), .ZN(n12696) );
  INV_X1 U15989 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20204) );
  INV_X1 U15990 ( .A(n12754), .ZN(n12749) );
  NAND2_X1 U15991 ( .A1(n12698), .A2(n12749), .ZN(n12703) );
  XNOR2_X1 U15992 ( .A(n12708), .B(n12707), .ZN(n12701) );
  INV_X1 U15993 ( .A(n20874), .ZN(n15857) );
  INV_X1 U15994 ( .A(n12699), .ZN(n12700) );
  AOI21_X1 U15995 ( .B1(n12701), .B2(n15857), .A(n12700), .ZN(n12702) );
  NAND2_X1 U15996 ( .A1(n12703), .A2(n12702), .ZN(n13133) );
  NAND2_X1 U15997 ( .A1(n13134), .A2(n13133), .ZN(n20197) );
  NAND2_X1 U15998 ( .A1(n12704), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12705) );
  NAND2_X1 U15999 ( .A1(n12708), .A2(n12707), .ZN(n12727) );
  INV_X1 U16000 ( .A(n12724), .ZN(n12709) );
  XNOR2_X1 U16001 ( .A(n12727), .B(n12709), .ZN(n12710) );
  NAND2_X1 U16002 ( .A1(n12710), .A2(n15857), .ZN(n12711) );
  NAND2_X1 U16003 ( .A1(n12712), .A2(n12711), .ZN(n13288) );
  NAND2_X1 U16004 ( .A1(n12713), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12714) );
  NAND2_X1 U16005 ( .A1(n12715), .A2(n12749), .ZN(n12719) );
  NAND2_X1 U16006 ( .A1(n12727), .A2(n12724), .ZN(n12716) );
  XNOR2_X1 U16007 ( .A(n12716), .B(n12725), .ZN(n12717) );
  NAND2_X1 U16008 ( .A1(n12717), .A2(n15857), .ZN(n12718) );
  NAND2_X1 U16009 ( .A1(n12719), .A2(n12718), .ZN(n12721) );
  XNOR2_X1 U16010 ( .A(n12721), .B(n12720), .ZN(n20155) );
  NAND2_X1 U16011 ( .A1(n12721), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12722) );
  NAND2_X1 U16012 ( .A1(n12723), .A2(n12749), .ZN(n12730) );
  AND2_X1 U16013 ( .A1(n12725), .A2(n12724), .ZN(n12726) );
  NAND2_X1 U16014 ( .A1(n12727), .A2(n12726), .ZN(n12734) );
  XNOR2_X1 U16015 ( .A(n12734), .B(n12735), .ZN(n12728) );
  NAND2_X1 U16016 ( .A1(n12728), .A2(n15857), .ZN(n12729) );
  NAND2_X1 U16017 ( .A1(n12730), .A2(n12729), .ZN(n12731) );
  INV_X1 U16018 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13801) );
  XNOR2_X1 U16019 ( .A(n12731), .B(n13801), .ZN(n16035) );
  NAND2_X1 U16020 ( .A1(n12731), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12732) );
  NAND3_X1 U16021 ( .A1(n12757), .A2(n12749), .A3(n12733), .ZN(n12739) );
  INV_X1 U16022 ( .A(n12734), .ZN(n12736) );
  NAND2_X1 U16023 ( .A1(n12736), .A2(n12735), .ZN(n12743) );
  XNOR2_X1 U16024 ( .A(n12743), .B(n12744), .ZN(n12737) );
  NAND2_X1 U16025 ( .A1(n12737), .A2(n15857), .ZN(n12738) );
  NAND2_X1 U16026 ( .A1(n16029), .A2(n16028), .ZN(n12740) );
  INV_X1 U16027 ( .A(n16029), .ZN(n12741) );
  NAND2_X1 U16028 ( .A1(n12741), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12742) );
  INV_X1 U16029 ( .A(n12743), .ZN(n12745) );
  NAND2_X1 U16030 ( .A1(n12745), .A2(n12744), .ZN(n12759) );
  XNOR2_X1 U16031 ( .A(n12759), .B(n12746), .ZN(n12747) );
  AND2_X1 U16032 ( .A1(n12747), .A2(n15857), .ZN(n12748) );
  AOI21_X1 U16033 ( .B1(n12750), .B2(n12749), .A(n12748), .ZN(n12752) );
  NAND2_X1 U16034 ( .A1(n12752), .A2(n12751), .ZN(n16023) );
  INV_X1 U16035 ( .A(n12752), .ZN(n12753) );
  NAND2_X1 U16036 ( .A1(n12753), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16022) );
  NOR3_X1 U16037 ( .A1(n12755), .A2(n12754), .A3(n12758), .ZN(n12756) );
  OR3_X1 U16038 ( .A1(n12759), .A2(n12758), .A3(n20874), .ZN(n12760) );
  INV_X1 U16039 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13731) );
  NAND2_X1 U16040 ( .A1(n13732), .A2(n13731), .ZN(n12761) );
  NAND2_X1 U16041 ( .A1(n13734), .A2(n12761), .ZN(n12764) );
  INV_X1 U16042 ( .A(n13732), .ZN(n12762) );
  NAND2_X1 U16043 ( .A1(n12762), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12763) );
  INV_X1 U16044 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13764) );
  NAND2_X1 U16045 ( .A1(n16013), .A2(n13764), .ZN(n12765) );
  INV_X1 U16046 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14992) );
  NAND2_X1 U16047 ( .A1(n9810), .A2(n14992), .ZN(n14823) );
  NAND2_X1 U16048 ( .A1(n12766), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12767) );
  NAND2_X1 U16049 ( .A1(n14823), .A2(n12767), .ZN(n14985) );
  OAI21_X1 U16050 ( .B1(n14858), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n14988), .ZN(n12768) );
  NAND2_X1 U16051 ( .A1(n9810), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13813) );
  INV_X1 U16052 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16081) );
  NAND2_X1 U16053 ( .A1(n12766), .A2(n16081), .ZN(n12769) );
  NAND2_X1 U16054 ( .A1(n13813), .A2(n12769), .ZN(n14848) );
  INV_X1 U16055 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12770) );
  NAND2_X1 U16056 ( .A1(n12766), .A2(n12770), .ZN(n15003) );
  NAND2_X1 U16057 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12771) );
  NAND2_X1 U16058 ( .A1(n12766), .A2(n12771), .ZN(n14845) );
  NAND2_X1 U16059 ( .A1(n15003), .A2(n14845), .ZN(n12772) );
  NOR2_X1 U16060 ( .A1(n14848), .A2(n12772), .ZN(n13812) );
  NAND2_X1 U16061 ( .A1(n16013), .A2(n21132), .ZN(n12773) );
  NAND2_X1 U16062 ( .A1(n13812), .A2(n12773), .ZN(n14820) );
  NAND2_X1 U16063 ( .A1(n14858), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14846) );
  INV_X1 U16064 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16102) );
  NAND2_X1 U16065 ( .A1(n16102), .A2(n16089), .ZN(n12774) );
  NAND2_X1 U16066 ( .A1(n14858), .A2(n12774), .ZN(n14843) );
  AND2_X1 U16067 ( .A1(n14846), .A2(n14843), .ZN(n13811) );
  NAND2_X1 U16068 ( .A1(n14858), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12775) );
  OAI21_X1 U16069 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n14858), .ZN(n12776) );
  NAND2_X1 U16070 ( .A1(n14858), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14822) );
  XNOR2_X1 U16071 ( .A(n16013), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14814) );
  NAND2_X1 U16072 ( .A1(n14815), .A2(n14814), .ZN(n14807) );
  INV_X1 U16073 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14953) );
  INV_X1 U16074 ( .A(n12777), .ZN(n14786) );
  NAND2_X1 U16075 ( .A1(n16055), .A2(n16045), .ZN(n14798) );
  OR4_X2 U16076 ( .A1(n14815), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A4(n14798), .ZN(n12778) );
  NAND2_X2 U16077 ( .A1(n12780), .A2(n14785), .ZN(n14726) );
  OR2_X2 U16078 ( .A1(n14726), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14761) );
  NAND2_X1 U16079 ( .A1(n14727), .A2(n14930), .ZN(n12779) );
  AND2_X1 U16081 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14928) );
  NAND2_X1 U16082 ( .A1(n14928), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14750) );
  NAND2_X1 U16083 ( .A1(n14726), .A2(n14750), .ZN(n12781) );
  NAND2_X1 U16084 ( .A1(n12780), .A2(n16013), .ZN(n14762) );
  AND2_X1 U16085 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14888) );
  INV_X1 U16086 ( .A(n14721), .ZN(n12783) );
  INV_X1 U16087 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14877) );
  NOR2_X1 U16088 ( .A1(n14858), .A2(n14877), .ZN(n12782) );
  NAND2_X1 U16089 ( .A1(n12783), .A2(n12782), .ZN(n14710) );
  NAND2_X1 U16090 ( .A1(n14710), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12786) );
  INV_X1 U16091 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14898) );
  INV_X1 U16092 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14732) );
  NAND2_X1 U16093 ( .A1(n14898), .A2(n14732), .ZN(n14890) );
  NOR2_X1 U16094 ( .A1(n14740), .A2(n10228), .ZN(n14722) );
  NAND2_X1 U16095 ( .A1(n14722), .A2(n14877), .ZN(n14711) );
  NAND2_X1 U16096 ( .A1(n14711), .A2(n12784), .ZN(n12785) );
  NAND2_X1 U16097 ( .A1(n12786), .A2(n12785), .ZN(n12788) );
  OR2_X1 U16098 ( .A1(n12790), .A2(n20781), .ZN(n12792) );
  NAND2_X1 U16099 ( .A1(n12791), .A2(n11773), .ZN(n13818) );
  NAND2_X1 U16100 ( .A1(n12792), .A2(n13818), .ZN(n13020) );
  NOR2_X1 U16101 ( .A1(n12793), .A2(n20781), .ZN(n12794) );
  NAND2_X1 U16102 ( .A1(n14392), .A2(n12794), .ZN(n13025) );
  OAI21_X1 U16103 ( .B1(n14395), .B2(n12795), .A(n13025), .ZN(n12796) );
  NAND2_X1 U16104 ( .A1(n12796), .A2(n14397), .ZN(n12797) );
  AND2_X1 U16105 ( .A1(n14704), .A2(n20264), .ZN(n12799) );
  NAND2_X1 U16106 ( .A1(n12800), .A2(n12799), .ZN(n12816) );
  INV_X1 U16107 ( .A(n13786), .ZN(n12801) );
  NOR4_X1 U16108 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12805) );
  NOR4_X1 U16109 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12804) );
  NOR4_X1 U16110 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12803) );
  NOR4_X1 U16111 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12802) );
  AND4_X1 U16112 ( .A1(n12805), .A2(n12804), .A3(n12803), .A4(n12802), .ZN(
        n12810) );
  NOR4_X1 U16113 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12808) );
  NOR4_X1 U16114 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12807) );
  NOR4_X1 U16115 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12806) );
  INV_X1 U16116 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20797) );
  AND4_X1 U16117 ( .A1(n12808), .A2(n12807), .A3(n12806), .A4(n20797), .ZN(
        n12809) );
  NAND2_X1 U16118 ( .A1(n12810), .A2(n12809), .ZN(n12811) );
  NOR2_X2 U16119 ( .A1(n13425), .A2(n14628), .ZN(n15987) );
  AOI22_X1 U16120 ( .A1(n15987), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15985), .ZN(n12812) );
  INV_X1 U16121 ( .A(n12812), .ZN(n12814) );
  INV_X1 U16122 ( .A(n14628), .ZN(n13411) );
  INV_X1 U16123 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19338) );
  NOR2_X1 U16124 ( .A1(n15992), .A2(n19338), .ZN(n12813) );
  NOR2_X1 U16125 ( .A1(n12814), .A2(n12813), .ZN(n12815) );
  NAND2_X1 U16126 ( .A1(n12816), .A2(n12815), .ZN(P1_U2873) );
  NOR2_X1 U16127 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12818) );
  NOR4_X1 U16128 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12817) );
  NAND4_X1 U16129 ( .A1(n12818), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n12817), .ZN(n12832) );
  NOR4_X1 U16130 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12821)
         );
  NAND2_X1 U16131 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(P1_W_R_N_REG_SCAN_IN), 
        .ZN(n12819) );
  NOR3_X1 U16132 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n12819), .ZN(n12820) );
  NAND3_X1 U16133 ( .A1(n14628), .A2(n12821), .A3(n12820), .ZN(U214) );
  NOR4_X1 U16134 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12825) );
  NOR4_X1 U16135 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_0__SCAN_IN), .ZN(n12824) );
  NOR4_X1 U16136 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12823) );
  NOR4_X1 U16137 ( .A1(P2_ADDRESS_REG_21__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12822) );
  NAND4_X1 U16138 ( .A1(n12825), .A2(n12824), .A3(n12823), .A4(n12822), .ZN(
        n12830) );
  NOR4_X1 U16139 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_7__SCAN_IN), .A4(
        P2_ADDRESS_REG_6__SCAN_IN), .ZN(n12828) );
  NOR4_X1 U16140 ( .A1(P2_ADDRESS_REG_12__SCAN_IN), .A2(
        P2_ADDRESS_REG_11__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_5__SCAN_IN), .ZN(n12827) );
  NOR4_X1 U16141 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n12826) );
  NAND4_X1 U16142 ( .A1(n12828), .A2(n12827), .A3(n12826), .A4(n21024), .ZN(
        n12829) );
  NOR2_X1 U16143 ( .A1(n14376), .A2(n12832), .ZN(n16493) );
  NAND2_X1 U16144 ( .A1(n16493), .A2(U214), .ZN(U212) );
  NOR3_X1 U16145 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16923) );
  NAND2_X1 U16146 ( .A1(n16923), .A2(n17263), .ZN(n16920) );
  NOR2_X1 U16147 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16920), .ZN(n16896) );
  INV_X1 U16148 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17257) );
  NAND2_X1 U16149 ( .A1(n16896), .A2(n17257), .ZN(n16889) );
  NOR2_X1 U16150 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16889), .ZN(n16872) );
  INV_X1 U16151 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16863) );
  NAND2_X1 U16152 ( .A1(n16872), .A2(n16863), .ZN(n16862) );
  INV_X1 U16153 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16846) );
  NAND2_X1 U16154 ( .A1(n16839), .A2(n16846), .ZN(n16830) );
  NAND2_X1 U16155 ( .A1(n16829), .A2(n16823), .ZN(n16815) );
  NAND2_X1 U16156 ( .A1(n16800), .A2(n16795), .ZN(n16794) );
  NAND2_X1 U16157 ( .A1(n16776), .A2(n16769), .ZN(n16767) );
  INV_X1 U16158 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17094) );
  NAND2_X1 U16159 ( .A1(n16755), .A2(n17094), .ZN(n16746) );
  INV_X1 U16160 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16721) );
  NAND2_X1 U16161 ( .A1(n16733), .A2(n16721), .ZN(n16719) );
  INV_X1 U16162 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17051) );
  NAND2_X1 U16163 ( .A1(n16705), .A2(n17051), .ZN(n16700) );
  INV_X1 U16164 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16679) );
  NAND2_X1 U16165 ( .A1(n16685), .A2(n16679), .ZN(n16678) );
  INV_X1 U16166 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16658) );
  NAND2_X1 U16167 ( .A1(n16663), .A2(n16658), .ZN(n16657) );
  NOR2_X1 U16168 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16657), .ZN(n16647) );
  NAND2_X1 U16169 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18809) );
  INV_X1 U16170 ( .A(n18809), .ZN(n18941) );
  NOR2_X1 U16171 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n18941), .ZN(n12837) );
  NAND2_X1 U16172 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18933), .ZN(n12836) );
  NOR3_X4 U16173 ( .A1(n12837), .A2(n12851), .A3(n12836), .ZN(n16954) );
  AOI211_X1 U16174 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16657), .A(n16647), .B(
        n16947), .ZN(n12856) );
  INV_X1 U16175 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21158) );
  NOR2_X1 U16176 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18806) );
  OAI211_X1 U16177 ( .C1(n18933), .C2(n18932), .A(n18809), .B(n16580), .ZN(
        n12850) );
  INV_X1 U16178 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18866) );
  INV_X1 U16179 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18862) );
  INV_X1 U16180 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18857) );
  INV_X1 U16181 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18855) );
  INV_X1 U16182 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18841) );
  INV_X1 U16183 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18836) );
  NAND3_X1 U16184 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16900) );
  NAND4_X1 U16185 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(P3_REIP_REG_5__SCAN_IN), .A4(P3_REIP_REG_4__SCAN_IN), .ZN(n16853)
         );
  NOR3_X1 U16186 ( .A1(n18836), .A2(n16900), .A3(n16853), .ZN(n16811) );
  INV_X1 U16187 ( .A(n16811), .ZN(n16824) );
  INV_X1 U16188 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18839) );
  NOR4_X1 U16189 ( .A1(n18841), .A2(n16824), .A3(n18839), .A4(n18837), .ZN(
        n16803) );
  AND2_X1 U16190 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16803), .ZN(n16790) );
  NAND3_X1 U16191 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16790), .ZN(n16722) );
  NAND3_X1 U16192 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16723) );
  NOR4_X1 U16193 ( .A1(n18857), .A2(n18855), .A3(n16722), .A4(n16723), .ZN(
        n16711) );
  NAND2_X1 U16194 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16711), .ZN(n16703) );
  NOR2_X1 U16195 ( .A1(n18862), .A2(n16703), .ZN(n16684) );
  NAND2_X1 U16196 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16684), .ZN(n16675) );
  NOR2_X1 U16197 ( .A1(n18866), .A2(n16675), .ZN(n16673) );
  NAND2_X1 U16198 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16673), .ZN(n12839) );
  NOR2_X1 U16199 ( .A1(n16943), .A2(n12839), .ZN(n16656) );
  NAND2_X1 U16200 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16656), .ZN(n16599) );
  INV_X2 U16201 ( .A(n16718), .ZN(n18235) );
  INV_X1 U16202 ( .A(n18660), .ZN(n18794) );
  NOR3_X1 U16203 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18936), .A3(n18794), 
        .ZN(n12838) );
  NOR4_X4 U16204 ( .A1(n18235), .A2(n18951), .A3(n16941), .A4(n12838), .ZN(
        n16950) );
  NOR3_X1 U16205 ( .A1(n16950), .A2(n12839), .A3(n21158), .ZN(n12840) );
  INV_X1 U16206 ( .A(n16950), .ZN(n16957) );
  NAND2_X1 U16207 ( .A1(n16943), .A2(n16957), .ZN(n16956) );
  AOI21_X1 U16208 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n12840), .A(n16902), 
        .ZN(n16645) );
  INV_X1 U16209 ( .A(n16645), .ZN(n12841) );
  AOI21_X1 U16210 ( .B1(n21158), .B2(n16599), .A(n12841), .ZN(n12855) );
  NOR2_X1 U16211 ( .A1(n17910), .A2(n17591), .ZN(n12844) );
  INV_X1 U16212 ( .A(n12844), .ZN(n12845) );
  NOR2_X1 U16213 ( .A1(n17592), .A2(n12845), .ZN(n17548) );
  NAND2_X1 U16214 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17548), .ZN(
        n16607) );
  OAI21_X1 U16215 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17548), .A(
        n16607), .ZN(n12842) );
  INV_X1 U16216 ( .A(n12842), .ZN(n17578) );
  INV_X1 U16217 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16653) );
  NAND2_X1 U16218 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12844), .ZN(
        n12843) );
  AOI21_X1 U16219 ( .B1(n16653), .B2(n12843), .A(n17548), .ZN(n17590) );
  INV_X1 U16220 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17604) );
  OAI22_X1 U16221 ( .A1(n17604), .A2(n12844), .B1(n12845), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17602) );
  INV_X1 U16222 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16693) );
  INV_X1 U16223 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12848) );
  NOR2_X1 U16224 ( .A1(n17910), .A2(n17673), .ZN(n17672) );
  INV_X1 U16225 ( .A(n17672), .ZN(n16729) );
  NOR2_X1 U16226 ( .A1(n17674), .A2(n16729), .ZN(n17636) );
  INV_X1 U16227 ( .A(n17636), .ZN(n16715) );
  NOR2_X1 U16228 ( .A1(n12848), .A2(n16715), .ZN(n12847) );
  NAND2_X1 U16229 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12847), .ZN(
        n12846) );
  NOR2_X1 U16230 ( .A1(n16693), .A2(n12846), .ZN(n17588) );
  OAI21_X1 U16231 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17588), .A(
        n12845), .ZN(n17625) );
  INV_X1 U16232 ( .A(n17625), .ZN(n16672) );
  AOI21_X1 U16233 ( .B1(n16693), .B2(n12846), .A(n17588), .ZN(n17638) );
  OAI21_X1 U16234 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12847), .A(
        n12846), .ZN(n17646) );
  INV_X1 U16235 ( .A(n17646), .ZN(n16696) );
  AOI21_X1 U16236 ( .B1(n12848), .B2(n16715), .A(n12847), .ZN(n17666) );
  NOR2_X1 U16237 ( .A1(n17910), .A2(n17712), .ZN(n17711) );
  NAND2_X1 U16238 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17711), .ZN(
        n16764) );
  NOR2_X1 U16239 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16764), .ZN(
        n16752) );
  AOI21_X1 U16240 ( .B1(n17636), .B2(n16752), .A(n16884), .ZN(n16707) );
  NOR2_X1 U16241 ( .A1(n17666), .A2(n16707), .ZN(n16706) );
  NOR2_X1 U16242 ( .A1(n16706), .A2(n16884), .ZN(n16695) );
  NOR2_X1 U16243 ( .A1(n16672), .A2(n9856), .ZN(n16671) );
  NOR2_X1 U16244 ( .A1(n16671), .A2(n16884), .ZN(n16665) );
  NOR2_X1 U16245 ( .A1(n17578), .A2(n12849), .ZN(n16608) );
  AOI211_X1 U16246 ( .C1(n17578), .C2(n12849), .A(n16608), .B(n18800), .ZN(
        n12854) );
  INV_X1 U16247 ( .A(n12850), .ZN(n18785) );
  AOI211_X4 U16248 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18933), .A(n18785), .B(
        n12851), .ZN(n16955) );
  AOI22_X1 U16249 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16939), .B1(
        n16955), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n12852) );
  INV_X1 U16250 ( .A(n12852), .ZN(n12853) );
  NAND2_X1 U16251 ( .A1(n10328), .A2(n12857), .ZN(n12858) );
  INV_X1 U16252 ( .A(n11340), .ZN(n15702) );
  NAND2_X1 U16253 ( .A1(n15702), .A2(n12969), .ZN(n19202) );
  INV_X1 U16254 ( .A(n19981), .ZN(n12861) );
  INV_X1 U16255 ( .A(n11546), .ZN(n12860) );
  OAI21_X1 U16256 ( .B1(n18957), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n12861), 
        .ZN(n12859) );
  OAI21_X1 U16257 ( .B1(n12861), .B2(n12860), .A(n12859), .ZN(P2_U3612) );
  OAI21_X1 U16258 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n12863), .A(
        n12862), .ZN(n16361) );
  INV_X1 U16259 ( .A(n16361), .ZN(n12866) );
  NAND2_X1 U16260 ( .A1(n15118), .A2(n16365), .ZN(n12864) );
  NAND2_X1 U16261 ( .A1(n12936), .A2(n12864), .ZN(n16368) );
  NAND2_X1 U16262 ( .A1(n19088), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16366) );
  OAI21_X1 U16263 ( .B1(n16292), .B2(n16368), .A(n16366), .ZN(n12865) );
  AOI21_X1 U16264 ( .B1(n16287), .B2(n12866), .A(n12865), .ZN(n12869) );
  OAI21_X1 U16265 ( .B1(n16299), .B2(n12867), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12868) );
  OAI211_X1 U16266 ( .C1(n16317), .C2(n10073), .A(n12869), .B(n12868), .ZN(
        P2_U3014) );
  AND2_X1 U16267 ( .A1(n20846), .A2(n16162), .ZN(n13495) );
  AOI21_X1 U16268 ( .B1(n12870), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13495), 
        .ZN(n12871) );
  NAND2_X1 U16269 ( .A1(n13114), .A2(n12871), .ZN(P1_U2801) );
  INV_X1 U16270 ( .A(n13539), .ZN(n18956) );
  AOI22_X1 U16271 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n12905), .B1(n13538), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12874) );
  NOR3_X1 U16272 ( .A1(n13539), .A2(n14294), .A3(n19976), .ZN(n12872) );
  CLKBUF_X1 U16273 ( .A(n12872), .Z(n12953) );
  AOI22_X1 U16274 ( .A1(n14372), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14376), .ZN(n19342) );
  INV_X1 U16275 ( .A(n19342), .ZN(n12873) );
  NAND2_X1 U16276 ( .A1(n12953), .A2(n12873), .ZN(n12875) );
  NAND2_X1 U16277 ( .A1(n12874), .A2(n12875), .ZN(P2_U2974) );
  AOI22_X1 U16278 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n12932), .B1(n13538), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12876) );
  NAND2_X1 U16279 ( .A1(n12876), .A2(n12875), .ZN(P2_U2959) );
  AOI22_X1 U16280 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n12932), .B1(n13538), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12877) );
  AOI22_X1 U16281 ( .A1(n14372), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14376), .ZN(n15273) );
  INV_X1 U16282 ( .A(n15273), .ZN(n19191) );
  NAND2_X1 U16283 ( .A1(n12953), .A2(n19191), .ZN(n12880) );
  NAND2_X1 U16284 ( .A1(n12877), .A2(n12880), .ZN(P2_U2957) );
  AOI22_X1 U16285 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n12905), .B1(n13538), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U16286 ( .A1(n14372), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14376), .ZN(n19320) );
  INV_X1 U16287 ( .A(n19320), .ZN(n13355) );
  NAND2_X1 U16288 ( .A1(n12953), .A2(n13355), .ZN(n12882) );
  NAND2_X1 U16289 ( .A1(n12878), .A2(n12882), .ZN(P2_U2970) );
  AOI22_X1 U16290 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n12932), .B1(n13538), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U16291 ( .A1(n14372), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14376), .ZN(n15288) );
  INV_X1 U16292 ( .A(n15288), .ZN(n13057) );
  NAND2_X1 U16293 ( .A1(n12953), .A2(n13057), .ZN(n12884) );
  NAND2_X1 U16294 ( .A1(n12879), .A2(n12884), .ZN(P2_U2968) );
  AOI22_X1 U16295 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n12905), .B1(n13538), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12881) );
  NAND2_X1 U16296 ( .A1(n12881), .A2(n12880), .ZN(P2_U2972) );
  AOI22_X1 U16297 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n12932), .B1(n13538), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12883) );
  NAND2_X1 U16298 ( .A1(n12883), .A2(n12882), .ZN(P2_U2955) );
  AOI22_X1 U16299 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n12932), .B1(n13538), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12885) );
  NAND2_X1 U16300 ( .A1(n12885), .A2(n12884), .ZN(P2_U2953) );
  AOI22_X1 U16301 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n12905), .B1(n13538), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12886) );
  OAI22_X1 U16302 ( .A1(n14376), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14372), .ZN(n12997) );
  INV_X1 U16303 ( .A(n12997), .ZN(n16235) );
  NAND2_X1 U16304 ( .A1(n12953), .A2(n16235), .ZN(n12887) );
  NAND2_X1 U16305 ( .A1(n12886), .A2(n12887), .ZN(P2_U2958) );
  AOI22_X1 U16306 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n12905), .B1(n13531), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12888) );
  NAND2_X1 U16307 ( .A1(n12888), .A2(n12887), .ZN(P2_U2973) );
  AOI22_X1 U16308 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n12905), .B1(n13538), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12892) );
  INV_X1 U16309 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12889) );
  OR2_X1 U16310 ( .A1(n14376), .A2(n12889), .ZN(n12891) );
  NAND2_X1 U16311 ( .A1(n14376), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12890) );
  NAND2_X1 U16312 ( .A1(n12891), .A2(n12890), .ZN(n15240) );
  NAND2_X1 U16313 ( .A1(n12953), .A2(n15240), .ZN(n12903) );
  NAND2_X1 U16314 ( .A1(n12892), .A2(n12903), .ZN(P2_U2978) );
  AOI22_X1 U16315 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n12905), .B1(n13531), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12895) );
  INV_X1 U16316 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16525) );
  OR2_X1 U16317 ( .A1(n14376), .A2(n16525), .ZN(n12894) );
  NAND2_X1 U16318 ( .A1(n14376), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U16319 ( .A1(n12894), .A2(n12893), .ZN(n15252) );
  NAND2_X1 U16320 ( .A1(n12953), .A2(n15252), .ZN(n12896) );
  NAND2_X1 U16321 ( .A1(n12895), .A2(n12896), .ZN(P2_U2976) );
  AOI22_X1 U16322 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n12905), .B1(n13531), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12897) );
  NAND2_X1 U16323 ( .A1(n12897), .A2(n12896), .ZN(P2_U2961) );
  AOI22_X1 U16324 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n12932), .B1(n13531), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12900) );
  INV_X1 U16325 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13166) );
  OR2_X1 U16326 ( .A1(n14376), .A2(n13166), .ZN(n12899) );
  NAND2_X1 U16327 ( .A1(n14376), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12898) );
  NAND2_X1 U16328 ( .A1(n12899), .A2(n12898), .ZN(n15228) );
  NAND2_X1 U16329 ( .A1(n12953), .A2(n15228), .ZN(n12901) );
  NAND2_X1 U16330 ( .A1(n12900), .A2(n12901), .ZN(P2_U2965) );
  AOI22_X1 U16331 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n12905), .B1(n13531), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12902) );
  NAND2_X1 U16332 ( .A1(n12902), .A2(n12901), .ZN(P2_U2980) );
  AOI22_X1 U16333 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n12932), .B1(n13538), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U16334 ( .A1(n12904), .A2(n12903), .ZN(P2_U2963) );
  AOI22_X1 U16335 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n12905), .B1(n13531), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12907) );
  OAI22_X1 U16336 ( .A1(n14376), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14372), .ZN(n12906) );
  INV_X1 U16337 ( .A(n12906), .ZN(n19314) );
  NAND2_X1 U16338 ( .A1(n12953), .A2(n19314), .ZN(n12910) );
  NAND2_X1 U16339 ( .A1(n12907), .A2(n12910), .ZN(P2_U2969) );
  AOI22_X1 U16340 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n12932), .B1(n13538), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12909) );
  OAI22_X1 U16341 ( .A1(n14376), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14372), .ZN(n12908) );
  INV_X1 U16342 ( .A(n12908), .ZN(n19326) );
  NAND2_X1 U16343 ( .A1(n12953), .A2(n19326), .ZN(n12912) );
  NAND2_X1 U16344 ( .A1(n12909), .A2(n12912), .ZN(P2_U2956) );
  AOI22_X1 U16345 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n12932), .B1(n13531), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12911) );
  NAND2_X1 U16346 ( .A1(n12911), .A2(n12910), .ZN(P2_U2954) );
  AOI22_X1 U16347 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n12932), .B1(n13531), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12913) );
  NAND2_X1 U16348 ( .A1(n12913), .A2(n12912), .ZN(P2_U2971) );
  INV_X1 U16349 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n19210) );
  INV_X1 U16350 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14629) );
  OR2_X1 U16351 ( .A1(n14376), .A2(n14629), .ZN(n12915) );
  NAND2_X1 U16352 ( .A1(n14376), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12914) );
  AND2_X1 U16353 ( .A1(n12915), .A2(n12914), .ZN(n14375) );
  INV_X1 U16354 ( .A(n14375), .ZN(n19178) );
  NAND2_X1 U16355 ( .A1(n12953), .A2(n19178), .ZN(n12924) );
  NAND2_X1 U16356 ( .A1(n12932), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12916) );
  OAI211_X1 U16357 ( .C1(n19210), .C2(n19201), .A(n12924), .B(n12916), .ZN(
        P2_U2966) );
  INV_X1 U16358 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19214) );
  INV_X1 U16359 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16520) );
  OR2_X1 U16360 ( .A1(n14376), .A2(n16520), .ZN(n12918) );
  NAND2_X1 U16361 ( .A1(n14376), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12917) );
  AND2_X1 U16362 ( .A1(n12918), .A2(n12917), .ZN(n15234) );
  INV_X1 U16363 ( .A(n15234), .ZN(n19181) );
  NAND2_X1 U16364 ( .A1(n12953), .A2(n19181), .ZN(n12928) );
  NAND2_X1 U16365 ( .A1(n12932), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12919) );
  OAI211_X1 U16366 ( .C1(n19214), .C2(n19201), .A(n12928), .B(n12919), .ZN(
        P2_U2964) );
  INV_X1 U16367 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19252) );
  INV_X1 U16368 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16527) );
  OR2_X1 U16369 ( .A1(n14376), .A2(n16527), .ZN(n12921) );
  NAND2_X1 U16370 ( .A1(n14376), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12920) );
  AND2_X1 U16371 ( .A1(n12921), .A2(n12920), .ZN(n15260) );
  INV_X1 U16372 ( .A(n15260), .ZN(n19187) );
  NAND2_X1 U16373 ( .A1(n12953), .A2(n19187), .ZN(n12926) );
  NAND2_X1 U16374 ( .A1(n12932), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12922) );
  OAI211_X1 U16375 ( .C1(n19252), .C2(n19201), .A(n12926), .B(n12922), .ZN(
        P2_U2975) );
  INV_X1 U16376 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19241) );
  NAND2_X1 U16377 ( .A1(n12932), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12923) );
  OAI211_X1 U16378 ( .C1(n19241), .C2(n19201), .A(n12924), .B(n12923), .ZN(
        P2_U2981) );
  INV_X1 U16379 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19222) );
  NAND2_X1 U16380 ( .A1(n12932), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12925) );
  OAI211_X1 U16381 ( .C1(n19222), .C2(n19201), .A(n12926), .B(n12925), .ZN(
        P2_U2960) );
  INV_X1 U16382 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19245) );
  NAND2_X1 U16383 ( .A1(n12932), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12927) );
  OAI211_X1 U16384 ( .C1(n19245), .C2(n19201), .A(n12928), .B(n12927), .ZN(
        P2_U2979) );
  INV_X1 U16385 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19249) );
  INV_X1 U16386 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16523) );
  OR2_X1 U16387 ( .A1(n14376), .A2(n16523), .ZN(n12930) );
  NAND2_X1 U16388 ( .A1(n14376), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12929) );
  NAND2_X1 U16389 ( .A1(n12930), .A2(n12929), .ZN(n19184) );
  NAND2_X1 U16390 ( .A1(n12953), .A2(n19184), .ZN(n12934) );
  NAND2_X1 U16391 ( .A1(n12932), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12931) );
  OAI211_X1 U16392 ( .C1(n19249), .C2(n19201), .A(n12934), .B(n12931), .ZN(
        P2_U2977) );
  INV_X1 U16393 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19218) );
  NAND2_X1 U16394 ( .A1(n12932), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12933) );
  OAI211_X1 U16395 ( .C1(n19218), .C2(n19201), .A(n12934), .B(n12933), .ZN(
        P2_U2962) );
  OAI21_X1 U16396 ( .B1(n13710), .B2(n12936), .A(n12935), .ZN(n12937) );
  XNOR2_X1 U16397 ( .A(n12937), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15687) );
  AND2_X1 U16398 ( .A1(n19088), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15685) );
  OAI21_X1 U16399 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12939), .A(
        n12938), .ZN(n15683) );
  OAI22_X1 U16400 ( .A1(n19282), .A2(n15683), .B1(n13705), .B2(n19288), .ZN(
        n12940) );
  AOI211_X1 U16401 ( .C1(n19276), .C2(n15687), .A(n15685), .B(n12940), .ZN(
        n12942) );
  NAND2_X1 U16402 ( .A1(n19274), .A2(n13705), .ZN(n12941) );
  OAI211_X1 U16403 ( .C1(n10619), .C2(n16317), .A(n12942), .B(n12941), .ZN(
        P2_U3013) );
  INV_X1 U16404 ( .A(n12943), .ZN(n12944) );
  AOI21_X1 U16405 ( .B1(n12946), .B2(n12945), .A(n12944), .ZN(n19302) );
  AOI21_X1 U16406 ( .B1(n13705), .B2(n13553), .A(n13443), .ZN(n13551) );
  AOI22_X1 U16407 ( .A1(n19302), .A2(n19276), .B1(n19274), .B2(n13551), .ZN(
        n12952) );
  OAI21_X1 U16408 ( .B1(n12949), .B2(n12948), .A(n12947), .ZN(n19294) );
  NAND2_X1 U16409 ( .A1(n19088), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19293) );
  OAI21_X1 U16410 ( .B1(n19282), .B2(n19294), .A(n19293), .ZN(n12950) );
  AOI21_X1 U16411 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16299), .A(
        n12950), .ZN(n12951) );
  OAI211_X1 U16412 ( .C1(n10655), .C2(n16317), .A(n12952), .B(n12951), .ZN(
        P2_U3012) );
  INV_X1 U16413 ( .A(n12953), .ZN(n12988) );
  OAI22_X1 U16414 ( .A1(n14376), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14372), .ZN(n13616) );
  INV_X1 U16415 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12954) );
  INV_X1 U16416 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19238) );
  OAI222_X1 U16417 ( .A1(n12988), .A2(n13616), .B1(n12954), .B2(n12989), .C1(
        n19201), .C2(n19238), .ZN(P2_U2952) );
  NAND2_X1 U16418 ( .A1(n13570), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12956) );
  AOI22_X1 U16419 ( .A1(n13146), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19924), .B2(n19958), .ZN(n12957) );
  NOR2_X1 U16420 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12960) );
  OAI21_X1 U16421 ( .B1(n11375), .B2(n12960), .A(n12959), .ZN(n12961) );
  MUX2_X1 U16422 ( .A(n10073), .B(n15119), .S(n15212), .Z(n12962) );
  OAI21_X1 U16423 ( .B1(n15219), .B2(n15124), .A(n12962), .ZN(P2_U2887) );
  NAND2_X1 U16424 ( .A1(n16402), .A2(n15743), .ZN(n12965) );
  AND2_X1 U16425 ( .A1(n11546), .A2(n19983), .ZN(n16389) );
  NAND2_X1 U16426 ( .A1(n11360), .A2(n16389), .ZN(n12963) );
  OR2_X1 U16427 ( .A1(n16398), .A2(n12963), .ZN(n12964) );
  NAND2_X1 U16428 ( .A1(n12965), .A2(n12964), .ZN(n15699) );
  NOR2_X1 U16429 ( .A1(n12967), .A2(n12966), .ZN(n12968) );
  NAND2_X1 U16430 ( .A1(n11367), .A2(n12972), .ZN(n12971) );
  INV_X1 U16431 ( .A(n11381), .ZN(n12978) );
  INV_X1 U16432 ( .A(n12973), .ZN(n12976) );
  INV_X1 U16433 ( .A(n12974), .ZN(n12975) );
  NAND2_X1 U16434 ( .A1(n12976), .A2(n12975), .ZN(n12977) );
  NAND2_X1 U16435 ( .A1(n12978), .A2(n12977), .ZN(n16359) );
  INV_X1 U16436 ( .A(n16359), .ZN(n12980) );
  AOI22_X1 U16437 ( .A1(n16246), .A2(n12980), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19190), .ZN(n12982) );
  NOR2_X1 U16438 ( .A1(n15124), .A2(n16359), .ZN(n13056) );
  INV_X1 U16439 ( .A(n13056), .ZN(n12979) );
  OAI211_X1 U16440 ( .C1(n19955), .C2(n12980), .A(n12979), .B(n19194), .ZN(
        n12981) );
  OAI211_X1 U16441 ( .C1(n13505), .C2(n13616), .A(n12982), .B(n12981), .ZN(
        P2_U2919) );
  INV_X1 U16442 ( .A(n20878), .ZN(n12984) );
  OAI21_X1 U16443 ( .B1(n13495), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n12984), 
        .ZN(n12983) );
  OAI21_X1 U16444 ( .B1(n12985), .B2(n12984), .A(n12983), .ZN(P1_U3487) );
  INV_X1 U16445 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12986) );
  OAI222_X1 U16446 ( .A1(n12987), .A2(n19201), .B1(n12986), .B2(n12989), .C1(
        n12988), .C2(n13616), .ZN(P2_U2967) );
  INV_X1 U16447 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12991) );
  INV_X1 U16448 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16449 ( .A1(n14372), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14376), .ZN(n13504) );
  OAI222_X1 U16450 ( .A1(n19201), .A2(n12991), .B1(n12990), .B2(n12989), .C1(
        n12988), .C2(n13504), .ZN(P2_U2982) );
  NAND2_X1 U16451 ( .A1(n13146), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12992) );
  XNOR2_X1 U16452 ( .A(n19958), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13743) );
  NAND2_X1 U16453 ( .A1(n13743), .A2(n19924), .ZN(n19606) );
  NAND2_X1 U16454 ( .A1(n12992), .A2(n19606), .ZN(n12993) );
  OR2_X1 U16455 ( .A1(n13036), .A2(n19313), .ZN(n13047) );
  MUX2_X1 U16456 ( .A(n10619), .B(n13706), .S(n15212), .Z(n12994) );
  OAI21_X1 U16457 ( .B1(n13715), .B2(n15219), .A(n12994), .ZN(P2_U2886) );
  XNOR2_X1 U16458 ( .A(n12996), .B(n12995), .ZN(n15677) );
  INV_X1 U16459 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19256) );
  OAI222_X1 U16460 ( .A1(n13505), .A2(n12997), .B1(n15677), .B2(n19200), .C1(
        n19256), .C2(n15286), .ZN(P2_U2913) );
  INV_X1 U16461 ( .A(n11939), .ZN(n20857) );
  AOI21_X1 U16462 ( .B1(n13779), .B2(n13786), .A(n12998), .ZN(n13005) );
  AND2_X1 U16463 ( .A1(n12999), .A2(n13794), .ZN(n13000) );
  NAND2_X1 U16464 ( .A1(n13001), .A2(n13000), .ZN(n13023) );
  INV_X1 U16465 ( .A(n13002), .ZN(n13003) );
  NAND2_X1 U16466 ( .A1(n13003), .A2(n12529), .ZN(n13004) );
  OAI211_X1 U16467 ( .C1(n20238), .C2(n13005), .A(n13023), .B(n13004), .ZN(
        n13797) );
  INV_X1 U16468 ( .A(n13006), .ZN(n13009) );
  NOR2_X1 U16469 ( .A1(n13007), .A2(n13667), .ZN(n13008) );
  NOR2_X1 U16470 ( .A1(n13009), .A2(n13008), .ZN(n13793) );
  AND2_X1 U16471 ( .A1(n13795), .A2(n13792), .ZN(n13011) );
  INV_X1 U16472 ( .A(n15858), .ZN(n13019) );
  NAND4_X1 U16473 ( .A1(n13793), .A2(n13011), .A3(n13019), .A4(n13010), .ZN(
        n13012) );
  NOR2_X1 U16474 ( .A1(n13797), .A2(n13012), .ZN(n13014) );
  AND3_X1 U16475 ( .A1(n12793), .A2(n13014), .A3(n13013), .ZN(n13098) );
  OAI22_X1 U16476 ( .A1(n20857), .A2(n13098), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13015), .ZN(n15835) );
  INV_X1 U16477 ( .A(n15835), .ZN(n13016) );
  OAI21_X1 U16478 ( .B1(n13016), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n16162), 
        .ZN(n13017) );
  NAND2_X1 U16479 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U16480 ( .A1(n13017), .A2(n13106), .B1(n13240), .B2(n13030), .ZN(
        n13032) );
  NAND2_X1 U16481 ( .A1(n12645), .A2(n11758), .ZN(n13802) );
  NAND2_X1 U16482 ( .A1(n15856), .A2(n20880), .ZN(n13018) );
  AOI21_X1 U16483 ( .B1(n13802), .B2(n13019), .A(n13018), .ZN(n13021) );
  OR2_X1 U16484 ( .A1(n13021), .A2(n13020), .ZN(n13027) );
  INV_X1 U16485 ( .A(n12645), .ZN(n14383) );
  NAND2_X1 U16486 ( .A1(n13023), .A2(n13022), .ZN(n13024) );
  NAND2_X1 U16487 ( .A1(n14383), .A2(n13024), .ZN(n13781) );
  OAI211_X1 U16488 ( .C1(n13667), .C2(n13779), .A(n13025), .B(n13781), .ZN(
        n13026) );
  AOI21_X1 U16489 ( .B1(n14388), .B2(n13027), .A(n13026), .ZN(n13028) );
  NAND2_X1 U16490 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16159) );
  INV_X1 U16491 ( .A(n16159), .ZN(n15864) );
  NAND2_X1 U16492 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15864), .ZN(n16163) );
  INV_X1 U16493 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20000) );
  OAI22_X1 U16494 ( .A1(n15838), .A2(n19992), .B1(n16163), .B2(n20000), .ZN(
        n16149) );
  AOI21_X1 U16495 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n16155), .A(n16149), 
        .ZN(n13067) );
  NOR2_X1 U16496 ( .A1(n13802), .A2(n13030), .ZN(n15834) );
  AOI22_X1 U16497 ( .A1(n15834), .A2(n19990), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13067), .ZN(n13031) );
  OAI21_X1 U16498 ( .B1(n13032), .B2(n13067), .A(n13031), .ZN(P1_U3474) );
  OAI21_X1 U16499 ( .B1(n13035), .B2(n13034), .A(n13033), .ZN(n19134) );
  OAI222_X1 U16500 ( .A1(n13505), .A2(n19342), .B1(n19134), .B2(n19200), .C1(
        n19254), .C2(n15286), .ZN(P2_U2912) );
  NAND2_X1 U16501 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19407) );
  NAND2_X1 U16502 ( .A1(n19407), .A2(n13038), .ZN(n13040) );
  NAND2_X1 U16503 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19724) );
  INV_X1 U16504 ( .A(n19724), .ZN(n13039) );
  NAND2_X1 U16505 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13039), .ZN(
        n13142) );
  NAND2_X1 U16506 ( .A1(n13040), .A2(n13142), .ZN(n13744) );
  NOR2_X1 U16507 ( .A1(n19722), .A2(n13744), .ZN(n13041) );
  AOI21_X1 U16508 ( .B1(n13146), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13041), .ZN(n13042) );
  NAND2_X1 U16509 ( .A1(n13046), .A2(n13045), .ZN(n13050) );
  NAND2_X1 U16510 ( .A1(n13048), .A2(n13047), .ZN(n13049) );
  MUX2_X1 U16511 ( .A(n10407), .B(n10655), .S(n15224), .Z(n13051) );
  OAI21_X1 U16512 ( .B1(n19938), .B2(n15219), .A(n13051), .ZN(P2_U2885) );
  XNOR2_X1 U16513 ( .A(n13053), .B(n13052), .ZN(n19948) );
  INV_X1 U16514 ( .A(n19948), .ZN(n13054) );
  NAND2_X1 U16515 ( .A1(n13715), .A2(n13054), .ZN(n13246) );
  OAI21_X1 U16516 ( .B1(n13715), .B2(n13054), .A(n13246), .ZN(n13055) );
  NOR2_X1 U16517 ( .A1(n13055), .A2(n13056), .ZN(n13248) );
  AOI21_X1 U16518 ( .B1(n13056), .B2(n13055), .A(n13248), .ZN(n13060) );
  AOI22_X1 U16519 ( .A1(n19192), .A2(n13057), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19190), .ZN(n13059) );
  NAND2_X1 U16520 ( .A1(n16246), .A2(n19948), .ZN(n13058) );
  OAI211_X1 U16521 ( .C1(n13060), .C2(n19171), .A(n13059), .B(n13058), .ZN(
        P2_U2918) );
  INV_X1 U16522 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13063) );
  OR2_X1 U16523 ( .A1(n12638), .A2(n11758), .ZN(n13823) );
  AOI21_X1 U16524 ( .B1(n13802), .B2(n13823), .A(n15880), .ZN(n13061) );
  NAND2_X1 U16525 ( .A1(n20104), .A2(n13794), .ZN(n13306) );
  NAND2_X1 U16526 ( .A1(n16155), .A2(n15864), .ZN(n20106) );
  INV_X2 U16527 ( .A(n20106), .ZN(n20121) );
  NOR2_X4 U16528 ( .A1(n20104), .A2(n20121), .ZN(n20112) );
  AOI22_X1 U16529 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13062) );
  OAI21_X1 U16530 ( .B1(n13063), .B2(n13306), .A(n13062), .ZN(P1_U2912) );
  AOI22_X1 U16531 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13064) );
  OAI21_X1 U16532 ( .B1(n14648), .B2(n13306), .A(n13064), .ZN(P1_U2910) );
  AOI22_X1 U16533 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13065) );
  OAI21_X1 U16534 ( .B1(n14638), .B2(n13306), .A(n13065), .ZN(P1_U2908) );
  AOI22_X1 U16535 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13066) );
  OAI21_X1 U16536 ( .B1(n14634), .B2(n13306), .A(n13066), .ZN(P1_U2907) );
  INV_X1 U16537 ( .A(n13067), .ZN(n16151) );
  INV_X1 U16538 ( .A(n13098), .ZN(n13227) );
  INV_X1 U16539 ( .A(n13069), .ZN(n13074) );
  INV_X1 U16540 ( .A(n13070), .ZN(n13073) );
  NAND3_X1 U16541 ( .A1(n13777), .A2(n13074), .A3(n13073), .ZN(n13071) );
  OAI21_X1 U16542 ( .B1(n13802), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13071), .ZN(n13072) );
  AOI21_X1 U16543 ( .B1(n20678), .B2(n13227), .A(n13072), .ZN(n15837) );
  INV_X1 U16544 ( .A(n19990), .ZN(n15016) );
  NOR2_X1 U16545 ( .A1(n15837), .A2(n15016), .ZN(n13077) );
  AOI22_X1 U16546 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20219), .B2(n12787), .ZN(
        n13108) );
  NAND3_X1 U16547 ( .A1(n13074), .A2(n13240), .A3(n13073), .ZN(n13075) );
  OAI21_X1 U16548 ( .B1(n13108), .B2(n13106), .A(n13075), .ZN(n13076) );
  OAI21_X1 U16549 ( .B1(n13077), .B2(n13076), .A(n16151), .ZN(n13078) );
  OAI21_X1 U16550 ( .B1(n16151), .B2(n13079), .A(n13078), .ZN(P1_U3473) );
  INV_X1 U16551 ( .A(n20159), .ZN(n20175) );
  NAND2_X1 U16552 ( .A1(n13081), .A2(n13080), .ZN(n13082) );
  NAND2_X1 U16553 ( .A1(n13083), .A2(n13082), .ZN(n14544) );
  NAND2_X1 U16554 ( .A1(n13084), .A2(n14805), .ZN(n13089) );
  INV_X2 U16555 ( .A(n20208), .ZN(n20164) );
  NAND2_X1 U16556 ( .A1(n20164), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20222) );
  INV_X1 U16557 ( .A(n20222), .ZN(n13088) );
  OAI21_X1 U16558 ( .B1(n13086), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13085), .ZN(n20221) );
  NOR2_X1 U16559 ( .A1(n19999), .A2(n20221), .ZN(n13087) );
  AOI211_X1 U16560 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13089), .A(
        n13088), .B(n13087), .ZN(n13090) );
  OAI21_X1 U16561 ( .B1(n20175), .B2(n14544), .A(n13090), .ZN(P1_U2999) );
  OR2_X1 U16562 ( .A1(n13092), .A2(n13091), .ZN(n13093) );
  NAND2_X1 U16563 ( .A1(n13126), .A2(n13093), .ZN(n20174) );
  XNOR2_X1 U16564 ( .A(n13666), .B(n14394), .ZN(n20209) );
  OAI22_X1 U16565 ( .A1(n20209), .A2(n14608), .B1(n14626), .B2(n13094), .ZN(
        n13095) );
  INV_X1 U16566 ( .A(n13095), .ZN(n13096) );
  OAI21_X1 U16567 ( .B1(n14627), .B2(n20174), .A(n13096), .ZN(P1_U2871) );
  INV_X1 U16568 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13111) );
  OR2_X1 U16569 ( .A1(n20612), .A2(n13098), .ZN(n13105) );
  INV_X1 U16570 ( .A(n13818), .ZN(n14384) );
  OR2_X1 U16571 ( .A1(n14385), .A2(n14384), .ZN(n13216) );
  XNOR2_X1 U16572 ( .A(n13070), .B(n13111), .ZN(n13107) );
  INV_X1 U16573 ( .A(n13107), .ZN(n13103) );
  XNOR2_X1 U16574 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13101) );
  NAND3_X1 U16575 ( .A1(n13777), .A2(n9890), .A3(n13107), .ZN(n13100) );
  OAI21_X1 U16576 ( .B1(n13802), .B2(n13101), .A(n13100), .ZN(n13102) );
  AOI21_X1 U16577 ( .B1(n13216), .B2(n13103), .A(n13102), .ZN(n13104) );
  NAND2_X1 U16578 ( .A1(n13105), .A2(n13104), .ZN(n13214) );
  INV_X1 U16579 ( .A(n13106), .ZN(n13109) );
  AOI222_X1 U16580 ( .A1(n13214), .A2(n19990), .B1(n13109), .B2(n13108), .C1(
        n13240), .C2(n13107), .ZN(n13110) );
  MUX2_X1 U16581 ( .A(n13111), .B(n13110), .S(n16151), .Z(n13112) );
  INV_X1 U16582 ( .A(n13112), .ZN(P1_U3472) );
  AND2_X2 U16583 ( .A1(n13176), .A2(n20238), .ZN(n20151) );
  INV_X2 U16584 ( .A(n13176), .ZN(n20150) );
  AOI22_X1 U16585 ( .A1(n20151), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13117) );
  NAND2_X1 U16586 ( .A1(n13176), .A2(n11758), .ZN(n13177) );
  INV_X1 U16587 ( .A(DATAI_4_), .ZN(n13116) );
  NAND2_X1 U16588 ( .A1(n14628), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13115) );
  OAI21_X1 U16589 ( .B1(n14628), .B2(n13116), .A(n13115), .ZN(n20250) );
  NAND2_X1 U16590 ( .A1(n20136), .A2(n20250), .ZN(n13121) );
  NAND2_X1 U16591 ( .A1(n13117), .A2(n13121), .ZN(P1_U2941) );
  AOI22_X1 U16592 ( .A1(n20151), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13120) );
  INV_X1 U16593 ( .A(DATAI_0_), .ZN(n13119) );
  NAND2_X1 U16594 ( .A1(n14628), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13118) );
  OAI21_X1 U16595 ( .B1(n14628), .B2(n13119), .A(n13118), .ZN(n13429) );
  NAND2_X1 U16596 ( .A1(n20136), .A2(n13429), .ZN(n13366) );
  NAND2_X1 U16597 ( .A1(n13120), .A2(n13366), .ZN(P1_U2937) );
  AOI22_X1 U16598 ( .A1(n20151), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13122) );
  NAND2_X1 U16599 ( .A1(n13122), .A2(n13121), .ZN(P1_U2956) );
  AOI22_X1 U16600 ( .A1(n20151), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13125) );
  INV_X1 U16601 ( .A(DATAI_7_), .ZN(n13124) );
  NAND2_X1 U16602 ( .A1(n14628), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13123) );
  OAI21_X1 U16603 ( .B1(n14628), .B2(n13124), .A(n13123), .ZN(n20270) );
  NAND2_X1 U16604 ( .A1(n20136), .A2(n20270), .ZN(n13359) );
  NAND2_X1 U16605 ( .A1(n13125), .A2(n13359), .ZN(P1_U2944) );
  NAND2_X1 U16606 ( .A1(n13127), .A2(n13126), .ZN(n13128) );
  INV_X1 U16607 ( .A(n20090), .ZN(n13427) );
  INV_X1 U16608 ( .A(n13130), .ZN(n20085) );
  INV_X1 U16609 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13131) );
  INV_X1 U16610 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20083) );
  OAI22_X1 U16611 ( .A1(n14805), .A2(n13131), .B1(n20208), .B2(n20083), .ZN(
        n13132) );
  AOI21_X1 U16612 ( .B1(n20085), .B2(n20171), .A(n13132), .ZN(n13136) );
  OR2_X1 U16613 ( .A1(n13134), .A2(n13133), .ZN(n20198) );
  NAND3_X1 U16614 ( .A1(n20198), .A2(n20197), .A3(n20169), .ZN(n13135) );
  OAI211_X1 U16615 ( .C1(n13427), .C2(n20175), .A(n13136), .B(n13135), .ZN(
        P1_U2997) );
  NAND2_X1 U16616 ( .A1(n15755), .A2(n13141), .ZN(n13148) );
  INV_X1 U16617 ( .A(n13142), .ZN(n13143) );
  NAND2_X1 U16618 ( .A1(n13143), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19773) );
  OAI211_X1 U16619 ( .C1(n13143), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19773), .B(n19924), .ZN(n13144) );
  INV_X1 U16620 ( .A(n13144), .ZN(n13145) );
  AOI21_X1 U16621 ( .B1(n13146), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13145), .ZN(n13147) );
  NOR2_X1 U16622 ( .A1(n13154), .A2(n15205), .ZN(n13155) );
  AOI21_X1 U16623 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n15205), .A(n13155), .ZN(
        n13156) );
  OAI21_X1 U16624 ( .B1(n19354), .B2(n15219), .A(n13156), .ZN(P2_U2884) );
  INV_X1 U16625 ( .A(n15252), .ZN(n13159) );
  INV_X1 U16626 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n21085) );
  OAI21_X1 U16627 ( .B1(n13643), .B2(n13158), .A(n13157), .ZN(n19120) );
  OAI222_X1 U16628 ( .A1(n13505), .A2(n13159), .B1(n15286), .B2(n21085), .C1(
        n19200), .C2(n19120), .ZN(P2_U2910) );
  INV_X1 U16629 ( .A(n20151), .ZN(n13178) );
  NAND2_X1 U16630 ( .A1(n14628), .A2(n12889), .ZN(n13160) );
  OAI21_X1 U16631 ( .B1(n14628), .B2(DATAI_11_), .A(n13160), .ZN(n14643) );
  INV_X1 U16632 ( .A(n14643), .ZN(n13161) );
  NAND2_X1 U16633 ( .A1(n20136), .A2(n13161), .ZN(n20144) );
  NAND2_X1 U16634 ( .A1(n20150), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13162) );
  OAI211_X1 U16635 ( .C1(n13178), .C2(n14642), .A(n20144), .B(n13162), .ZN(
        P1_U2948) );
  INV_X1 U16636 ( .A(DATAI_12_), .ZN(n13163) );
  MUX2_X1 U16637 ( .A(n13163), .B(n16520), .S(n14628), .Z(n14707) );
  INV_X1 U16638 ( .A(n14707), .ZN(n13164) );
  NAND2_X1 U16639 ( .A1(n20136), .A2(n13164), .ZN(n20146) );
  NAND2_X1 U16640 ( .A1(n20150), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13165) );
  OAI211_X1 U16641 ( .C1(n13178), .C2(n14638), .A(n20146), .B(n13165), .ZN(
        P1_U2949) );
  INV_X1 U16642 ( .A(DATAI_13_), .ZN(n13167) );
  MUX2_X1 U16643 ( .A(n13167), .B(n13166), .S(n14628), .Z(n14703) );
  INV_X1 U16644 ( .A(n14703), .ZN(n13168) );
  NAND2_X1 U16645 ( .A1(n20136), .A2(n13168), .ZN(n20148) );
  NAND2_X1 U16646 ( .A1(n20150), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13169) );
  OAI211_X1 U16647 ( .C1(n13178), .C2(n14634), .A(n20148), .B(n13169), .ZN(
        P1_U2950) );
  INV_X1 U16648 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13173) );
  NOR2_X1 U16649 ( .A1(n13171), .A2(n13170), .ZN(n13172) );
  OR2_X1 U16650 ( .A1(n13284), .A2(n13172), .ZN(n20196) );
  OAI222_X1 U16651 ( .A1(n13427), .A2(n14627), .B1(n14626), .B2(n13173), .C1(
        n20196), .C2(n14608), .ZN(P1_U2870) );
  INV_X1 U16652 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14698) );
  INV_X1 U16653 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13174) );
  NOR2_X1 U16654 ( .A1(n13411), .A2(n13174), .ZN(n13175) );
  AOI21_X1 U16655 ( .B1(DATAI_15_), .B2(n13411), .A(n13175), .ZN(n14699) );
  INV_X1 U16656 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20100) );
  OAI222_X1 U16657 ( .A1(n13178), .A2(n14698), .B1(n13177), .B2(n14699), .C1(
        n13176), .C2(n20100), .ZN(P1_U2967) );
  INV_X1 U16658 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14539) );
  OR2_X1 U16659 ( .A1(n13179), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13180) );
  NAND2_X1 U16660 ( .A1(n13181), .A2(n13180), .ZN(n20225) );
  OAI222_X1 U16661 ( .A1(n14544), .A2(n14627), .B1(n14539), .B2(n14626), .C1(
        n14608), .C2(n20225), .ZN(P1_U2872) );
  NAND2_X1 U16662 ( .A1(n13182), .A2(n13183), .ZN(n13184) );
  INV_X1 U16663 ( .A(n16338), .ZN(n13196) );
  NAND2_X1 U16664 ( .A1(n13570), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13185) );
  AND2_X1 U16665 ( .A1(n13186), .A2(n13185), .ZN(n13187) );
  AND2_X1 U16666 ( .A1(n14288), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13197) );
  AND2_X1 U16667 ( .A1(n14065), .A2(n13197), .ZN(n13189) );
  NAND2_X1 U16668 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13311) );
  NOR2_X1 U16669 ( .A1(n19348), .A2(n13311), .ZN(n13190) );
  AND2_X1 U16670 ( .A1(n13189), .A2(n13190), .ZN(n13193) );
  AND2_X1 U16671 ( .A1(n13192), .A2(n13190), .ZN(n13191) );
  AND2_X1 U16672 ( .A1(n13191), .A2(n13197), .ZN(n13206) );
  NAND2_X1 U16673 ( .A1(n14065), .A2(n13206), .ZN(n13260) );
  OAI211_X1 U16674 ( .C1(n13193), .C2(n13192), .A(n13260), .B(n15199), .ZN(
        n13195) );
  NAND2_X1 U16675 ( .A1(n15212), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13194) );
  OAI211_X1 U16676 ( .C1(n13196), .C2(n15205), .A(n13195), .B(n13194), .ZN(
        P2_U2879) );
  OR2_X1 U16677 ( .A1(n14065), .A2(n13197), .ZN(n13198) );
  NAND2_X1 U16678 ( .A1(n14065), .A2(n13197), .ZN(n13312) );
  NAND2_X1 U16679 ( .A1(n13198), .A2(n13312), .ZN(n19193) );
  NAND2_X1 U16680 ( .A1(n15212), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n13204) );
  INV_X1 U16681 ( .A(n13200), .ZN(n13201) );
  NAND2_X1 U16682 ( .A1(n10423), .A2(n13201), .ZN(n13202) );
  AND2_X1 U16683 ( .A1(n13202), .A2(n13269), .ZN(n19279) );
  NAND2_X1 U16684 ( .A1(n19279), .A2(n15224), .ZN(n13203) );
  OAI211_X1 U16685 ( .C1(n19193), .C2(n15219), .A(n13204), .B(n13203), .ZN(
        P2_U2883) );
  INV_X1 U16686 ( .A(n13261), .ZN(n13205) );
  NOR2_X1 U16687 ( .A1(n13260), .A2(n13205), .ZN(n13209) );
  AND2_X1 U16688 ( .A1(n13208), .A2(n13261), .ZN(n13207) );
  AND2_X1 U16689 ( .A1(n13207), .A2(n13206), .ZN(n13328) );
  NAND2_X1 U16690 ( .A1(n14065), .A2(n13328), .ZN(n13330) );
  OAI211_X1 U16691 ( .C1(n13209), .C2(n13208), .A(n15199), .B(n13330), .ZN(
        n13213) );
  OR2_X1 U16692 ( .A1(n13264), .A2(n13210), .ZN(n13211) );
  NAND2_X1 U16693 ( .A1(n13326), .A2(n13211), .ZN(n16285) );
  INV_X1 U16694 ( .A(n16285), .ZN(n19110) );
  NAND2_X1 U16695 ( .A1(n19110), .A2(n15224), .ZN(n13212) );
  OAI211_X1 U16696 ( .C1(n15224), .C2(n10009), .A(n13213), .B(n13212), .ZN(
        P2_U2877) );
  NOR2_X1 U16697 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16162), .ZN(n13232) );
  MUX2_X1 U16698 ( .A(n13214), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15838), .Z(n15841) );
  AOI22_X1 U16699 ( .A1(n13232), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15841), .B2(n16162), .ZN(n13234) );
  MUX2_X1 U16700 ( .A(n13215), .B(n11619), .S(n13070), .Z(n13217) );
  OAI21_X1 U16701 ( .B1(n13218), .B2(n13217), .A(n13216), .ZN(n13225) );
  AOI21_X1 U16702 ( .B1(n13070), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n15019), .ZN(n13219) );
  NOR2_X1 U16703 ( .A1(n11792), .A2(n13219), .ZN(n15013) );
  NAND3_X1 U16704 ( .A1(n13777), .A2(n9890), .A3(n15013), .ZN(n13224) );
  INV_X1 U16705 ( .A(n13802), .ZN(n13831) );
  NAND2_X1 U16706 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13220) );
  INV_X1 U16707 ( .A(n13220), .ZN(n13221) );
  MUX2_X1 U16708 ( .A(n13221), .B(n13220), .S(n15019), .Z(n13222) );
  NAND2_X1 U16709 ( .A1(n13831), .A2(n13222), .ZN(n13223) );
  NAND3_X1 U16710 ( .A1(n13225), .A2(n13224), .A3(n13223), .ZN(n13226) );
  AOI21_X1 U16711 ( .B1(n20476), .B2(n13227), .A(n13226), .ZN(n15017) );
  MUX2_X1 U16712 ( .A(n15017), .B(n11619), .S(n15838), .Z(n13228) );
  AOI22_X1 U16713 ( .A1(n13232), .A2(n15019), .B1(n16162), .B2(n15844), .ZN(
        n13233) );
  INV_X1 U16714 ( .A(n20365), .ZN(n20611) );
  XNOR2_X1 U16715 ( .A(n13229), .B(n11963), .ZN(n20071) );
  NOR2_X1 U16716 ( .A1(n20071), .A2(n12793), .ZN(n16148) );
  OAI21_X1 U16717 ( .B1(n15838), .B2(n16148), .A(n16162), .ZN(n13230) );
  AOI21_X1 U16718 ( .B1(n15838), .B2(n11963), .A(n13230), .ZN(n13231) );
  AOI21_X1 U16719 ( .B1(n13232), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13231), .ZN(n13236) );
  OAI21_X1 U16720 ( .B1(n13234), .B2(n13233), .A(n13236), .ZN(n15853) );
  NAND2_X1 U16721 ( .A1(n13236), .A2(n13069), .ZN(n13237) );
  NAND2_X1 U16722 ( .A1(n15853), .A2(n13237), .ZN(n15865) );
  NAND2_X1 U16723 ( .A1(n15865), .A2(n20000), .ZN(n13239) );
  INV_X1 U16724 ( .A(n16163), .ZN(n13238) );
  NAND2_X1 U16725 ( .A1(n13239), .A2(n13238), .ZN(n13241) );
  OAI21_X1 U16726 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(
        P1_STATE2_REG_1__SCAN_IN), .A(n16155), .ZN(n20875) );
  AND2_X1 U16727 ( .A1(n20615), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20858) );
  AND2_X1 U16728 ( .A1(n9817), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20332) );
  AOI21_X1 U16729 ( .B1(n20481), .B2(n20332), .A(n20859), .ZN(n20720) );
  OAI21_X1 U16730 ( .B1(n20481), .B2(n20332), .A(n20720), .ZN(n13243) );
  OAI21_X1 U16731 ( .B1(n20858), .B2(n20612), .A(n13243), .ZN(n13244) );
  NAND2_X1 U16732 ( .A1(n20864), .A2(n13244), .ZN(n13245) );
  OAI21_X1 U16733 ( .B1(n20864), .B2(n11859), .A(n13245), .ZN(P1_U3476) );
  INV_X1 U16734 ( .A(n13246), .ZN(n13247) );
  NOR2_X1 U16735 ( .A1(n13248), .A2(n13247), .ZN(n13256) );
  NAND2_X1 U16736 ( .A1(n13250), .A2(n13249), .ZN(n13253) );
  INV_X1 U16737 ( .A(n13251), .ZN(n13252) );
  NAND2_X1 U16738 ( .A1(n13253), .A2(n13252), .ZN(n19940) );
  INV_X1 U16739 ( .A(n19940), .ZN(n13254) );
  NAND2_X1 U16740 ( .A1(n19938), .A2(n13254), .ZN(n13346) );
  OAI21_X1 U16741 ( .B1(n19938), .B2(n13254), .A(n13346), .ZN(n13255) );
  NOR2_X1 U16742 ( .A1(n13256), .A2(n13255), .ZN(n13348) );
  AOI21_X1 U16743 ( .B1(n13256), .B2(n13255), .A(n13348), .ZN(n13259) );
  AOI22_X1 U16744 ( .A1(n19192), .A2(n19314), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19190), .ZN(n13258) );
  NAND2_X1 U16745 ( .A1(n19940), .A2(n16246), .ZN(n13257) );
  OAI211_X1 U16746 ( .C1(n13259), .C2(n19171), .A(n13258), .B(n13257), .ZN(
        P2_U2917) );
  XOR2_X1 U16747 ( .A(n13261), .B(n13260), .Z(n13267) );
  AND2_X1 U16748 ( .A1(n13263), .A2(n13262), .ZN(n13265) );
  OR2_X1 U16749 ( .A1(n13265), .A2(n13264), .ZN(n19119) );
  MUX2_X1 U16750 ( .A(n19119), .B(n10008), .S(n15212), .Z(n13266) );
  OAI21_X1 U16751 ( .B1(n13267), .B2(n15219), .A(n13266), .ZN(P2_U2878) );
  XOR2_X1 U16752 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13312), .Z(n13273)
         );
  AND2_X1 U16753 ( .A1(n13269), .A2(n13268), .ZN(n13271) );
  OR2_X1 U16754 ( .A1(n13271), .A2(n13270), .ZN(n19152) );
  MUX2_X1 U16755 ( .A(n19152), .B(n10429), .S(n15212), .Z(n13272) );
  OAI21_X1 U16756 ( .B1(n13273), .B2(n15219), .A(n13272), .ZN(P2_U2882) );
  INV_X1 U16757 ( .A(n15240), .ZN(n13277) );
  OAI21_X1 U16758 ( .B1(n13276), .B2(n13275), .A(n13274), .ZN(n15639) );
  INV_X1 U16759 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19247) );
  OAI222_X1 U16760 ( .A1(n13505), .A2(n13277), .B1(n15639), .B2(n19200), .C1(
        n19247), .C2(n15286), .ZN(P2_U2908) );
  OR3_X1 U16761 ( .A1(n9817), .A2(n20859), .A3(n20847), .ZN(n20396) );
  INV_X1 U16762 ( .A(n20396), .ZN(n20853) );
  INV_X1 U16763 ( .A(n9817), .ZN(n13278) );
  NAND2_X1 U16764 ( .A1(n20846), .A2(n20847), .ZN(n20609) );
  OAI22_X1 U16765 ( .A1(n13278), .A2(n20609), .B1(n20613), .B2(n20858), .ZN(
        n13279) );
  OAI21_X1 U16766 ( .B1(n20853), .B2(n13279), .A(n20864), .ZN(n13280) );
  OAI21_X1 U16767 ( .B1(n20864), .B2(n20539), .A(n13280), .ZN(P1_U3477) );
  XOR2_X1 U16768 ( .A(n13281), .B(n13282), .Z(n13292) );
  OR2_X1 U16769 ( .A1(n13284), .A2(n13283), .ZN(n13285) );
  NAND2_X1 U16770 ( .A1(n13320), .A2(n13285), .ZN(n13683) );
  INV_X1 U16771 ( .A(n13683), .ZN(n20185) );
  AOI22_X1 U16772 ( .A1(n14614), .A2(n20185), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14612), .ZN(n13286) );
  OAI21_X1 U16773 ( .B1(n13690), .B2(n14627), .A(n13286), .ZN(P1_U2869) );
  OAI21_X1 U16774 ( .B1(n13289), .B2(n13288), .A(n13287), .ZN(n20187) );
  INV_X1 U16775 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13687) );
  NOR2_X1 U16776 ( .A1(n20208), .A2(n13687), .ZN(n20184) );
  AOI21_X1 U16777 ( .B1(n20165), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20184), .ZN(n13290) );
  OAI21_X1 U16778 ( .B1(n20163), .B2(n13679), .A(n13290), .ZN(n13291) );
  AOI21_X1 U16779 ( .B1(n13292), .B2(n20159), .A(n13291), .ZN(n13293) );
  OAI21_X1 U16780 ( .B1(n20187), .B2(n19999), .A(n13293), .ZN(P1_U2996) );
  INV_X1 U16781 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14676) );
  AOI22_X1 U16782 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13294) );
  OAI21_X1 U16783 ( .B1(n14676), .B2(n13306), .A(n13294), .ZN(P1_U2916) );
  INV_X1 U16784 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21096) );
  AOI22_X1 U16785 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13295) );
  OAI21_X1 U16786 ( .B1(n21096), .B2(n13306), .A(n13295), .ZN(P1_U2915) );
  AOI22_X1 U16787 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13296) );
  OAI21_X1 U16788 ( .B1(n14666), .B2(n13306), .A(n13296), .ZN(P1_U2914) );
  AOI22_X1 U16789 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13297) );
  OAI21_X1 U16790 ( .B1(n14660), .B2(n13306), .A(n13297), .ZN(P1_U2913) );
  AOI22_X1 U16791 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13298) );
  OAI21_X1 U16792 ( .B1(n14653), .B2(n13306), .A(n13298), .ZN(P1_U2911) );
  AOI22_X1 U16793 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13299) );
  OAI21_X1 U16794 ( .B1(n14642), .B2(n13306), .A(n13299), .ZN(P1_U2909) );
  AOI22_X1 U16795 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13300) );
  OAI21_X1 U16796 ( .B1(n12201), .B2(n13306), .A(n13300), .ZN(P1_U2918) );
  INV_X1 U16797 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14693) );
  AOI22_X1 U16798 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13301) );
  OAI21_X1 U16799 ( .B1(n14693), .B2(n13306), .A(n13301), .ZN(P1_U2920) );
  AOI22_X1 U16800 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13302) );
  OAI21_X1 U16801 ( .B1(n14686), .B2(n13306), .A(n13302), .ZN(P1_U2919) );
  INV_X1 U16802 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U16803 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13303) );
  OAI21_X1 U16804 ( .B1(n13304), .B2(n13306), .A(n13303), .ZN(P1_U2906) );
  INV_X1 U16805 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13307) );
  AOI22_X1 U16806 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13305) );
  OAI21_X1 U16807 ( .B1(n13307), .B2(n13306), .A(n13305), .ZN(P1_U2917) );
  OR2_X1 U16808 ( .A1(n13270), .A2(n13309), .ZN(n13310) );
  NAND2_X1 U16809 ( .A1(n13308), .A2(n13310), .ZN(n16316) );
  INV_X1 U16810 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13525) );
  NOR2_X1 U16811 ( .A1(n13312), .A2(n13525), .ZN(n13313) );
  OR2_X1 U16812 ( .A1(n13312), .A2(n13311), .ZN(n13341) );
  OAI211_X1 U16813 ( .C1(n13313), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15199), .B(n13341), .ZN(n13315) );
  NAND2_X1 U16814 ( .A1(n15212), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13314) );
  OAI211_X1 U16815 ( .C1(n16316), .C2(n15205), .A(n13315), .B(n13314), .ZN(
        P2_U2881) );
  AOI21_X1 U16816 ( .B1(n13318), .B2(n13317), .A(n13316), .ZN(n20158) );
  INV_X1 U16817 ( .A(n20158), .ZN(n13428) );
  NAND2_X1 U16818 ( .A1(n13320), .A2(n13319), .ZN(n13321) );
  NAND2_X1 U16819 ( .A1(n13338), .A2(n13321), .ZN(n20178) );
  INV_X1 U16820 ( .A(n20178), .ZN(n13322) );
  AOI22_X1 U16821 ( .A1(n14614), .A2(n13322), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14612), .ZN(n13323) );
  OAI21_X1 U16822 ( .B1(n13428), .B2(n14627), .A(n13323), .ZN(P1_U2868) );
  NAND2_X1 U16823 ( .A1(n13326), .A2(n13325), .ZN(n13327) );
  AND2_X1 U16824 ( .A1(n13324), .A2(n13327), .ZN(n19095) );
  NOR2_X1 U16825 ( .A1(n15224), .A2(n10449), .ZN(n13333) );
  INV_X1 U16826 ( .A(n13331), .ZN(n13329) );
  AND2_X1 U16827 ( .A1(n13329), .A2(n13328), .ZN(n13391) );
  AND2_X1 U16828 ( .A1(n14065), .A2(n13391), .ZN(n13394) );
  AOI211_X1 U16829 ( .C1(n13331), .C2(n13330), .A(n15219), .B(n13394), .ZN(
        n13332) );
  AOI211_X1 U16830 ( .C1(n19095), .C2(n15224), .A(n13333), .B(n13332), .ZN(
        n13334) );
  INV_X1 U16831 ( .A(n13334), .ZN(P2_U2876) );
  OR2_X1 U16832 ( .A1(n13316), .A2(n13336), .ZN(n13337) );
  AND2_X1 U16833 ( .A1(n13335), .A2(n13337), .ZN(n20063) );
  INV_X1 U16834 ( .A(n20063), .ZN(n13430) );
  INV_X1 U16835 ( .A(n13400), .ZN(n13454) );
  AOI21_X1 U16836 ( .B1(n13339), .B2(n13338), .A(n13454), .ZN(n20055) );
  AOI22_X1 U16837 ( .A1(n14614), .A2(n20055), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14612), .ZN(n13340) );
  OAI21_X1 U16838 ( .B1(n13430), .B2(n14627), .A(n13340), .ZN(P1_U2867) );
  XOR2_X1 U16839 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13341), .Z(n13345)
         );
  NAND2_X1 U16840 ( .A1(n13308), .A2(n13342), .ZN(n13343) );
  NAND2_X1 U16841 ( .A1(n13182), .A2(n13343), .ZN(n19135) );
  MUX2_X1 U16842 ( .A(n10847), .B(n19135), .S(n15224), .Z(n13344) );
  OAI21_X1 U16843 ( .B1(n13345), .B2(n15219), .A(n13344), .ZN(P2_U2880) );
  INV_X1 U16844 ( .A(n13346), .ZN(n13347) );
  NOR2_X1 U16845 ( .A1(n13348), .A2(n13347), .ZN(n13354) );
  OR2_X1 U16846 ( .A1(n13350), .A2(n13349), .ZN(n13352) );
  NAND2_X1 U16847 ( .A1(n13352), .A2(n13351), .ZN(n19932) );
  XNOR2_X1 U16848 ( .A(n19354), .B(n19932), .ZN(n13353) );
  NOR2_X1 U16849 ( .A1(n13354), .A2(n13353), .ZN(n13434) );
  AOI21_X1 U16850 ( .B1(n13354), .B2(n13353), .A(n13434), .ZN(n13358) );
  AOI22_X1 U16851 ( .A1(n19192), .A2(n13355), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19190), .ZN(n13357) );
  INV_X1 U16852 ( .A(n19932), .ZN(n16349) );
  NAND2_X1 U16853 ( .A1(n16349), .A2(n16246), .ZN(n13356) );
  OAI211_X1 U16854 ( .C1(n13358), .C2(n19171), .A(n13357), .B(n13356), .ZN(
        P2_U2916) );
  AOI22_X1 U16855 ( .A1(n20151), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13360) );
  NAND2_X1 U16856 ( .A1(n13360), .A2(n13359), .ZN(P1_U2959) );
  AOI22_X1 U16857 ( .A1(n20151), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13363) );
  INV_X1 U16858 ( .A(DATAI_6_), .ZN(n13362) );
  NAND2_X1 U16859 ( .A1(n14628), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13361) );
  OAI21_X1 U16860 ( .B1(n14628), .B2(n13362), .A(n13361), .ZN(n20259) );
  NAND2_X1 U16861 ( .A1(n20136), .A2(n20259), .ZN(n13364) );
  NAND2_X1 U16862 ( .A1(n13363), .A2(n13364), .ZN(P1_U2958) );
  AOI22_X1 U16863 ( .A1(n20151), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13365) );
  NAND2_X1 U16864 ( .A1(n13365), .A2(n13364), .ZN(P1_U2943) );
  AOI22_X1 U16865 ( .A1(n20151), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13367) );
  NAND2_X1 U16866 ( .A1(n13367), .A2(n13366), .ZN(P1_U2952) );
  AOI22_X1 U16867 ( .A1(n20151), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13370) );
  INV_X1 U16868 ( .A(DATAI_3_), .ZN(n13369) );
  NAND2_X1 U16869 ( .A1(n14628), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13368) );
  OAI21_X1 U16870 ( .B1(n14628), .B2(n13369), .A(n13368), .ZN(n20246) );
  NAND2_X1 U16871 ( .A1(n20136), .A2(n20246), .ZN(n13386) );
  NAND2_X1 U16872 ( .A1(n13370), .A2(n13386), .ZN(P1_U2955) );
  AOI22_X1 U16873 ( .A1(n20151), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13373) );
  INV_X1 U16874 ( .A(DATAI_2_), .ZN(n13372) );
  NAND2_X1 U16875 ( .A1(n14628), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13371) );
  OAI21_X1 U16876 ( .B1(n14628), .B2(n13372), .A(n13371), .ZN(n20242) );
  NAND2_X1 U16877 ( .A1(n20136), .A2(n20242), .ZN(n13384) );
  NAND2_X1 U16878 ( .A1(n13373), .A2(n13384), .ZN(P1_U2954) );
  AOI22_X1 U16879 ( .A1(n20151), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13376) );
  INV_X1 U16880 ( .A(DATAI_1_), .ZN(n13375) );
  NAND2_X1 U16881 ( .A1(n14628), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13374) );
  OAI21_X1 U16882 ( .B1(n14628), .B2(n13375), .A(n13374), .ZN(n20239) );
  NAND2_X1 U16883 ( .A1(n20136), .A2(n20239), .ZN(n13380) );
  NAND2_X1 U16884 ( .A1(n13376), .A2(n13380), .ZN(P1_U2953) );
  AOI22_X1 U16885 ( .A1(n20151), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13379) );
  INV_X1 U16886 ( .A(DATAI_5_), .ZN(n13378) );
  NAND2_X1 U16887 ( .A1(n14628), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13377) );
  OAI21_X1 U16888 ( .B1(n14628), .B2(n13378), .A(n13377), .ZN(n20255) );
  NAND2_X1 U16889 ( .A1(n20136), .A2(n20255), .ZN(n13382) );
  NAND2_X1 U16890 ( .A1(n13379), .A2(n13382), .ZN(P1_U2942) );
  AOI22_X1 U16891 ( .A1(n20151), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U16892 ( .A1(n13381), .A2(n13380), .ZN(P1_U2938) );
  AOI22_X1 U16893 ( .A1(n20151), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13383) );
  NAND2_X1 U16894 ( .A1(n13383), .A2(n13382), .ZN(P1_U2957) );
  AOI22_X1 U16895 ( .A1(n20151), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13385) );
  NAND2_X1 U16896 ( .A1(n13385), .A2(n13384), .ZN(P1_U2939) );
  AOI22_X1 U16897 ( .A1(n20151), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U16898 ( .A1(n13387), .A2(n13386), .ZN(P1_U2940) );
  AND2_X1 U16899 ( .A1(n13324), .A2(n13389), .ZN(n13390) );
  NOR2_X1 U16900 ( .A1(n13388), .A2(n13390), .ZN(n19081) );
  INV_X1 U16901 ( .A(n19081), .ZN(n13397) );
  AND2_X1 U16902 ( .A1(n14065), .A2(n13466), .ZN(n13457) );
  INV_X1 U16903 ( .A(n13457), .ZN(n13392) );
  OAI211_X1 U16904 ( .C1(n13394), .C2(n13393), .A(n13392), .B(n15199), .ZN(
        n13396) );
  NAND2_X1 U16905 ( .A1(n15212), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13395) );
  OAI211_X1 U16906 ( .C1(n13397), .C2(n15205), .A(n13396), .B(n13395), .ZN(
        P2_U2875) );
  AOI21_X1 U16907 ( .B1(n13399), .B2(n13335), .A(n12027), .ZN(n20051) );
  INV_X1 U16908 ( .A(n20051), .ZN(n13431) );
  XNOR2_X1 U16909 ( .A(n13400), .B(n13453), .ZN(n16131) );
  AOI22_X1 U16910 ( .A1(n14614), .A2(n16131), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14612), .ZN(n13401) );
  OAI21_X1 U16911 ( .B1(n13431), .B2(n14627), .A(n13401), .ZN(P1_U2866) );
  INV_X1 U16912 ( .A(n20481), .ZN(n20848) );
  NAND2_X1 U16913 ( .A1(n20481), .A2(n13402), .ZN(n20676) );
  AOI21_X1 U16914 ( .B1(n20292), .B2(n20775), .A(n20847), .ZN(n13404) );
  NOR2_X1 U16915 ( .A1(n13404), .A2(n20859), .ZN(n13406) );
  INV_X1 U16916 ( .A(n20612), .ZN(n20088) );
  OR2_X1 U16917 ( .A1(n20476), .A2(n20088), .ZN(n20335) );
  OR2_X1 U16918 ( .A1(n20335), .A2(n20678), .ZN(n13409) );
  NAND2_X1 U16919 ( .A1(n13408), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20673) );
  NAND2_X1 U16920 ( .A1(n20269), .A2(n20673), .ZN(n20480) );
  NOR2_X1 U16921 ( .A1(n20536), .A2(n20477), .ZN(n13407) );
  NOR3_X1 U16922 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20281) );
  INV_X1 U16923 ( .A(n20281), .ZN(n20278) );
  NOR2_X1 U16924 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20278), .ZN(
        n20268) );
  OAI22_X1 U16925 ( .A1(n13407), .A2(n20715), .B1(n20268), .B2(n20615), .ZN(
        n13405) );
  AOI211_X1 U16926 ( .C1(n13406), .C2(n13409), .A(n20480), .B(n13405), .ZN(
        n20263) );
  INV_X1 U16927 ( .A(n13406), .ZN(n13410) );
  INV_X1 U16928 ( .A(n13407), .ZN(n20366) );
  NOR2_X1 U16929 ( .A1(n13408), .A2(n20715), .ZN(n20538) );
  INV_X1 U16930 ( .A(n20538), .ZN(n20479) );
  NAND2_X1 U16931 ( .A1(n13429), .A2(n20269), .ZN(n20548) );
  NAND2_X1 U16932 ( .A1(n20159), .A2(n14628), .ZN(n20236) );
  NAND2_X1 U16933 ( .A1(n13411), .A2(n20159), .ZN(n20235) );
  NOR2_X1 U16934 ( .A1(n20775), .A2(n20727), .ZN(n13415) );
  INV_X1 U16935 ( .A(n20265), .ZN(n13412) );
  NAND2_X1 U16936 ( .A1(n13412), .A2(n13794), .ZN(n20275) );
  INV_X1 U16937 ( .A(n20268), .ZN(n13413) );
  AOI22_X1 U16938 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20267), .B1(DATAI_16_), 
        .B2(n20266), .ZN(n20649) );
  OAI22_X1 U16939 ( .A1(n20275), .A2(n13413), .B1(n20649), .B2(n20292), .ZN(
        n13414) );
  AOI211_X1 U16940 ( .C1(n20271), .C2(n20717), .A(n13415), .B(n13414), .ZN(
        n13416) );
  OAI21_X1 U16941 ( .B1(n20263), .B2(n13417), .A(n13416), .ZN(P1_U3033) );
  INV_X1 U16942 ( .A(n15228), .ZN(n13421) );
  INV_X1 U16943 ( .A(n13418), .ZN(n13419) );
  OAI21_X1 U16944 ( .B1(n15616), .B2(n13420), .A(n13419), .ZN(n19073) );
  INV_X1 U16945 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19243) );
  OAI222_X1 U16946 ( .A1(n13505), .A2(n13421), .B1(n19073), .B2(n19200), .C1(
        n19243), .C2(n15286), .ZN(P2_U2906) );
  NAND2_X1 U16947 ( .A1(n20254), .A2(n12524), .ZN(n13423) );
  AND2_X1 U16948 ( .A1(n13786), .A2(n13423), .ZN(n13422) );
  INV_X1 U16949 ( .A(n13423), .ZN(n13424) );
  INV_X1 U16950 ( .A(n20242), .ZN(n13426) );
  OAI222_X1 U16951 ( .A1(n13427), .A2(n14708), .B1(n14706), .B2(n13426), .C1(
        n14704), .C2(n11927), .ZN(P1_U2902) );
  INV_X1 U16952 ( .A(n20250), .ZN(n14677) );
  INV_X1 U16953 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20117) );
  OAI222_X1 U16954 ( .A1(n13428), .A2(n14708), .B1(n14677), .B2(n14706), .C1(
        n14704), .C2(n20117), .ZN(P1_U2900) );
  INV_X1 U16955 ( .A(n20239), .ZN(n14687) );
  OAI222_X1 U16956 ( .A1(n20174), .A2(n14708), .B1(n14687), .B2(n14706), .C1(
        n14704), .C2(n11931), .ZN(P1_U2903) );
  INV_X1 U16957 ( .A(n13429), .ZN(n14694) );
  INV_X1 U16958 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20124) );
  OAI222_X1 U16959 ( .A1(n14544), .A2(n14708), .B1(n14694), .B2(n14706), .C1(
        n14704), .C2(n20124), .ZN(P1_U2904) );
  INV_X1 U16960 ( .A(n20255), .ZN(n14672) );
  OAI222_X1 U16961 ( .A1(n13430), .A2(n14708), .B1(n14672), .B2(n14706), .C1(
        n14704), .C2(n11989), .ZN(P1_U2899) );
  INV_X1 U16962 ( .A(n20246), .ZN(n14682) );
  OAI222_X1 U16963 ( .A1(n13690), .A2(n14708), .B1(n14682), .B2(n14706), .C1(
        n14704), .C2(n11920), .ZN(P1_U2901) );
  INV_X1 U16964 ( .A(n20259), .ZN(n14667) );
  OAI222_X1 U16965 ( .A1(n13431), .A2(n14708), .B1(n14667), .B2(n14706), .C1(
        n20114), .C2(n14704), .ZN(P1_U2898) );
  XNOR2_X1 U16966 ( .A(n13351), .B(n13432), .ZN(n13658) );
  INV_X1 U16967 ( .A(n19354), .ZN(n19928) );
  NOR2_X1 U16968 ( .A1(n19928), .A2(n16349), .ZN(n13433) );
  OAI21_X1 U16969 ( .B1(n13434), .B2(n13433), .A(n13658), .ZN(n19196) );
  XNOR2_X1 U16970 ( .A(n19196), .B(n19193), .ZN(n13435) );
  NAND2_X1 U16971 ( .A1(n13435), .A2(n19194), .ZN(n13437) );
  AOI22_X1 U16972 ( .A1(n19192), .A2(n19326), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19190), .ZN(n13436) );
  OAI211_X1 U16973 ( .C1(n13658), .C2(n19170), .A(n13437), .B(n13436), .ZN(
        P2_U2915) );
  XNOR2_X1 U16974 ( .A(n13439), .B(n13438), .ZN(n16351) );
  XNOR2_X1 U16975 ( .A(n13440), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13441) );
  XNOR2_X1 U16976 ( .A(n13442), .B(n13441), .ZN(n16353) );
  NAND2_X1 U16977 ( .A1(n16353), .A2(n19276), .ZN(n13447) );
  INV_X1 U16978 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21048) );
  NAND2_X1 U16979 ( .A1(n19088), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16347) );
  OAI21_X1 U16980 ( .B1(n19288), .B2(n21048), .A(n16347), .ZN(n13445) );
  OAI21_X1 U16981 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13443), .A(
        n13623), .ZN(n13624) );
  NOR2_X1 U16982 ( .A1(n16314), .A2(n13624), .ZN(n13444) );
  AOI211_X1 U16983 ( .C1(n19278), .C2(n15755), .A(n13445), .B(n13444), .ZN(
        n13446) );
  OAI211_X1 U16984 ( .C1(n16351), .C2(n19282), .A(n13447), .B(n13446), .ZN(
        P2_U3011) );
  INV_X1 U16985 ( .A(n13449), .ZN(n13450) );
  AOI21_X1 U16986 ( .B1(n13451), .B2(n13398), .A(n13450), .ZN(n20039) );
  INV_X1 U16987 ( .A(n20039), .ZN(n13463) );
  AOI21_X1 U16988 ( .B1(n13454), .B2(n13453), .A(n13452), .ZN(n13455) );
  OR2_X1 U16989 ( .A1(n13455), .A2(n13695), .ZN(n20034) );
  INV_X1 U16990 ( .A(n20034), .ZN(n16125) );
  AOI22_X1 U16991 ( .A1(n14614), .A2(n16125), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14612), .ZN(n13456) );
  OAI21_X1 U16992 ( .B1(n13463), .B2(n14627), .A(n13456), .ZN(P1_U2865) );
  XNOR2_X1 U16993 ( .A(n13457), .B(n13467), .ZN(n13462) );
  NOR2_X1 U16994 ( .A1(n13388), .A2(n13459), .ZN(n13460) );
  OR2_X1 U16995 ( .A1(n13458), .A2(n13460), .ZN(n19069) );
  INV_X1 U16996 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n21127) );
  MUX2_X1 U16997 ( .A(n19069), .B(n21127), .S(n15212), .Z(n13461) );
  OAI21_X1 U16998 ( .B1(n13462), .B2(n15219), .A(n13461), .ZN(P2_U2874) );
  INV_X1 U16999 ( .A(n20270), .ZN(n14661) );
  OAI222_X1 U17000 ( .A1(n13463), .A2(n14708), .B1(n14661), .B2(n14706), .C1(
        n14704), .C2(n12024), .ZN(P1_U2897) );
  OR2_X1 U17001 ( .A1(n13458), .A2(n13464), .ZN(n13465) );
  AND2_X1 U17002 ( .A1(n15217), .A2(n13465), .ZN(n19057) );
  INV_X1 U17003 ( .A(n19057), .ZN(n13474) );
  AND2_X1 U17004 ( .A1(n14065), .A2(n13469), .ZN(n13471) );
  INV_X1 U17005 ( .A(n13468), .ZN(n13470) );
  NAND2_X1 U17006 ( .A1(n14065), .A2(n14062), .ZN(n15220) );
  OAI211_X1 U17007 ( .C1(n13471), .C2(n13470), .A(n15199), .B(n15220), .ZN(
        n13473) );
  NAND2_X1 U17008 ( .A1(n15212), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13472) );
  OAI211_X1 U17009 ( .C1(n13474), .C2(n15205), .A(n13473), .B(n13472), .ZN(
        P2_U2873) );
  NAND2_X1 U17010 ( .A1(n13476), .A2(n13475), .ZN(n13477) );
  XNOR2_X1 U17011 ( .A(n13477), .B(n13482), .ZN(n19283) );
  INV_X1 U17012 ( .A(n13478), .ZN(n13479) );
  XNOR2_X1 U17013 ( .A(n13480), .B(n13479), .ZN(n19277) );
  INV_X1 U17014 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19868) );
  INV_X2 U17015 ( .A(n19088), .ZN(n19131) );
  NOR2_X1 U17016 ( .A1(n19868), .A2(n19131), .ZN(n13481) );
  AOI221_X1 U17017 ( .B1(n13594), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n13586), .C2(n13482), .A(n13481), .ZN(n13484) );
  NAND2_X1 U17018 ( .A1(n19279), .A2(n16339), .ZN(n13483) );
  OAI211_X1 U17019 ( .C1(n16360), .C2(n13658), .A(n13484), .B(n13483), .ZN(
        n13485) );
  AOI21_X1 U17020 ( .B1(n19303), .B2(n19277), .A(n13485), .ZN(n13486) );
  OAI21_X1 U17021 ( .B1(n19295), .B2(n19283), .A(n13486), .ZN(P2_U3042) );
  AOI21_X1 U17022 ( .B1(n13488), .B2(n13449), .A(n13487), .ZN(n13489) );
  INV_X1 U17023 ( .A(n13489), .ZN(n13741) );
  INV_X1 U17024 ( .A(DATAI_8_), .ZN(n13490) );
  MUX2_X1 U17025 ( .A(n13490), .B(n16527), .S(n14628), .Z(n20125) );
  INV_X1 U17026 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13491) );
  OAI222_X1 U17027 ( .A1(n13741), .A2(n14708), .B1(n20125), .B2(n14706), .C1(
        n13491), .C2(n14704), .ZN(P1_U2896) );
  INV_X1 U17028 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13492) );
  XNOR2_X1 U17029 ( .A(n13695), .B(n13694), .ZN(n13494) );
  OAI222_X1 U17030 ( .A1(n14627), .A2(n13741), .B1(n13492), .B2(n14626), .C1(
        n14608), .C2(n13494), .ZN(P1_U2864) );
  NAND2_X1 U17031 ( .A1(n20054), .A2(n20079), .ZN(n20060) );
  NOR2_X1 U17032 ( .A1(n13493), .A2(n20060), .ZN(n14480) );
  NOR2_X1 U17033 ( .A1(n20062), .A2(n14480), .ZN(n20028) );
  INV_X1 U17034 ( .A(n13494), .ZN(n16111) );
  AOI22_X1 U17035 ( .A1(n20056), .A2(n16111), .B1(n20081), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n13496) );
  NAND2_X1 U17036 ( .A1(n20079), .A2(n13495), .ZN(n20022) );
  OAI211_X1 U17037 ( .C1(n20025), .C2(n13736), .A(n13496), .B(n20022), .ZN(
        n13497) );
  AOI21_X1 U17038 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n20028), .A(n13497), .ZN(
        n13502) );
  NAND4_X1 U17039 ( .A1(n20084), .A2(n20054), .A3(P1_REIP_REG_6__SCAN_IN), 
        .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n20037) );
  NOR2_X1 U17040 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20037), .ZN(n13500) );
  AOI22_X1 U17041 ( .A1(n13500), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n13738), 
        .B2(n20086), .ZN(n13501) );
  OAI211_X1 U17042 ( .C1(n13741), .C2(n15945), .A(n13502), .B(n13501), .ZN(
        P1_U2832) );
  OAI21_X1 U17043 ( .B1(n15587), .B2(n13503), .A(n15107), .ZN(n19046) );
  OAI222_X1 U17044 ( .A1(n13505), .A2(n13504), .B1(n19046), .B2(n19200), .C1(
        n12991), .C2(n15286), .ZN(P2_U2904) );
  NAND2_X1 U17045 ( .A1(n19834), .A2(n19373), .ZN(n13506) );
  NAND2_X1 U17046 ( .A1(n13506), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13507) );
  NAND2_X1 U17047 ( .A1(n13507), .A2(n19924), .ZN(n13522) );
  NAND2_X1 U17048 ( .A1(n19935), .A2(n13038), .ZN(n19406) );
  INV_X1 U17049 ( .A(n19406), .ZN(n13508) );
  NAND2_X1 U17050 ( .A1(n13508), .A2(n19950), .ZN(n19357) );
  NOR2_X1 U17051 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19357), .ZN(
        n19341) );
  INV_X1 U17052 ( .A(n19341), .ZN(n13516) );
  AND2_X1 U17053 ( .A1(n19773), .A2(n13516), .ZN(n13521) );
  INV_X1 U17054 ( .A(n13521), .ZN(n13509) );
  OR2_X1 U17055 ( .A1(n13522), .A2(n13509), .ZN(n13513) );
  INV_X1 U17056 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19975) );
  OAI21_X1 U17057 ( .B1(n13519), .B2(n19975), .A(n19951), .ZN(n13511) );
  NAND2_X1 U17058 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19206) );
  AOI21_X1 U17059 ( .B1(n13516), .B2(n13511), .A(n9793), .ZN(n13512) );
  AOI22_X1 U17060 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19343), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19344), .ZN(n19818) );
  INV_X1 U17061 ( .A(n19818), .ZN(n19753) );
  INV_X1 U17062 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16509) );
  INV_X1 U17063 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18285) );
  OAI22_X2 U17064 ( .A1(n16509), .A2(n19337), .B1(n18285), .B2(n19335), .ZN(
        n19813) );
  INV_X1 U17065 ( .A(n19813), .ZN(n13517) );
  NAND2_X1 U17066 ( .A1(n13515), .A2(n19319), .ZN(n19370) );
  OAI22_X1 U17067 ( .A1(n13517), .A2(n19373), .B1(n13516), .B2(n19370), .ZN(
        n13518) );
  AOI21_X1 U17068 ( .B1(n19814), .B2(n19753), .A(n13518), .ZN(n13524) );
  OAI21_X1 U17069 ( .B1(n13519), .B2(n19341), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13520) );
  NOR2_X2 U17070 ( .A1(n15273), .A2(n9793), .ZN(n19812) );
  NAND2_X1 U17071 ( .A1(n19345), .A2(n19812), .ZN(n13523) );
  OAI211_X1 U17072 ( .C1(n19349), .C2(n13525), .A(n13524), .B(n13523), .ZN(
        P2_U3053) );
  INV_X1 U17073 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14050) );
  AOI22_X1 U17074 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20977), .ZN(n15115) );
  AOI22_X1 U17075 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13705), .B2(n20977), .ZN(
        n13703) );
  NAND2_X1 U17076 ( .A1(n15115), .A2(n13703), .ZN(n13702) );
  NOR2_X1 U17077 ( .A1(n13551), .A2(n13702), .ZN(n13625) );
  NOR2_X1 U17078 ( .A1(n19147), .A2(n13625), .ZN(n13528) );
  XNOR2_X1 U17079 ( .A(n13528), .B(n13624), .ZN(n13529) );
  NAND4_X1 U17080 ( .A1(n19975), .A2(n20977), .A3(n10593), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19840) );
  NAND2_X1 U17081 ( .A1(n13529), .A2(n19154), .ZN(n13549) );
  NAND2_X1 U17082 ( .A1(n16388), .A2(n10593), .ZN(n16410) );
  INV_X1 U17083 ( .A(n16410), .ZN(n13530) );
  AND2_X1 U17084 ( .A1(n19981), .A2(n10376), .ZN(n13536) );
  NAND2_X1 U17085 ( .A1(n10593), .A2(n19983), .ZN(n13541) );
  INV_X1 U17086 ( .A(n13541), .ZN(n13532) );
  INV_X1 U17087 ( .A(n19837), .ZN(n18961) );
  NOR2_X1 U17088 ( .A1(n19951), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19510) );
  INV_X1 U17089 ( .A(n19510), .ZN(n19836) );
  NOR2_X1 U17090 ( .A1(n18961), .A2(n19836), .ZN(n16414) );
  NOR2_X1 U17091 ( .A1(n16414), .A2(n19154), .ZN(n13533) );
  NAND2_X1 U17092 ( .A1(n19131), .A2(n13533), .ZN(n13534) );
  AND2_X1 U17093 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13541), .ZN(n13535) );
  NOR2_X1 U17094 ( .A1(n19142), .A2(n13537), .ZN(n13545) );
  NAND2_X1 U17095 ( .A1(n13538), .A2(n16410), .ZN(n16166) );
  NOR2_X1 U17096 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13539), .ZN(n13540) );
  NAND2_X1 U17097 ( .A1(n13541), .A2(n13540), .ZN(n13542) );
  INV_X1 U17098 ( .A(n19128), .ZN(n19143) );
  INV_X1 U17099 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19866) );
  OAI22_X1 U17100 ( .A1(n19143), .A2(n13543), .B1(n19866), .B2(n19133), .ZN(
        n13544) );
  AOI211_X1 U17101 ( .C1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n19138), .A(
        n13545), .B(n13544), .ZN(n13546) );
  OAI21_X1 U17102 ( .B1(n10627), .B2(n19151), .A(n13546), .ZN(n13547) );
  AOI21_X1 U17103 ( .B1(n16349), .B2(n19089), .A(n13547), .ZN(n13548) );
  OAI211_X1 U17104 ( .C1(n19354), .C2(n18958), .A(n13549), .B(n13548), .ZN(
        P2_U2852) );
  NAND2_X1 U17105 ( .A1(n19075), .A2(n13702), .ZN(n13550) );
  XNOR2_X1 U17106 ( .A(n13551), .B(n13550), .ZN(n13559) );
  INV_X1 U17107 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19864) );
  OAI22_X1 U17108 ( .A1(n19142), .A2(n13552), .B1(n19864), .B2(n19133), .ZN(
        n13555) );
  OAI22_X1 U17109 ( .A1(n19143), .A2(n10407), .B1(n13553), .B2(n19158), .ZN(
        n13554) );
  AOI211_X1 U17110 ( .C1(n19089), .C2(n19940), .A(n13555), .B(n13554), .ZN(
        n13557) );
  NAND2_X1 U17111 ( .A1(n10645), .A2(n19109), .ZN(n13556) );
  OAI211_X1 U17112 ( .C1(n19938), .C2(n18958), .A(n13557), .B(n13556), .ZN(
        n13558) );
  AOI21_X1 U17113 ( .B1(n13559), .B2(n19154), .A(n13558), .ZN(n13560) );
  INV_X1 U17114 ( .A(n13560), .ZN(P2_U2853) );
  OR2_X1 U17115 ( .A1(n19354), .A2(n10593), .ZN(n19689) );
  NAND2_X1 U17116 ( .A1(n13038), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19607) );
  INV_X1 U17117 ( .A(n19607), .ZN(n19539) );
  NAND2_X1 U17118 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19539), .ZN(
        n13566) );
  OAI21_X1 U17119 ( .B1(n19689), .B2(n13742), .A(n13566), .ZN(n13565) );
  INV_X1 U17120 ( .A(n19407), .ZN(n13561) );
  NAND2_X1 U17121 ( .A1(n13561), .A2(n19539), .ZN(n19637) );
  AND2_X1 U17122 ( .A1(n19637), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13562) );
  AND2_X1 U17123 ( .A1(n19637), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13563) );
  NOR3_X1 U17124 ( .A1(n9793), .A2(n13569), .A3(n13563), .ZN(n13564) );
  NAND2_X1 U17125 ( .A1(n13565), .A2(n13564), .ZN(n19654) );
  INV_X1 U17126 ( .A(n19654), .ZN(n19641) );
  NAND2_X1 U17127 ( .A1(n16235), .A2(n19777), .ZN(n19760) );
  INV_X1 U17128 ( .A(n13566), .ZN(n13567) );
  AOI21_X1 U17129 ( .B1(n19951), .B2(n13567), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13568) );
  INV_X1 U17130 ( .A(n19819), .ZN(n13574) );
  INV_X1 U17131 ( .A(n19720), .ZN(n13571) );
  INV_X1 U17132 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n21113) );
  OAI22_X2 U17133 ( .A1(n21113), .A2(n19337), .B1(n14378), .B2(n19335), .ZN(
        n19821) );
  AOI22_X1 U17134 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19344), .B1(
        BUF1_REG_22__SCAN_IN), .B2(n19343), .ZN(n19824) );
  INV_X1 U17135 ( .A(n19824), .ZN(n19757) );
  AOI22_X1 U17136 ( .A1(n19653), .A2(n19821), .B1(n19681), .B2(n19757), .ZN(
        n13573) );
  OAI21_X1 U17137 ( .B1(n13574), .B2(n19637), .A(n13573), .ZN(n13575) );
  AOI21_X1 U17138 ( .B1(n19820), .B2(n19652), .A(n13575), .ZN(n13576) );
  OAI21_X1 U17139 ( .B1(n19641), .B2(n13577), .A(n13576), .ZN(P2_U3142) );
  NOR2_X2 U17140 ( .A1(n15288), .A2(n9793), .ZN(n19788) );
  NOR2_X2 U17141 ( .A1(n14294), .A2(n19339), .ZN(n19787) );
  INV_X1 U17142 ( .A(n19787), .ZN(n13579) );
  INV_X1 U17143 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16503) );
  INV_X1 U17144 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18271) );
  OAI22_X2 U17145 ( .A1(n16503), .A2(n19337), .B1(n18271), .B2(n19335), .ZN(
        n19789) );
  AOI22_X1 U17146 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19343), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19344), .ZN(n19792) );
  INV_X1 U17147 ( .A(n19792), .ZN(n19737) );
  AOI22_X1 U17148 ( .A1(n19653), .A2(n19789), .B1(n19681), .B2(n19737), .ZN(
        n13578) );
  OAI21_X1 U17149 ( .B1(n13579), .B2(n19637), .A(n13578), .ZN(n13580) );
  AOI21_X1 U17150 ( .B1(n19652), .B2(n19788), .A(n13580), .ZN(n13581) );
  OAI21_X1 U17151 ( .B1(n19641), .B2(n13582), .A(n13581), .ZN(P2_U3137) );
  XNOR2_X1 U17152 ( .A(n13584), .B(n13583), .ZN(n13609) );
  OAI211_X1 U17153 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n13586), .B(n13585), .ZN(n13592) );
  XNOR2_X1 U17154 ( .A(n13588), .B(n13587), .ZN(n19199) );
  INV_X1 U17155 ( .A(n19199), .ZN(n13590) );
  INV_X1 U17156 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13589) );
  NOR2_X1 U17157 ( .A1(n19131), .A2(n13589), .ZN(n13603) );
  AOI21_X1 U17158 ( .B1(n19301), .B2(n13590), .A(n13603), .ZN(n13591) );
  OAI211_X1 U17159 ( .C1(n19296), .C2(n19152), .A(n13592), .B(n13591), .ZN(
        n13593) );
  AOI21_X1 U17160 ( .B1(n13594), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13593), .ZN(n13601) );
  NAND2_X1 U17161 ( .A1(n13596), .A2(n13595), .ZN(n13606) );
  OAI21_X1 U17162 ( .B1(n13599), .B2(n13598), .A(n13597), .ZN(n13605) );
  NAND3_X1 U17163 ( .A1(n13606), .A2(n16337), .A3(n13605), .ZN(n13600) );
  OAI211_X1 U17164 ( .C1(n13609), .C2(n16369), .A(n13601), .B(n13600), .ZN(
        P2_U3041) );
  INV_X1 U17165 ( .A(n19152), .ZN(n13604) );
  INV_X1 U17166 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19159) );
  OAI21_X1 U17167 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13622), .A(
        n13621), .ZN(n19149) );
  OAI22_X1 U17168 ( .A1(n19288), .A2(n19159), .B1(n16314), .B2(n19149), .ZN(
        n13602) );
  AOI211_X1 U17169 ( .C1(n13604), .C2(n19278), .A(n13603), .B(n13602), .ZN(
        n13608) );
  NAND3_X1 U17170 ( .A1(n13606), .A2(n16310), .A3(n13605), .ZN(n13607) );
  OAI211_X1 U17171 ( .C1(n13609), .C2(n16292), .A(n13608), .B(n13607), .ZN(
        P2_U3009) );
  NOR2_X1 U17172 ( .A1(n19606), .A2(n19406), .ZN(n13611) );
  AOI221_X1 U17173 ( .B1(n19401), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19430), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n13611), .ZN(n13615) );
  INV_X1 U17174 ( .A(n13617), .ZN(n13612) );
  AOI21_X1 U17175 ( .B1(n13612), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U17176 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19958), .ZN(
        n19604) );
  NOR2_X1 U17177 ( .A1(n19604), .A2(n19406), .ZN(n19399) );
  NOR2_X1 U17178 ( .A1(n13613), .A2(n19399), .ZN(n13614) );
  INV_X1 U17179 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14158) );
  INV_X1 U17180 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n21083) );
  INV_X1 U17181 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18263) );
  OAI22_X2 U17182 ( .A1(n21083), .A2(n19337), .B1(n18263), .B2(n19335), .ZN(
        n19783) );
  AOI22_X1 U17183 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19344), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19343), .ZN(n19786) );
  INV_X1 U17184 ( .A(n19786), .ZN(n19727) );
  AOI22_X1 U17185 ( .A1(n19430), .A2(n19783), .B1(n19401), .B2(n19727), .ZN(
        n13620) );
  INV_X1 U17186 ( .A(n13616), .ZN(n19165) );
  NAND2_X1 U17187 ( .A1(n19165), .A2(n19777), .ZN(n19736) );
  OAI21_X1 U17188 ( .B1(n13617), .B2(n19399), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13618) );
  OAI21_X1 U17189 ( .B1(n19406), .B2(n19606), .A(n13618), .ZN(n19400) );
  NOR2_X2 U17190 ( .A1(n16397), .A2(n19339), .ZN(n19774) );
  AOI22_X1 U17191 ( .A1(n19775), .A2(n19400), .B1(n19774), .B2(n19399), .ZN(
        n13619) );
  OAI211_X1 U17192 ( .C1(n19405), .C2(n14158), .A(n13620), .B(n13619), .ZN(
        P2_U3064) );
  AOI21_X1 U17193 ( .B1(n16323), .B2(n13621), .A(n13639), .ZN(n16315) );
  AOI21_X1 U17194 ( .B1(n19287), .B2(n13623), .A(n13622), .ZN(n19273) );
  NAND2_X1 U17195 ( .A1(n13625), .A2(n13624), .ZN(n13654) );
  NOR2_X1 U17196 ( .A1(n19273), .A2(n13654), .ZN(n19146) );
  NAND2_X1 U17197 ( .A1(n19146), .A2(n19149), .ZN(n13636) );
  NAND2_X1 U17198 ( .A1(n19075), .A2(n13636), .ZN(n13626) );
  XNOR2_X1 U17199 ( .A(n16315), .B(n13626), .ZN(n13627) );
  NAND2_X1 U17200 ( .A1(n13627), .A2(n19154), .ZN(n13634) );
  INV_X1 U17201 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19870) );
  OAI21_X1 U17202 ( .B1(n19870), .B2(n19133), .A(n19131), .ZN(n13628) );
  AOI21_X1 U17203 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19138), .A(
        n13628), .ZN(n13629) );
  OAI21_X1 U17204 ( .B1(n19150), .B2(n15677), .A(n13629), .ZN(n13632) );
  NOR2_X1 U17205 ( .A1(n19142), .A2(n13630), .ZN(n13631) );
  AOI211_X1 U17206 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19128), .A(n13632), .B(
        n13631), .ZN(n13633) );
  OAI211_X1 U17207 ( .C1(n16316), .C2(n19151), .A(n13634), .B(n13633), .ZN(
        P2_U2849) );
  OAI21_X1 U17208 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13637), .A(
        n15027), .ZN(n16313) );
  NOR2_X1 U17209 ( .A1(n16315), .A2(n13636), .ZN(n19125) );
  OAI21_X1 U17210 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13639), .A(
        n13638), .ZN(n19127) );
  NAND2_X1 U17211 ( .A1(n19125), .A2(n19127), .ZN(n15024) );
  NAND2_X1 U17212 ( .A1(n19075), .A2(n15024), .ZN(n13640) );
  XOR2_X1 U17213 ( .A(n16313), .B(n13640), .Z(n13641) );
  NAND2_X1 U17214 ( .A1(n13641), .A2(n19154), .ZN(n13653) );
  INV_X1 U17215 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13650) );
  NAND2_X1 U17216 ( .A1(n13642), .A2(n19129), .ZN(n13649) );
  AOI21_X1 U17217 ( .B1(n13644), .B2(n13033), .A(n13643), .ZN(n13645) );
  INV_X1 U17218 ( .A(n13645), .ZN(n19189) );
  AOI22_X1 U17219 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19138), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19128), .ZN(n13646) );
  OAI211_X1 U17220 ( .C1(n19150), .C2(n19189), .A(n13646), .B(n19131), .ZN(
        n13647) );
  INV_X1 U17221 ( .A(n13647), .ZN(n13648) );
  OAI211_X1 U17222 ( .C1(n19133), .C2(n13650), .A(n13649), .B(n13648), .ZN(
        n13651) );
  AOI21_X1 U17223 ( .B1(n16338), .B2(n19109), .A(n13651), .ZN(n13652) );
  NAND2_X1 U17224 ( .A1(n13653), .A2(n13652), .ZN(P2_U2847) );
  AND2_X1 U17225 ( .A1(n19075), .A2(n13654), .ZN(n13656) );
  AOI21_X1 U17226 ( .B1(n19273), .B2(n13656), .A(n19840), .ZN(n13655) );
  OAI21_X1 U17227 ( .B1(n19273), .B2(n13656), .A(n13655), .ZN(n13664) );
  INV_X1 U17228 ( .A(n19133), .ZN(n19145) );
  AOI22_X1 U17229 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19138), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19128), .ZN(n13657) );
  OAI211_X1 U17230 ( .C1(n19150), .C2(n13658), .A(n13657), .B(n19131), .ZN(
        n13659) );
  AOI21_X1 U17231 ( .B1(n19145), .B2(P2_REIP_REG_4__SCAN_IN), .A(n13659), .ZN(
        n13660) );
  OAI21_X1 U17232 ( .B1(n13661), .B2(n19142), .A(n13660), .ZN(n13662) );
  AOI21_X1 U17233 ( .B1(n19279), .B2(n19109), .A(n13662), .ZN(n13663) );
  OAI211_X1 U17234 ( .C1(n18958), .C2(n19193), .A(n13664), .B(n13663), .ZN(
        P2_U2851) );
  NAND2_X1 U17235 ( .A1(n13669), .A2(n11773), .ZN(n13665) );
  NAND2_X1 U17236 ( .A1(n15945), .A2(n13665), .ZN(n20091) );
  INV_X1 U17237 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20796) );
  AOI22_X1 U17238 ( .A1(n20796), .A2(n20084), .B1(n20056), .B2(n13666), .ZN(
        n13676) );
  NAND2_X1 U17239 ( .A1(n20081), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n13674) );
  INV_X1 U17240 ( .A(n13667), .ZN(n13668) );
  NAND2_X1 U17241 ( .A1(n13669), .A2(n13668), .ZN(n20072) );
  INV_X1 U17242 ( .A(n20072), .ZN(n20089) );
  NAND2_X1 U17243 ( .A1(n20089), .A2(n20678), .ZN(n13673) );
  INV_X1 U17244 ( .A(n20079), .ZN(n13670) );
  AOI22_X1 U17245 ( .A1(n20087), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13670), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13672) );
  NAND2_X1 U17246 ( .A1(n20086), .A2(n20170), .ZN(n13671) );
  AND4_X1 U17247 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13675) );
  OAI211_X1 U17248 ( .C1(n14545), .C2(n20174), .A(n13676), .B(n13675), .ZN(
        P1_U2839) );
  NAND2_X1 U17249 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n13677) );
  OR2_X1 U17250 ( .A1(n20080), .A2(n13677), .ZN(n20073) );
  INV_X1 U17251 ( .A(n20073), .ZN(n13688) );
  OAI221_X1 U17252 ( .B1(n20080), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n20080), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n20079), .ZN(n13678) );
  AOI22_X1 U17253 ( .A1(n20087), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13678), .ZN(n13682) );
  INV_X1 U17254 ( .A(n13679), .ZN(n13680) );
  NAND2_X1 U17255 ( .A1(n20086), .A2(n13680), .ZN(n13681) );
  OAI211_X1 U17256 ( .C1(n20098), .C2(n13683), .A(n13682), .B(n13681), .ZN(
        n13686) );
  INV_X1 U17257 ( .A(n20476), .ZN(n20850) );
  OAI22_X1 U17258 ( .A1(n13684), .A2(n20043), .B1(n20072), .B2(n20850), .ZN(
        n13685) );
  AOI211_X1 U17259 ( .C1(n13688), .C2(n13687), .A(n13686), .B(n13685), .ZN(
        n13689) );
  OAI21_X1 U17260 ( .B1(n14545), .B2(n13690), .A(n13689), .ZN(P1_U2837) );
  NOR2_X1 U17261 ( .A1(n13487), .A2(n13692), .ZN(n13693) );
  OR2_X1 U17262 ( .A1(n13691), .A2(n13693), .ZN(n20017) );
  INV_X1 U17263 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13699) );
  NAND2_X1 U17264 ( .A1(n13695), .A2(n13694), .ZN(n13697) );
  NAND2_X1 U17265 ( .A1(n13697), .A2(n13696), .ZN(n13698) );
  NAND2_X1 U17266 ( .A1(n13698), .A2(n13721), .ZN(n20020) );
  OAI222_X1 U17267 ( .A1(n20017), .A2(n14627), .B1(n13699), .B2(n14626), .C1(
        n20020), .C2(n14608), .ZN(P1_U2863) );
  INV_X1 U17268 ( .A(DATAI_9_), .ZN(n13700) );
  MUX2_X1 U17269 ( .A(n13700), .B(n16525), .S(n14628), .Z(n20128) );
  INV_X1 U17270 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13701) );
  OAI222_X1 U17271 ( .A1(n20017), .A2(n14708), .B1(n20128), .B2(n14706), .C1(
        n13701), .C2(n14704), .ZN(P1_U2895) );
  NAND2_X1 U17272 ( .A1(n19147), .A2(n19154), .ZN(n19102) );
  OAI211_X1 U17273 ( .C1(n15115), .C2(n13703), .A(n19075), .B(n13702), .ZN(
        n15716) );
  OAI22_X1 U17274 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19102), .B1(
        n15716), .B2(n19840), .ZN(n13704) );
  INV_X1 U17275 ( .A(n13704), .ZN(n13714) );
  OAI22_X1 U17276 ( .A1(n19143), .A2(n13706), .B1(n13705), .B2(n19158), .ZN(
        n13707) );
  AOI21_X1 U17277 ( .B1(n19145), .B2(P2_REIP_REG_1__SCAN_IN), .A(n13707), .ZN(
        n13709) );
  NAND2_X1 U17278 ( .A1(n19089), .A2(n19948), .ZN(n13708) );
  OAI211_X1 U17279 ( .C1(n19142), .C2(n13710), .A(n13709), .B(n13708), .ZN(
        n13711) );
  AOI21_X1 U17280 ( .B1(n19109), .B2(n13712), .A(n13711), .ZN(n13713) );
  OAI211_X1 U17281 ( .C1(n13715), .C2(n18958), .A(n13714), .B(n13713), .ZN(
        P2_U2854) );
  OR2_X1 U17282 ( .A1(n13691), .A2(n13717), .ZN(n13718) );
  NAND2_X1 U17283 ( .A1(n13716), .A2(n13718), .ZN(n14864) );
  INV_X1 U17284 ( .A(n13719), .ZN(n14861) );
  NAND2_X1 U17285 ( .A1(n13721), .A2(n13720), .ZN(n13722) );
  NAND2_X1 U17286 ( .A1(n13772), .A2(n13722), .ZN(n16097) );
  AOI21_X1 U17287 ( .B1(n20087), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20069), .ZN(n13726) );
  INV_X1 U17288 ( .A(n14480), .ZN(n13723) );
  NOR2_X1 U17289 ( .A1(n14525), .A2(n13723), .ZN(n13724) );
  OR2_X1 U17290 ( .A1(n13724), .A2(n20062), .ZN(n14529) );
  INV_X1 U17291 ( .A(n14529), .ZN(n15981) );
  AOI22_X1 U17292 ( .A1(n15981), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_EBX_REG_10__SCAN_IN), .B2(n20081), .ZN(n13725) );
  OAI211_X1 U17293 ( .C1(n20098), .C2(n16097), .A(n13726), .B(n13725), .ZN(
        n13729) );
  INV_X1 U17294 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20806) );
  NAND2_X1 U17295 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .ZN(n13727) );
  INV_X1 U17296 ( .A(n20027), .ZN(n14524) );
  NOR3_X1 U17297 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20806), .A3(n14524), 
        .ZN(n13728) );
  AOI211_X1 U17298 ( .C1(n20086), .C2(n14861), .A(n13729), .B(n13728), .ZN(
        n13730) );
  OAI21_X1 U17299 ( .B1(n15945), .B2(n14864), .A(n13730), .ZN(P1_U2830) );
  XNOR2_X1 U17300 ( .A(n13732), .B(n13731), .ZN(n13733) );
  XNOR2_X1 U17301 ( .A(n13734), .B(n13733), .ZN(n16119) );
  NAND2_X1 U17302 ( .A1(n16119), .A2(n20169), .ZN(n13740) );
  INV_X1 U17303 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13735) );
  NOR2_X1 U17304 ( .A1(n20208), .A2(n13735), .ZN(n16110) );
  NOR2_X1 U17305 ( .A1(n14805), .A2(n13736), .ZN(n13737) );
  AOI211_X1 U17306 ( .C1(n20171), .C2(n13738), .A(n16110), .B(n13737), .ZN(
        n13739) );
  OAI211_X1 U17307 ( .C1(n20175), .C2(n13741), .A(n13740), .B(n13739), .ZN(
        P1_U2991) );
  OAI21_X1 U17308 ( .B1(n19449), .B2(n19475), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13747) );
  NOR2_X1 U17309 ( .A1(n13744), .A2(n13743), .ZN(n19657) );
  NAND2_X1 U17310 ( .A1(n19657), .A2(n19935), .ZN(n13750) );
  INV_X1 U17311 ( .A(n13745), .ZN(n13748) );
  NAND3_X1 U17312 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19935), .A3(
        n19950), .ZN(n19458) );
  NOR2_X1 U17313 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19458), .ZN(
        n19447) );
  AOI211_X1 U17314 ( .C1(n13748), .C2(n19951), .A(n19447), .B(n19924), .ZN(
        n13746) );
  OAI21_X1 U17315 ( .B1(n13748), .B2(n19447), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13749) );
  INV_X1 U17316 ( .A(n19447), .ZN(n13755) );
  AOI22_X1 U17317 ( .A1(n19475), .A2(n19813), .B1(n19449), .B2(n19753), .ZN(
        n13751) );
  OAI21_X1 U17318 ( .B1(n19370), .B2(n13755), .A(n13751), .ZN(n13752) );
  AOI21_X1 U17319 ( .B1(n19448), .B2(n19812), .A(n13752), .ZN(n13753) );
  OAI21_X1 U17320 ( .B1(n19452), .B2(n14296), .A(n13753), .ZN(P2_U3085) );
  INV_X1 U17321 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13759) );
  INV_X1 U17322 ( .A(n19774), .ZN(n13756) );
  AOI22_X1 U17323 ( .A1(n19475), .A2(n19783), .B1(n19449), .B2(n19727), .ZN(
        n13754) );
  OAI21_X1 U17324 ( .B1(n13756), .B2(n13755), .A(n13754), .ZN(n13757) );
  AOI21_X1 U17325 ( .B1(n19775), .B2(n19448), .A(n13757), .ZN(n13758) );
  OAI21_X1 U17326 ( .B1(n19452), .B2(n13759), .A(n13758), .ZN(P2_U3080) );
  INV_X1 U17327 ( .A(DATAI_10_), .ZN(n13760) );
  MUX2_X1 U17328 ( .A(n13760), .B(n16523), .S(n14628), .Z(n20131) );
  INV_X1 U17329 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13761) );
  OAI222_X1 U17330 ( .A1(n14864), .A2(n14708), .B1(n20131), .B2(n14706), .C1(
        n13761), .C2(n14704), .ZN(P1_U2894) );
  INV_X1 U17331 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13762) );
  OAI222_X1 U17332 ( .A1(n16097), .A2(n14608), .B1(n14626), .B2(n13762), .C1(
        n14864), .C2(n14627), .ZN(P1_U2862) );
  MUX2_X1 U17333 ( .A(n13764), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n16013), .Z(n13765) );
  XNOR2_X1 U17334 ( .A(n13763), .B(n13765), .ZN(n16103) );
  OAI22_X1 U17335 ( .A1(n14805), .A2(n20024), .B1(n20208), .B2(n20806), .ZN(
        n13767) );
  NOR2_X1 U17336 ( .A1(n20017), .A2(n20175), .ZN(n13766) );
  AOI211_X1 U17337 ( .C1(n20171), .C2(n20018), .A(n13767), .B(n13766), .ZN(
        n13768) );
  OAI21_X1 U17338 ( .B1(n16103), .B2(n19999), .A(n13768), .ZN(P1_U2990) );
  NAND2_X1 U17339 ( .A1(n13716), .A2(n13770), .ZN(n13771) );
  NAND2_X1 U17340 ( .A1(n13769), .A2(n13771), .ZN(n14521) );
  XOR2_X1 U17341 ( .A(n14520), .B(n14521), .Z(n16018) );
  INV_X1 U17342 ( .A(n16018), .ZN(n13776) );
  AOI21_X1 U17343 ( .B1(n13773), .B2(n13772), .A(n14623), .ZN(n16083) );
  AOI22_X1 U17344 ( .A1(n14614), .A2(n16083), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14612), .ZN(n13774) );
  OAI21_X1 U17345 ( .B1(n13776), .B2(n14627), .A(n13774), .ZN(P1_U2861) );
  OAI222_X1 U17346 ( .A1(n13776), .A2(n14708), .B1(n14643), .B2(n14706), .C1(
        n13775), .C2(n14704), .ZN(P1_U2893) );
  NAND2_X1 U17347 ( .A1(n13777), .A2(n11758), .ZN(n13782) );
  NAND2_X1 U17348 ( .A1(n11758), .A2(n15880), .ZN(n13778) );
  NAND4_X1 U17349 ( .A1(n13779), .A2(n14392), .A3(n20880), .A4(n13778), .ZN(
        n13780) );
  OAI211_X1 U17350 ( .C1(n14388), .C2(n13782), .A(n13781), .B(n13780), .ZN(
        n13783) );
  NAND2_X1 U17351 ( .A1(n13783), .A2(n14397), .ZN(n13791) );
  NAND3_X1 U17352 ( .A1(n15858), .A2(n20880), .A3(n13785), .ZN(n13787) );
  NAND3_X1 U17353 ( .A1(n13787), .A2(n13794), .A3(n13786), .ZN(n13788) );
  NAND3_X1 U17354 ( .A1(n13789), .A2(n13784), .A3(n13788), .ZN(n13790) );
  NOR2_X1 U17355 ( .A1(n20164), .A2(n13832), .ZN(n20220) );
  OAI211_X1 U17356 ( .C1(n13795), .C2(n13794), .A(n13793), .B(n13792), .ZN(
        n13796) );
  NOR2_X1 U17357 ( .A1(n13797), .A2(n13796), .ZN(n13799) );
  AND2_X1 U17358 ( .A1(n13799), .A2(n13798), .ZN(n13803) );
  INV_X1 U17359 ( .A(n13803), .ZN(n13800) );
  NAND2_X1 U17360 ( .A1(n13832), .A2(n13800), .ZN(n14973) );
  NOR2_X1 U17361 ( .A1(n14973), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20227) );
  NAND2_X1 U17362 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20176) );
  NOR2_X1 U17363 ( .A1(n13801), .A2(n20176), .ZN(n16117) );
  NAND3_X1 U17364 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n16117), .ZN(n16091) );
  AND2_X1 U17365 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16123) );
  NAND4_X1 U17366 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16123), .ZN(n13805) );
  NOR2_X1 U17367 ( .A1(n16091), .A2(n13805), .ZN(n16074) );
  NOR3_X1 U17368 ( .A1(n16089), .A2(n12770), .A3(n16081), .ZN(n13949) );
  NAND2_X1 U17369 ( .A1(n13803), .A2(n13802), .ZN(n13804) );
  NAND2_X1 U17370 ( .A1(n13832), .A2(n13804), .ZN(n13946) );
  AOI21_X1 U17371 ( .B1(n16074), .B2(n13949), .A(n13946), .ZN(n13807) );
  INV_X1 U17372 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20233) );
  OAI21_X1 U17373 ( .B1(n20233), .B2(n20219), .A(n20204), .ZN(n20194) );
  NAND2_X1 U17374 ( .A1(n16117), .A2(n20194), .ZN(n16134) );
  NOR2_X1 U17375 ( .A1(n13805), .A2(n16134), .ZN(n16086) );
  AND2_X1 U17376 ( .A1(n13949), .A2(n16086), .ZN(n13833) );
  NOR2_X1 U17377 ( .A1(n16116), .A2(n13833), .ZN(n13806) );
  NOR2_X1 U17378 ( .A1(n13807), .A2(n13806), .ZN(n13808) );
  INV_X1 U17379 ( .A(n16082), .ZN(n14977) );
  NOR2_X1 U17380 ( .A1(n20208), .A2(n13809), .ZN(n13830) );
  AND2_X1 U17381 ( .A1(n13810), .A2(n13811), .ZN(n14821) );
  INV_X1 U17382 ( .A(n13812), .ZN(n13814) );
  OAI21_X1 U17383 ( .B1(n14821), .B2(n13814), .A(n13813), .ZN(n13816) );
  XNOR2_X1 U17384 ( .A(n16013), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13815) );
  XNOR2_X1 U17385 ( .A(n13816), .B(n13815), .ZN(n16007) );
  INV_X1 U17386 ( .A(n13817), .ZN(n13821) );
  OAI21_X1 U17387 ( .B1(n13825), .B2(n20249), .A(n13818), .ZN(n13819) );
  NOR2_X1 U17388 ( .A1(n15847), .A2(n13819), .ZN(n13820) );
  NAND2_X1 U17389 ( .A1(n13821), .A2(n13820), .ZN(n13822) );
  OAI21_X1 U17390 ( .B1(n13825), .B2(n13824), .A(n13823), .ZN(n13826) );
  NAND2_X1 U17391 ( .A1(n9897), .A2(n13827), .ZN(n13828) );
  NAND2_X1 U17392 ( .A1(n14512), .A2(n13828), .ZN(n15961) );
  OAI22_X1 U17393 ( .A1(n16007), .A2(n16049), .B1(n20224), .B2(n15961), .ZN(
        n13829) );
  AOI211_X1 U17394 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n14977), .A(
        n13830), .B(n13829), .ZN(n13835) );
  NAND2_X1 U17395 ( .A1(n13832), .A2(n13831), .ZN(n20231) );
  NAND2_X1 U17396 ( .A1(n20233), .A2(n20231), .ZN(n20207) );
  NAND2_X1 U17397 ( .A1(n16114), .A2(n20207), .ZN(n20193) );
  NOR3_X1 U17398 ( .A1(n20204), .A2(n20219), .A3(n20193), .ZN(n16118) );
  INV_X1 U17399 ( .A(n16135), .ZN(n16142) );
  NAND3_X1 U17400 ( .A1(n16142), .A2(n21132), .A3(n13833), .ZN(n13834) );
  NAND2_X1 U17401 ( .A1(n13835), .A2(n13834), .ZN(P1_U3017) );
  AND2_X1 U17402 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16996) );
  NOR2_X2 U17403 ( .A1(n18730), .A2(n13838), .ZN(n15791) );
  NAND2_X1 U17404 ( .A1(n18297), .A2(n17284), .ZN(n17278) );
  INV_X2 U17405 ( .A(n17281), .ZN(n17275) );
  INV_X1 U17406 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17283) );
  INV_X1 U17407 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17277) );
  NOR2_X1 U17408 ( .A1(n17283), .A2(n17277), .ZN(n17271) );
  AND2_X1 U17409 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17271), .ZN(n17262) );
  NAND3_X1 U17410 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17262), .ZN(n15772) );
  NOR2_X2 U17411 ( .A1(n13841), .A2(n15772), .ZN(n17258) );
  NAND3_X1 U17412 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .ZN(n15771) );
  INV_X1 U17413 ( .A(n15771), .ZN(n13842) );
  NOR3_X2 U17414 ( .A1(n17227), .A2(n16823), .A3(n17208), .ZN(n17189) );
  AND2_X1 U17415 ( .A1(n18297), .A2(n17083), .ZN(n17066) );
  NAND2_X1 U17416 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17027), .ZN(n17014) );
  NAND2_X1 U17417 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17017), .ZN(n17008) );
  NAND2_X1 U17418 ( .A1(n17275), .A2(n17008), .ZN(n17006) );
  OAI21_X1 U17419 ( .B1(n16996), .B2(n17278), .A(n17006), .ZN(n17000) );
  AOI22_X1 U17420 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13843) );
  OAI21_X1 U17421 ( .B1(n9842), .B2(n17264), .A(n13843), .ZN(n13853) );
  AOI22_X1 U17422 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13850) );
  OAI22_X1 U17423 ( .A1(n11037), .A2(n18500), .B1(n17072), .B2(n17170), .ZN(
        n13848) );
  AOI22_X1 U17424 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17425 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U17426 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13844) );
  NAND3_X1 U17427 ( .A1(n13846), .A2(n13845), .A3(n13844), .ZN(n13847) );
  AOI211_X1 U17428 ( .C1(n9806), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n13848), .B(n13847), .ZN(n13849) );
  OAI211_X1 U17429 ( .C1(n17177), .C2(n13851), .A(n13850), .B(n13849), .ZN(
        n13852) );
  AOI211_X1 U17430 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n13853), .B(n13852), .ZN(n17004) );
  AOI22_X1 U17431 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13854) );
  OAI21_X1 U17432 ( .B1(n17072), .B2(n17193), .A(n13854), .ZN(n13864) );
  INV_X1 U17433 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13862) );
  AOI22_X1 U17434 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13861) );
  AOI22_X1 U17435 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13855) );
  OAI21_X1 U17436 ( .B1(n11037), .B2(n18494), .A(n13855), .ZN(n13859) );
  INV_X1 U17437 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18598) );
  AOI22_X1 U17438 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13857) );
  AOI22_X1 U17439 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17235), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13856) );
  OAI211_X1 U17440 ( .C1(n17246), .C2(n18598), .A(n13857), .B(n13856), .ZN(
        n13858) );
  AOI211_X1 U17441 ( .C1(n17216), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n13859), .B(n13858), .ZN(n13860) );
  OAI211_X1 U17442 ( .C1(n10244), .C2(n13862), .A(n13861), .B(n13860), .ZN(
        n13863) );
  AOI211_X1 U17443 ( .C1(n11226), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n13864), .B(n13863), .ZN(n17015) );
  AOI22_X1 U17444 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13865) );
  OAI21_X1 U17445 ( .B1(n17151), .B2(n21045), .A(n13865), .ZN(n13874) );
  AOI22_X1 U17446 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U17447 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13866) );
  OAI21_X1 U17448 ( .B1(n11037), .B2(n18489), .A(n13866), .ZN(n13870) );
  AOI22_X1 U17449 ( .A1(n11011), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13868) );
  AOI22_X1 U17450 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13867) );
  OAI211_X1 U17451 ( .C1(n17246), .C2(n18593), .A(n13868), .B(n13867), .ZN(
        n13869) );
  AOI211_X1 U17452 ( .C1(n17216), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n13870), .B(n13869), .ZN(n13871) );
  OAI211_X1 U17453 ( .C1(n11054), .C2(n18304), .A(n13872), .B(n13871), .ZN(
        n13873) );
  AOI211_X1 U17454 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n13874), .B(n13873), .ZN(n17025) );
  AOI22_X1 U17455 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17105), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13875) );
  OAI21_X1 U17456 ( .B1(n10227), .B2(n18618), .A(n13875), .ZN(n13884) );
  AOI22_X1 U17457 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n9812), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13882) );
  INV_X1 U17458 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21080) );
  AOI22_X1 U17459 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9801), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13876) );
  OAI21_X1 U17460 ( .B1(n21080), .B2(n11037), .A(n13876), .ZN(n13880) );
  AOI22_X1 U17461 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13878) );
  AOI22_X1 U17462 ( .A1(n17236), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n11051), .ZN(n13877) );
  OAI211_X1 U17463 ( .C1(n16981), .C2(n11056), .A(n13878), .B(n13877), .ZN(
        n13879) );
  AOI211_X1 U17464 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n13880), .B(n13879), .ZN(n13881) );
  OAI211_X1 U17465 ( .C1(n11054), .C2(n17252), .A(n13882), .B(n13881), .ZN(
        n13883) );
  AOI211_X1 U17466 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n13884), .B(n13883), .ZN(n17024) );
  NOR2_X1 U17467 ( .A1(n17025), .A2(n17024), .ZN(n17020) );
  AOI22_X1 U17468 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U17469 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U17470 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13892) );
  OAI22_X1 U17471 ( .A1(n11037), .A2(n20981), .B1(n17246), .B2(n21111), .ZN(
        n13890) );
  AOI22_X1 U17472 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U17473 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13887) );
  AOI22_X1 U17474 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13886) );
  NAND2_X1 U17475 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13885) );
  NAND4_X1 U17476 ( .A1(n13888), .A2(n13887), .A3(n13886), .A4(n13885), .ZN(
        n13889) );
  AOI211_X1 U17477 ( .C1(n17195), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n13890), .B(n13889), .ZN(n13891) );
  NAND4_X1 U17478 ( .A1(n13894), .A2(n13893), .A3(n13892), .A4(n13891), .ZN(
        n17019) );
  NAND2_X1 U17479 ( .A1(n17020), .A2(n17019), .ZN(n17018) );
  NOR2_X1 U17480 ( .A1(n17015), .A2(n17018), .ZN(n17011) );
  AOI22_X1 U17481 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13904) );
  AOI22_X1 U17482 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13903) );
  AOI22_X1 U17483 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13902) );
  OAI22_X1 U17484 ( .A1(n11037), .A2(n18497), .B1(n9841), .B2(n17176), .ZN(
        n13900) );
  AOI22_X1 U17485 ( .A1(n9801), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13898) );
  AOI22_X1 U17486 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17487 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13896) );
  NAND2_X1 U17488 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n13895) );
  NAND4_X1 U17489 ( .A1(n13898), .A2(n13897), .A3(n13896), .A4(n13895), .ZN(
        n13899) );
  AOI211_X1 U17490 ( .C1(n17236), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n13900), .B(n13899), .ZN(n13901) );
  NAND4_X1 U17491 ( .A1(n13904), .A2(n13903), .A3(n13902), .A4(n13901), .ZN(
        n17010) );
  NAND2_X1 U17492 ( .A1(n17011), .A2(n17010), .ZN(n17009) );
  NOR2_X1 U17493 ( .A1(n17004), .A2(n17009), .ZN(n17003) );
  AOI22_X1 U17494 ( .A1(n17236), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13916) );
  AOI22_X1 U17495 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U17496 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13907) );
  OAI211_X1 U17497 ( .C1(n11056), .C2(n21130), .A(n13908), .B(n13907), .ZN(
        n13914) );
  AOI22_X1 U17498 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U17499 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U17500 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13910) );
  NAND2_X1 U17501 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13909) );
  NAND4_X1 U17502 ( .A1(n13912), .A2(n13911), .A3(n13910), .A4(n13909), .ZN(
        n13913) );
  AOI211_X1 U17503 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n13914), .B(n13913), .ZN(n13915) );
  OAI211_X1 U17504 ( .C1(n11054), .C2(n15760), .A(n13916), .B(n13915), .ZN(
        n16997) );
  XOR2_X1 U17505 ( .A(n17003), .B(n16997), .Z(n17299) );
  AOI22_X1 U17506 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17000), .B1(n17281), 
        .B2(n17299), .ZN(n13919) );
  INV_X1 U17507 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n13917) );
  INV_X1 U17508 ( .A(n17008), .ZN(n17013) );
  NAND3_X1 U17509 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n13917), .A3(n17013), 
        .ZN(n13918) );
  NAND2_X1 U17510 ( .A1(n13919), .A2(n13918), .ZN(P3_U2675) );
  NAND2_X1 U17511 ( .A1(n14021), .A2(n14017), .ZN(n13926) );
  NAND2_X1 U17512 ( .A1(n13923), .A2(n13922), .ZN(n14023) );
  NAND2_X1 U17513 ( .A1(n14024), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13924) );
  AOI21_X1 U17514 ( .B1(n15056), .B2(n10931), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14020) );
  INV_X1 U17515 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14039) );
  NOR2_X1 U17516 ( .A1(n14020), .A2(n9855), .ZN(n13925) );
  XNOR2_X1 U17517 ( .A(n13926), .B(n13925), .ZN(n15305) );
  AOI22_X1 U17518 ( .A1(n14030), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n13928) );
  NAND2_X1 U17519 ( .A1(n14031), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13927) );
  OAI211_X1 U17520 ( .C1(n10424), .C2(n14039), .A(n13928), .B(n13927), .ZN(
        n13929) );
  AOI211_X1 U17521 ( .C1(n16364), .C2(n13932), .A(n14039), .B(n14001), .ZN(
        n14048) );
  AOI21_X1 U17522 ( .B1(n14051), .B2(n14049), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13933) );
  NOR2_X1 U17523 ( .A1(n14048), .A2(n13933), .ZN(n13943) );
  AOI22_X1 U17524 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n13936) );
  NAND2_X1 U17525 ( .A1(n14043), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13935) );
  NAND2_X1 U17526 ( .A1(n13936), .A2(n13935), .ZN(n13938) );
  NAND2_X1 U17527 ( .A1(n13937), .A2(n13938), .ZN(n14047) );
  INV_X1 U17528 ( .A(n13937), .ZN(n13940) );
  INV_X1 U17529 ( .A(n13938), .ZN(n13939) );
  NAND2_X1 U17530 ( .A1(n13940), .A2(n13939), .ZN(n13941) );
  NAND2_X1 U17531 ( .A1(n19088), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15298) );
  OAI21_X1 U17532 ( .B1(n16360), .B2(n15054), .A(n15298), .ZN(n13942) );
  XNOR2_X1 U17533 ( .A(n14040), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15302) );
  NAND2_X1 U17534 ( .A1(n15302), .A2(n16337), .ZN(n13944) );
  OAI211_X1 U17535 ( .C1(n15305), .C2(n16369), .A(n13945), .B(n13944), .ZN(
        P2_U3016) );
  NAND2_X1 U17536 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13951) );
  NOR2_X1 U17537 ( .A1(n14990), .A2(n14992), .ZN(n16057) );
  NAND2_X1 U17538 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n16057), .ZN(
        n16047) );
  INV_X1 U17539 ( .A(n16047), .ZN(n14949) );
  NAND3_X1 U17540 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n14949), .ZN(n14978) );
  NOR3_X1 U17541 ( .A1(n14970), .A2(n16045), .A3(n14978), .ZN(n13952) );
  NAND2_X1 U17542 ( .A1(n16082), .A2(n13952), .ZN(n13947) );
  NAND2_X1 U17543 ( .A1(n20218), .A2(n20215), .ZN(n13948) );
  AOI21_X1 U17544 ( .B1(n16095), .B2(n13951), .A(n14963), .ZN(n14927) );
  OAI21_X1 U17545 ( .B1(n14928), .B2(n20215), .A(n14927), .ZN(n14922) );
  NAND2_X1 U17546 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13955) );
  NOR2_X1 U17547 ( .A1(n14922), .A2(n13955), .ZN(n14887) );
  INV_X1 U17548 ( .A(n13948), .ZN(n14886) );
  AOI21_X1 U17549 ( .B1(n14887), .B2(n14888), .A(n14886), .ZN(n14883) );
  AOI211_X1 U17550 ( .C1(n14877), .C2(n16095), .A(n12784), .B(n14883), .ZN(
        n14869) );
  NOR3_X1 U17551 ( .A1(n14869), .A2(n14886), .A3(n12787), .ZN(n13958) );
  NAND2_X1 U17552 ( .A1(n20206), .A2(n16086), .ZN(n14972) );
  INV_X1 U17553 ( .A(n13949), .ZN(n13950) );
  INV_X1 U17554 ( .A(n16074), .ZN(n15000) );
  NOR2_X1 U17555 ( .A1(n15000), .A2(n20193), .ZN(n14998) );
  NAND2_X1 U17556 ( .A1(n14998), .A2(n13949), .ZN(n14929) );
  OAI21_X1 U17557 ( .B1(n14972), .B2(n13950), .A(n14929), .ZN(n14948) );
  INV_X1 U17558 ( .A(n13951), .ZN(n14951) );
  AND2_X1 U17559 ( .A1(n13952), .A2(n14951), .ZN(n13953) );
  NAND2_X1 U17560 ( .A1(n14948), .A2(n13953), .ZN(n14937) );
  INV_X1 U17561 ( .A(n14928), .ZN(n13954) );
  NOR2_X1 U17562 ( .A1(n14909), .A2(n13955), .ZN(n14899) );
  NAND3_X1 U17563 ( .A1(n14899), .A2(n14888), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14870) );
  NOR3_X1 U17564 ( .A1(n14870), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12784), .ZN(n13956) );
  NAND2_X1 U17565 ( .A1(n13964), .A2(n13962), .ZN(n13960) );
  NAND2_X1 U17566 ( .A1(n10248), .A2(n13961), .ZN(n13990) );
  INV_X1 U17567 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14002) );
  AOI21_X1 U17568 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(n13965) );
  NOR2_X1 U17569 ( .A1(n13989), .A2(n13965), .ZN(n13968) );
  XOR2_X1 U17570 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n13966), .Z(
        n13967) );
  XNOR2_X1 U17571 ( .A(n13968), .B(n13967), .ZN(n13988) );
  XNOR2_X1 U17572 ( .A(n9840), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13986) );
  AOI21_X1 U17573 ( .B1(n13969), .B2(n13998), .A(n9852), .ZN(n15059) );
  INV_X1 U17574 ( .A(n15059), .ZN(n15134) );
  AOI21_X1 U17575 ( .B1(n13970), .B2(n9857), .A(n11541), .ZN(n15233) );
  INV_X1 U17576 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19907) );
  NOR2_X1 U17577 ( .A1(n19131), .A2(n19907), .ZN(n13982) );
  NOR3_X1 U17578 ( .A1(n13973), .A2(n13972), .A3(n13971), .ZN(n13974) );
  AOI211_X1 U17579 ( .C1(n19301), .C2(n15233), .A(n13982), .B(n13974), .ZN(
        n13976) );
  NAND2_X1 U17580 ( .A1(n14001), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13975) );
  OAI211_X1 U17581 ( .C1(n15134), .C2(n19296), .A(n13976), .B(n13975), .ZN(
        n13977) );
  AOI21_X1 U17582 ( .B1(n13986), .B2(n16337), .A(n13977), .ZN(n13978) );
  OAI21_X1 U17583 ( .B1(n13988), .B2(n16369), .A(n13978), .ZN(P2_U3018) );
  NAND2_X1 U17584 ( .A1(n14008), .A2(n13979), .ZN(n13980) );
  NAND2_X1 U17585 ( .A1(n13981), .A2(n13980), .ZN(n15063) );
  NAND2_X1 U17586 ( .A1(n15059), .A2(n19278), .ZN(n13984) );
  AOI21_X1 U17587 ( .B1(n16299), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n13982), .ZN(n13983) );
  OAI211_X1 U17588 ( .C1(n16314), .C2(n15063), .A(n13984), .B(n13983), .ZN(
        n13985) );
  AOI21_X1 U17589 ( .B1(n13986), .B2(n16287), .A(n13985), .ZN(n13987) );
  OAI21_X1 U17590 ( .B1(n13988), .B2(n16292), .A(n13987), .ZN(P2_U2986) );
  NAND2_X1 U17591 ( .A1(n13990), .A2(n14002), .ZN(n14007) );
  NAND2_X1 U17592 ( .A1(n14007), .A2(n19303), .ZN(n14006) );
  NAND2_X1 U17593 ( .A1(n13991), .A2(n13992), .ZN(n13993) );
  NAND2_X1 U17594 ( .A1(n9857), .A2(n13993), .ZN(n16189) );
  INV_X1 U17595 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19906) );
  NOR2_X1 U17596 ( .A1(n19131), .A2(n19906), .ZN(n14009) );
  AOI21_X1 U17597 ( .B1(n14002), .B2(n14049), .A(n14009), .ZN(n13994) );
  OAI21_X1 U17598 ( .B1(n16360), .B2(n16189), .A(n13994), .ZN(n14000) );
  NAND2_X1 U17599 ( .A1(n15144), .A2(n13996), .ZN(n13997) );
  NAND2_X1 U17600 ( .A1(n13998), .A2(n13997), .ZN(n16190) );
  NOR2_X1 U17601 ( .A1(n16190), .A2(n19296), .ZN(n13999) );
  AOI211_X1 U17602 ( .C1(n14001), .C2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14000), .B(n13999), .ZN(n14005) );
  INV_X1 U17603 ( .A(n15310), .ZN(n14003) );
  NAND2_X1 U17604 ( .A1(n14003), .A2(n14002), .ZN(n14013) );
  NAND3_X1 U17605 ( .A1(n14013), .A2(n16337), .A3(n9840), .ZN(n14004) );
  OAI211_X1 U17606 ( .C1(n13989), .C2(n14006), .A(n14005), .B(n14004), .ZN(
        P2_U3019) );
  NAND2_X1 U17607 ( .A1(n14007), .A2(n19276), .ZN(n14016) );
  AOI21_X1 U17608 ( .B1(n16186), .B2(n15048), .A(n9929), .ZN(n15049) );
  INV_X1 U17609 ( .A(n14009), .ZN(n14010) );
  OAI21_X1 U17610 ( .B1(n19288), .B2(n16186), .A(n14010), .ZN(n14012) );
  NOR2_X1 U17611 ( .A1(n16190), .A2(n16317), .ZN(n14011) );
  AOI211_X1 U17612 ( .C1(n19274), .C2(n15049), .A(n14012), .B(n14011), .ZN(
        n14015) );
  NAND3_X1 U17613 ( .A1(n14013), .A2(n16310), .A3(n9840), .ZN(n14014) );
  OAI211_X1 U17614 ( .C1(n13989), .C2(n14016), .A(n14015), .B(n14014), .ZN(
        P2_U2987) );
  INV_X1 U17615 ( .A(n14017), .ZN(n14018) );
  INV_X1 U17616 ( .A(n14022), .ZN(n14026) );
  NOR2_X1 U17617 ( .A1(n14023), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14025) );
  MUX2_X1 U17618 ( .A(n14026), .B(n14025), .S(n14024), .Z(n16165) );
  NAND2_X1 U17619 ( .A1(n16165), .A2(n10931), .ZN(n14027) );
  XNOR2_X1 U17620 ( .A(n14027), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14028) );
  XNOR2_X1 U17621 ( .A(n14029), .B(n14028), .ZN(n14061) );
  AOI22_X1 U17622 ( .A1(n14030), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14033) );
  NAND2_X1 U17623 ( .A1(n14031), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14032) );
  OAI211_X1 U17624 ( .C1(n10424), .C2(n14050), .A(n14033), .B(n14032), .ZN(
        n14034) );
  NAND2_X1 U17625 ( .A1(n19088), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14052) );
  NAND2_X1 U17626 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14036) );
  OAI211_X1 U17627 ( .C1(n16314), .C2(n14037), .A(n14052), .B(n14036), .ZN(
        n14038) );
  AOI21_X1 U17628 ( .B1(n16171), .B2(n19278), .A(n14038), .ZN(n14042) );
  NAND2_X1 U17629 ( .A1(n14058), .A2(n16310), .ZN(n14041) );
  OAI211_X1 U17630 ( .C1(n14061), .C2(n16292), .A(n14042), .B(n14041), .ZN(
        P2_U2983) );
  NAND2_X1 U17631 ( .A1(n14043), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14045) );
  AOI22_X1 U17632 ( .A1(n11516), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n13934), .B2(P2_EAX_REG_31__SCAN_IN), .ZN(n14044) );
  AND2_X1 U17633 ( .A1(n14045), .A2(n14044), .ZN(n14046) );
  NOR3_X1 U17634 ( .A1(n14048), .A2(n15446), .A3(n14050), .ZN(n14055) );
  NAND4_X1 U17635 ( .A1(n14051), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14050), .A4(n14049), .ZN(n14053) );
  NAND2_X1 U17636 ( .A1(n14053), .A2(n14052), .ZN(n14054) );
  OAI211_X1 U17637 ( .C1(n14061), .C2(n16369), .A(n14060), .B(n14059), .ZN(
        P2_U3015) );
  INV_X1 U17638 ( .A(n15221), .ZN(n14063) );
  AOI22_X1 U17639 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14069) );
  AOI22_X1 U17640 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14068) );
  AOI22_X1 U17641 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14067) );
  AOI22_X1 U17642 ( .A1(n14142), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14066) );
  NAND4_X1 U17643 ( .A1(n14069), .A2(n14068), .A3(n14067), .A4(n14066), .ZN(
        n14075) );
  AOI22_X1 U17644 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14073) );
  AOI22_X1 U17645 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14072) );
  AOI22_X1 U17646 ( .A1(n10669), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14071) );
  AOI22_X1 U17647 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14070) );
  NAND4_X1 U17648 ( .A1(n14073), .A2(n14072), .A3(n14071), .A4(n14070), .ZN(
        n14074) );
  AOI22_X1 U17649 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14079) );
  AOI22_X1 U17650 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U17651 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14077) );
  AOI22_X1 U17652 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14142), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14076) );
  NAND4_X1 U17653 ( .A1(n14079), .A2(n14078), .A3(n14077), .A4(n14076), .ZN(
        n14085) );
  AOI22_X1 U17654 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14151), .ZN(n14083) );
  AOI22_X1 U17655 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17656 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U17657 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14080) );
  NAND4_X1 U17658 ( .A1(n14083), .A2(n14082), .A3(n14081), .A4(n14080), .ZN(
        n14084) );
  INV_X1 U17659 ( .A(n15197), .ZN(n14097) );
  AOI22_X1 U17660 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14089) );
  AOI22_X1 U17661 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14088) );
  AOI22_X1 U17662 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14087) );
  AOI22_X1 U17663 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14142), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14086) );
  NAND4_X1 U17664 ( .A1(n14089), .A2(n14088), .A3(n14087), .A4(n14086), .ZN(
        n14095) );
  AOI22_X1 U17665 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n14151), .ZN(n14093) );
  AOI22_X1 U17666 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U17667 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U17668 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14090) );
  NAND4_X1 U17669 ( .A1(n14093), .A2(n14092), .A3(n14091), .A4(n14090), .ZN(
        n14094) );
  NOR2_X1 U17670 ( .A1(n14095), .A2(n14094), .ZN(n15198) );
  NAND2_X1 U17671 ( .A1(n14097), .A2(n14096), .ZN(n15193) );
  INV_X1 U17672 ( .A(n15193), .ZN(n14109) );
  AOI22_X1 U17673 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14101) );
  AOI22_X1 U17674 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14100) );
  AOI22_X1 U17675 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14099) );
  AOI22_X1 U17676 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n14142), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14098) );
  NAND4_X1 U17677 ( .A1(n14101), .A2(n14100), .A3(n14099), .A4(n14098), .ZN(
        n14107) );
  AOI22_X1 U17678 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n14151), .ZN(n14105) );
  AOI22_X1 U17679 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U17680 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14103) );
  AOI22_X1 U17681 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14102) );
  NAND4_X1 U17682 ( .A1(n14105), .A2(n14104), .A3(n14103), .A4(n14102), .ZN(
        n14106) );
  NOR2_X1 U17683 ( .A1(n14107), .A2(n14106), .ZN(n15194) );
  NAND2_X1 U17684 ( .A1(n14109), .A2(n14108), .ZN(n15182) );
  AOI22_X1 U17685 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U17686 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14112) );
  AOI22_X1 U17687 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U17688 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14142), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14110) );
  NAND4_X1 U17689 ( .A1(n14113), .A2(n14112), .A3(n14111), .A4(n14110), .ZN(
        n14119) );
  AOI22_X1 U17690 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n14151), .ZN(n14117) );
  AOI22_X1 U17691 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14116) );
  AOI22_X1 U17692 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14115) );
  AOI22_X1 U17693 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14114) );
  NAND4_X1 U17694 ( .A1(n14117), .A2(n14116), .A3(n14115), .A4(n14114), .ZN(
        n14118) );
  NOR2_X1 U17695 ( .A1(n14119), .A2(n14118), .ZN(n15183) );
  AOI22_X1 U17696 ( .A1(n11447), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U17697 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17698 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17699 ( .A1(n14142), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14120) );
  NAND4_X1 U17700 ( .A1(n14123), .A2(n14122), .A3(n14121), .A4(n14120), .ZN(
        n14129) );
  AOI22_X1 U17701 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14151), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14127) );
  AOI22_X1 U17702 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U17703 ( .A1(n10669), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U17704 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14124) );
  NAND4_X1 U17705 ( .A1(n14127), .A2(n14126), .A3(n14125), .A4(n14124), .ZN(
        n14128) );
  AOI22_X1 U17706 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11447), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14134) );
  AOI22_X1 U17707 ( .A1(n14141), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14133) );
  AOI22_X1 U17708 ( .A1(n10678), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14132) );
  AOI22_X1 U17709 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14142), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14131) );
  NAND4_X1 U17710 ( .A1(n14134), .A2(n14133), .A3(n14132), .A4(n14131), .ZN(
        n14140) );
  AOI22_X1 U17711 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n14151), .ZN(n14138) );
  AOI22_X1 U17712 ( .A1(n10685), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10573), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U17713 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14136) );
  AOI22_X1 U17714 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14135) );
  NAND4_X1 U17715 ( .A1(n14138), .A2(n14137), .A3(n14136), .A4(n14135), .ZN(
        n14139) );
  NOR2_X1 U17716 ( .A1(n14140), .A2(n14139), .ZN(n15175) );
  AOI22_X1 U17717 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11447), .B1(
        n10678), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U17718 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14141), .B1(
        n14130), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U17719 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n14142), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14145) );
  AOI22_X1 U17720 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10676), .B1(
        n10684), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14144) );
  NAND4_X1 U17721 ( .A1(n14147), .A2(n14146), .A3(n14145), .A4(n14144), .ZN(
        n14157) );
  INV_X1 U17722 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14149) );
  INV_X1 U17723 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14148) );
  OAI22_X1 U17724 ( .A1(n14149), .A2(n10668), .B1(n10738), .B2(n14148), .ZN(
        n14150) );
  INV_X1 U17725 ( .A(n14150), .ZN(n14155) );
  AOI22_X1 U17726 ( .A1(n10573), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14151), .ZN(n14154) );
  AOI22_X1 U17727 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10669), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17728 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10759), .B1(
        n10565), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14152) );
  NAND4_X1 U17729 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        n14156) );
  NOR2_X1 U17730 ( .A1(n14157), .A2(n14156), .ZN(n14200) );
  INV_X1 U17731 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19310) );
  INV_X1 U17732 ( .A(n14353), .ZN(n14270) );
  OAI22_X1 U17733 ( .A1(n14272), .A2(n19310), .B1(n14270), .B2(n14158), .ZN(
        n14163) );
  INV_X1 U17734 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14161) );
  INV_X1 U17735 ( .A(n14351), .ZN(n15745) );
  INV_X1 U17736 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14160) );
  OAI22_X1 U17737 ( .A1(n14159), .A2(n14161), .B1(n15745), .B2(n14160), .ZN(
        n14162) );
  NOR2_X1 U17738 ( .A1(n14163), .A2(n14162), .ZN(n14166) );
  AOI22_X1 U17739 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14165) );
  AOI22_X1 U17740 ( .A1(n14354), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14164) );
  XNOR2_X1 U17741 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14348) );
  NAND4_X1 U17742 ( .A1(n14166), .A2(n14165), .A3(n14164), .A4(n14348), .ZN(
        n14176) );
  INV_X1 U17743 ( .A(n14354), .ZN(n14330) );
  INV_X1 U17744 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14167) );
  INV_X1 U17745 ( .A(n14357), .ZN(n14328) );
  INV_X1 U17746 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19584) );
  OAI22_X1 U17747 ( .A1(n14330), .A2(n14167), .B1(n14328), .B2(n19584), .ZN(
        n14171) );
  INV_X1 U17748 ( .A(n14359), .ZN(n14334) );
  INV_X1 U17749 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14169) );
  INV_X1 U17750 ( .A(n14358), .ZN(n14332) );
  INV_X1 U17751 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14168) );
  OAI22_X1 U17752 ( .A1(n14334), .A2(n14169), .B1(n14332), .B2(n14168), .ZN(
        n14170) );
  NOR2_X1 U17753 ( .A1(n14171), .A2(n14170), .ZN(n14174) );
  INV_X1 U17754 ( .A(n14348), .ZN(n14360) );
  AOI22_X1 U17755 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14173) );
  AOI22_X1 U17756 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14172) );
  NAND4_X1 U17757 ( .A1(n14174), .A2(n14360), .A3(n14173), .A4(n14172), .ZN(
        n14175) );
  NAND2_X1 U17758 ( .A1(n14176), .A2(n14175), .ZN(n14205) );
  NOR2_X1 U17759 ( .A1(n19970), .A2(n14205), .ZN(n14177) );
  XOR2_X1 U17760 ( .A(n14200), .B(n14177), .Z(n14206) );
  INV_X1 U17761 ( .A(n14205), .ZN(n14201) );
  NAND2_X1 U17762 ( .A1(n14294), .A2(n14201), .ZN(n15163) );
  INV_X1 U17763 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14180) );
  OAI22_X1 U17764 ( .A1(n14330), .A2(n14181), .B1(n14332), .B2(n14180), .ZN(
        n14185) );
  INV_X1 U17765 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14182) );
  OAI22_X1 U17766 ( .A1(n14334), .A2(n14183), .B1(n14328), .B2(n14182), .ZN(
        n14184) );
  NOR2_X1 U17767 ( .A1(n14185), .A2(n14184), .ZN(n14188) );
  AOI22_X1 U17768 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14187) );
  AOI22_X1 U17769 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14186) );
  NAND4_X1 U17770 ( .A1(n14188), .A2(n14187), .A3(n14186), .A4(n14348), .ZN(
        n14199) );
  INV_X1 U17771 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14190) );
  OAI22_X1 U17772 ( .A1(n14330), .A2(n14190), .B1(n14332), .B2(n14189), .ZN(
        n14194) );
  INV_X1 U17773 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14192) );
  OAI22_X1 U17774 ( .A1(n14334), .A2(n14192), .B1(n14328), .B2(n14191), .ZN(
        n14193) );
  NOR2_X1 U17775 ( .A1(n14194), .A2(n14193), .ZN(n14197) );
  AOI22_X1 U17776 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U17777 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14195) );
  NAND4_X1 U17778 ( .A1(n14197), .A2(n14360), .A3(n14196), .A4(n14195), .ZN(
        n14198) );
  NAND2_X1 U17779 ( .A1(n14199), .A2(n14198), .ZN(n14208) );
  INV_X1 U17780 ( .A(n14200), .ZN(n14202) );
  NAND2_X1 U17781 ( .A1(n14202), .A2(n14201), .ZN(n14209) );
  XOR2_X1 U17782 ( .A(n14208), .B(n14209), .Z(n14203) );
  NAND2_X1 U17783 ( .A1(n14203), .A2(n14288), .ZN(n15156) );
  INV_X1 U17784 ( .A(n14208), .ZN(n14204) );
  NAND2_X1 U17785 ( .A1(n19970), .A2(n14204), .ZN(n15159) );
  NOR3_X1 U17786 ( .A1(n14206), .A2(n14205), .A3(n15159), .ZN(n14207) );
  NOR2_X1 U17787 ( .A1(n14209), .A2(n14208), .ZN(n14230) );
  INV_X1 U17788 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14211) );
  INV_X1 U17789 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14210) );
  OAI22_X1 U17790 ( .A1(n14272), .A2(n14211), .B1(n14270), .B2(n14210), .ZN(
        n14215) );
  INV_X1 U17791 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14213) );
  OAI22_X1 U17792 ( .A1(n14275), .A2(n14213), .B1(n15745), .B2(n14212), .ZN(
        n14214) );
  NOR2_X1 U17793 ( .A1(n14215), .A2(n14214), .ZN(n14218) );
  AOI22_X1 U17794 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14217) );
  AOI22_X1 U17795 ( .A1(n14354), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14216) );
  NAND4_X1 U17796 ( .A1(n14218), .A2(n14217), .A3(n14216), .A4(n14348), .ZN(
        n14229) );
  INV_X1 U17797 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14220) );
  INV_X1 U17798 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14219) );
  OAI22_X1 U17799 ( .A1(n14272), .A2(n14220), .B1(n14270), .B2(n14219), .ZN(
        n14224) );
  INV_X1 U17800 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14222) );
  OAI22_X1 U17801 ( .A1(n14275), .A2(n14222), .B1(n15745), .B2(n14221), .ZN(
        n14223) );
  NOR2_X1 U17802 ( .A1(n14224), .A2(n14223), .ZN(n14227) );
  AOI22_X1 U17803 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14226) );
  AOI22_X1 U17804 ( .A1(n14354), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14225) );
  NAND4_X1 U17805 ( .A1(n14227), .A2(n14360), .A3(n14226), .A4(n14225), .ZN(
        n14228) );
  AND2_X1 U17806 ( .A1(n14229), .A2(n14228), .ZN(n14231) );
  NAND2_X1 U17807 ( .A1(n14230), .A2(n14231), .ZN(n14285) );
  OAI211_X1 U17808 ( .C1(n14230), .C2(n14231), .A(n14285), .B(n14288), .ZN(
        n14234) );
  INV_X1 U17809 ( .A(n14231), .ZN(n14232) );
  NOR2_X1 U17810 ( .A1(n14316), .A2(n14232), .ZN(n15151) );
  NAND2_X1 U17811 ( .A1(n15152), .A2(n15151), .ZN(n15150) );
  INV_X1 U17812 ( .A(n14233), .ZN(n14236) );
  OAI22_X1 U17813 ( .A1(n14330), .A2(n14239), .B1(n14332), .B2(n14238), .ZN(
        n14243) );
  INV_X1 U17814 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14240) );
  OAI22_X1 U17815 ( .A1(n14334), .A2(n14241), .B1(n14328), .B2(n14240), .ZN(
        n14242) );
  NOR2_X1 U17816 ( .A1(n14243), .A2(n14242), .ZN(n14246) );
  AOI22_X1 U17817 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14245) );
  AOI22_X1 U17818 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14244) );
  NAND4_X1 U17819 ( .A1(n14246), .A2(n14245), .A3(n14244), .A4(n14348), .ZN(
        n14257) );
  INV_X1 U17820 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14248) );
  OAI22_X1 U17821 ( .A1(n14330), .A2(n14248), .B1(n14332), .B2(n14247), .ZN(
        n14252) );
  OAI22_X1 U17822 ( .A1(n14334), .A2(n14250), .B1(n14328), .B2(n14249), .ZN(
        n14251) );
  NOR2_X1 U17823 ( .A1(n14252), .A2(n14251), .ZN(n14255) );
  AOI22_X1 U17824 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14254) );
  AOI22_X1 U17825 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14253) );
  NAND4_X1 U17826 ( .A1(n14255), .A2(n14360), .A3(n14254), .A4(n14253), .ZN(
        n14256) );
  AND2_X1 U17827 ( .A1(n14257), .A2(n14256), .ZN(n14283) );
  XNOR2_X1 U17828 ( .A(n14285), .B(n14283), .ZN(n14258) );
  NAND2_X1 U17829 ( .A1(n14294), .A2(n14283), .ZN(n15146) );
  INV_X1 U17830 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19331) );
  OAI22_X1 U17831 ( .A1(n14272), .A2(n19331), .B1(n14270), .B2(n14261), .ZN(
        n14265) );
  INV_X1 U17832 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14263) );
  INV_X1 U17833 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14262) );
  OAI22_X1 U17834 ( .A1(n14275), .A2(n14263), .B1(n15745), .B2(n14262), .ZN(
        n14264) );
  NOR2_X1 U17835 ( .A1(n14265), .A2(n14264), .ZN(n14268) );
  AOI22_X1 U17836 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14267) );
  AOI22_X1 U17837 ( .A1(n14354), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14266) );
  NAND4_X1 U17838 ( .A1(n14268), .A2(n14267), .A3(n14266), .A4(n14348), .ZN(
        n14282) );
  INV_X1 U17839 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14271) );
  OAI22_X1 U17840 ( .A1(n14272), .A2(n14271), .B1(n14270), .B2(n14269), .ZN(
        n14277) );
  INV_X1 U17841 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14274) );
  INV_X1 U17842 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14273) );
  OAI22_X1 U17843 ( .A1(n14275), .A2(n14274), .B1(n15745), .B2(n14273), .ZN(
        n14276) );
  NOR2_X1 U17844 ( .A1(n14277), .A2(n14276), .ZN(n14280) );
  AOI22_X1 U17845 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14279) );
  AOI22_X1 U17846 ( .A1(n14354), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14278) );
  NAND4_X1 U17847 ( .A1(n14280), .A2(n14360), .A3(n14279), .A4(n14278), .ZN(
        n14281) );
  NAND2_X1 U17848 ( .A1(n14282), .A2(n14281), .ZN(n14286) );
  INV_X1 U17849 ( .A(n14286), .ZN(n14293) );
  INV_X1 U17850 ( .A(n14283), .ZN(n14284) );
  INV_X1 U17851 ( .A(n14287), .ZN(n14289) );
  OR2_X1 U17852 ( .A1(n14287), .A2(n14286), .ZN(n15131) );
  OAI211_X1 U17853 ( .C1(n14293), .C2(n14289), .A(n14288), .B(n15131), .ZN(
        n14291) );
  NOR2_X1 U17854 ( .A1(n14290), .A2(n14291), .ZN(n14315) );
  NAND2_X1 U17855 ( .A1(n14294), .A2(n14293), .ZN(n15137) );
  OAI22_X1 U17856 ( .A1(n14330), .A2(n14296), .B1(n14332), .B2(n14295), .ZN(
        n14300) );
  INV_X1 U17857 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14297) );
  OAI22_X1 U17858 ( .A1(n14334), .A2(n14298), .B1(n14328), .B2(n14297), .ZN(
        n14299) );
  NOR2_X1 U17859 ( .A1(n14300), .A2(n14299), .ZN(n14303) );
  AOI22_X1 U17860 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14302) );
  AOI22_X1 U17861 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14301) );
  NAND4_X1 U17862 ( .A1(n14303), .A2(n14302), .A3(n14301), .A4(n14348), .ZN(
        n14314) );
  INV_X1 U17863 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14305) );
  OAI22_X1 U17864 ( .A1(n14330), .A2(n14305), .B1(n14332), .B2(n14304), .ZN(
        n14309) );
  OAI22_X1 U17865 ( .A1(n14334), .A2(n14307), .B1(n14328), .B2(n14306), .ZN(
        n14308) );
  NOR2_X1 U17866 ( .A1(n14309), .A2(n14308), .ZN(n14312) );
  AOI22_X1 U17867 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14311) );
  AOI22_X1 U17868 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14310) );
  NAND4_X1 U17869 ( .A1(n14312), .A2(n14360), .A3(n14311), .A4(n14310), .ZN(
        n14313) );
  AND2_X1 U17870 ( .A1(n14314), .A2(n14313), .ZN(n15132) );
  NAND2_X1 U17871 ( .A1(n14316), .A2(n15132), .ZN(n14317) );
  NOR2_X1 U17872 ( .A1(n15131), .A2(n14317), .ZN(n14343) );
  OAI22_X1 U17873 ( .A1(n14330), .A2(n14319), .B1(n14332), .B2(n14318), .ZN(
        n14323) );
  INV_X1 U17874 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14320) );
  OAI22_X1 U17875 ( .A1(n14334), .A2(n14321), .B1(n14328), .B2(n14320), .ZN(
        n14322) );
  NOR2_X1 U17876 ( .A1(n14323), .A2(n14322), .ZN(n14326) );
  AOI22_X1 U17877 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14325) );
  AOI22_X1 U17878 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14324) );
  NAND4_X1 U17879 ( .A1(n14326), .A2(n14325), .A3(n14324), .A4(n14348), .ZN(
        n14341) );
  INV_X1 U17880 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14329) );
  OAI22_X1 U17881 ( .A1(n14330), .A2(n14329), .B1(n14328), .B2(n14327), .ZN(
        n14336) );
  OAI22_X1 U17882 ( .A1(n14334), .A2(n14333), .B1(n14332), .B2(n14331), .ZN(
        n14335) );
  NOR2_X1 U17883 ( .A1(n14336), .A2(n14335), .ZN(n14339) );
  AOI22_X1 U17884 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U17885 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14337) );
  NAND4_X1 U17886 ( .A1(n14339), .A2(n14360), .A3(n14338), .A4(n14337), .ZN(
        n14340) );
  AND2_X1 U17887 ( .A1(n14341), .A2(n14340), .ZN(n14342) );
  NAND2_X1 U17888 ( .A1(n14343), .A2(n14342), .ZN(n14344) );
  OAI21_X1 U17889 ( .B1(n14343), .B2(n14342), .A(n14344), .ZN(n15128) );
  INV_X1 U17890 ( .A(n14344), .ZN(n14345) );
  AOI22_X1 U17891 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14347) );
  AOI22_X1 U17892 ( .A1(n14354), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14346) );
  NAND2_X1 U17893 ( .A1(n14347), .A2(n14346), .ZN(n14366) );
  AOI22_X1 U17894 ( .A1(n9807), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14350) );
  AOI22_X1 U17895 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14349) );
  NAND3_X1 U17896 ( .A1(n14350), .A2(n14349), .A3(n14348), .ZN(n14365) );
  AOI22_X1 U17897 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14356) );
  AOI22_X1 U17898 ( .A1(n14354), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14355) );
  NAND2_X1 U17899 ( .A1(n14356), .A2(n14355), .ZN(n14364) );
  AOI22_X1 U17900 ( .A1(n10543), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14357), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U17901 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14361) );
  NAND3_X1 U17902 ( .A1(n14362), .A2(n14361), .A3(n14360), .ZN(n14363) );
  OAI22_X1 U17903 ( .A1(n14366), .A2(n14365), .B1(n14364), .B2(n14363), .ZN(
        n14367) );
  XNOR2_X1 U17904 ( .A(n14368), .B(n14367), .ZN(n14382) );
  NOR2_X1 U17905 ( .A1(n15058), .A2(n15205), .ZN(n14369) );
  AOI21_X1 U17906 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15205), .A(n14369), .ZN(
        n14370) );
  OAI21_X1 U17907 ( .B1(n14382), .B2(n15219), .A(n14370), .ZN(P2_U2857) );
  NAND2_X1 U17908 ( .A1(n14371), .A2(n14372), .ZN(n14373) );
  OR2_X1 U17909 ( .A1(n19190), .A2(n14373), .ZN(n19160) );
  OR2_X1 U17910 ( .A1(n19190), .A2(n14374), .ZN(n15287) );
  OAI22_X1 U17911 ( .A1(n14375), .A2(n15287), .B1(n15286), .B2(n19210), .ZN(
        n14380) );
  NAND2_X1 U17912 ( .A1(n14371), .A2(n14376), .ZN(n14377) );
  INV_X1 U17913 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14378) );
  OAI22_X1 U17914 ( .A1(n15292), .A2(n14378), .B1(n19170), .B2(n15054), .ZN(
        n14379) );
  AOI211_X1 U17915 ( .C1(n19168), .C2(BUF1_REG_30__SCAN_IN), .A(n14380), .B(
        n14379), .ZN(n14381) );
  OAI21_X1 U17916 ( .B1(n14382), .B2(n19171), .A(n14381), .ZN(P2_U2889) );
  OAI22_X1 U17917 ( .A1(n14388), .A2(n12638), .B1(n14392), .B2(n14383), .ZN(
        n14390) );
  NOR2_X1 U17918 ( .A1(n15847), .A2(n14384), .ZN(n14387) );
  NAND2_X1 U17919 ( .A1(n14388), .A2(n14385), .ZN(n14386) );
  OAI21_X1 U17920 ( .B1(n14388), .B2(n14387), .A(n14386), .ZN(n14389) );
  NOR2_X1 U17921 ( .A1(n14390), .A2(n14389), .ZN(n15849) );
  INV_X1 U17922 ( .A(n15849), .ZN(n14398) );
  AOI21_X1 U17923 ( .B1(n14392), .B2(n12645), .A(n14391), .ZN(n14393) );
  AOI21_X1 U17924 ( .B1(n15862), .B2(n14395), .A(n14393), .ZN(n19991) );
  NAND3_X1 U17925 ( .A1(n14395), .A2(n14394), .A3(n15880), .ZN(n14396) );
  NAND2_X1 U17926 ( .A1(n14396), .A2(n20880), .ZN(n20877) );
  NAND2_X1 U17927 ( .A1(n19991), .A2(n20877), .ZN(n15851) );
  AND2_X1 U17928 ( .A1(n15851), .A2(n14397), .ZN(n20001) );
  MUX2_X1 U17929 ( .A(P1_MORE_REG_SCAN_IN), .B(n14398), .S(n20001), .Z(
        P1_U3484) );
  NAND2_X1 U17930 ( .A1(n14716), .A2(n20050), .ZN(n14407) );
  INV_X1 U17931 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20833) );
  INV_X1 U17932 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14399) );
  OAI21_X1 U17933 ( .B1(n14415), .B2(n20833), .A(n14399), .ZN(n14405) );
  NOR2_X1 U17934 ( .A1(n20043), .A2(n14400), .ZN(n14403) );
  OAI22_X1 U17935 ( .A1(n14401), .A2(n20025), .B1(n20078), .B2(n14714), .ZN(
        n14402) );
  AOI211_X1 U17936 ( .C1(n14405), .C2(n14404), .A(n14403), .B(n14402), .ZN(
        n14406) );
  OAI211_X1 U17937 ( .C1(n20098), .C2(n14867), .A(n14407), .B(n14406), .ZN(
        P1_U2810) );
  NAND2_X1 U17938 ( .A1(n14421), .A2(n14408), .ZN(n14409) );
  NAND2_X1 U17939 ( .A1(n14410), .A2(n14409), .ZN(n14881) );
  INV_X1 U17940 ( .A(n14725), .ZN(n14413) );
  NAND2_X1 U17941 ( .A1(n14413), .A2(n20050), .ZN(n14418) );
  AOI22_X1 U17942 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20087), .B1(
        n20081), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n14414) );
  OAI221_X1 U17943 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14415), .C1(n20833), 
        .C2(n14428), .A(n14414), .ZN(n14416) );
  AOI21_X1 U17944 ( .B1(n20086), .B2(n14720), .A(n14416), .ZN(n14417) );
  OAI211_X1 U17945 ( .C1(n20098), .C2(n14881), .A(n14418), .B(n14417), .ZN(
        P1_U2811) );
  OR2_X1 U17946 ( .A1(n14436), .A2(n14419), .ZN(n14420) );
  NAND2_X1 U17947 ( .A1(n14421), .A2(n14420), .ZN(n14893) );
  INV_X1 U17948 ( .A(n14422), .ZN(n14425) );
  INV_X1 U17949 ( .A(n14423), .ZN(n14424) );
  NAND2_X1 U17950 ( .A1(n14737), .A2(n20050), .ZN(n14434) );
  OAI22_X1 U17951 ( .A1(n14426), .A2(n20025), .B1(n20078), .B2(n14735), .ZN(
        n14432) );
  INV_X1 U17952 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14430) );
  NAND3_X1 U17953 ( .A1(n20084), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14427), 
        .ZN(n14429) );
  AOI21_X1 U17954 ( .B1(n14430), .B2(n14429), .A(n14428), .ZN(n14431) );
  AOI211_X1 U17955 ( .C1(n20081), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14432), .B(
        n14431), .ZN(n14433) );
  OAI211_X1 U17956 ( .C1(n20098), .C2(n14893), .A(n14434), .B(n14433), .ZN(
        P1_U2812) );
  AND2_X1 U17957 ( .A1(n14449), .A2(n14435), .ZN(n14437) );
  OR2_X1 U17958 ( .A1(n14437), .A2(n14436), .ZN(n14902) );
  AOI21_X1 U17959 ( .B1(n14439), .B2(n14438), .A(n14423), .ZN(n14744) );
  NAND2_X1 U17960 ( .A1(n14744), .A2(n20050), .ZN(n14446) );
  NAND2_X1 U17961 ( .A1(n20084), .A2(n14440), .ZN(n14458) );
  NAND2_X1 U17962 ( .A1(n14458), .A2(n20079), .ZN(n14461) );
  INV_X1 U17963 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14550) );
  INV_X1 U17964 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20828) );
  NAND2_X1 U17965 ( .A1(n14441), .A2(n20828), .ZN(n14443) );
  AOI22_X1 U17966 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20087), .B1(
        n20086), .B2(n14747), .ZN(n14442) );
  OAI211_X1 U17967 ( .C1(n14550), .C2(n20043), .A(n14443), .B(n14442), .ZN(
        n14444) );
  AOI21_X1 U17968 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14461), .A(n14444), 
        .ZN(n14445) );
  OAI211_X1 U17969 ( .C1(n20098), .C2(n14902), .A(n14446), .B(n14445), .ZN(
        P1_U2813) );
  NAND2_X1 U17970 ( .A1(n14556), .A2(n14447), .ZN(n14448) );
  NAND2_X1 U17971 ( .A1(n14449), .A2(n14448), .ZN(n14910) );
  INV_X1 U17972 ( .A(n14438), .ZN(n14452) );
  AOI21_X1 U17973 ( .B1(n14453), .B2(n14450), .A(n14452), .ZN(n14759) );
  NAND2_X1 U17974 ( .A1(n14759), .A2(n20050), .ZN(n14463) );
  INV_X1 U17975 ( .A(n14454), .ZN(n14459) );
  OAI22_X1 U17976 ( .A1(n14455), .A2(n20025), .B1(n20078), .B2(n14757), .ZN(
        n14456) );
  AOI21_X1 U17977 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(n20081), .A(n14456), .ZN(
        n14457) );
  OAI21_X1 U17978 ( .B1(n14459), .B2(n14458), .A(n14457), .ZN(n14460) );
  AOI21_X1 U17979 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n14461), .A(n14460), 
        .ZN(n14462) );
  OAI211_X1 U17980 ( .C1(n20098), .C2(n14910), .A(n14463), .B(n14462), .ZN(
        P1_U2814) );
  INV_X1 U17981 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14476) );
  INV_X1 U17982 ( .A(n14464), .ZN(n15903) );
  NAND2_X1 U17983 ( .A1(n20079), .A2(n15903), .ZN(n14469) );
  NAND2_X1 U17984 ( .A1(n20031), .A2(n14469), .ZN(n15896) );
  AOI21_X1 U17985 ( .B1(n14466), .B2(n9847), .A(n14465), .ZN(n14783) );
  NAND2_X1 U17986 ( .A1(n14783), .A2(n20050), .ZN(n14475) );
  AND2_X1 U17987 ( .A1(n9874), .A2(n14467), .ZN(n14468) );
  NOR2_X1 U17988 ( .A1(n14565), .A2(n14468), .ZN(n14938) );
  NAND3_X1 U17989 ( .A1(n20084), .A2(n14470), .A3(n14469), .ZN(n14472) );
  AOI22_X1 U17990 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20087), .B1(
        n20086), .B2(n14779), .ZN(n14471) );
  OAI211_X1 U17991 ( .C1(n21069), .C2(n20043), .A(n14472), .B(n14471), .ZN(
        n14473) );
  AOI21_X1 U17992 ( .B1(n14938), .B2(n20056), .A(n14473), .ZN(n14474) );
  OAI211_X1 U17993 ( .C1(n14476), .C2(n15896), .A(n14475), .B(n14474), .ZN(
        P1_U2817) );
  OAI21_X1 U17994 ( .B1(n14477), .B2(n14479), .A(n14478), .ZN(n14803) );
  NAND3_X1 U17995 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .ZN(n14482) );
  NAND2_X1 U17996 ( .A1(n14495), .A2(n14480), .ZN(n14510) );
  OR2_X1 U17997 ( .A1(n14481), .A2(n14510), .ZN(n14497) );
  NOR2_X1 U17998 ( .A1(n14482), .A2(n14497), .ZN(n14483) );
  NOR2_X1 U17999 ( .A1(n14483), .A2(n20062), .ZN(n15928) );
  NOR2_X1 U18000 ( .A1(n20080), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15914) );
  AOI22_X1 U18001 ( .A1(n14483), .A2(n15914), .B1(n20081), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n14484) );
  OAI21_X1 U18002 ( .B1(n14793), .B2(n20025), .A(n14484), .ZN(n14485) );
  AOI21_X1 U18003 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15928), .A(n14485), 
        .ZN(n14489) );
  INV_X1 U18004 ( .A(n14582), .ZN(n14486) );
  AOI21_X1 U18005 ( .B1(n14487), .B2(n14486), .A(n10165), .ZN(n14959) );
  AOI22_X1 U18006 ( .A1(n14959), .A2(n20056), .B1(n14795), .B2(n20086), .ZN(
        n14488) );
  OAI211_X1 U18007 ( .C1(n14803), .C2(n15945), .A(n14489), .B(n14488), .ZN(
        P1_U2819) );
  INV_X1 U18008 ( .A(n14492), .ZN(n14493) );
  AOI21_X1 U18009 ( .B1(n14494), .B2(n14490), .A(n14493), .ZN(n14829) );
  INV_X1 U18010 ( .A(n14829), .ZN(n14692) );
  NAND2_X1 U18011 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14496) );
  NAND2_X1 U18012 ( .A1(n14495), .A2(n20027), .ZN(n15954) );
  NOR2_X1 U18013 ( .A1(n14496), .A2(n15954), .ZN(n15912) );
  AND2_X1 U18014 ( .A1(n14497), .A2(n20031), .ZN(n15941) );
  OAI21_X1 U18015 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15912), .A(n15941), 
        .ZN(n14505) );
  OR2_X1 U18016 ( .A1(n14604), .A2(n14498), .ZN(n14499) );
  AND2_X1 U18017 ( .A1(n14499), .A2(n14598), .ZN(n16059) );
  INV_X1 U18018 ( .A(n14827), .ZN(n14500) );
  AOI22_X1 U18019 ( .A1(P1_EBX_REG_17__SCAN_IN), .A2(n20081), .B1(n20086), 
        .B2(n14500), .ZN(n14501) );
  OAI211_X1 U18020 ( .C1(n20025), .C2(n14502), .A(n14501), .B(n20022), .ZN(
        n14503) );
  AOI21_X1 U18021 ( .B1(n20056), .B2(n16059), .A(n14503), .ZN(n14504) );
  OAI211_X1 U18022 ( .C1(n14692), .C2(n15945), .A(n14505), .B(n14504), .ZN(
        P1_U2823) );
  OAI21_X1 U18023 ( .B1(n14506), .B2(n14509), .A(n14508), .ZN(n14836) );
  INV_X1 U18024 ( .A(n14838), .ZN(n14518) );
  INV_X1 U18025 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20813) );
  NAND2_X1 U18026 ( .A1(n20031), .A2(n14510), .ZN(n15965) );
  AOI21_X1 U18027 ( .B1(n20087), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20069), .ZN(n14515) );
  NAND2_X1 U18028 ( .A1(n14512), .A2(n14511), .ZN(n14513) );
  AND2_X1 U18029 ( .A1(n14603), .A2(n14513), .ZN(n16066) );
  AOI22_X1 U18030 ( .A1(n20056), .A2(n16066), .B1(n20081), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14514) );
  OAI211_X1 U18031 ( .C1(n20813), .C2(n15965), .A(n14515), .B(n14514), .ZN(
        n14517) );
  NOR2_X1 U18032 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15954), .ZN(n14516) );
  AOI211_X1 U18033 ( .C1(n20086), .C2(n14518), .A(n14517), .B(n14516), .ZN(
        n14519) );
  OAI21_X1 U18034 ( .B1(n14836), .B2(n15945), .A(n14519), .ZN(P1_U2825) );
  OR2_X1 U18035 ( .A1(n14521), .A2(n14520), .ZN(n14522) );
  NAND2_X1 U18036 ( .A1(n14522), .A2(n13769), .ZN(n14617) );
  NOR2_X1 U18037 ( .A1(n14525), .A2(n14524), .ZN(n15980) );
  NAND2_X1 U18038 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14528) );
  NOR2_X1 U18039 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14528), .ZN(n14537) );
  OR2_X1 U18040 ( .A1(n14625), .A2(n14526), .ZN(n14527) );
  NAND2_X1 U18041 ( .A1(n9897), .A2(n14527), .ZN(n16071) );
  INV_X1 U18042 ( .A(n14850), .ZN(n14534) );
  INV_X1 U18043 ( .A(n14528), .ZN(n14530) );
  OAI21_X1 U18044 ( .B1(n20062), .B2(n14530), .A(n14529), .ZN(n15972) );
  AOI22_X1 U18045 ( .A1(n20081), .A2(P1_EBX_REG_13__SCAN_IN), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n15972), .ZN(n14531) );
  OAI211_X1 U18046 ( .C1(n20025), .C2(n14532), .A(n14531), .B(n20022), .ZN(
        n14533) );
  AOI21_X1 U18047 ( .B1(n20086), .B2(n14534), .A(n14533), .ZN(n14535) );
  OAI21_X1 U18048 ( .B1(n20098), .B2(n16071), .A(n14535), .ZN(n14536) );
  AOI21_X1 U18049 ( .B1(n15980), .B2(n14537), .A(n14536), .ZN(n14538) );
  OAI21_X1 U18050 ( .B1(n14854), .B2(n15945), .A(n14538), .ZN(P1_U2827) );
  OAI22_X1 U18051 ( .A1(n20098), .A2(n20225), .B1(n20043), .B2(n14539), .ZN(
        n14540) );
  AOI21_X1 U18052 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n20031), .A(n14540), .ZN(
        n14543) );
  NAND2_X1 U18053 ( .A1(n20025), .A2(n20078), .ZN(n14541) );
  AOI22_X1 U18054 ( .A1(n20089), .A2(n11939), .B1(n14541), .B2(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14542) );
  OAI211_X1 U18055 ( .C1(n14545), .C2(n14544), .A(n14543), .B(n14542), .ZN(
        P1_U2840) );
  OAI22_X1 U18056 ( .A1(n14546), .A2(n14608), .B1(n14626), .B2(n12670), .ZN(
        P1_U2841) );
  OAI222_X1 U18057 ( .A1(n14627), .A2(n14725), .B1(n14547), .B2(n14626), .C1(
        n14881), .C2(n14608), .ZN(P1_U2843) );
  INV_X1 U18058 ( .A(n14737), .ZN(n14549) );
  INV_X1 U18059 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14548) );
  OAI222_X1 U18060 ( .A1(n14627), .A2(n14549), .B1(n14548), .B2(n14626), .C1(
        n14893), .C2(n14608), .ZN(P1_U2844) );
  INV_X1 U18061 ( .A(n14744), .ZN(n14647) );
  OAI222_X1 U18062 ( .A1(n14627), .A2(n14647), .B1(n14626), .B2(n14550), .C1(
        n14902), .C2(n14608), .ZN(P1_U2845) );
  INV_X1 U18063 ( .A(n14759), .ZN(n14652) );
  INV_X1 U18064 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14551) );
  OAI222_X1 U18065 ( .A1(n14627), .A2(n14652), .B1(n14626), .B2(n14551), .C1(
        n14910), .C2(n14608), .ZN(P1_U2846) );
  OAI21_X1 U18066 ( .B1(n14552), .B2(n14553), .A(n14450), .ZN(n15893) );
  OR2_X1 U18067 ( .A1(n14562), .A2(n14554), .ZN(n14555) );
  NAND2_X1 U18068 ( .A1(n14556), .A2(n14555), .ZN(n15892) );
  OAI22_X1 U18069 ( .A1(n15892), .A2(n14608), .B1(n14557), .B2(n14626), .ZN(
        n14558) );
  INV_X1 U18070 ( .A(n14558), .ZN(n14559) );
  OAI21_X1 U18071 ( .B1(n15893), .B2(n14627), .A(n14559), .ZN(P1_U2847) );
  NOR2_X1 U18072 ( .A1(n14465), .A2(n14560), .ZN(n14561) );
  OR2_X1 U18073 ( .A1(n14552), .A2(n14561), .ZN(n14774) );
  INV_X1 U18074 ( .A(n14562), .ZN(n14563) );
  OAI21_X1 U18075 ( .B1(n14565), .B2(n14564), .A(n14563), .ZN(n15907) );
  INV_X1 U18076 ( .A(n15907), .ZN(n14926) );
  AOI22_X1 U18077 ( .A1(n14926), .A2(n14614), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14612), .ZN(n14566) );
  OAI21_X1 U18078 ( .B1(n14774), .B2(n14627), .A(n14566), .ZN(P1_U2848) );
  INV_X1 U18079 ( .A(n14783), .ZN(n14665) );
  AOI22_X1 U18080 ( .A1(n14938), .A2(n14614), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14612), .ZN(n14567) );
  OAI21_X1 U18081 ( .B1(n14665), .B2(n14627), .A(n14567), .ZN(P1_U2849) );
  NAND2_X1 U18082 ( .A1(n14478), .A2(n14568), .ZN(n14569) );
  NAND2_X1 U18083 ( .A1(n14571), .A2(n14570), .ZN(n14572) );
  NAND2_X1 U18084 ( .A1(n9874), .A2(n14572), .ZN(n15924) );
  OAI22_X1 U18085 ( .A1(n15924), .A2(n14608), .B1(n14573), .B2(n14626), .ZN(
        n14574) );
  AOI21_X1 U18086 ( .B1(n15922), .B2(n14584), .A(n14574), .ZN(n14575) );
  INV_X1 U18087 ( .A(n14575), .ZN(P1_U2850) );
  AOI22_X1 U18088 ( .A1(n14959), .A2(n14614), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14612), .ZN(n14576) );
  OAI21_X1 U18089 ( .B1(n14803), .B2(n14627), .A(n14576), .ZN(P1_U2851) );
  NOR2_X1 U18090 ( .A1(n14577), .A2(n14578), .ZN(n14579) );
  OR2_X1 U18091 ( .A1(n14477), .A2(n14579), .ZN(n14681) );
  NOR2_X1 U18092 ( .A1(n14590), .A2(n14580), .ZN(n14581) );
  OR2_X1 U18093 ( .A1(n14582), .A2(n14581), .ZN(n15931) );
  OAI22_X1 U18094 ( .A1(n15931), .A2(n14608), .B1(n15925), .B2(n14626), .ZN(
        n14583) );
  AOI21_X1 U18095 ( .B1(n15994), .B2(n14584), .A(n14583), .ZN(n14585) );
  INV_X1 U18096 ( .A(n14585), .ZN(P1_U2852) );
  INV_X1 U18097 ( .A(n14577), .ZN(n14587) );
  OAI21_X1 U18098 ( .B1(n14588), .B2(n14586), .A(n14587), .ZN(n15935) );
  AND2_X1 U18099 ( .A1(n9873), .A2(n14589), .ZN(n14591) );
  OR2_X1 U18100 ( .A1(n14591), .A2(n14590), .ZN(n16040) );
  OAI22_X1 U18101 ( .A1(n16040), .A2(n14608), .B1(n14592), .B2(n14626), .ZN(
        n14593) );
  INV_X1 U18102 ( .A(n14593), .ZN(n14594) );
  OAI21_X1 U18103 ( .B1(n15935), .B2(n14627), .A(n14594), .ZN(P1_U2853) );
  AND2_X1 U18104 ( .A1(n14492), .A2(n14595), .ZN(n14596) );
  OR2_X1 U18105 ( .A1(n14596), .A2(n14586), .ZN(n15946) );
  INV_X1 U18106 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14600) );
  NAND2_X1 U18107 ( .A1(n14598), .A2(n14597), .ZN(n14599) );
  NAND2_X1 U18108 ( .A1(n9873), .A2(n14599), .ZN(n16048) );
  OAI222_X1 U18109 ( .A1(n15946), .A2(n14627), .B1(n14600), .B2(n14626), .C1(
        n16048), .C2(n14608), .ZN(P1_U2854) );
  AOI22_X1 U18110 ( .A1(n16059), .A2(n14614), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14612), .ZN(n14601) );
  OAI21_X1 U18111 ( .B1(n14692), .B2(n14627), .A(n14601), .ZN(P1_U2855) );
  AND2_X1 U18112 ( .A1(n14603), .A2(n14602), .ZN(n14605) );
  OR2_X1 U18113 ( .A1(n14605), .A2(n14604), .ZN(n15951) );
  INV_X1 U18114 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21014) );
  AOI21_X1 U18115 ( .B1(n14606), .B2(n14508), .A(n10211), .ZN(n15998) );
  INV_X1 U18116 ( .A(n15998), .ZN(n14607) );
  OAI222_X1 U18117 ( .A1(n15951), .A2(n14608), .B1(n14626), .B2(n21014), .C1(
        n14607), .C2(n14627), .ZN(P1_U2856) );
  AOI22_X1 U18118 ( .A1(n14614), .A2(n16066), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14612), .ZN(n14609) );
  OAI21_X1 U18119 ( .B1(n14836), .B2(n14627), .A(n14609), .ZN(P1_U2857) );
  INV_X1 U18120 ( .A(n14610), .ZN(n14611) );
  AOI21_X1 U18121 ( .B1(n14611), .B2(n9876), .A(n14506), .ZN(n16004) );
  INV_X1 U18122 ( .A(n16004), .ZN(n14701) );
  INV_X1 U18123 ( .A(n15961), .ZN(n14613) );
  AOI22_X1 U18124 ( .A1(n14614), .A2(n14613), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14612), .ZN(n14615) );
  OAI21_X1 U18125 ( .B1(n14701), .B2(n14627), .A(n14615), .ZN(P1_U2858) );
  INV_X1 U18126 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14616) );
  OAI222_X1 U18127 ( .A1(n16071), .A2(n14608), .B1(n14616), .B2(n14626), .C1(
        n14854), .C2(n14627), .ZN(P1_U2859) );
  INV_X1 U18128 ( .A(n14617), .ZN(n14621) );
  INV_X1 U18129 ( .A(n14618), .ZN(n14620) );
  AOI21_X1 U18130 ( .B1(n14621), .B2(n14620), .A(n14619), .ZN(n16008) );
  INV_X1 U18131 ( .A(n16008), .ZN(n14709) );
  INV_X1 U18132 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15968) );
  NOR2_X1 U18133 ( .A1(n14623), .A2(n14622), .ZN(n14624) );
  OR2_X1 U18134 ( .A1(n14625), .A2(n14624), .ZN(n15969) );
  OAI222_X1 U18135 ( .A1(n14709), .A2(n14627), .B1(n15968), .B2(n14626), .C1(
        n15969), .C2(n14608), .ZN(P1_U2860) );
  NAND2_X1 U18136 ( .A1(n14716), .A2(n15988), .ZN(n14633) );
  INV_X1 U18137 ( .A(DATAI_14_), .ZN(n14630) );
  MUX2_X1 U18138 ( .A(n14630), .B(n14629), .S(n14628), .Z(n20134) );
  OAI22_X1 U18139 ( .A1(n15984), .A2(n20134), .B1(n13304), .B2(n14704), .ZN(
        n14631) );
  AOI21_X1 U18140 ( .B1(n15987), .B2(DATAI_30_), .A(n14631), .ZN(n14632) );
  OAI211_X1 U18141 ( .C1(n15992), .C2(n21113), .A(n14633), .B(n14632), .ZN(
        P1_U2874) );
  OAI22_X1 U18142 ( .A1(n15984), .A2(n14703), .B1(n14634), .B2(n14704), .ZN(
        n14635) );
  AOI21_X1 U18143 ( .B1(n15987), .B2(DATAI_29_), .A(n14635), .ZN(n14637) );
  NAND2_X1 U18144 ( .A1(n14689), .A2(BUF1_REG_29__SCAN_IN), .ZN(n14636) );
  OAI211_X1 U18145 ( .C1(n14725), .C2(n14708), .A(n14637), .B(n14636), .ZN(
        P1_U2875) );
  INV_X1 U18146 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16497) );
  NAND2_X1 U18147 ( .A1(n14737), .A2(n15988), .ZN(n14641) );
  OAI22_X1 U18148 ( .A1(n15984), .A2(n14707), .B1(n14638), .B2(n14704), .ZN(
        n14639) );
  AOI21_X1 U18149 ( .B1(n15987), .B2(DATAI_28_), .A(n14639), .ZN(n14640) );
  OAI211_X1 U18150 ( .C1(n15992), .C2(n16497), .A(n14641), .B(n14640), .ZN(
        P1_U2876) );
  OAI22_X1 U18151 ( .A1(n15984), .A2(n14643), .B1(n14642), .B2(n14704), .ZN(
        n14644) );
  AOI21_X1 U18152 ( .B1(n15987), .B2(DATAI_27_), .A(n14644), .ZN(n14646) );
  NAND2_X1 U18153 ( .A1(n14689), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14645) );
  OAI211_X1 U18154 ( .C1(n14647), .C2(n14708), .A(n14646), .B(n14645), .ZN(
        P1_U2877) );
  OAI22_X1 U18155 ( .A1(n15984), .A2(n20131), .B1(n14648), .B2(n14704), .ZN(
        n14649) );
  AOI21_X1 U18156 ( .B1(n15987), .B2(DATAI_26_), .A(n14649), .ZN(n14651) );
  NAND2_X1 U18157 ( .A1(n14689), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14650) );
  OAI211_X1 U18158 ( .C1(n14652), .C2(n14708), .A(n14651), .B(n14650), .ZN(
        P1_U2878) );
  OAI22_X1 U18159 ( .A1(n15984), .A2(n20128), .B1(n14653), .B2(n14704), .ZN(
        n14654) );
  AOI21_X1 U18160 ( .B1(n15987), .B2(DATAI_25_), .A(n14654), .ZN(n14656) );
  NAND2_X1 U18161 ( .A1(n14689), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14655) );
  OAI211_X1 U18162 ( .C1(n15893), .C2(n14708), .A(n14656), .B(n14655), .ZN(
        P1_U2879) );
  OAI22_X1 U18163 ( .A1(n15984), .A2(n20125), .B1(n13063), .B2(n14704), .ZN(
        n14657) );
  AOI21_X1 U18164 ( .B1(n15987), .B2(DATAI_24_), .A(n14657), .ZN(n14659) );
  NAND2_X1 U18165 ( .A1(n14689), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14658) );
  OAI211_X1 U18166 ( .C1(n14774), .C2(n14708), .A(n14659), .B(n14658), .ZN(
        P1_U2880) );
  OAI22_X1 U18167 ( .A1(n15984), .A2(n14661), .B1(n14660), .B2(n14704), .ZN(
        n14662) );
  AOI21_X1 U18168 ( .B1(n15987), .B2(DATAI_23_), .A(n14662), .ZN(n14664) );
  NAND2_X1 U18169 ( .A1(n14689), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14663) );
  OAI211_X1 U18170 ( .C1(n14665), .C2(n14708), .A(n14664), .B(n14663), .ZN(
        P1_U2881) );
  INV_X1 U18171 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14671) );
  NAND2_X1 U18172 ( .A1(n15922), .A2(n15988), .ZN(n14670) );
  OAI22_X1 U18173 ( .A1(n15984), .A2(n14667), .B1(n14666), .B2(n14704), .ZN(
        n14668) );
  AOI21_X1 U18174 ( .B1(n15987), .B2(DATAI_22_), .A(n14668), .ZN(n14669) );
  OAI211_X1 U18175 ( .C1(n15992), .C2(n14671), .A(n14670), .B(n14669), .ZN(
        P1_U2882) );
  OAI22_X1 U18176 ( .A1(n15984), .A2(n14672), .B1(n21096), .B2(n14704), .ZN(
        n14673) );
  AOI21_X1 U18177 ( .B1(n15987), .B2(DATAI_21_), .A(n14673), .ZN(n14675) );
  NAND2_X1 U18178 ( .A1(n14689), .A2(BUF1_REG_21__SCAN_IN), .ZN(n14674) );
  OAI211_X1 U18179 ( .C1(n14803), .C2(n14708), .A(n14675), .B(n14674), .ZN(
        P1_U2883) );
  OAI22_X1 U18180 ( .A1(n15984), .A2(n14677), .B1(n14676), .B2(n14704), .ZN(
        n14678) );
  AOI21_X1 U18181 ( .B1(n15987), .B2(DATAI_20_), .A(n14678), .ZN(n14680) );
  NAND2_X1 U18182 ( .A1(n14689), .A2(BUF1_REG_20__SCAN_IN), .ZN(n14679) );
  OAI211_X1 U18183 ( .C1(n14681), .C2(n14708), .A(n14680), .B(n14679), .ZN(
        P1_U2884) );
  OAI22_X1 U18184 ( .A1(n15984), .A2(n14682), .B1(n13307), .B2(n14704), .ZN(
        n14683) );
  AOI21_X1 U18185 ( .B1(n15987), .B2(DATAI_19_), .A(n14683), .ZN(n14685) );
  NAND2_X1 U18186 ( .A1(n14689), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14684) );
  OAI211_X1 U18187 ( .C1(n15935), .C2(n14708), .A(n14685), .B(n14684), .ZN(
        P1_U2885) );
  OAI22_X1 U18188 ( .A1(n15984), .A2(n14687), .B1(n14686), .B2(n14704), .ZN(
        n14688) );
  AOI21_X1 U18189 ( .B1(n15987), .B2(DATAI_17_), .A(n14688), .ZN(n14691) );
  NAND2_X1 U18190 ( .A1(n14689), .A2(BUF1_REG_17__SCAN_IN), .ZN(n14690) );
  OAI211_X1 U18191 ( .C1(n14692), .C2(n14708), .A(n14691), .B(n14690), .ZN(
        P1_U2887) );
  NAND2_X1 U18192 ( .A1(n15998), .A2(n15988), .ZN(n14697) );
  OAI22_X1 U18193 ( .A1(n15984), .A2(n14694), .B1(n14693), .B2(n14704), .ZN(
        n14695) );
  AOI21_X1 U18194 ( .B1(n15987), .B2(DATAI_16_), .A(n14695), .ZN(n14696) );
  OAI211_X1 U18195 ( .C1(n15992), .C2(n21083), .A(n14697), .B(n14696), .ZN(
        P1_U2888) );
  OAI222_X1 U18196 ( .A1(n14836), .A2(n14708), .B1(n14706), .B2(n14699), .C1(
        n14704), .C2(n14698), .ZN(P1_U2889) );
  INV_X1 U18197 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14700) );
  OAI222_X1 U18198 ( .A1(n14701), .A2(n14708), .B1(n20134), .B2(n14706), .C1(
        n14700), .C2(n14704), .ZN(P1_U2890) );
  OAI222_X1 U18199 ( .A1(n14854), .A2(n14708), .B1(n14703), .B2(n14706), .C1(
        n14702), .C2(n14704), .ZN(P1_U2891) );
  OAI222_X1 U18200 ( .A1(n14709), .A2(n14708), .B1(n14707), .B2(n14706), .C1(
        n14705), .C2(n14704), .ZN(P1_U2892) );
  NAND2_X1 U18201 ( .A1(n14711), .A2(n14710), .ZN(n14712) );
  XNOR2_X1 U18202 ( .A(n14712), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14875) );
  NAND2_X1 U18203 ( .A1(n20164), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14868) );
  NAND2_X1 U18204 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14713) );
  OAI211_X1 U18205 ( .C1(n20163), .C2(n14714), .A(n14868), .B(n14713), .ZN(
        n14715) );
  AOI21_X1 U18206 ( .B1(n14716), .B2(n20159), .A(n14715), .ZN(n14717) );
  OAI21_X1 U18207 ( .B1(n14875), .B2(n19999), .A(n14717), .ZN(P1_U2969) );
  NOR2_X1 U18208 ( .A1(n20208), .A2(n20833), .ZN(n14878) );
  NOR2_X1 U18209 ( .A1(n14805), .A2(n14718), .ZN(n14719) );
  AOI211_X1 U18210 ( .C1(n14720), .C2(n20171), .A(n14878), .B(n14719), .ZN(
        n14724) );
  NAND2_X1 U18211 ( .A1(n14876), .A2(n20169), .ZN(n14723) );
  OAI211_X1 U18212 ( .C1(n14725), .C2(n20175), .A(n14724), .B(n14723), .ZN(
        P1_U2970) );
  INV_X1 U18213 ( .A(n14726), .ZN(n14770) );
  INV_X1 U18214 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14907) );
  NAND3_X1 U18215 ( .A1(n14727), .A2(n14907), .A3(n14898), .ZN(n14728) );
  OR4_X1 U18216 ( .A1(n14729), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A4(n14728), .ZN(n14731) );
  NAND3_X1 U18217 ( .A1(n14729), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14730) );
  MUX2_X1 U18218 ( .A(n14731), .B(n14730), .S(n16013), .Z(n14733) );
  XNOR2_X1 U18219 ( .A(n14733), .B(n14732), .ZN(n14896) );
  NAND2_X1 U18220 ( .A1(n20164), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14892) );
  NAND2_X1 U18221 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14734) );
  OAI211_X1 U18222 ( .C1(n20163), .C2(n14735), .A(n14892), .B(n14734), .ZN(
        n14736) );
  AOI21_X1 U18223 ( .B1(n14737), .B2(n20159), .A(n14736), .ZN(n14738) );
  OAI21_X1 U18224 ( .B1(n19999), .B2(n14896), .A(n14738), .ZN(P1_U2971) );
  INV_X1 U18225 ( .A(n14739), .ZN(n14742) );
  INV_X1 U18226 ( .A(n14740), .ZN(n14741) );
  MUX2_X1 U18227 ( .A(n14742), .B(n14741), .S(n14858), .Z(n14743) );
  XNOR2_X1 U18228 ( .A(n14743), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14906) );
  NAND2_X1 U18229 ( .A1(n14744), .A2(n20159), .ZN(n14749) );
  NOR2_X1 U18230 ( .A1(n20208), .A2(n20828), .ZN(n14897) );
  INV_X1 U18231 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14745) );
  NOR2_X1 U18232 ( .A1(n14805), .A2(n14745), .ZN(n14746) );
  AOI211_X1 U18233 ( .C1(n20171), .C2(n14747), .A(n14897), .B(n14746), .ZN(
        n14748) );
  OAI211_X1 U18234 ( .C1(n14906), .C2(n19999), .A(n14749), .B(n14748), .ZN(
        P1_U2972) );
  INV_X1 U18235 ( .A(n14750), .ZN(n14908) );
  NAND2_X1 U18236 ( .A1(n14726), .A2(n14908), .ZN(n14751) );
  NAND2_X1 U18237 ( .A1(n14751), .A2(n12766), .ZN(n14752) );
  NAND2_X1 U18238 ( .A1(n14753), .A2(n14752), .ZN(n14754) );
  XNOR2_X1 U18239 ( .A(n14754), .B(n14907), .ZN(n14918) );
  INV_X1 U18240 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14755) );
  NOR2_X1 U18241 ( .A1(n20208), .A2(n14755), .ZN(n14911) );
  AOI21_X1 U18242 ( .B1(n20165), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14911), .ZN(n14756) );
  OAI21_X1 U18243 ( .B1(n20163), .B2(n14757), .A(n14756), .ZN(n14758) );
  AOI21_X1 U18244 ( .B1(n14759), .B2(n20159), .A(n14758), .ZN(n14760) );
  OAI21_X1 U18245 ( .B1(n19999), .B2(n14918), .A(n14760), .ZN(P1_U2973) );
  MUX2_X1 U18246 ( .A(n14761), .B(n14930), .S(n16013), .Z(n14764) );
  NAND2_X1 U18247 ( .A1(n14762), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14771) );
  AND2_X1 U18248 ( .A1(n14771), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14763) );
  NOR2_X1 U18249 ( .A1(n14764), .A2(n14763), .ZN(n14765) );
  XNOR2_X1 U18250 ( .A(n14765), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14924) );
  INV_X1 U18251 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14766) );
  NAND2_X1 U18252 ( .A1(n20164), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14919) );
  OAI21_X1 U18253 ( .B1(n14805), .B2(n14766), .A(n14919), .ZN(n14768) );
  NOR2_X1 U18254 ( .A1(n15893), .A2(n20175), .ZN(n14767) );
  AOI211_X1 U18255 ( .C1(n20171), .C2(n15895), .A(n14768), .B(n14767), .ZN(
        n14769) );
  OAI21_X1 U18256 ( .B1(n19999), .B2(n14924), .A(n14769), .ZN(P1_U2974) );
  NAND2_X1 U18257 ( .A1(n14771), .A2(n14770), .ZN(n14772) );
  MUX2_X1 U18258 ( .A(n14772), .B(n14771), .S(n12766), .Z(n14773) );
  XNOR2_X1 U18259 ( .A(n14773), .B(n14930), .ZN(n14936) );
  INV_X1 U18260 ( .A(n14774), .ZN(n15909) );
  NOR2_X1 U18261 ( .A1(n20208), .A2(n20822), .ZN(n14925) );
  AOI21_X1 U18262 ( .B1(n20165), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14925), .ZN(n14775) );
  OAI21_X1 U18263 ( .B1(n20163), .B2(n15911), .A(n14775), .ZN(n14776) );
  AOI21_X1 U18264 ( .B1(n15909), .B2(n20159), .A(n14776), .ZN(n14777) );
  OAI21_X1 U18265 ( .B1(n19999), .B2(n14936), .A(n14777), .ZN(P1_U2975) );
  XNOR2_X1 U18266 ( .A(n12766), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14778) );
  XNOR2_X1 U18267 ( .A(n14726), .B(n14778), .ZN(n14945) );
  NAND2_X1 U18268 ( .A1(n20171), .A2(n14779), .ZN(n14780) );
  NAND2_X1 U18269 ( .A1(n20164), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14939) );
  OAI211_X1 U18270 ( .C1(n14805), .C2(n14781), .A(n14780), .B(n14939), .ZN(
        n14782) );
  AOI21_X1 U18271 ( .B1(n14783), .B2(n20159), .A(n14782), .ZN(n14784) );
  OAI21_X1 U18272 ( .B1(n14945), .B2(n19999), .A(n14784), .ZN(P1_U2976) );
  NAND2_X1 U18273 ( .A1(n14786), .A2(n14785), .ZN(n14787) );
  XNOR2_X1 U18274 ( .A(n14787), .B(n14952), .ZN(n14957) );
  NAND2_X1 U18275 ( .A1(n15922), .A2(n20159), .ZN(n14791) );
  INV_X1 U18276 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14788) );
  NOR2_X1 U18277 ( .A1(n20208), .A2(n14788), .ZN(n14946) );
  NOR2_X1 U18278 ( .A1(n14805), .A2(n15916), .ZN(n14789) );
  AOI211_X1 U18279 ( .C1(n20171), .C2(n15918), .A(n14946), .B(n14789), .ZN(
        n14790) );
  OAI211_X1 U18280 ( .C1(n14957), .C2(n19999), .A(n14791), .B(n14790), .ZN(
        P1_U2977) );
  INV_X1 U18281 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14792) );
  NOR2_X1 U18282 ( .A1(n20208), .A2(n14792), .ZN(n14962) );
  NOR2_X1 U18283 ( .A1(n14805), .A2(n14793), .ZN(n14794) );
  AOI211_X1 U18284 ( .C1(n20171), .C2(n14795), .A(n14962), .B(n14794), .ZN(
        n14802) );
  INV_X1 U18285 ( .A(n14796), .ZN(n14797) );
  NOR2_X1 U18286 ( .A1(n14797), .A2(n14858), .ZN(n14969) );
  OR3_X1 U18287 ( .A1(n14815), .A2(n16013), .A3(n14798), .ZN(n14967) );
  NOR2_X1 U18288 ( .A1(n14967), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14799) );
  AOI21_X1 U18289 ( .B1(n14969), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14799), .ZN(n14800) );
  XNOR2_X1 U18290 ( .A(n14800), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14958) );
  NAND2_X1 U18291 ( .A1(n14958), .A2(n20169), .ZN(n14801) );
  OAI211_X1 U18292 ( .C1(n14803), .C2(n20175), .A(n14802), .B(n14801), .ZN(
        P1_U2978) );
  INV_X1 U18293 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14804) );
  OAI22_X1 U18294 ( .A1(n14805), .A2(n15934), .B1(n20208), .B2(n14804), .ZN(
        n14806) );
  AOI21_X1 U18295 ( .B1(n20171), .B2(n15938), .A(n14806), .ZN(n14812) );
  OAI21_X1 U18296 ( .B1(n12766), .B2(n16055), .A(n14813), .ZN(n14810) );
  XNOR2_X1 U18297 ( .A(n16013), .B(n16045), .ZN(n14809) );
  XNOR2_X1 U18298 ( .A(n14810), .B(n14809), .ZN(n16042) );
  NAND2_X1 U18299 ( .A1(n16042), .A2(n20169), .ZN(n14811) );
  OAI211_X1 U18300 ( .C1(n15935), .C2(n20175), .A(n14812), .B(n14811), .ZN(
        P1_U2980) );
  OAI21_X1 U18301 ( .B1(n14815), .B2(n14814), .A(n14813), .ZN(n16050) );
  INV_X1 U18302 ( .A(n15946), .ZN(n15989) );
  AOI22_X1 U18303 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14816) );
  OAI21_X1 U18304 ( .B1(n20163), .B2(n15943), .A(n14816), .ZN(n14817) );
  AOI21_X1 U18305 ( .B1(n15989), .B2(n20159), .A(n14817), .ZN(n14818) );
  OAI21_X1 U18306 ( .B1(n19999), .B2(n16050), .A(n14818), .ZN(P1_U2981) );
  NAND2_X1 U18307 ( .A1(n14988), .A2(n14823), .ZN(n14824) );
  OAI21_X1 U18308 ( .B1(n14821), .B2(n14820), .A(n14819), .ZN(n14832) );
  INV_X1 U18309 ( .A(n14822), .ZN(n14833) );
  NOR2_X1 U18310 ( .A1(n14832), .A2(n14833), .ZN(n14831) );
  MUX2_X1 U18311 ( .A(n14824), .B(n14823), .S(n14831), .Z(n14825) );
  XOR2_X1 U18312 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n14825), .Z(
        n16058) );
  AOI22_X1 U18313 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n14826) );
  OAI21_X1 U18314 ( .B1(n20163), .B2(n14827), .A(n14826), .ZN(n14828) );
  AOI21_X1 U18315 ( .B1(n14829), .B2(n20159), .A(n14828), .ZN(n14830) );
  OAI21_X1 U18316 ( .B1(n16058), .B2(n19999), .A(n14830), .ZN(P1_U2982) );
  INV_X1 U18317 ( .A(n14831), .ZN(n14986) );
  OAI21_X1 U18318 ( .B1(n14835), .B2(n14833), .A(n14832), .ZN(n14834) );
  OAI21_X1 U18319 ( .B1(n14986), .B2(n14835), .A(n14834), .ZN(n16067) );
  INV_X1 U18320 ( .A(n16067), .ZN(n14842) );
  INV_X1 U18321 ( .A(n14836), .ZN(n14840) );
  AOI22_X1 U18322 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14837) );
  OAI21_X1 U18323 ( .B1(n20163), .B2(n14838), .A(n14837), .ZN(n14839) );
  AOI21_X1 U18324 ( .B1(n14840), .B2(n20159), .A(n14839), .ZN(n14841) );
  OAI21_X1 U18325 ( .B1(n14842), .B2(n19999), .A(n14841), .ZN(P1_U2984) );
  INV_X1 U18326 ( .A(n13810), .ZN(n16014) );
  INV_X1 U18327 ( .A(n14843), .ZN(n14844) );
  AOI21_X1 U18328 ( .B1(n16014), .B2(n14845), .A(n14844), .ZN(n15002) );
  NAND3_X1 U18329 ( .A1(n15002), .A2(n15003), .A3(n14846), .ZN(n15004) );
  NAND2_X1 U18330 ( .A1(n15004), .A2(n15003), .ZN(n14847) );
  XOR2_X1 U18331 ( .A(n14848), .B(n14847), .Z(n16078) );
  NAND2_X1 U18332 ( .A1(n16078), .A2(n20169), .ZN(n14853) );
  INV_X1 U18333 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14849) );
  NOR2_X1 U18334 ( .A1(n20208), .A2(n14849), .ZN(n16072) );
  NOR2_X1 U18335 ( .A1(n20163), .A2(n14850), .ZN(n14851) );
  AOI211_X1 U18336 ( .C1(n20165), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16072), .B(n14851), .ZN(n14852) );
  OAI211_X1 U18337 ( .C1(n20175), .C2(n14854), .A(n14853), .B(n14852), .ZN(
        P1_U2986) );
  NAND2_X1 U18338 ( .A1(n14855), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14857) );
  XNOR2_X1 U18339 ( .A(n13810), .B(n16102), .ZN(n14856) );
  MUX2_X1 U18340 ( .A(n14857), .B(n14856), .S(n16013), .Z(n14860) );
  INV_X1 U18341 ( .A(n14855), .ZN(n14859) );
  NAND3_X1 U18342 ( .A1(n14859), .A2(n14858), .A3(n16102), .ZN(n16015) );
  NAND2_X1 U18343 ( .A1(n14860), .A2(n16015), .ZN(n16100) );
  AOI22_X1 U18344 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14863) );
  NAND2_X1 U18345 ( .A1(n20171), .A2(n14861), .ZN(n14862) );
  OAI211_X1 U18346 ( .C1(n14864), .C2(n20175), .A(n14863), .B(n14862), .ZN(
        n14865) );
  AOI21_X1 U18347 ( .B1(n16100), .B2(n20169), .A(n14865), .ZN(n14866) );
  INV_X1 U18348 ( .A(n14866), .ZN(P1_U2989) );
  INV_X1 U18349 ( .A(n14867), .ZN(n14873) );
  INV_X1 U18350 ( .A(n14868), .ZN(n14872) );
  AOI21_X1 U18351 ( .B1(n12784), .B2(n14870), .A(n14869), .ZN(n14871) );
  AOI211_X1 U18352 ( .C1(n20186), .C2(n14873), .A(n14872), .B(n14871), .ZN(
        n14874) );
  OAI21_X1 U18353 ( .B1(n14875), .B2(n16049), .A(n14874), .ZN(P1_U3001) );
  INV_X1 U18354 ( .A(n14876), .ZN(n14885) );
  NAND3_X1 U18355 ( .A1(n14899), .A2(n14888), .A3(n14877), .ZN(n14880) );
  INV_X1 U18356 ( .A(n14878), .ZN(n14879) );
  OAI211_X1 U18357 ( .C1(n14881), .C2(n20224), .A(n14880), .B(n14879), .ZN(
        n14882) );
  AOI21_X1 U18358 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14883), .A(
        n14882), .ZN(n14884) );
  OAI21_X1 U18359 ( .B1(n14885), .B2(n16049), .A(n14884), .ZN(P1_U3002) );
  NOR2_X1 U18360 ( .A1(n14887), .A2(n14886), .ZN(n14904) );
  INV_X1 U18361 ( .A(n14888), .ZN(n14889) );
  NAND3_X1 U18362 ( .A1(n14899), .A2(n14890), .A3(n14889), .ZN(n14891) );
  OAI211_X1 U18363 ( .C1(n14893), .C2(n20224), .A(n14892), .B(n14891), .ZN(
        n14894) );
  AOI21_X1 U18364 ( .B1(n14904), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14894), .ZN(n14895) );
  OAI21_X1 U18365 ( .B1(n14896), .B2(n16049), .A(n14895), .ZN(P1_U3003) );
  INV_X1 U18366 ( .A(n14897), .ZN(n14901) );
  NAND2_X1 U18367 ( .A1(n14899), .A2(n14898), .ZN(n14900) );
  OAI211_X1 U18368 ( .C1(n14902), .C2(n20224), .A(n14901), .B(n14900), .ZN(
        n14903) );
  AOI21_X1 U18369 ( .B1(n14904), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14903), .ZN(n14905) );
  OAI21_X1 U18370 ( .B1(n14906), .B2(n16049), .A(n14905), .ZN(P1_U3004) );
  NAND2_X1 U18371 ( .A1(n14908), .A2(n14907), .ZN(n14915) );
  NOR2_X1 U18372 ( .A1(n14909), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14920) );
  OAI21_X1 U18373 ( .B1(n14922), .B2(n14920), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14914) );
  INV_X1 U18374 ( .A(n14910), .ZN(n14912) );
  AOI21_X1 U18375 ( .B1(n14912), .B2(n20186), .A(n14911), .ZN(n14913) );
  OAI211_X1 U18376 ( .C1(n14937), .C2(n14915), .A(n14914), .B(n14913), .ZN(
        n14916) );
  INV_X1 U18377 ( .A(n14916), .ZN(n14917) );
  OAI21_X1 U18378 ( .B1(n14918), .B2(n16049), .A(n14917), .ZN(P1_U3005) );
  OAI21_X1 U18379 ( .B1(n15892), .B2(n20224), .A(n14919), .ZN(n14921) );
  AOI211_X1 U18380 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n14922), .A(
        n14921), .B(n14920), .ZN(n14923) );
  OAI21_X1 U18381 ( .B1(n14924), .B2(n16049), .A(n14923), .ZN(P1_U3006) );
  AOI21_X1 U18382 ( .B1(n14926), .B2(n20186), .A(n14925), .ZN(n14935) );
  INV_X1 U18383 ( .A(n14927), .ZN(n14943) );
  AOI21_X1 U18384 ( .B1(n14929), .B2(n16116), .A(n14928), .ZN(n14933) );
  OAI21_X1 U18385 ( .B1(n14937), .B2(n14931), .A(n14930), .ZN(n14932) );
  OAI21_X1 U18386 ( .B1(n14943), .B2(n14933), .A(n14932), .ZN(n14934) );
  OAI211_X1 U18387 ( .C1(n14936), .C2(n16049), .A(n14935), .B(n14934), .ZN(
        P1_U3007) );
  NOR2_X1 U18388 ( .A1(n14937), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14942) );
  INV_X1 U18389 ( .A(n14938), .ZN(n14940) );
  OAI21_X1 U18390 ( .B1(n14940), .B2(n20224), .A(n14939), .ZN(n14941) );
  AOI211_X1 U18391 ( .C1(n14943), .C2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14942), .B(n14941), .ZN(n14944) );
  OAI21_X1 U18392 ( .B1(n14945), .B2(n16049), .A(n14944), .ZN(P1_U3008) );
  INV_X1 U18393 ( .A(n14946), .ZN(n14947) );
  OAI21_X1 U18394 ( .B1(n15924), .B2(n20224), .A(n14947), .ZN(n14955) );
  NAND2_X1 U18395 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14948), .ZN(
        n16070) );
  NAND3_X1 U18396 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14949), .A3(
        n16056), .ZN(n16046) );
  INV_X1 U18397 ( .A(n16046), .ZN(n14950) );
  NAND3_X1 U18398 ( .A1(n14950), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14966) );
  AOI211_X1 U18399 ( .C1(n14953), .C2(n14952), .A(n14951), .B(n14966), .ZN(
        n14954) );
  AOI211_X1 U18400 ( .C1(n14963), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n14955), .B(n14954), .ZN(n14956) );
  OAI21_X1 U18401 ( .B1(n14957), .B2(n16049), .A(n14956), .ZN(P1_U3009) );
  NAND2_X1 U18402 ( .A1(n14958), .A2(n20228), .ZN(n14965) );
  INV_X1 U18403 ( .A(n14959), .ZN(n14960) );
  NOR2_X1 U18404 ( .A1(n14960), .A2(n20224), .ZN(n14961) );
  AOI211_X1 U18405 ( .C1(n14963), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14962), .B(n14961), .ZN(n14964) );
  OAI211_X1 U18406 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n14966), .A(
        n14965), .B(n14964), .ZN(P1_U3010) );
  INV_X1 U18407 ( .A(n14967), .ZN(n14968) );
  OR2_X1 U18408 ( .A1(n14969), .A2(n14968), .ZN(n14971) );
  XNOR2_X1 U18409 ( .A(n14971), .B(n14970), .ZN(n15993) );
  INV_X1 U18410 ( .A(n15993), .ZN(n14984) );
  INV_X1 U18411 ( .A(n14972), .ZN(n14976) );
  NOR2_X1 U18412 ( .A1(n20233), .A2(n14973), .ZN(n14975) );
  NOR2_X1 U18413 ( .A1(n16089), .A2(n12770), .ZN(n14974) );
  OAI221_X1 U18414 ( .B1(n14976), .B2(n16074), .C1(n14976), .C2(n14975), .A(
        n14974), .ZN(n16075) );
  AOI21_X1 U18415 ( .B1(n16095), .B2(n14978), .A(n14977), .ZN(n16044) );
  OAI221_X1 U18416 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16075), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n20231), .A(n16044), .ZN(
        n14982) );
  INV_X1 U18417 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14979) );
  OAI22_X1 U18418 ( .A1(n15931), .A2(n20224), .B1(n20208), .B2(n14979), .ZN(
        n14981) );
  NOR3_X1 U18419 ( .A1(n16046), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n16045), .ZN(n14980) );
  AOI211_X1 U18420 ( .C1(n14982), .C2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14981), .B(n14980), .ZN(n14983) );
  OAI21_X1 U18421 ( .B1(n14984), .B2(n16049), .A(n14983), .ZN(P1_U3011) );
  INV_X1 U18422 ( .A(n14985), .ZN(n14987) );
  OAI22_X1 U18423 ( .A1(n14989), .A2(n14988), .B1(n14987), .B2(n14986), .ZN(
        n15999) );
  NAND2_X1 U18424 ( .A1(n15999), .A2(n20228), .ZN(n14997) );
  AOI21_X1 U18425 ( .B1(n14990), .B2(n14992), .A(n16057), .ZN(n14995) );
  INV_X1 U18426 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14993) );
  OAI21_X1 U18427 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n20215), .A(
        n16082), .ZN(n16065) );
  INV_X1 U18428 ( .A(n16065), .ZN(n14991) );
  OAI22_X1 U18429 ( .A1(n20208), .A2(n14993), .B1(n14992), .B2(n14991), .ZN(
        n14994) );
  AOI21_X1 U18430 ( .B1(n14995), .B2(n16056), .A(n14994), .ZN(n14996) );
  OAI211_X1 U18431 ( .C1(n20224), .C2(n15951), .A(n14997), .B(n14996), .ZN(
        P1_U3015) );
  INV_X1 U18432 ( .A(n14998), .ZN(n15001) );
  AOI21_X1 U18433 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16086), .A(
        n16116), .ZN(n14999) );
  INV_X1 U18434 ( .A(n20218), .ZN(n16112) );
  AOI211_X1 U18435 ( .C1(n16114), .C2(n15000), .A(n14999), .B(n16112), .ZN(
        n16090) );
  OAI21_X1 U18436 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15001), .A(
        n16090), .ZN(n15010) );
  NAND3_X1 U18437 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16086), .A3(
        n12770), .ZN(n15008) );
  INV_X1 U18438 ( .A(n15002), .ZN(n15007) );
  OAI21_X1 U18439 ( .B1(n12770), .B2(n16013), .A(n15003), .ZN(n15006) );
  INV_X1 U18440 ( .A(n15004), .ZN(n15005) );
  AOI21_X1 U18441 ( .B1(n15007), .B2(n15006), .A(n15005), .ZN(n16012) );
  OAI22_X1 U18442 ( .A1(n16135), .A2(n15008), .B1(n16012), .B2(n16049), .ZN(
        n15009) );
  AOI21_X1 U18443 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15010), .A(
        n15009), .ZN(n15012) );
  NAND2_X1 U18444 ( .A1(n20164), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15011) );
  OAI211_X1 U18445 ( .C1(n20224), .C2(n15969), .A(n15012), .B(n15011), .ZN(
        P1_U3019) );
  INV_X1 U18446 ( .A(n15013), .ZN(n15015) );
  OAI22_X1 U18447 ( .A1(n15017), .A2(n15016), .B1(n15015), .B2(n15014), .ZN(
        n15018) );
  MUX2_X1 U18448 ( .A(n15019), .B(n15018), .S(n16151), .Z(P1_U3469) );
  INV_X1 U18449 ( .A(n15020), .ZN(n16181) );
  AOI21_X1 U18450 ( .B1(n15321), .B2(n15045), .A(n15046), .ZN(n15324) );
  INV_X1 U18451 ( .A(n15324), .ZN(n16217) );
  AOI21_X1 U18452 ( .B1(n15339), .B2(n15041), .A(n15043), .ZN(n15341) );
  INV_X1 U18453 ( .A(n15341), .ZN(n18996) );
  INV_X1 U18454 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15021) );
  XNOR2_X1 U18455 ( .A(n15039), .B(n15021), .ZN(n15379) );
  AND2_X1 U18456 ( .A1(n15034), .A2(n15398), .ZN(n15022) );
  OR2_X1 U18457 ( .A1(n15022), .A2(n15037), .ZN(n15104) );
  INV_X1 U18458 ( .A(n15104), .ZN(n15396) );
  OR2_X1 U18459 ( .A1(n15032), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15023) );
  NAND2_X1 U18460 ( .A1(n15036), .A2(n15023), .ZN(n15419) );
  INV_X1 U18461 ( .A(n15419), .ZN(n19053) );
  OAI21_X1 U18462 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15029), .A(
        n15031), .ZN(n16271) );
  INV_X1 U18463 ( .A(n16271), .ZN(n19076) );
  OAI21_X1 U18464 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n15026), .A(
        n15030), .ZN(n19108) );
  INV_X1 U18465 ( .A(n19108), .ZN(n15028) );
  INV_X1 U18466 ( .A(n16313), .ZN(n15025) );
  NOR2_X1 U18467 ( .A1(n15025), .A2(n15024), .ZN(n19114) );
  AOI21_X1 U18468 ( .B1(n16298), .B2(n15027), .A(n15026), .ZN(n16290) );
  INV_X1 U18469 ( .A(n16290), .ZN(n19115) );
  NAND2_X1 U18470 ( .A1(n19114), .A2(n19115), .ZN(n19106) );
  NOR2_X1 U18471 ( .A1(n15028), .A2(n19106), .ZN(n19098) );
  AOI21_X1 U18472 ( .B1(n19085), .B2(n15030), .A(n15029), .ZN(n16272) );
  INV_X1 U18473 ( .A(n16272), .ZN(n19101) );
  NAND2_X1 U18474 ( .A1(n19098), .A2(n19101), .ZN(n19074) );
  NOR2_X1 U18475 ( .A1(n19076), .A2(n19074), .ZN(n19063) );
  AND2_X1 U18476 ( .A1(n15031), .A2(n15429), .ZN(n15033) );
  OR2_X1 U18477 ( .A1(n15033), .A2(n15032), .ZN(n19068) );
  NAND2_X1 U18478 ( .A1(n19063), .A2(n19068), .ZN(n19052) );
  NOR2_X1 U18479 ( .A1(n19053), .A2(n19052), .ZN(n19040) );
  INV_X1 U18480 ( .A(n15034), .ZN(n15035) );
  AOI21_X1 U18481 ( .B1(n15409), .B2(n15036), .A(n15035), .ZN(n15407) );
  INV_X1 U18482 ( .A(n15407), .ZN(n19041) );
  NAND2_X1 U18483 ( .A1(n19040), .A2(n19041), .ZN(n15102) );
  NOR2_X1 U18484 ( .A1(n15396), .A2(n15102), .ZN(n19036) );
  NOR2_X1 U18485 ( .A1(n15037), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15038) );
  OR2_X1 U18486 ( .A1(n15039), .A2(n15038), .ZN(n19035) );
  NAND2_X1 U18487 ( .A1(n19036), .A2(n19035), .ZN(n15086) );
  NOR2_X1 U18488 ( .A1(n15379), .A2(n15086), .ZN(n19011) );
  AOI21_X1 U18489 ( .B1(n15039), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15040) );
  OR2_X1 U18490 ( .A1(n15042), .A2(n15040), .ZN(n19013) );
  NAND2_X1 U18491 ( .A1(n19011), .A2(n19013), .ZN(n19001) );
  OAI21_X1 U18492 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15042), .A(
        n15041), .ZN(n15353) );
  INV_X1 U18493 ( .A(n15353), .ZN(n19004) );
  OAI21_X1 U18494 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n15043), .A(
        n15044), .ZN(n16265) );
  NAND2_X1 U18495 ( .A1(n15829), .A2(n16265), .ZN(n15828) );
  NAND2_X1 U18496 ( .A1(n19075), .A2(n15828), .ZN(n16230) );
  AOI21_X1 U18497 ( .B1(n9925), .B2(n15044), .A(n9877), .ZN(n16251) );
  INV_X1 U18498 ( .A(n16251), .ZN(n16231) );
  OAI21_X1 U18499 ( .B1(n9877), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15045), .ZN(n15334) );
  OR2_X1 U18500 ( .A1(n15046), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15047) );
  NAND2_X1 U18501 ( .A1(n15048), .A2(n15047), .ZN(n16206) );
  NAND2_X1 U18502 ( .A1(n19075), .A2(n16204), .ZN(n16193) );
  INV_X1 U18503 ( .A(n15049), .ZN(n16194) );
  XNOR2_X1 U18504 ( .A(n15050), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15299) );
  OAI211_X1 U18505 ( .C1(n15051), .C2(n15299), .A(n19154), .B(n16174), .ZN(
        n15057) );
  AOI22_X1 U18506 ( .A1(n19128), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19145), .ZN(n15052) );
  INV_X1 U18507 ( .A(n15052), .ZN(n15055) );
  INV_X1 U18508 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15053) );
  NAND2_X1 U18509 ( .A1(n15059), .A2(n19109), .ZN(n15069) );
  OAI22_X1 U18510 ( .A1(n19143), .A2(n10506), .B1(n19907), .B2(n19133), .ZN(
        n15061) );
  NOR2_X1 U18511 ( .A1(n19158), .A2(n13979), .ZN(n15060) );
  AOI211_X1 U18512 ( .C1(n15233), .C2(n19089), .A(n15061), .B(n15060), .ZN(
        n15068) );
  OAI211_X1 U18513 ( .C1(n15064), .C2(n15063), .A(n19154), .B(n15062), .ZN(
        n15067) );
  NAND2_X1 U18514 ( .A1(n15065), .A2(n19129), .ZN(n15066) );
  NAND4_X1 U18515 ( .A1(n15069), .A2(n15068), .A3(n15067), .A4(n15066), .ZN(
        P2_U2827) );
  INV_X1 U18516 ( .A(n15070), .ZN(n15071) );
  OAI21_X1 U18517 ( .B1(n15166), .B2(n15072), .A(n15071), .ZN(n15468) );
  NAND2_X1 U18518 ( .A1(n15267), .A2(n15073), .ZN(n15074) );
  NAND2_X1 U18519 ( .A1(n15253), .A2(n15074), .ZN(n15475) );
  INV_X1 U18520 ( .A(n15475), .ZN(n15079) );
  INV_X1 U18521 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19899) );
  AOI22_X1 U18522 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19138), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n19128), .ZN(n15075) );
  OAI21_X1 U18523 ( .B1(n19899), .B2(n19133), .A(n15075), .ZN(n15078) );
  AOI211_X1 U18524 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n15076), .A(n19142), .B(
        n16220), .ZN(n15077) );
  AOI211_X1 U18525 ( .C1(n19089), .C2(n15079), .A(n15078), .B(n15077), .ZN(
        n15083) );
  OAI211_X1 U18526 ( .C1(n15081), .C2(n15334), .A(n19154), .B(n15080), .ZN(
        n15082) );
  OAI211_X1 U18527 ( .C1(n15468), .C2(n19151), .A(n15083), .B(n15082), .ZN(
        P2_U2831) );
  OR2_X1 U18528 ( .A1(n15206), .A2(n15084), .ZN(n15085) );
  NAND2_X1 U18529 ( .A1(n15191), .A2(n15085), .ZN(n15549) );
  INV_X1 U18530 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15378) );
  INV_X1 U18531 ( .A(n15086), .ZN(n15096) );
  OAI211_X1 U18532 ( .C1(n15096), .C2(n19147), .A(n19154), .B(n15379), .ZN(
        n15093) );
  NAND2_X1 U18533 ( .A1(n15289), .A2(n15088), .ZN(n15089) );
  AND2_X1 U18534 ( .A1(n15280), .A2(n15089), .ZN(n16245) );
  AOI22_X1 U18535 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19138), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19128), .ZN(n15090) );
  NAND2_X1 U18536 ( .A1(n19131), .A2(n15090), .ZN(n15091) );
  AOI21_X1 U18537 ( .B1(n19089), .B2(n16245), .A(n15091), .ZN(n15092) );
  OAI211_X1 U18538 ( .C1(n15378), .C2(n19133), .A(n15093), .B(n15092), .ZN(
        n15094) );
  AOI21_X1 U18539 ( .B1(n15095), .B2(n19129), .A(n15094), .ZN(n15099) );
  NAND2_X1 U18540 ( .A1(n19154), .A2(n19075), .ZN(n16175) );
  NOR2_X1 U18541 ( .A1(n15096), .A2(n16175), .ZN(n19034) );
  INV_X1 U18542 ( .A(n15379), .ZN(n15097) );
  NAND2_X1 U18543 ( .A1(n19034), .A2(n15097), .ZN(n15098) );
  OAI211_X1 U18544 ( .C1(n15549), .C2(n19151), .A(n15099), .B(n15098), .ZN(
        P2_U2837) );
  NAND2_X1 U18545 ( .A1(n15215), .A2(n15100), .ZN(n15101) );
  NAND2_X1 U18546 ( .A1(n9878), .A2(n15101), .ZN(n15395) );
  NAND2_X1 U18547 ( .A1(n19075), .A2(n15102), .ZN(n15103) );
  XOR2_X1 U18548 ( .A(n15104), .B(n15103), .Z(n15105) );
  NAND2_X1 U18549 ( .A1(n15105), .A2(n19154), .ZN(n15114) );
  AND2_X1 U18550 ( .A1(n15107), .A2(n15106), .ZN(n15108) );
  OR2_X1 U18551 ( .A1(n15108), .A2(n9879), .ZN(n19169) );
  AOI22_X1 U18552 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19138), .B1(
        P2_EBX_REG_16__SCAN_IN), .B2(n19128), .ZN(n15109) );
  OAI211_X1 U18553 ( .C1(n19150), .C2(n19169), .A(n15109), .B(n19131), .ZN(
        n15112) );
  NOR2_X1 U18554 ( .A1(n15110), .A2(n19142), .ZN(n15111) );
  AOI211_X1 U18555 ( .C1(n19145), .C2(P2_REIP_REG_16__SCAN_IN), .A(n15112), 
        .B(n15111), .ZN(n15113) );
  OAI211_X1 U18556 ( .C1(n19151), .C2(n15395), .A(n15114), .B(n15113), .ZN(
        P2_U2839) );
  NOR2_X1 U18557 ( .A1(n19147), .A2(n15115), .ZN(n15696) );
  NAND2_X1 U18558 ( .A1(n15696), .A2(n19154), .ZN(n15123) );
  INV_X1 U18559 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18982) );
  OR2_X1 U18560 ( .A1(n19150), .A2(n16359), .ZN(n15117) );
  INV_X1 U18561 ( .A(n19102), .ZN(n19028) );
  OAI21_X1 U18562 ( .B1(n19138), .B2(n19028), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15116) );
  OAI211_X1 U18563 ( .C1(n19133), .C2(n18982), .A(n15117), .B(n15116), .ZN(
        n15121) );
  OAI22_X1 U18564 ( .A1(n19143), .A2(n15119), .B1(n19142), .B2(n15118), .ZN(
        n15120) );
  AOI211_X1 U18565 ( .C1(n15695), .C2(n19109), .A(n15121), .B(n15120), .ZN(
        n15122) );
  OAI211_X1 U18566 ( .C1(n15124), .C2(n18958), .A(n15123), .B(n15122), .ZN(
        P2_U2855) );
  MUX2_X1 U18567 ( .A(n16171), .B(P2_EBX_REG_31__SCAN_IN), .S(n15212), .Z(
        P2_U2856) );
  INV_X1 U18568 ( .A(n15126), .ZN(n15227) );
  NAND2_X1 U18569 ( .A1(n15127), .A2(n15128), .ZN(n15226) );
  NAND3_X1 U18570 ( .A1(n15227), .A2(n15199), .A3(n15226), .ZN(n15130) );
  NAND2_X1 U18571 ( .A1(n15212), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15129) );
  OAI211_X1 U18572 ( .C1(n15212), .C2(n15125), .A(n15130), .B(n15129), .ZN(
        P2_U2858) );
  NAND2_X1 U18573 ( .A1(n9802), .A2(n15131), .ZN(n15133) );
  XNOR2_X1 U18574 ( .A(n15133), .B(n15132), .ZN(n15238) );
  NOR2_X1 U18575 ( .A1(n15134), .A2(n15205), .ZN(n15135) );
  AOI21_X1 U18576 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15205), .A(n15135), .ZN(
        n15136) );
  OAI21_X1 U18577 ( .B1(n15238), .B2(n15219), .A(n15136), .ZN(P2_U2859) );
  AOI21_X1 U18578 ( .B1(n15138), .B2(n15137), .A(n9868), .ZN(n15239) );
  NAND2_X1 U18579 ( .A1(n15239), .A2(n15199), .ZN(n15140) );
  NAND2_X1 U18580 ( .A1(n15212), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15139) );
  OAI211_X1 U18581 ( .C1(n15212), .C2(n16190), .A(n15140), .B(n15139), .ZN(
        P2_U2860) );
  NAND2_X1 U18582 ( .A1(n15141), .A2(n15142), .ZN(n15143) );
  NAND2_X1 U18583 ( .A1(n15144), .A2(n15143), .ZN(n16200) );
  AOI21_X1 U18584 ( .B1(n15147), .B2(n15146), .A(n15145), .ZN(n15245) );
  NAND2_X1 U18585 ( .A1(n15245), .A2(n15199), .ZN(n15149) );
  NAND2_X1 U18586 ( .A1(n15212), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15148) );
  OAI211_X1 U18587 ( .C1(n16200), .C2(n15205), .A(n15149), .B(n15148), .ZN(
        P2_U2861) );
  OAI21_X1 U18588 ( .B1(n15152), .B2(n15151), .A(n15150), .ZN(n15259) );
  OAI21_X1 U18589 ( .B1(n15070), .B2(n15153), .A(n15141), .ZN(n16212) );
  NOR2_X1 U18590 ( .A1(n16212), .A2(n15205), .ZN(n15154) );
  AOI21_X1 U18591 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15205), .A(n15154), .ZN(
        n15155) );
  OAI21_X1 U18592 ( .B1(n15259), .B2(n15219), .A(n15155), .ZN(P2_U2862) );
  AOI21_X1 U18593 ( .B1(n15157), .B2(n15156), .A(n9883), .ZN(n15158) );
  XOR2_X1 U18594 ( .A(n15159), .B(n15158), .Z(n15265) );
  NOR2_X1 U18595 ( .A1(n15468), .A2(n15205), .ZN(n15160) );
  AOI21_X1 U18596 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15205), .A(n15160), .ZN(
        n15161) );
  OAI21_X1 U18597 ( .B1(n15265), .B2(n15219), .A(n15161), .ZN(P2_U2863) );
  AOI21_X1 U18598 ( .B1(n15164), .B2(n15163), .A(n15162), .ZN(n15266) );
  NAND2_X1 U18599 ( .A1(n15266), .A2(n15199), .ZN(n15169) );
  AND2_X1 U18600 ( .A1(n15172), .A2(n15165), .ZN(n15167) );
  NAND2_X1 U18601 ( .A1(n9875), .A2(n15224), .ZN(n15168) );
  OAI211_X1 U18602 ( .C1(n15224), .C2(n10489), .A(n15169), .B(n15168), .ZN(
        P2_U2864) );
  NAND2_X1 U18603 ( .A1(n11604), .A2(n15170), .ZN(n15171) );
  NAND2_X1 U18604 ( .A1(n15172), .A2(n15171), .ZN(n16260) );
  INV_X1 U18605 ( .A(n14178), .ZN(n15174) );
  AOI21_X1 U18606 ( .B1(n15175), .B2(n15173), .A(n15174), .ZN(n16237) );
  NAND2_X1 U18607 ( .A1(n16237), .A2(n15199), .ZN(n15177) );
  NAND2_X1 U18608 ( .A1(n15212), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15176) );
  OAI211_X1 U18609 ( .C1(n16260), .C2(n15205), .A(n15177), .B(n15176), .ZN(
        P2_U2865) );
  OAI21_X1 U18610 ( .B1(n15178), .B2(n15179), .A(n15173), .ZN(n15277) );
  MUX2_X1 U18611 ( .A(n18989), .B(n15180), .S(n15212), .Z(n15181) );
  OAI21_X1 U18612 ( .B1(n15277), .B2(n15219), .A(n15181), .ZN(P2_U2866) );
  AND2_X1 U18613 ( .A1(n15182), .A2(n15183), .ZN(n15184) );
  NOR2_X1 U18614 ( .A1(n15178), .A2(n15184), .ZN(n16241) );
  NAND2_X1 U18615 ( .A1(n16241), .A2(n15199), .ZN(n15188) );
  AND2_X1 U18616 ( .A1(n9819), .A2(n15185), .ZN(n15186) );
  NOR2_X1 U18617 ( .A1(n11605), .A2(n15186), .ZN(n19006) );
  NAND2_X1 U18618 ( .A1(n19006), .A2(n15224), .ZN(n15187) );
  OAI211_X1 U18619 ( .C1(n15224), .C2(n15189), .A(n15188), .B(n15187), .ZN(
        P2_U2867) );
  NAND2_X1 U18620 ( .A1(n15191), .A2(n15190), .ZN(n15192) );
  NAND2_X1 U18621 ( .A1(n9819), .A2(n15192), .ZN(n19021) );
  AOI21_X1 U18622 ( .B1(n15194), .B2(n15193), .A(n10089), .ZN(n15278) );
  NAND2_X1 U18623 ( .A1(n15278), .A2(n15199), .ZN(n15196) );
  NAND2_X1 U18624 ( .A1(n15212), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15195) );
  OAI211_X1 U18625 ( .C1(n19021), .C2(n15205), .A(n15196), .B(n15195), .ZN(
        P2_U2868) );
  AOI21_X1 U18626 ( .B1(n15198), .B2(n15203), .A(n14109), .ZN(n16247) );
  NAND2_X1 U18627 ( .A1(n16247), .A2(n15199), .ZN(n15201) );
  NAND2_X1 U18628 ( .A1(n15205), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15200) );
  OAI211_X1 U18629 ( .C1(n15549), .C2(n15205), .A(n15201), .B(n15200), .ZN(
        P2_U2869) );
  OAI21_X1 U18630 ( .B1(n15202), .B2(n15204), .A(n15203), .ZN(n15296) );
  NAND2_X1 U18631 ( .A1(n15205), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15209) );
  AOI21_X1 U18632 ( .B1(n15207), .B2(n9878), .A(n15206), .ZN(n19033) );
  NAND2_X1 U18633 ( .A1(n19033), .A2(n15224), .ZN(n15208) );
  OAI211_X1 U18634 ( .C1(n15296), .C2(n15219), .A(n15209), .B(n15208), .ZN(
        P2_U2870) );
  NOR2_X1 U18635 ( .A1(n9881), .A2(n15210), .ZN(n15211) );
  OR2_X1 U18636 ( .A1(n15202), .A2(n15211), .ZN(n19172) );
  MUX2_X1 U18637 ( .A(n15395), .B(n15213), .S(n15212), .Z(n15214) );
  OAI21_X1 U18638 ( .B1(n19172), .B2(n15219), .A(n15214), .ZN(P2_U2871) );
  INV_X1 U18639 ( .A(n15215), .ZN(n15216) );
  AOI21_X1 U18640 ( .B1(n15218), .B2(n15217), .A(n15216), .ZN(n19045) );
  NOR2_X1 U18641 ( .A1(n15224), .A2(n10462), .ZN(n15223) );
  AOI211_X1 U18642 ( .C1(n15221), .C2(n15220), .A(n15219), .B(n9881), .ZN(
        n15222) );
  AOI211_X1 U18643 ( .C1(n19045), .C2(n15224), .A(n15223), .B(n15222), .ZN(
        n15225) );
  INV_X1 U18644 ( .A(n15225), .ZN(P2_U2872) );
  NAND3_X1 U18645 ( .A1(n15227), .A2(n19194), .A3(n15226), .ZN(n15232) );
  INV_X1 U18646 ( .A(n15287), .ZN(n19166) );
  AOI22_X1 U18647 ( .A1(n19167), .A2(BUF2_REG_29__SCAN_IN), .B1(n19166), .B2(
        n15228), .ZN(n15231) );
  INV_X1 U18648 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19212) );
  OAI22_X1 U18649 ( .A1(n16177), .A2(n19170), .B1(n15286), .B2(n19212), .ZN(
        n15229) );
  AOI21_X1 U18650 ( .B1(n19168), .B2(BUF1_REG_29__SCAN_IN), .A(n15229), .ZN(
        n15230) );
  NAND3_X1 U18651 ( .A1(n15232), .A2(n15231), .A3(n15230), .ZN(P2_U2890) );
  AOI22_X1 U18652 ( .A1(n19167), .A2(BUF2_REG_28__SCAN_IN), .B1(n16246), .B2(
        n15233), .ZN(n15237) );
  OAI22_X1 U18653 ( .A1(n15234), .A2(n15287), .B1(n15286), .B2(n19214), .ZN(
        n15235) );
  AOI21_X1 U18654 ( .B1(n19168), .B2(BUF1_REG_28__SCAN_IN), .A(n15235), .ZN(
        n15236) );
  OAI211_X1 U18655 ( .C1(n15238), .C2(n19171), .A(n15237), .B(n15236), .ZN(
        P2_U2891) );
  INV_X1 U18656 ( .A(n15239), .ZN(n15244) );
  AOI22_X1 U18657 ( .A1(n19167), .A2(BUF2_REG_27__SCAN_IN), .B1(n19166), .B2(
        n15240), .ZN(n15243) );
  INV_X1 U18658 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19216) );
  OAI22_X1 U18659 ( .A1(n16189), .A2(n19170), .B1(n15286), .B2(n19216), .ZN(
        n15241) );
  AOI21_X1 U18660 ( .B1(n19168), .B2(BUF1_REG_27__SCAN_IN), .A(n15241), .ZN(
        n15242) );
  OAI211_X1 U18661 ( .C1(n15244), .C2(n19171), .A(n15243), .B(n15242), .ZN(
        P2_U2892) );
  INV_X1 U18662 ( .A(n15245), .ZN(n15251) );
  AOI22_X1 U18663 ( .A1(n19167), .A2(BUF2_REG_26__SCAN_IN), .B1(n19166), .B2(
        n19184), .ZN(n15250) );
  OAI21_X1 U18664 ( .B1(n15247), .B2(n15246), .A(n13991), .ZN(n16201) );
  OAI22_X1 U18665 ( .A1(n16201), .A2(n19170), .B1(n15286), .B2(n19218), .ZN(
        n15248) );
  AOI21_X1 U18666 ( .B1(n19168), .B2(BUF1_REG_26__SCAN_IN), .A(n15248), .ZN(
        n15249) );
  OAI211_X1 U18667 ( .C1(n15251), .C2(n19171), .A(n15250), .B(n15249), .ZN(
        P2_U2893) );
  AOI22_X1 U18668 ( .A1(n19167), .A2(BUF2_REG_25__SCAN_IN), .B1(n19166), .B2(
        n15252), .ZN(n15258) );
  XOR2_X1 U18669 ( .A(n15254), .B(n15253), .Z(n16213) );
  INV_X1 U18670 ( .A(n16213), .ZN(n15255) );
  INV_X1 U18671 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19220) );
  OAI22_X1 U18672 ( .A1(n15255), .A2(n19170), .B1(n15286), .B2(n19220), .ZN(
        n15256) );
  AOI21_X1 U18673 ( .B1(n19168), .B2(BUF1_REG_25__SCAN_IN), .A(n15256), .ZN(
        n15257) );
  OAI211_X1 U18674 ( .C1(n15259), .C2(n19171), .A(n15258), .B(n15257), .ZN(
        P2_U2894) );
  OAI22_X1 U18675 ( .A1(n15260), .A2(n15287), .B1(n15286), .B2(n19222), .ZN(
        n15263) );
  INV_X1 U18676 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n15261) );
  OAI22_X1 U18677 ( .A1(n15292), .A2(n15261), .B1(n19170), .B2(n15475), .ZN(
        n15262) );
  AOI211_X1 U18678 ( .C1(n19168), .C2(BUF1_REG_24__SCAN_IN), .A(n15263), .B(
        n15262), .ZN(n15264) );
  OAI21_X1 U18679 ( .B1(n15265), .B2(n19171), .A(n15264), .ZN(P2_U2895) );
  INV_X1 U18680 ( .A(n15266), .ZN(n15272) );
  OAI21_X1 U18681 ( .B1(n15504), .B2(n15268), .A(n15267), .ZN(n16234) );
  INV_X1 U18682 ( .A(n16234), .ZN(n15488) );
  AOI22_X1 U18683 ( .A1(n19167), .A2(BUF2_REG_23__SCAN_IN), .B1(n16246), .B2(
        n15488), .ZN(n15271) );
  INV_X1 U18684 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19224) );
  OAI22_X1 U18685 ( .A1(n19342), .A2(n15287), .B1(n15286), .B2(n19224), .ZN(
        n15269) );
  AOI21_X1 U18686 ( .B1(n19168), .B2(BUF1_REG_23__SCAN_IN), .A(n15269), .ZN(
        n15270) );
  OAI211_X1 U18687 ( .C1(n15272), .C2(n19171), .A(n15271), .B(n15270), .ZN(
        P2_U2896) );
  OAI22_X1 U18688 ( .A1(n15273), .A2(n15287), .B1(n15286), .B2(n19228), .ZN(
        n15275) );
  OAI22_X1 U18689 ( .A1(n19170), .A2(n18999), .B1(n15292), .B2(n18285), .ZN(
        n15274) );
  AOI211_X1 U18690 ( .C1(n19168), .C2(BUF1_REG_21__SCAN_IN), .A(n15275), .B(
        n15274), .ZN(n15276) );
  OAI21_X1 U18691 ( .B1(n15277), .B2(n19171), .A(n15276), .ZN(P2_U2898) );
  INV_X1 U18692 ( .A(n15278), .ZN(n15285) );
  NAND2_X1 U18693 ( .A1(n15280), .A2(n15279), .ZN(n15281) );
  AND2_X1 U18694 ( .A1(n15516), .A2(n15281), .ZN(n19019) );
  AOI22_X1 U18695 ( .A1(n19167), .A2(BUF2_REG_19__SCAN_IN), .B1(n16246), .B2(
        n19019), .ZN(n15284) );
  INV_X1 U18696 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19232) );
  OAI22_X1 U18697 ( .A1(n19320), .A2(n15287), .B1(n15286), .B2(n19232), .ZN(
        n15282) );
  AOI21_X1 U18698 ( .B1(n19168), .B2(BUF1_REG_19__SCAN_IN), .A(n15282), .ZN(
        n15283) );
  OAI211_X1 U18699 ( .C1(n15285), .C2(n19171), .A(n15284), .B(n15283), .ZN(
        P2_U2900) );
  INV_X1 U18700 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n21133) );
  OAI22_X1 U18701 ( .A1(n15288), .A2(n15287), .B1(n15286), .B2(n21133), .ZN(
        n15294) );
  INV_X1 U18702 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15291) );
  OAI21_X1 U18703 ( .B1(n9879), .B2(n15290), .A(n15289), .ZN(n19039) );
  OAI22_X1 U18704 ( .A1(n15292), .A2(n15291), .B1(n19170), .B2(n19039), .ZN(
        n15293) );
  AOI211_X1 U18705 ( .C1(n19168), .C2(BUF1_REG_17__SCAN_IN), .A(n15294), .B(
        n15293), .ZN(n15295) );
  OAI21_X1 U18706 ( .B1(n15296), .B2(n19171), .A(n15295), .ZN(P2_U2902) );
  NAND2_X1 U18707 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15297) );
  OAI211_X1 U18708 ( .C1(n16314), .C2(n15299), .A(n15298), .B(n15297), .ZN(
        n15300) );
  AOI21_X1 U18709 ( .B1(n15301), .B2(n19278), .A(n15300), .ZN(n15304) );
  NAND2_X1 U18710 ( .A1(n15302), .A2(n16310), .ZN(n15303) );
  OAI211_X1 U18711 ( .C1(n15305), .C2(n16292), .A(n15304), .B(n15303), .ZN(
        P2_U2984) );
  NOR2_X1 U18712 ( .A1(n15306), .A2(n15319), .ZN(n15307) );
  XOR2_X1 U18713 ( .A(n15308), .B(n15307), .Z(n15457) );
  AOI21_X1 U18714 ( .B1(n15311), .B2(n15309), .A(n15310), .ZN(n15455) );
  NOR2_X1 U18715 ( .A1(n16200), .A2(n16317), .ZN(n15314) );
  NAND2_X1 U18716 ( .A1(n19088), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15449) );
  NAND2_X1 U18717 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15312) );
  OAI211_X1 U18718 ( .C1(n16314), .C2(n16206), .A(n15449), .B(n15312), .ZN(
        n15313) );
  AOI211_X1 U18719 ( .C1(n15455), .C2(n16287), .A(n15314), .B(n15313), .ZN(
        n15315) );
  OAI21_X1 U18720 ( .B1(n15457), .B2(n16292), .A(n15315), .ZN(P2_U2988) );
  INV_X1 U18721 ( .A(n15306), .ZN(n15320) );
  OAI21_X1 U18722 ( .B1(n15317), .B2(n15319), .A(n15316), .ZN(n15318) );
  OAI21_X1 U18723 ( .B1(n15320), .B2(n15319), .A(n15318), .ZN(n15467) );
  NAND2_X1 U18724 ( .A1(n19088), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15458) );
  OAI21_X1 U18725 ( .B1(n19288), .B2(n15321), .A(n15458), .ZN(n15323) );
  NOR2_X1 U18726 ( .A1(n16212), .A2(n16317), .ZN(n15322) );
  AOI211_X1 U18727 ( .C1(n19274), .C2(n15324), .A(n15323), .B(n15322), .ZN(
        n15328) );
  INV_X1 U18728 ( .A(n15332), .ZN(n15326) );
  NAND2_X1 U18729 ( .A1(n15326), .A2(n15325), .ZN(n15464) );
  NAND3_X1 U18730 ( .A1(n15464), .A2(n16310), .A3(n15309), .ZN(n15327) );
  OAI211_X1 U18731 ( .C1(n15467), .C2(n16292), .A(n15328), .B(n15327), .ZN(
        P2_U2989) );
  XNOR2_X1 U18732 ( .A(n15329), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15330) );
  XNOR2_X1 U18733 ( .A(n15331), .B(n15330), .ZN(n15482) );
  AOI21_X1 U18734 ( .B1(n15474), .B2(n15493), .A(n15332), .ZN(n15479) );
  NOR2_X1 U18735 ( .A1(n15468), .A2(n16317), .ZN(n15336) );
  AOI22_X1 U18736 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19088), .ZN(n15333) );
  OAI21_X1 U18737 ( .B1(n16314), .B2(n15334), .A(n15333), .ZN(n15335) );
  AOI211_X1 U18738 ( .C1(n15479), .C2(n16310), .A(n15336), .B(n15335), .ZN(
        n15337) );
  OAI21_X1 U18739 ( .B1(n15482), .B2(n16292), .A(n15337), .ZN(P2_U2990) );
  OAI21_X1 U18740 ( .B1(n19288), .B2(n15339), .A(n15338), .ZN(n15340) );
  AOI21_X1 U18741 ( .B1(n19274), .B2(n15341), .A(n15340), .ZN(n15342) );
  OAI21_X1 U18742 ( .B1(n18989), .B2(n16317), .A(n15342), .ZN(n15343) );
  AOI21_X1 U18743 ( .B1(n15344), .B2(n16310), .A(n15343), .ZN(n15345) );
  OAI21_X1 U18744 ( .B1(n15346), .B2(n16292), .A(n15345), .ZN(P2_U2993) );
  NAND2_X1 U18745 ( .A1(n15347), .A2(n10234), .ZN(n15351) );
  NAND2_X1 U18746 ( .A1(n15349), .A2(n15348), .ZN(n15350) );
  XNOR2_X1 U18747 ( .A(n15351), .B(n15350), .ZN(n15533) );
  NAND2_X1 U18748 ( .A1(n19088), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15518) );
  NAND2_X1 U18749 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15352) );
  OAI211_X1 U18750 ( .C1(n16314), .C2(n15353), .A(n15518), .B(n15352), .ZN(
        n15355) );
  XNOR2_X1 U18751 ( .A(n15361), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15530) );
  NOR2_X1 U18752 ( .A1(n15530), .A2(n19282), .ZN(n15354) );
  AOI211_X1 U18753 ( .C1(n19278), .C2(n19006), .A(n15355), .B(n15354), .ZN(
        n15356) );
  OAI21_X1 U18754 ( .B1(n15533), .B2(n16292), .A(n15356), .ZN(P2_U2994) );
  INV_X1 U18755 ( .A(n15369), .ZN(n15357) );
  NOR2_X1 U18756 ( .A1(n15370), .A2(n15357), .ZN(n15360) );
  XNOR2_X1 U18757 ( .A(n15360), .B(n10229), .ZN(n15543) );
  AOI21_X1 U18758 ( .B1(n15534), .B2(n15375), .A(n15361), .ZN(n15541) );
  INV_X1 U18759 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n21177) );
  NOR2_X1 U18760 ( .A1(n19131), .A2(n21177), .ZN(n15536) );
  NOR2_X1 U18761 ( .A1(n19013), .A2(n16314), .ZN(n15362) );
  AOI211_X1 U18762 ( .C1(n16299), .C2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15536), .B(n15362), .ZN(n15363) );
  OAI21_X1 U18763 ( .B1(n19021), .B2(n16317), .A(n15363), .ZN(n15364) );
  AOI21_X1 U18764 ( .B1(n15541), .B2(n16287), .A(n15364), .ZN(n15365) );
  OAI21_X1 U18765 ( .B1(n15543), .B2(n16292), .A(n15365), .ZN(P2_U2995) );
  AOI21_X1 U18766 ( .B1(n15369), .B2(n15367), .A(n15366), .ZN(n15368) );
  AOI21_X1 U18767 ( .B1(n15370), .B2(n15369), .A(n15368), .ZN(n15553) );
  INV_X1 U18768 ( .A(n15644), .ZN(n15372) );
  INV_X1 U18769 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15636) );
  INV_X1 U18770 ( .A(n15590), .ZN(n15373) );
  INV_X1 U18771 ( .A(n15525), .ZN(n15374) );
  NAND2_X1 U18772 ( .A1(n15386), .A2(n15374), .ZN(n15387) );
  INV_X1 U18773 ( .A(n15375), .ZN(n15376) );
  AOI21_X1 U18774 ( .B1(n15387), .B2(n15377), .A(n15376), .ZN(n15551) );
  NOR2_X1 U18775 ( .A1(n19131), .A2(n15378), .ZN(n15545) );
  AOI21_X1 U18776 ( .B1(n16299), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15545), .ZN(n15381) );
  NAND2_X1 U18777 ( .A1(n15379), .A2(n19274), .ZN(n15380) );
  OAI211_X1 U18778 ( .C1(n15549), .C2(n16317), .A(n15381), .B(n15380), .ZN(
        n15382) );
  AOI21_X1 U18779 ( .B1(n15551), .B2(n16287), .A(n15382), .ZN(n15383) );
  OAI21_X1 U18780 ( .B1(n15553), .B2(n16292), .A(n15383), .ZN(P2_U2996) );
  XOR2_X1 U18781 ( .A(n15385), .B(n15384), .Z(n15564) );
  INV_X1 U18782 ( .A(n15386), .ZN(n15406) );
  NAND2_X1 U18783 ( .A1(n15556), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15558) );
  INV_X1 U18784 ( .A(n15558), .ZN(n15388) );
  OAI211_X1 U18785 ( .C1(n15388), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16310), .B(n15387), .ZN(n15392) );
  NAND2_X1 U18786 ( .A1(n19088), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15554) );
  NAND2_X1 U18787 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15389) );
  OAI211_X1 U18788 ( .C1(n16314), .C2(n19035), .A(n15554), .B(n15389), .ZN(
        n15390) );
  AOI21_X1 U18789 ( .B1(n19033), .B2(n19278), .A(n15390), .ZN(n15391) );
  OAI211_X1 U18790 ( .C1(n15564), .C2(n16292), .A(n15392), .B(n15391), .ZN(
        P2_U2997) );
  XNOR2_X1 U18791 ( .A(n15394), .B(n15393), .ZN(n15573) );
  OAI211_X1 U18792 ( .C1(n15556), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15558), .B(n16287), .ZN(n15401) );
  INV_X1 U18793 ( .A(n15395), .ZN(n15569) );
  NAND2_X1 U18794 ( .A1(n19274), .A2(n15396), .ZN(n15397) );
  NAND2_X1 U18795 ( .A1(n19088), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15565) );
  OAI211_X1 U18796 ( .C1(n19288), .C2(n15398), .A(n15397), .B(n15565), .ZN(
        n15399) );
  AOI21_X1 U18797 ( .B1(n15569), .B2(n19278), .A(n15399), .ZN(n15400) );
  OAI211_X1 U18798 ( .C1(n15573), .C2(n16292), .A(n15401), .B(n15400), .ZN(
        P2_U2998) );
  NAND2_X1 U18799 ( .A1(n15403), .A2(n15402), .ZN(n15405) );
  XOR2_X1 U18800 ( .A(n15405), .B(n15404), .Z(n15584) );
  AOI21_X1 U18801 ( .B1(n15578), .B2(n15406), .A(n15556), .ZN(n15574) );
  NAND2_X1 U18802 ( .A1(n15574), .A2(n16287), .ZN(n15412) );
  NAND2_X1 U18803 ( .A1(n19274), .A2(n15407), .ZN(n15408) );
  NAND2_X1 U18804 ( .A1(n19088), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15576) );
  OAI211_X1 U18805 ( .C1(n19288), .C2(n15409), .A(n15408), .B(n15576), .ZN(
        n15410) );
  AOI21_X1 U18806 ( .B1(n19045), .B2(n19278), .A(n15410), .ZN(n15411) );
  OAI211_X1 U18807 ( .C1(n15584), .C2(n16292), .A(n15412), .B(n15411), .ZN(
        P2_U2999) );
  NAND2_X1 U18808 ( .A1(n15414), .A2(n15413), .ZN(n15415) );
  XNOR2_X1 U18809 ( .A(n15416), .B(n15415), .ZN(n15596) );
  AOI21_X1 U18810 ( .B1(n15588), .B2(n15417), .A(n15386), .ZN(n15598) );
  NAND2_X1 U18811 ( .A1(n15598), .A2(n16310), .ZN(n15422) );
  AOI22_X1 U18812 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19088), .ZN(n15418) );
  OAI21_X1 U18813 ( .B1(n16314), .B2(n15419), .A(n15418), .ZN(n15420) );
  AOI21_X1 U18814 ( .B1(n19057), .B2(n19278), .A(n15420), .ZN(n15421) );
  OAI211_X1 U18815 ( .C1(n16292), .C2(n15596), .A(n15422), .B(n15421), .ZN(
        P2_U3000) );
  NAND2_X1 U18816 ( .A1(n15425), .A2(n15424), .ZN(n15426) );
  XNOR2_X1 U18817 ( .A(n15423), .B(n15426), .ZN(n15609) );
  NAND2_X1 U18818 ( .A1(n15625), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15428) );
  INV_X1 U18819 ( .A(n15417), .ZN(n15427) );
  AOI21_X1 U18820 ( .B1(n10895), .B2(n15428), .A(n15427), .ZN(n15600) );
  NAND2_X1 U18821 ( .A1(n15600), .A2(n16287), .ZN(n15434) );
  INV_X1 U18822 ( .A(n19069), .ZN(n15432) );
  INV_X1 U18823 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n21209) );
  OAI22_X1 U18824 ( .A1(n19288), .A2(n15429), .B1(n21209), .B2(n19131), .ZN(
        n15431) );
  NOR2_X1 U18825 ( .A1(n16314), .A2(n19068), .ZN(n15430) );
  AOI211_X1 U18826 ( .C1(n15432), .C2(n19278), .A(n15431), .B(n15430), .ZN(
        n15433) );
  OAI211_X1 U18827 ( .C1(n16292), .C2(n15609), .A(n15434), .B(n15433), .ZN(
        P2_U3001) );
  NAND2_X1 U18828 ( .A1(n15435), .A2(n15436), .ZN(n16301) );
  INV_X1 U18829 ( .A(n16300), .ZN(n15438) );
  AND2_X1 U18830 ( .A1(n16300), .A2(n15436), .ZN(n15437) );
  OAI22_X1 U18831 ( .A1(n16301), .A2(n15438), .B1(n15437), .B2(n15435), .ZN(
        n15667) );
  OR2_X1 U18832 ( .A1(n15440), .A2(n15439), .ZN(n15659) );
  NAND3_X1 U18833 ( .A1(n15659), .A2(n15658), .A3(n16310), .ZN(n15445) );
  INV_X1 U18834 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15441) );
  OAI22_X1 U18835 ( .A1(n19288), .A2(n15441), .B1(n16314), .B2(n19127), .ZN(
        n15443) );
  NOR2_X1 U18836 ( .A1(n19135), .A2(n16317), .ZN(n15442) );
  AOI211_X1 U18837 ( .C1(n19088), .C2(P2_REIP_REG_7__SCAN_IN), .A(n15443), .B(
        n15442), .ZN(n15444) );
  OAI211_X1 U18838 ( .C1(n16292), .C2(n15667), .A(n15445), .B(n15444), .ZN(
        P2_U3007) );
  AOI21_X1 U18839 ( .B1(n15447), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15446), .ZN(n15463) );
  NOR2_X1 U18840 ( .A1(n16360), .A2(n16201), .ZN(n15452) );
  NAND2_X1 U18841 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15469), .ZN(
        n15460) );
  OAI21_X1 U18842 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15448), .ZN(n15450) );
  OAI21_X1 U18843 ( .B1(n15460), .B2(n15450), .A(n15449), .ZN(n15451) );
  AOI211_X1 U18844 ( .C1(n15463), .C2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15452), .B(n15451), .ZN(n15453) );
  OAI21_X1 U18845 ( .B1(n16200), .B2(n19296), .A(n15453), .ZN(n15454) );
  AOI21_X1 U18846 ( .B1(n15455), .B2(n16337), .A(n15454), .ZN(n15456) );
  OAI21_X1 U18847 ( .B1(n15457), .B2(n16369), .A(n15456), .ZN(P2_U3020) );
  NAND2_X1 U18848 ( .A1(n19301), .A2(n16213), .ZN(n15459) );
  OAI211_X1 U18849 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15460), .A(
        n15459), .B(n15458), .ZN(n15462) );
  NOR2_X1 U18850 ( .A1(n16212), .A2(n19296), .ZN(n15461) );
  AOI211_X1 U18851 ( .C1(n15463), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15462), .B(n15461), .ZN(n15466) );
  NAND3_X1 U18852 ( .A1(n15464), .A2(n16337), .A3(n15309), .ZN(n15465) );
  OAI211_X1 U18853 ( .C1(n15467), .C2(n16369), .A(n15466), .B(n15465), .ZN(
        P2_U3021) );
  INV_X1 U18854 ( .A(n15468), .ZN(n15478) );
  INV_X1 U18855 ( .A(n15469), .ZN(n15473) );
  AOI21_X1 U18856 ( .B1(n15471), .B2(n15470), .A(n15474), .ZN(n15472) );
  AOI21_X1 U18857 ( .B1(n15474), .B2(n15473), .A(n15472), .ZN(n15477) );
  OAI22_X1 U18858 ( .A1(n16360), .A2(n15475), .B1(n19899), .B2(n19131), .ZN(
        n15476) );
  AOI211_X1 U18859 ( .C1(n15478), .C2(n16339), .A(n15477), .B(n15476), .ZN(
        n15481) );
  NAND2_X1 U18860 ( .A1(n15479), .A2(n16337), .ZN(n15480) );
  OAI211_X1 U18861 ( .C1(n15482), .C2(n16369), .A(n15481), .B(n15480), .ZN(
        P2_U3022) );
  XNOR2_X1 U18862 ( .A(n15483), .B(n15484), .ZN(n16253) );
  NAND2_X1 U18863 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15485), .ZN(
        n15507) );
  AOI211_X1 U18864 ( .C1(n20965), .C2(n10999), .A(n15486), .B(n15507), .ZN(
        n15492) );
  INV_X1 U18865 ( .A(n15510), .ZN(n15490) );
  NOR2_X1 U18866 ( .A1(n19897), .A2(n19131), .ZN(n15487) );
  AOI21_X1 U18867 ( .B1(n19301), .B2(n15488), .A(n15487), .ZN(n15489) );
  OAI21_X1 U18868 ( .B1(n15490), .B2(n20965), .A(n15489), .ZN(n15491) );
  AOI211_X1 U18869 ( .C1(n9875), .C2(n16339), .A(n15492), .B(n15491), .ZN(
        n15496) );
  OR2_X1 U18870 ( .A1(n15511), .A2(n10999), .ZN(n16258) );
  NAND2_X1 U18871 ( .A1(n16258), .A2(n20965), .ZN(n15494) );
  NAND2_X1 U18872 ( .A1(n15494), .A2(n15493), .ZN(n16252) );
  OR2_X1 U18873 ( .A1(n16252), .A2(n19295), .ZN(n15495) );
  OAI211_X1 U18874 ( .C1(n16253), .C2(n16369), .A(n15496), .B(n15495), .ZN(
        P2_U3023) );
  NAND2_X1 U18875 ( .A1(n15499), .A2(n15498), .ZN(n15500) );
  XNOR2_X1 U18876 ( .A(n15497), .B(n15500), .ZN(n16262) );
  INV_X1 U18877 ( .A(n16262), .ZN(n15514) );
  NOR2_X1 U18878 ( .A1(n15502), .A2(n15501), .ZN(n15503) );
  OR2_X1 U18879 ( .A1(n15504), .A2(n15503), .ZN(n15826) );
  INV_X1 U18880 ( .A(n15826), .ZN(n16236) );
  NAND2_X1 U18881 ( .A1(n19301), .A2(n16236), .ZN(n15506) );
  INV_X1 U18882 ( .A(n19131), .ZN(n19275) );
  NAND2_X1 U18883 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19275), .ZN(n15505) );
  OAI211_X1 U18884 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15507), .A(
        n15506), .B(n15505), .ZN(n15509) );
  NOR2_X1 U18885 ( .A1(n16260), .A2(n19296), .ZN(n15508) );
  AOI211_X1 U18886 ( .C1(n15510), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15509), .B(n15508), .ZN(n15513) );
  NAND2_X1 U18887 ( .A1(n15511), .A2(n10999), .ZN(n16257) );
  NAND3_X1 U18888 ( .A1(n16258), .A2(n16257), .A3(n16337), .ZN(n15512) );
  OAI211_X1 U18889 ( .C1(n15514), .C2(n16369), .A(n15513), .B(n15512), .ZN(
        P2_U3024) );
  AND2_X1 U18890 ( .A1(n15516), .A2(n15515), .ZN(n15517) );
  NOR2_X1 U18891 ( .A1(n11609), .A2(n15517), .ZN(n19005) );
  NAND2_X1 U18892 ( .A1(n19301), .A2(n19005), .ZN(n15519) );
  OAI211_X1 U18893 ( .C1(n15520), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15519), .B(n15518), .ZN(n15529) );
  INV_X1 U18894 ( .A(n15523), .ZN(n15521) );
  OAI21_X1 U18895 ( .B1(n15522), .B2(n15562), .A(n15649), .ZN(n15615) );
  AOI21_X1 U18896 ( .B1(n15521), .B2(n16364), .A(n15615), .ZN(n15579) );
  OAI21_X1 U18897 ( .B1(n15562), .B2(n15374), .A(n15579), .ZN(n15546) );
  NAND2_X1 U18898 ( .A1(n15652), .A2(n15522), .ZN(n15591) );
  INV_X1 U18899 ( .A(n15591), .ZN(n15524) );
  NAND2_X1 U18900 ( .A1(n15524), .A2(n15523), .ZN(n15555) );
  NOR3_X1 U18901 ( .A1(n15555), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15525), .ZN(n15544) );
  NOR2_X1 U18902 ( .A1(n15546), .A2(n15544), .ZN(n15535) );
  NAND3_X1 U18903 ( .A1(n15652), .A2(n15526), .A3(n15534), .ZN(n15537) );
  AOI21_X1 U18904 ( .B1(n15535), .B2(n15537), .A(n15527), .ZN(n15528) );
  AOI211_X1 U18905 ( .C1(n19006), .C2(n16339), .A(n15529), .B(n15528), .ZN(
        n15532) );
  OR2_X1 U18906 ( .A1(n15530), .A2(n19295), .ZN(n15531) );
  OAI211_X1 U18907 ( .C1(n15533), .C2(n16369), .A(n15532), .B(n15531), .ZN(
        P2_U3026) );
  NOR2_X1 U18908 ( .A1(n15535), .A2(n15534), .ZN(n15540) );
  AOI21_X1 U18909 ( .B1(n19301), .B2(n19019), .A(n15536), .ZN(n15538) );
  OAI211_X1 U18910 ( .C1(n19021), .C2(n19296), .A(n15538), .B(n15537), .ZN(
        n15539) );
  AOI211_X1 U18911 ( .C1(n15541), .C2(n16337), .A(n15540), .B(n15539), .ZN(
        n15542) );
  OAI21_X1 U18912 ( .B1(n15543), .B2(n16369), .A(n15542), .ZN(P2_U3027) );
  AOI211_X1 U18913 ( .C1(n19301), .C2(n16245), .A(n15545), .B(n15544), .ZN(
        n15548) );
  NAND2_X1 U18914 ( .A1(n15546), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15547) );
  OAI211_X1 U18915 ( .C1(n15549), .C2(n19296), .A(n15548), .B(n15547), .ZN(
        n15550) );
  AOI21_X1 U18916 ( .B1(n15551), .B2(n16337), .A(n15550), .ZN(n15552) );
  OAI21_X1 U18917 ( .B1(n15553), .B2(n16369), .A(n15552), .ZN(P2_U3028) );
  OAI21_X1 U18918 ( .B1(n16360), .B2(n19039), .A(n15554), .ZN(n15557) );
  INV_X1 U18919 ( .A(n15555), .ZN(n15575) );
  INV_X1 U18920 ( .A(n15559), .ZN(n15560) );
  NOR2_X1 U18921 ( .A1(n15562), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15563) );
  OAI21_X1 U18922 ( .B1(n16360), .B2(n19169), .A(n15565), .ZN(n15568) );
  NOR2_X1 U18923 ( .A1(n15566), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15567) );
  AOI211_X1 U18924 ( .C1(n16339), .C2(n15569), .A(n15568), .B(n15567), .ZN(
        n15572) );
  NAND2_X1 U18925 ( .A1(n15570), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15571) );
  OAI211_X1 U18926 ( .C1(n16369), .C2(n15573), .A(n15572), .B(n15571), .ZN(
        P2_U3030) );
  NAND2_X1 U18927 ( .A1(n15574), .A2(n16337), .ZN(n15583) );
  NAND2_X1 U18928 ( .A1(n15575), .A2(n15578), .ZN(n15577) );
  OAI211_X1 U18929 ( .C1(n16360), .C2(n19046), .A(n15577), .B(n15576), .ZN(
        n15581) );
  NOR2_X1 U18930 ( .A1(n15579), .A2(n15578), .ZN(n15580) );
  AOI211_X1 U18931 ( .C1(n19045), .C2(n16339), .A(n15581), .B(n15580), .ZN(
        n15582) );
  OAI211_X1 U18932 ( .C1(n15584), .C2(n16369), .A(n15583), .B(n15582), .ZN(
        P2_U3031) );
  NOR2_X1 U18933 ( .A1(n13418), .A2(n15585), .ZN(n15586) );
  NOR2_X1 U18934 ( .A1(n15587), .A2(n15586), .ZN(n19177) );
  INV_X1 U18935 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19881) );
  NOR2_X1 U18936 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15591), .ZN(
        n15603) );
  NOR2_X1 U18937 ( .A1(n15591), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15619) );
  OR2_X1 U18938 ( .A1(n15615), .A2(n15619), .ZN(n15606) );
  NOR2_X1 U18939 ( .A1(n15603), .A2(n15606), .ZN(n15589) );
  OAI22_X1 U18940 ( .A1(n19131), .A2(n19881), .B1(n15589), .B2(n15588), .ZN(
        n15593) );
  NOR3_X1 U18941 ( .A1(n15591), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15590), .ZN(n15592) );
  AOI211_X1 U18942 ( .C1(n19301), .C2(n19177), .A(n15593), .B(n15592), .ZN(
        n15595) );
  NAND2_X1 U18943 ( .A1(n19057), .A2(n16339), .ZN(n15594) );
  OAI211_X1 U18944 ( .C1(n15596), .C2(n16369), .A(n15595), .B(n15594), .ZN(
        n15597) );
  AOI21_X1 U18945 ( .B1(n15598), .B2(n16337), .A(n15597), .ZN(n15599) );
  INV_X1 U18946 ( .A(n15599), .ZN(P2_U3032) );
  NAND2_X1 U18947 ( .A1(n15600), .A2(n16337), .ZN(n15608) );
  NOR2_X1 U18948 ( .A1(n21209), .A2(n19131), .ZN(n15602) );
  NOR2_X1 U18949 ( .A1(n16360), .A2(n19073), .ZN(n15601) );
  AOI211_X1 U18950 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15603), .A(
        n15602), .B(n15601), .ZN(n15604) );
  OAI21_X1 U18951 ( .B1(n19069), .B2(n19296), .A(n15604), .ZN(n15605) );
  AOI21_X1 U18952 ( .B1(n15606), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15605), .ZN(n15607) );
  OAI211_X1 U18953 ( .C1(n15609), .C2(n16369), .A(n15608), .B(n15607), .ZN(
        P2_U3033) );
  XNOR2_X1 U18954 ( .A(n15625), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16266) );
  INV_X1 U18955 ( .A(n15611), .ZN(n15613) );
  NAND2_X1 U18956 ( .A1(n15613), .A2(n15612), .ZN(n15614) );
  XNOR2_X1 U18957 ( .A(n15610), .B(n15614), .ZN(n16268) );
  INV_X1 U18958 ( .A(n15615), .ZN(n15622) );
  AOI21_X1 U18959 ( .B1(n15617), .B2(n13274), .A(n15616), .ZN(n19080) );
  INV_X1 U18960 ( .A(n19080), .ZN(n19183) );
  NAND2_X1 U18961 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19275), .ZN(n15618) );
  OAI21_X1 U18962 ( .B1(n16360), .B2(n19183), .A(n15618), .ZN(n15620) );
  AOI211_X1 U18963 ( .C1(n19081), .C2(n16339), .A(n15620), .B(n15619), .ZN(
        n15621) );
  OAI21_X1 U18964 ( .B1(n15622), .B2(n10874), .A(n15621), .ZN(n15623) );
  AOI21_X1 U18965 ( .B1(n16268), .B2(n19303), .A(n15623), .ZN(n15624) );
  OAI21_X1 U18966 ( .B1(n16266), .B2(n19295), .A(n15624), .ZN(P2_U3034) );
  INV_X1 U18967 ( .A(n15625), .ZN(n15626) );
  OAI21_X1 U18968 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n9843), .A(
        n15626), .ZN(n16274) );
  AND2_X1 U18969 ( .A1(n16281), .A2(n15645), .ZN(n15628) );
  NAND2_X1 U18970 ( .A1(n15627), .A2(n15628), .ZN(n15633) );
  INV_X1 U18971 ( .A(n15629), .ZN(n15630) );
  NOR2_X1 U18972 ( .A1(n15631), .A2(n15630), .ZN(n15632) );
  XNOR2_X1 U18973 ( .A(n15633), .B(n15632), .ZN(n16273) );
  OAI21_X1 U18974 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15634), .A(
        n15649), .ZN(n16328) );
  INV_X1 U18975 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19876) );
  NOR2_X1 U18976 ( .A1(n19876), .A2(n19131), .ZN(n15638) );
  NAND2_X1 U18977 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15652), .ZN(
        n16325) );
  AOI211_X1 U18978 ( .C1(n16278), .C2(n15636), .A(n15635), .B(n16325), .ZN(
        n15637) );
  AOI211_X1 U18979 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16328), .A(
        n15638), .B(n15637), .ZN(n15641) );
  INV_X1 U18980 ( .A(n15639), .ZN(n19090) );
  AOI22_X1 U18981 ( .A1(n19095), .A2(n16339), .B1(n19301), .B2(n19090), .ZN(
        n15640) );
  OAI211_X1 U18982 ( .C1(n16273), .C2(n16369), .A(n15641), .B(n15640), .ZN(
        n15642) );
  INV_X1 U18983 ( .A(n15642), .ZN(n15643) );
  OAI21_X1 U18984 ( .B1(n16274), .B2(n19295), .A(n15643), .ZN(P2_U3035) );
  OAI21_X1 U18985 ( .B1(n15371), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15644), .ZN(n16293) );
  INV_X1 U18986 ( .A(n15645), .ZN(n16279) );
  OR2_X1 U18987 ( .A1(n16279), .A2(n15646), .ZN(n15647) );
  XNOR2_X1 U18988 ( .A(n15648), .B(n15647), .ZN(n16291) );
  INV_X1 U18989 ( .A(n15649), .ZN(n15651) );
  INV_X1 U18990 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19873) );
  NOR2_X1 U18991 ( .A1(n19873), .A2(n19131), .ZN(n15650) );
  AOI221_X1 U18992 ( .B1(n15652), .B2(n21028), .C1(n15651), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15650), .ZN(n15655) );
  OAI22_X1 U18993 ( .A1(n19120), .A2(n16360), .B1(n19296), .B2(n19119), .ZN(
        n15653) );
  INV_X1 U18994 ( .A(n15653), .ZN(n15654) );
  OAI211_X1 U18995 ( .C1(n16291), .C2(n16369), .A(n15655), .B(n15654), .ZN(
        n15656) );
  INV_X1 U18996 ( .A(n15656), .ZN(n15657) );
  OAI21_X1 U18997 ( .B1(n16293), .B2(n19295), .A(n15657), .ZN(P2_U3037) );
  NAND3_X1 U18998 ( .A1(n15659), .A2(n15658), .A3(n16337), .ZN(n15666) );
  INV_X1 U18999 ( .A(n19134), .ZN(n15660) );
  AOI22_X1 U19000 ( .A1(n19301), .A2(n15660), .B1(n19088), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n15661) );
  OAI21_X1 U19001 ( .B1(n19135), .B2(n19296), .A(n15661), .ZN(n15663) );
  NOR2_X1 U19002 ( .A1(n16334), .A2(n15664), .ZN(n15662) );
  AOI211_X1 U19003 ( .C1(n16342), .C2(n15664), .A(n15663), .B(n15662), .ZN(
        n15665) );
  OAI211_X1 U19004 ( .C1(n15667), .C2(n16369), .A(n15666), .B(n15665), .ZN(
        P2_U3039) );
  XOR2_X1 U19005 ( .A(n15668), .B(n15670), .Z(n16320) );
  INV_X1 U19006 ( .A(n16320), .ZN(n15682) );
  OAI21_X1 U19007 ( .B1(n15672), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15671), .ZN(n16318) );
  INV_X1 U19008 ( .A(n16318), .ZN(n15680) );
  NAND2_X1 U19009 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19275), .ZN(n15673) );
  OAI221_X1 U19010 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15676), .C1(
        n15675), .C2(n15674), .A(n15673), .ZN(n15679) );
  OAI22_X1 U19011 ( .A1(n16316), .A2(n19296), .B1(n16360), .B2(n15677), .ZN(
        n15678) );
  AOI211_X1 U19012 ( .C1(n15680), .C2(n16337), .A(n15679), .B(n15678), .ZN(
        n15681) );
  OAI21_X1 U19013 ( .B1(n16369), .B2(n15682), .A(n15681), .ZN(P2_U3040) );
  INV_X1 U19014 ( .A(n16358), .ZN(n15686) );
  OAI22_X1 U19015 ( .A1(n19295), .A2(n15683), .B1(n10619), .B2(n19296), .ZN(
        n15684) );
  AOI211_X1 U19016 ( .C1(n15686), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15685), .B(n15684), .ZN(n15690) );
  AOI22_X1 U19017 ( .A1(n19303), .A2(n15687), .B1(n19301), .B2(n19948), .ZN(
        n15689) );
  OAI211_X1 U19018 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16364), .B(n19306), .ZN(n15688) );
  NAND3_X1 U19019 ( .A1(n15690), .A2(n15689), .A3(n15688), .ZN(P2_U3045) );
  INV_X1 U19020 ( .A(n16413), .ZN(n15756) );
  INV_X1 U19021 ( .A(n15719), .ZN(n19926) );
  INV_X1 U19022 ( .A(n15715), .ZN(n15754) );
  INV_X1 U19023 ( .A(n11361), .ZN(n15692) );
  NAND2_X1 U19024 ( .A1(n15692), .A2(n15691), .ZN(n15712) );
  MUX2_X1 U19025 ( .A(n15748), .B(n15712), .S(n15693), .Z(n15694) );
  AOI21_X1 U19026 ( .B1(n15695), .B2(n15754), .A(n15694), .ZN(n16373) );
  AOI21_X1 U19027 ( .B1(n19147), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n15696), .ZN(n15717) );
  INV_X1 U19028 ( .A(n15717), .ZN(n15697) );
  OAI222_X1 U19029 ( .A1(n15756), .A2(n15698), .B1(n19926), .B2(n16373), .C1(
        n16419), .C2(n15697), .ZN(n15708) );
  NOR2_X1 U19030 ( .A1(n20977), .A2(n19206), .ZN(n15883) );
  INV_X1 U19031 ( .A(n15699), .ZN(n15706) );
  AND2_X1 U19032 ( .A1(n15701), .A2(n15700), .ZN(n15705) );
  NAND2_X1 U19033 ( .A1(n15702), .A2(n16388), .ZN(n15703) );
  OR2_X1 U19034 ( .A1(n19203), .A2(n15703), .ZN(n15704) );
  OAI22_X1 U19035 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19951), .B1(n16404), 
        .B2(n18965), .ZN(n15707) );
  MUX2_X1 U19036 ( .A(n15708), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15795), .Z(P2_U3601) );
  NOR2_X1 U19037 ( .A1(n15709), .A2(n15724), .ZN(n15713) );
  AOI22_X1 U19038 ( .A1(n15713), .A2(n15712), .B1(n15748), .B2(n15711), .ZN(
        n15714) );
  OAI21_X1 U19039 ( .B1(n10619), .B2(n15715), .A(n15714), .ZN(n16372) );
  OAI21_X1 U19040 ( .B1(n19075), .B2(n10357), .A(n15716), .ZN(n15737) );
  INV_X1 U19041 ( .A(n15737), .ZN(n15718) );
  NOR2_X1 U19042 ( .A1(n15717), .A2(n16419), .ZN(n15736) );
  AOI222_X1 U19043 ( .A1(n16372), .A2(n15719), .B1(n16413), .B2(n19944), .C1(
        n15718), .C2(n15736), .ZN(n15721) );
  NAND2_X1 U19044 ( .A1(n15795), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15720) );
  OAI21_X1 U19045 ( .B1(n15721), .B2(n15795), .A(n15720), .ZN(P2_U3600) );
  INV_X1 U19046 ( .A(n15722), .ZN(n15723) );
  NAND2_X1 U19047 ( .A1(n15748), .A2(n15723), .ZN(n15742) );
  INV_X1 U19048 ( .A(n15744), .ZN(n16399) );
  INV_X1 U19049 ( .A(n15724), .ZN(n15726) );
  NAND2_X1 U19050 ( .A1(n15726), .A2(n15725), .ZN(n15746) );
  NAND2_X1 U19051 ( .A1(n15745), .A2(n15746), .ZN(n15729) );
  OAI21_X1 U19052 ( .B1(n16399), .B2(n15743), .A(n15729), .ZN(n15732) );
  NAND2_X1 U19053 ( .A1(n15728), .A2(n15727), .ZN(n15740) );
  INV_X1 U19054 ( .A(n15729), .ZN(n15730) );
  NAND2_X1 U19055 ( .A1(n15740), .A2(n15730), .ZN(n15731) );
  OAI211_X1 U19056 ( .C1(n15742), .C2(n15733), .A(n15732), .B(n15731), .ZN(
        n15734) );
  AOI21_X1 U19057 ( .B1(n10645), .B2(n15754), .A(n15734), .ZN(n16371) );
  OAI22_X1 U19058 ( .A1(n19938), .A2(n15756), .B1(n16371), .B2(n19926), .ZN(
        n15735) );
  AOI21_X1 U19059 ( .B1(n15737), .B2(n15736), .A(n15735), .ZN(n15738) );
  MUX2_X1 U19060 ( .A(n15738), .B(n16370), .S(n15795), .Z(n15739) );
  INV_X1 U19061 ( .A(n15739), .ZN(P2_U3599) );
  NAND2_X1 U19062 ( .A1(n15740), .A2(n15745), .ZN(n15741) );
  NAND3_X1 U19063 ( .A1(n15742), .A2(n15741), .A3(n15746), .ZN(n15752) );
  INV_X1 U19064 ( .A(n15743), .ZN(n16401) );
  NAND3_X1 U19065 ( .A1(n16401), .A2(n15745), .A3(n15744), .ZN(n15747) );
  NAND2_X1 U19066 ( .A1(n15747), .A2(n15746), .ZN(n15750) );
  NAND2_X1 U19067 ( .A1(n15748), .A2(n15722), .ZN(n15749) );
  NAND2_X1 U19068 ( .A1(n15750), .A2(n15749), .ZN(n15751) );
  MUX2_X1 U19069 ( .A(n15752), .B(n15751), .S(n16379), .Z(n15753) );
  AOI21_X1 U19070 ( .B1(n15755), .B2(n15754), .A(n15753), .ZN(n16382) );
  OAI22_X1 U19071 ( .A1(n19354), .A2(n15756), .B1(n16382), .B2(n19926), .ZN(
        n15757) );
  MUX2_X1 U19072 ( .A(n15757), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15795), .Z(P2_U3596) );
  INV_X1 U19073 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18503) );
  AOI22_X1 U19074 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15758) );
  OAI21_X1 U19075 ( .B1(n17186), .B2(n18503), .A(n15758), .ZN(n15769) );
  INV_X1 U19076 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15767) );
  AOI22_X1 U19077 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15766) );
  AOI22_X1 U19078 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15759) );
  OAI21_X1 U19079 ( .B1(n11076), .B2(n15760), .A(n15759), .ZN(n15764) );
  INV_X1 U19080 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17261) );
  AOI22_X1 U19081 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U19082 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15761) );
  OAI211_X1 U19083 ( .C1(n11056), .C2(n17261), .A(n15762), .B(n15761), .ZN(
        n15763) );
  AOI211_X1 U19084 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n15764), .B(n15763), .ZN(n15765) );
  OAI211_X1 U19085 ( .C1(n17177), .C2(n15767), .A(n15766), .B(n15765), .ZN(
        n15768) );
  AOI211_X1 U19086 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n15769), .B(n15768), .ZN(n17380) );
  NAND2_X1 U19087 ( .A1(n17275), .A2(n15770), .ZN(n17173) );
  INV_X1 U19088 ( .A(n17173), .ZN(n17155) );
  NAND2_X1 U19089 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17155), .ZN(n15776) );
  NOR2_X1 U19090 ( .A1(n16823), .A2(n17208), .ZN(n15774) );
  NOR2_X1 U19091 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17278), .ZN(n17154) );
  NOR4_X1 U19092 ( .A1(n16846), .A2(n17249), .A3(n15772), .A4(n15771), .ZN(
        n15773) );
  NAND4_X1 U19093 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n15774), .A3(n17154), 
        .A4(n15773), .ZN(n15775) );
  OAI211_X1 U19094 ( .C1(n17380), .C2(n17275), .A(n15776), .B(n15775), .ZN(
        P3_U2690) );
  NOR2_X1 U19095 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18626), .ZN(
        n18301) );
  NOR3_X1 U19096 ( .A1(n21022), .A2(n18936), .A3(n18948), .ZN(n15778) );
  INV_X1 U19097 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16897) );
  NAND2_X1 U19098 ( .A1(n15793), .A2(n16897), .ZN(n15777) );
  OR2_X1 U19099 ( .A1(n17237), .A2(n15777), .ZN(n18249) );
  INV_X1 U19100 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18250) );
  INV_X1 U19101 ( .A(n15778), .ZN(n18890) );
  NOR2_X1 U19102 ( .A1(n18250), .A2(n18890), .ZN(n15792) );
  AOI211_X1 U19103 ( .C1(n15778), .C2(n18249), .A(n18625), .B(n15792), .ZN(
        n15779) );
  NOR2_X1 U19104 ( .A1(n18301), .A2(n15779), .ZN(n18255) );
  INV_X1 U19105 ( .A(n18564), .ZN(n18622) );
  INV_X1 U19106 ( .A(n15779), .ZN(n18260) );
  INV_X1 U19107 ( .A(n17816), .ZN(n18252) );
  OAI22_X1 U19108 ( .A1(n18938), .A2(n18252), .B1(n18765), .B2(n18626), .ZN(
        n18256) );
  NAND3_X1 U19109 ( .A1(n18767), .A2(n18260), .A3(n18256), .ZN(n15780) );
  OAI221_X1 U19110 ( .B1(n18767), .B2(n18255), .C1(n18767), .C2(n18622), .A(
        n15780), .ZN(P3_U2864) );
  INV_X1 U19111 ( .A(n17481), .ZN(n15782) );
  NAND2_X1 U19112 ( .A1(n15810), .A2(n18809), .ZN(n15784) );
  NOR2_X1 U19113 ( .A1(n15784), .A2(n17442), .ZN(n15790) );
  INV_X1 U19114 ( .A(n15785), .ZN(n15786) );
  OAI211_X1 U19115 ( .C1(n15789), .C2(n15788), .A(n15787), .B(n15786), .ZN(
        n15803) );
  NOR4_X2 U19116 ( .A1(n15888), .A2(n15791), .A3(n15790), .A4(n15803), .ZN(
        n18770) );
  INV_X1 U19117 ( .A(n18770), .ZN(n18758) );
  NOR2_X1 U19118 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18626), .ZN(n18267) );
  INV_X1 U19119 ( .A(n18917), .ZN(n18914) );
  AOI21_X1 U19120 ( .B1(n15793), .B2(n16897), .A(n18747), .ZN(n18732) );
  NAND3_X1 U19121 ( .A1(n18914), .A2(n18949), .A3(n18732), .ZN(n15794) );
  OAI21_X1 U19122 ( .B1(n18914), .B2(n16897), .A(n15794), .ZN(P3_U3284) );
  INV_X1 U19123 ( .A(n15795), .ZN(n15799) );
  NOR4_X1 U19124 ( .A1(n15796), .A2(n11312), .A3(n16391), .A4(n19926), .ZN(
        n15797) );
  NAND2_X1 U19125 ( .A1(n15799), .A2(n15797), .ZN(n15798) );
  OAI21_X1 U19126 ( .B1(n15799), .B2(n11329), .A(n15798), .ZN(P2_U3595) );
  INV_X1 U19127 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16443) );
  NOR2_X1 U19128 ( .A1(n11132), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16484) );
  AOI21_X1 U19129 ( .B1(n15800), .B2(n16470), .A(n16484), .ZN(n15801) );
  XOR2_X1 U19130 ( .A(n16443), .B(n15801), .Z(n16457) );
  INV_X1 U19131 ( .A(n18728), .ZN(n15805) );
  AOI211_X1 U19132 ( .C1(n18282), .C2(n15802), .A(n9796), .B(n18730), .ZN(
        n15804) );
  AOI21_X1 U19133 ( .B1(n18272), .B2(n9796), .A(n18932), .ZN(n15808) );
  AOI21_X1 U19134 ( .B1(n15808), .B2(n15807), .A(n18941), .ZN(n16581) );
  NAND3_X1 U19135 ( .A1(n15810), .A2(n16581), .A3(n15809), .ZN(n15811) );
  INV_X1 U19136 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17928) );
  NOR2_X1 U19137 ( .A1(n18739), .A2(n18220), .ZN(n18127) );
  INV_X1 U19138 ( .A(n18127), .ZN(n17982) );
  NAND2_X1 U19139 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18151) );
  NOR2_X1 U19140 ( .A1(n21098), .A2(n18151), .ZN(n18029) );
  NAND3_X1 U19141 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18173) );
  NOR2_X1 U19142 ( .A1(n18216), .A2(n20976), .ZN(n18191) );
  INV_X1 U19143 ( .A(n18191), .ZN(n18212) );
  NOR2_X1 U19144 ( .A1(n18173), .A2(n18212), .ZN(n18044) );
  NAND2_X1 U19145 ( .A1(n18029), .A2(n18044), .ZN(n18072) );
  NOR2_X1 U19146 ( .A1(n18913), .A2(n18072), .ZN(n18135) );
  NAND2_X1 U19147 ( .A1(n16426), .A2(n18135), .ZN(n18047) );
  NOR2_X1 U19148 ( .A1(n17632), .A2(n18047), .ZN(n17998) );
  NAND2_X1 U19149 ( .A1(n16482), .A2(n17998), .ZN(n17979) );
  OR2_X1 U19150 ( .A1(n16428), .A2(n17928), .ZN(n16483) );
  OAI21_X1 U19151 ( .B1(n17979), .B2(n16483), .A(n18759), .ZN(n15814) );
  INV_X1 U19152 ( .A(n16427), .ZN(n17946) );
  AOI21_X1 U19153 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18193) );
  NOR2_X1 U19154 ( .A1(n18193), .A2(n18173), .ZN(n18148) );
  NAND2_X1 U19155 ( .A1(n18148), .A2(n18029), .ZN(n18070) );
  NOR2_X1 U19156 ( .A1(n18031), .A2(n18070), .ZN(n18021) );
  NAND2_X1 U19157 ( .A1(n17946), .A2(n18021), .ZN(n17967) );
  OAI21_X1 U19158 ( .B1(n16428), .B2(n17967), .A(n18220), .ZN(n17925) );
  INV_X1 U19159 ( .A(n16464), .ZN(n15820) );
  NOR2_X1 U19160 ( .A1(n18031), .A2(n18072), .ZN(n18020) );
  INV_X1 U19161 ( .A(n18020), .ZN(n17984) );
  OAI21_X1 U19162 ( .B1(n15820), .B2(n17984), .A(n18739), .ZN(n15813) );
  NAND4_X1 U19163 ( .A1(n18224), .A2(n15814), .A3(n17925), .A4(n15813), .ZN(
        n15874) );
  AOI21_X1 U19164 ( .B1(n17928), .B2(n17982), .A(n15874), .ZN(n16473) );
  NAND2_X1 U19165 ( .A1(n18149), .A2(n17551), .ZN(n15816) );
  NAND2_X1 U19166 ( .A1(n18113), .A2(n18224), .ZN(n18175) );
  NAND2_X1 U19167 ( .A1(n17410), .A2(n18242), .ZN(n18088) );
  OAI22_X1 U19168 ( .A1(n18175), .A2(n16436), .B1(n18088), .B2(n16437), .ZN(
        n15815) );
  INV_X1 U19169 ( .A(n15815), .ZN(n15876) );
  OAI221_X1 U19170 ( .B1(n18140), .B2(n16473), .C1(n18235), .C2(n15816), .A(
        n15876), .ZN(n15817) );
  AOI22_X1 U19171 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15817), .B1(
        n18140), .B2(P3_REIP_REG_29__SCAN_IN), .ZN(n15823) );
  INV_X1 U19172 ( .A(n15818), .ZN(n18727) );
  NAND2_X1 U19173 ( .A1(n17410), .A2(n18727), .ZN(n18092) );
  AOI22_X1 U19174 ( .A1(n18113), .A2(n16425), .B1(n15819), .B2(n18111), .ZN(
        n18030) );
  INV_X1 U19175 ( .A(n18759), .ZN(n18749) );
  OAI21_X1 U19176 ( .B1(n18749), .B2(n18913), .A(n18761), .ZN(n18215) );
  AOI22_X1 U19177 ( .A1(n18220), .A2(n18021), .B1(n18020), .B2(n18215), .ZN(
        n17948) );
  OAI21_X1 U19178 ( .B1(n18030), .B2(n18031), .A(n17948), .ZN(n17987) );
  NAND2_X1 U19179 ( .A1(n18224), .A2(n17987), .ZN(n16481) );
  NOR2_X1 U19180 ( .A1(n15820), .A2(n16481), .ZN(n17921) );
  NAND3_X1 U19181 ( .A1(n15821), .A2(n17921), .A3(n16443), .ZN(n15822) );
  OAI211_X1 U19182 ( .C1(n16457), .C2(n18161), .A(n15823), .B(n15822), .ZN(
        P3_U2833) );
  AOI22_X1 U19183 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19145), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19128), .ZN(n15833) );
  INV_X1 U19184 ( .A(n15824), .ZN(n15825) );
  AOI22_X1 U19185 ( .A1(n15825), .A2(n19129), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19138), .ZN(n15832) );
  OAI22_X1 U19186 ( .A1(n16260), .A2(n19151), .B1(n15826), .B2(n19150), .ZN(
        n15827) );
  INV_X1 U19187 ( .A(n15827), .ZN(n15831) );
  OAI211_X1 U19188 ( .C1(n16265), .C2(n15829), .A(n19154), .B(n15828), .ZN(
        n15830) );
  NAND4_X1 U19189 ( .A1(n15833), .A2(n15832), .A3(n15831), .A4(n15830), .ZN(
        P2_U2833) );
  NOR3_X1 U19190 ( .A1(n15835), .A2(n15834), .A3(n20863), .ZN(n15836) );
  NAND2_X1 U19191 ( .A1(n15836), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15840) );
  OAI22_X1 U19192 ( .A1(n15838), .A2(n15837), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15836), .ZN(n15839) );
  NAND2_X1 U19193 ( .A1(n15840), .A2(n15839), .ZN(n15843) );
  INV_X1 U19194 ( .A(n15841), .ZN(n15842) );
  AOI222_X1 U19195 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15843), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15842), .C1(n15843), 
        .C2(n15842), .ZN(n15845) );
  AOI222_X1 U19196 ( .A1(n15845), .A2(n20574), .B1(n15845), .B2(n15844), .C1(
        n20574), .C2(n15844), .ZN(n15846) );
  NOR2_X1 U19197 ( .A1(n15846), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n15854) );
  NOR2_X1 U19198 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15850) );
  INV_X1 U19199 ( .A(n15847), .ZN(n15848) );
  OAI211_X1 U19200 ( .C1(n15851), .C2(n15850), .A(n15849), .B(n15848), .ZN(
        n15852) );
  NOR3_X1 U19201 ( .A1(n15854), .A2(n15853), .A3(n15852), .ZN(n15870) );
  NAND4_X1 U19202 ( .A1(n15858), .A2(n15857), .A3(n15856), .A4(n15855), .ZN(
        n15860) );
  OAI21_X1 U19203 ( .B1(n20777), .B2(n20880), .A(n20778), .ZN(n15859) );
  AND2_X1 U19204 ( .A1(n15860), .A2(n15859), .ZN(n16158) );
  OAI221_X1 U19205 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15870), 
        .A(n16158), .ZN(n16164) );
  NOR2_X1 U19206 ( .A1(n15862), .A2(n15861), .ZN(n15863) );
  NOR2_X1 U19207 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15863), .ZN(n15868) );
  AOI21_X1 U19208 ( .B1(n20615), .B2(n20880), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n16152) );
  NAND2_X1 U19209 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20880), .ZN(n16154) );
  AND2_X1 U19210 ( .A1(n15865), .A2(n15864), .ZN(n20861) );
  AOI21_X1 U19211 ( .B1(n16152), .B2(n16154), .A(n20861), .ZN(n15866) );
  NAND2_X1 U19212 ( .A1(n16164), .A2(n15866), .ZN(n15867) );
  AOI22_X1 U19213 ( .A1(n16164), .A2(n15868), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15867), .ZN(n15869) );
  OAI21_X1 U19214 ( .B1(n15870), .B2(n19992), .A(n15869), .ZN(P1_U3161) );
  AOI21_X1 U19215 ( .B1(n15872), .B2(n11132), .A(n15871), .ZN(n15873) );
  XOR2_X1 U19216 ( .A(n15873), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16440) );
  NOR2_X1 U19217 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16458), .ZN(
        n16435) );
  OAI221_X1 U19218 ( .B1(n15874), .B2(n18149), .C1(n15874), .C2(n16458), .A(
        n16718), .ZN(n16460) );
  INV_X1 U19219 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15875) );
  AOI21_X1 U19220 ( .B1(n15876), .B2(n16460), .A(n15875), .ZN(n15877) );
  AOI21_X1 U19221 ( .B1(n17921), .B2(n16435), .A(n15877), .ZN(n15878) );
  NAND2_X1 U19222 ( .A1(n18140), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16432) );
  OAI211_X1 U19223 ( .C1(n16440), .C2(n18161), .A(n15878), .B(n16432), .ZN(
        P3_U2832) );
  INV_X1 U19224 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21079) );
  NOR2_X1 U19225 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21079), .ZN(n20788) );
  INV_X1 U19226 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20790) );
  NOR2_X1 U19227 ( .A1(n21063), .A2(n20790), .ZN(n20787) );
  NAND2_X1 U19228 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n15879) );
  AOI22_X1 U19229 ( .A1(HOLD), .A2(n20788), .B1(n20787), .B2(n15879), .ZN(
        n15881) );
  OAI211_X1 U19230 ( .C1(n20880), .C2(n21079), .A(n15881), .B(n15880), .ZN(
        P1_U3195) );
  AND2_X1 U19231 ( .A1(n20112), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19232 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15882) );
  NOR3_X1 U19233 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20977), .A3(n19983), 
        .ZN(n16415) );
  NOR4_X1 U19234 ( .A1(n19977), .A2(n15882), .A3(n16415), .A4(n15883), .ZN(
        P2_U3178) );
  INV_X1 U19235 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18968) );
  INV_X1 U19236 ( .A(n15883), .ZN(n16423) );
  INV_X1 U19237 ( .A(n19964), .ZN(n15884) );
  OAI221_X1 U19238 ( .B1(n18968), .B2(n16423), .C1(n15884), .C2(n16423), .A(
        n9793), .ZN(n19956) );
  NOR2_X1 U19239 ( .A1(n15885), .A2(n19956), .ZN(P2_U3047) );
  NAND2_X1 U19240 ( .A1(n18297), .A2(n17429), .ZN(n17372) );
  INV_X1 U19241 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17511) );
  AOI22_X1 U19242 ( .A1(n17435), .A2(BUF2_REG_0__SCAN_IN), .B1(n17434), .B2(
        n15890), .ZN(n15891) );
  OAI221_X1 U19243 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17372), .C1(n17511), 
        .C2(n17429), .A(n15891), .ZN(P3_U2735) );
  AOI22_X1 U19244 ( .A1(n20081), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20087), .ZN(n15901) );
  OAI22_X1 U19245 ( .A1(n15893), .A2(n15945), .B1(n15892), .B2(n20098), .ZN(
        n15894) );
  AOI21_X1 U19246 ( .B1(n15895), .B2(n20086), .A(n15894), .ZN(n15900) );
  NOR2_X1 U19247 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20080), .ZN(n15902) );
  INV_X1 U19248 ( .A(n15896), .ZN(n15904) );
  OAI21_X1 U19249 ( .B1(n15902), .B2(n15904), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15899) );
  INV_X1 U19250 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20825) );
  NAND3_X1 U19251 ( .A1(n20084), .A2(n15897), .A3(n20825), .ZN(n15898) );
  NAND4_X1 U19252 ( .A1(n15901), .A2(n15900), .A3(n15899), .A4(n15898), .ZN(
        P1_U2815) );
  AOI22_X1 U19253 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15904), .B1(n15903), 
        .B2(n15902), .ZN(n15906) );
  AOI22_X1 U19254 ( .A1(n20081), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20087), .ZN(n15905) );
  OAI211_X1 U19255 ( .C1(n15907), .C2(n20098), .A(n15906), .B(n15905), .ZN(
        n15908) );
  AOI21_X1 U19256 ( .B1(n15909), .B2(n20050), .A(n15908), .ZN(n15910) );
  OAI21_X1 U19257 ( .B1(n15911), .B2(n20078), .A(n15910), .ZN(P1_U2816) );
  NAND2_X1 U19258 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n15912), .ZN(n15950) );
  NOR3_X1 U19259 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15913), .A3(n15950), 
        .ZN(n15921) );
  OAI21_X1 U19260 ( .B1(n15928), .B2(n15914), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15915) );
  OAI21_X1 U19261 ( .B1(n20025), .B2(n15916), .A(n15915), .ZN(n15917) );
  AOI21_X1 U19262 ( .B1(n15918), .B2(n20086), .A(n15917), .ZN(n15919) );
  OAI21_X1 U19263 ( .B1(n20043), .B2(n14573), .A(n15919), .ZN(n15920) );
  AOI211_X1 U19264 ( .C1(n15922), .C2(n20050), .A(n15921), .B(n15920), .ZN(
        n15923) );
  OAI21_X1 U19265 ( .B1(n20098), .B2(n15924), .A(n15923), .ZN(P1_U2818) );
  OAI22_X1 U19266 ( .A1(n15925), .A2(n20043), .B1(n20078), .B2(n15997), .ZN(
        n15926) );
  AOI21_X1 U19267 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20087), .A(
        n15926), .ZN(n15930) );
  NAND2_X1 U19268 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15932) );
  OAI21_X1 U19269 ( .B1(n15932), .B2(n15950), .A(n14979), .ZN(n15927) );
  AOI22_X1 U19270 ( .A1(n15994), .A2(n20050), .B1(n15928), .B2(n15927), .ZN(
        n15929) );
  OAI211_X1 U19271 ( .C1(n20098), .C2(n15931), .A(n15930), .B(n15929), .ZN(
        P1_U2820) );
  OAI21_X1 U19272 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15932), .ZN(n15940) );
  AOI22_X1 U19273 ( .A1(n15941), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n20081), 
        .B2(P1_EBX_REG_19__SCAN_IN), .ZN(n15933) );
  OAI211_X1 U19274 ( .C1(n20025), .C2(n15934), .A(n15933), .B(n20022), .ZN(
        n15937) );
  OAI22_X1 U19275 ( .A1(n15935), .A2(n15945), .B1(n20098), .B2(n16040), .ZN(
        n15936) );
  AOI211_X1 U19276 ( .C1(n15938), .C2(n20086), .A(n15937), .B(n15936), .ZN(
        n15939) );
  OAI21_X1 U19277 ( .B1(n15950), .B2(n15940), .A(n15939), .ZN(P1_U2821) );
  AOI22_X1 U19278 ( .A1(n15941), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n20081), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n15942) );
  OAI21_X1 U19279 ( .B1(n15943), .B2(n20078), .A(n15942), .ZN(n15944) );
  AOI211_X1 U19280 ( .C1(n20087), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20069), .B(n15944), .ZN(n15949) );
  OAI22_X1 U19281 ( .A1(n15946), .A2(n15945), .B1(n20098), .B2(n16048), .ZN(
        n15947) );
  INV_X1 U19282 ( .A(n15947), .ZN(n15948) );
  OAI211_X1 U19283 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15950), .A(n15949), 
        .B(n15948), .ZN(P1_U2822) );
  OAI22_X1 U19284 ( .A1(n20098), .A2(n15951), .B1(n20043), .B2(n21014), .ZN(
        n15952) );
  AOI211_X1 U19285 ( .C1(n20087), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20069), .B(n15952), .ZN(n15957) );
  XNOR2_X1 U19286 ( .A(P1_REIP_REG_16__SCAN_IN), .B(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15953) );
  OAI22_X1 U19287 ( .A1(n15954), .A2(n15953), .B1(n15965), .B2(n14993), .ZN(
        n15955) );
  AOI21_X1 U19288 ( .B1(n15998), .B2(n20050), .A(n15955), .ZN(n15956) );
  OAI211_X1 U19289 ( .C1(n16002), .C2(n20078), .A(n15957), .B(n15956), .ZN(
        P1_U2824) );
  INV_X1 U19290 ( .A(n15958), .ZN(n15959) );
  AOI21_X1 U19291 ( .B1(n15959), .B2(n15980), .A(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n15966) );
  OAI22_X1 U19292 ( .A1(n15961), .A2(n20098), .B1(n20043), .B2(n15960), .ZN(
        n15962) );
  AOI211_X1 U19293 ( .C1(n20087), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20069), .B(n15962), .ZN(n15964) );
  AOI22_X1 U19294 ( .A1(n16004), .A2(n20050), .B1(n20086), .B2(n16003), .ZN(
        n15963) );
  OAI211_X1 U19295 ( .C1(n15966), .C2(n15965), .A(n15964), .B(n15963), .ZN(
        P1_U2826) );
  NAND2_X1 U19296 ( .A1(n20087), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15967) );
  OAI211_X1 U19297 ( .C1(n20043), .C2(n15968), .A(n15967), .B(n20022), .ZN(
        n15971) );
  NOR2_X1 U19298 ( .A1(n20098), .A2(n15969), .ZN(n15970) );
  NOR2_X1 U19299 ( .A1(n15971), .A2(n15970), .ZN(n15975) );
  AOI22_X1 U19300 ( .A1(n16009), .A2(n20086), .B1(n20050), .B2(n16008), .ZN(
        n15974) );
  OAI221_X1 U19301 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(P1_REIP_REG_11__SCAN_IN), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n15980), .A(n15972), .ZN(n15973) );
  NAND3_X1 U19302 ( .A1(n15975), .A2(n15974), .A3(n15973), .ZN(P1_U2828) );
  INV_X1 U19303 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15979) );
  INV_X1 U19304 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15977) );
  AOI22_X1 U19305 ( .A1(n20056), .A2(n16083), .B1(n20081), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15976) );
  OAI211_X1 U19306 ( .C1(n20025), .C2(n15977), .A(n15976), .B(n20022), .ZN(
        n15978) );
  AOI221_X1 U19307 ( .B1(n15981), .B2(P1_REIP_REG_11__SCAN_IN), .C1(n15980), 
        .C2(n15979), .A(n15978), .ZN(n15983) );
  NAND2_X1 U19308 ( .A1(n20050), .A2(n16018), .ZN(n15982) );
  OAI211_X1 U19309 ( .C1(n20078), .C2(n16021), .A(n15983), .B(n15982), .ZN(
        P1_U2829) );
  INV_X1 U19310 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n19315) );
  INV_X1 U19311 ( .A(n15984), .ZN(n15986) );
  AOI22_X1 U19312 ( .A1(n15986), .A2(n20242), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n15985), .ZN(n15991) );
  AOI22_X1 U19313 ( .A1(n15989), .A2(n15988), .B1(n15987), .B2(DATAI_18_), 
        .ZN(n15990) );
  OAI211_X1 U19314 ( .C1(n15992), .C2(n19315), .A(n15991), .B(n15990), .ZN(
        P1_U2886) );
  AOI22_X1 U19315 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15996) );
  AOI22_X1 U19316 ( .A1(n15994), .A2(n20159), .B1(n20169), .B2(n15993), .ZN(
        n15995) );
  OAI211_X1 U19317 ( .C1(n20163), .C2(n15997), .A(n15996), .B(n15995), .ZN(
        P1_U2979) );
  AOI22_X1 U19318 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16001) );
  AOI22_X1 U19319 ( .A1(n15999), .A2(n20169), .B1(n20159), .B2(n15998), .ZN(
        n16000) );
  OAI211_X1 U19320 ( .C1(n20163), .C2(n16002), .A(n16001), .B(n16000), .ZN(
        P1_U2983) );
  AOI22_X1 U19321 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16006) );
  AOI22_X1 U19322 ( .A1(n16004), .A2(n20159), .B1(n20171), .B2(n16003), .ZN(
        n16005) );
  OAI211_X1 U19323 ( .C1(n16007), .C2(n19999), .A(n16006), .B(n16005), .ZN(
        P1_U2985) );
  AOI22_X1 U19324 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16011) );
  AOI22_X1 U19325 ( .A1(n20171), .A2(n16009), .B1(n20159), .B2(n16008), .ZN(
        n16010) );
  OAI211_X1 U19326 ( .C1(n16012), .C2(n19999), .A(n16011), .B(n16010), .ZN(
        P1_U2987) );
  AOI22_X1 U19327 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16020) );
  NAND3_X1 U19328 ( .A1(n16014), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n12766), .ZN(n16016) );
  NAND2_X1 U19329 ( .A1(n16016), .A2(n16015), .ZN(n16017) );
  XNOR2_X1 U19330 ( .A(n16017), .B(n16089), .ZN(n16084) );
  AOI22_X1 U19331 ( .A1(n20169), .A2(n16084), .B1(n20159), .B2(n16018), .ZN(
        n16019) );
  OAI211_X1 U19332 ( .C1(n20163), .C2(n16021), .A(n16020), .B(n16019), .ZN(
        P1_U2988) );
  AOI22_X1 U19333 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16027) );
  NAND2_X1 U19334 ( .A1(n16023), .A2(n16022), .ZN(n16024) );
  XNOR2_X1 U19335 ( .A(n16025), .B(n16024), .ZN(n16126) );
  AOI22_X1 U19336 ( .A1(n16126), .A2(n20169), .B1(n20159), .B2(n20039), .ZN(
        n16026) );
  OAI211_X1 U19337 ( .C1(n20163), .C2(n20041), .A(n16027), .B(n16026), .ZN(
        P1_U2992) );
  AOI22_X1 U19338 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16033) );
  XNOR2_X1 U19339 ( .A(n16029), .B(n16028), .ZN(n16030) );
  XNOR2_X1 U19340 ( .A(n16031), .B(n16030), .ZN(n16137) );
  AOI22_X1 U19341 ( .A1(n16137), .A2(n20169), .B1(n20159), .B2(n20051), .ZN(
        n16032) );
  OAI211_X1 U19342 ( .C1(n20163), .C2(n20053), .A(n16033), .B(n16032), .ZN(
        P1_U2993) );
  AOI22_X1 U19343 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16039) );
  OAI21_X1 U19344 ( .B1(n16036), .B2(n16035), .A(n16034), .ZN(n16037) );
  INV_X1 U19345 ( .A(n16037), .ZN(n16143) );
  AOI22_X1 U19346 ( .A1(n16143), .A2(n20169), .B1(n20159), .B2(n20063), .ZN(
        n16038) );
  OAI211_X1 U19347 ( .C1(n20163), .C2(n20066), .A(n16039), .B(n16038), .ZN(
        P1_U2994) );
  OAI22_X1 U19348 ( .A1(n16040), .A2(n20224), .B1(n14804), .B2(n20208), .ZN(
        n16041) );
  AOI21_X1 U19349 ( .B1(n20228), .B2(n16042), .A(n16041), .ZN(n16043) );
  OAI221_X1 U19350 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16046), 
        .C1(n16045), .C2(n16044), .A(n16043), .ZN(P1_U3012) );
  AOI21_X1 U19351 ( .B1(n16095), .B2(n16047), .A(n16065), .ZN(n16064) );
  NOR2_X1 U19352 ( .A1(n16047), .A2(n16070), .ZN(n16052) );
  OAI22_X1 U19353 ( .A1(n16050), .A2(n16049), .B1(n20224), .B2(n16048), .ZN(
        n16051) );
  AOI21_X1 U19354 ( .B1(n16052), .B2(n16055), .A(n16051), .ZN(n16054) );
  NAND2_X1 U19355 ( .A1(n20164), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16053) );
  OAI211_X1 U19356 ( .C1(n16064), .C2(n16055), .A(n16054), .B(n16053), .ZN(
        P1_U3013) );
  AOI21_X1 U19357 ( .B1(n16057), .B2(n16056), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16063) );
  INV_X1 U19358 ( .A(n16058), .ZN(n16060) );
  AOI22_X1 U19359 ( .A1(n16060), .A2(n20228), .B1(n20186), .B2(n16059), .ZN(
        n16062) );
  NAND2_X1 U19360 ( .A1(n20164), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16061) );
  OAI211_X1 U19361 ( .C1(n16064), .C2(n16063), .A(n16062), .B(n16061), .ZN(
        P1_U3014) );
  AOI22_X1 U19362 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16065), .B1(
        n20164), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16069) );
  AOI22_X1 U19363 ( .A1(n16067), .A2(n20228), .B1(n20186), .B2(n16066), .ZN(
        n16068) );
  OAI211_X1 U19364 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16070), .A(
        n16069), .B(n16068), .ZN(P1_U3016) );
  INV_X1 U19365 ( .A(n16071), .ZN(n16073) );
  AOI21_X1 U19366 ( .B1(n20186), .B2(n16073), .A(n16072), .ZN(n16080) );
  NAND3_X1 U19367 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n16074), .ZN(n16076) );
  OAI21_X1 U19368 ( .B1(n16076), .B2(n20231), .A(n16075), .ZN(n16077) );
  AOI22_X1 U19369 ( .A1(n16078), .A2(n20228), .B1(n16081), .B2(n16077), .ZN(
        n16079) );
  OAI211_X1 U19370 ( .C1(n16082), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        P1_U3018) );
  AOI22_X1 U19371 ( .A1(n20186), .A2(n16083), .B1(n20164), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16088) );
  NOR2_X1 U19372 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16135), .ZN(
        n16085) );
  AOI22_X1 U19373 ( .A1(n16086), .A2(n16085), .B1(n20228), .B2(n16084), .ZN(
        n16087) );
  OAI211_X1 U19374 ( .C1(n16090), .C2(n16089), .A(n16088), .B(n16087), .ZN(
        P1_U3020) );
  INV_X1 U19375 ( .A(n16091), .ZN(n16093) );
  NOR2_X1 U19376 ( .A1(n16114), .A2(n16134), .ZN(n16092) );
  OAI211_X1 U19377 ( .C1(n16093), .C2(n16092), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16123), .ZN(n16094) );
  AOI21_X1 U19378 ( .B1(n16095), .B2(n16094), .A(n16112), .ZN(n16109) );
  NOR3_X1 U19379 ( .A1(n16135), .A2(n16134), .A3(n16028), .ZN(n16124) );
  NAND2_X1 U19380 ( .A1(n16123), .A2(n16124), .ZN(n16104) );
  AOI221_X1 U19381 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16102), .C2(n13764), .A(
        n16104), .ZN(n16099) );
  INV_X1 U19382 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n16096) );
  OAI22_X1 U19383 ( .A1(n20224), .A2(n16097), .B1(n16096), .B2(n20208), .ZN(
        n16098) );
  AOI211_X1 U19384 ( .C1(n16100), .C2(n20228), .A(n16099), .B(n16098), .ZN(
        n16101) );
  OAI21_X1 U19385 ( .B1(n16102), .B2(n16109), .A(n16101), .ZN(P1_U3021) );
  INV_X1 U19386 ( .A(n16103), .ZN(n16107) );
  NOR2_X1 U19387 ( .A1(n16104), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16106) );
  OAI22_X1 U19388 ( .A1(n20224), .A2(n20020), .B1(n20806), .B2(n20208), .ZN(
        n16105) );
  AOI211_X1 U19389 ( .C1(n16107), .C2(n20228), .A(n16106), .B(n16105), .ZN(
        n16108) );
  OAI21_X1 U19390 ( .B1(n13764), .B2(n16109), .A(n16108), .ZN(P1_U3022) );
  OAI21_X1 U19391 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16124), .ZN(n16122) );
  AOI21_X1 U19392 ( .B1(n20186), .B2(n16111), .A(n16110), .ZN(n16121) );
  NOR2_X1 U19393 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20176), .ZN(
        n16141) );
  NAND2_X1 U19394 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16113) );
  AOI21_X1 U19395 ( .B1(n16114), .B2(n16113), .A(n16112), .ZN(n20203) );
  OAI21_X1 U19396 ( .B1(n20194), .B2(n16116), .A(n20203), .ZN(n20189) );
  AOI21_X1 U19397 ( .B1(n16114), .B2(n20176), .A(n20189), .ZN(n16115) );
  OAI21_X1 U19398 ( .B1(n16117), .B2(n16116), .A(n16115), .ZN(n16144) );
  AOI21_X1 U19399 ( .B1(n16118), .B2(n16141), .A(n16144), .ZN(n16140) );
  OAI21_X1 U19400 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n20215), .A(
        n16140), .ZN(n16127) );
  AOI22_X1 U19401 ( .A1(n20228), .A2(n16119), .B1(n16127), .B2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16120) );
  OAI211_X1 U19402 ( .C1(n16123), .C2(n16122), .A(n16121), .B(n16120), .ZN(
        P1_U3023) );
  INV_X1 U19403 ( .A(n16124), .ZN(n16130) );
  AOI22_X1 U19404 ( .A1(n20186), .A2(n16125), .B1(n20164), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16129) );
  AOI22_X1 U19405 ( .A1(n16127), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20228), .B2(n16126), .ZN(n16128) );
  OAI211_X1 U19406 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16130), .A(
        n16129), .B(n16128), .ZN(P1_U3024) );
  INV_X1 U19407 ( .A(n16131), .ZN(n20044) );
  INV_X1 U19408 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n16132) );
  OAI22_X1 U19409 ( .A1(n20224), .A2(n20044), .B1(n20208), .B2(n16132), .ZN(
        n16133) );
  INV_X1 U19410 ( .A(n16133), .ZN(n16139) );
  NOR2_X1 U19411 ( .A1(n16135), .A2(n16134), .ZN(n16136) );
  AOI22_X1 U19412 ( .A1(n16137), .A2(n20228), .B1(n16136), .B2(n16028), .ZN(
        n16138) );
  OAI211_X1 U19413 ( .C1(n16140), .C2(n16028), .A(n16139), .B(n16138), .ZN(
        P1_U3025) );
  INV_X1 U19414 ( .A(n16141), .ZN(n16147) );
  NAND2_X1 U19415 ( .A1(n20194), .A2(n16142), .ZN(n20192) );
  AOI22_X1 U19416 ( .A1(n20186), .A2(n20055), .B1(n20164), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16146) );
  AOI22_X1 U19417 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16144), .B1(
        n16143), .B2(n20228), .ZN(n16145) );
  OAI211_X1 U19418 ( .C1(n16147), .C2(n20192), .A(n16146), .B(n16145), .ZN(
        P1_U3026) );
  NAND3_X1 U19419 ( .A1(n16149), .A2(n19990), .A3(n16148), .ZN(n16150) );
  OAI21_X1 U19420 ( .B1(n16151), .B2(n11963), .A(n16150), .ZN(P1_U3468) );
  INV_X1 U19421 ( .A(n16164), .ZN(n16153) );
  OR3_X1 U19422 ( .A1(n16155), .A2(n16153), .A3(n16152), .ZN(n16161) );
  NOR3_X1 U19423 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n16155), .A3(n16154), 
        .ZN(n16157) );
  NOR2_X1 U19424 ( .A1(n16157), .A2(n16156), .ZN(n20779) );
  AOI21_X1 U19425 ( .B1(n20779), .B2(n16159), .A(n16158), .ZN(n16160) );
  AOI21_X1 U19426 ( .B1(n16162), .B2(n16161), .A(n16160), .ZN(P1_U3162) );
  OAI221_X1 U19427 ( .B1(n20615), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20615), 
        .C2(n16164), .A(n16163), .ZN(P1_U3466) );
  INV_X1 U19428 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19914) );
  INV_X1 U19429 ( .A(n16165), .ZN(n16168) );
  INV_X1 U19430 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16167) );
  OAI222_X1 U19431 ( .A1(n19133), .A2(n19914), .B1(n19142), .B2(n16168), .C1(
        n16167), .C2(n16166), .ZN(n16169) );
  AOI21_X1 U19432 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19138), .A(
        n16169), .ZN(n16173) );
  INV_X1 U19433 ( .A(n19161), .ZN(n16170) );
  AOI22_X1 U19434 ( .A1(n16171), .A2(n19109), .B1(n19089), .B2(n16170), .ZN(
        n16172) );
  OAI211_X1 U19435 ( .C1(n16175), .C2(n16174), .A(n16173), .B(n16172), .ZN(
        P2_U2824) );
  AOI22_X1 U19436 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19145), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19128), .ZN(n16185) );
  AOI22_X1 U19437 ( .A1(n16176), .A2(n19129), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19138), .ZN(n16184) );
  OAI22_X1 U19438 ( .A1(n15125), .A2(n19151), .B1(n16177), .B2(n19150), .ZN(
        n16178) );
  INV_X1 U19439 ( .A(n16178), .ZN(n16183) );
  OAI211_X1 U19440 ( .C1(n16181), .C2(n16180), .A(n19154), .B(n16179), .ZN(
        n16182) );
  NAND4_X1 U19441 ( .A1(n16185), .A2(n16184), .A3(n16183), .A4(n16182), .ZN(
        P2_U2826) );
  AOI22_X1 U19442 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n19145), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n19128), .ZN(n16198) );
  OAI22_X1 U19443 ( .A1(n16187), .A2(n19142), .B1(n19158), .B2(n16186), .ZN(
        n16188) );
  INV_X1 U19444 ( .A(n16188), .ZN(n16197) );
  OAI22_X1 U19445 ( .A1(n16190), .A2(n19151), .B1(n16189), .B2(n19150), .ZN(
        n16191) );
  INV_X1 U19446 ( .A(n16191), .ZN(n16196) );
  OAI211_X1 U19447 ( .C1(n16194), .C2(n16193), .A(n19154), .B(n16192), .ZN(
        n16195) );
  NAND4_X1 U19448 ( .A1(n16198), .A2(n16197), .A3(n16196), .A4(n16195), .ZN(
        P2_U2828) );
  AOI22_X1 U19449 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19145), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19128), .ZN(n16210) );
  AOI22_X1 U19450 ( .A1(n16199), .A2(n19129), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19138), .ZN(n16209) );
  INV_X1 U19451 ( .A(n16200), .ZN(n16203) );
  INV_X1 U19452 ( .A(n16201), .ZN(n16202) );
  AOI22_X1 U19453 ( .A1(n16203), .A2(n19109), .B1(n16202), .B2(n19089), .ZN(
        n16208) );
  OAI211_X1 U19454 ( .C1(n16206), .C2(n16205), .A(n19154), .B(n16204), .ZN(
        n16207) );
  NAND4_X1 U19455 ( .A1(n16210), .A2(n16209), .A3(n16208), .A4(n16207), .ZN(
        P2_U2829) );
  INV_X1 U19456 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19901) );
  OAI22_X1 U19457 ( .A1(n19143), .A2(n16219), .B1(n19901), .B2(n19133), .ZN(
        n16211) );
  AOI21_X1 U19458 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19138), .A(
        n16211), .ZN(n16224) );
  INV_X1 U19459 ( .A(n16212), .ZN(n16214) );
  AOI22_X1 U19460 ( .A1(n16214), .A2(n19109), .B1(n19089), .B2(n16213), .ZN(
        n16223) );
  OAI211_X1 U19461 ( .C1(n16217), .C2(n16216), .A(n19154), .B(n16215), .ZN(
        n16222) );
  OAI211_X1 U19462 ( .C1(n16220), .C2(n16219), .A(n16218), .B(n19129), .ZN(
        n16221) );
  NAND4_X1 U19463 ( .A1(n16224), .A2(n16223), .A3(n16222), .A4(n16221), .ZN(
        P2_U2830) );
  OAI22_X1 U19464 ( .A1(n19143), .A2(n10489), .B1(n19897), .B2(n19133), .ZN(
        n16225) );
  AOI21_X1 U19465 ( .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19138), .A(
        n16225), .ZN(n16226) );
  OAI21_X1 U19466 ( .B1(n16227), .B2(n19142), .A(n16226), .ZN(n16228) );
  AOI21_X1 U19467 ( .B1(n9875), .B2(n19109), .A(n16228), .ZN(n16233) );
  OAI211_X1 U19468 ( .C1(n16231), .C2(n16230), .A(n19154), .B(n16229), .ZN(
        n16232) );
  OAI211_X1 U19469 ( .C1(n19150), .C2(n16234), .A(n16233), .B(n16232), .ZN(
        P2_U2832) );
  AOI22_X1 U19470 ( .A1(n19166), .A2(n16235), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19190), .ZN(n16240) );
  AOI22_X1 U19471 ( .A1(n19168), .A2(BUF1_REG_22__SCAN_IN), .B1(n19167), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16239) );
  AOI22_X1 U19472 ( .A1(n16237), .A2(n19194), .B1(n16246), .B2(n16236), .ZN(
        n16238) );
  NAND3_X1 U19473 ( .A1(n16240), .A2(n16239), .A3(n16238), .ZN(P2_U2897) );
  AOI22_X1 U19474 ( .A1(n19166), .A2(n19326), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19190), .ZN(n16244) );
  AOI22_X1 U19475 ( .A1(n19168), .A2(BUF1_REG_20__SCAN_IN), .B1(n19167), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16243) );
  AOI22_X1 U19476 ( .A1(n16241), .A2(n19194), .B1(n16246), .B2(n19005), .ZN(
        n16242) );
  NAND3_X1 U19477 ( .A1(n16244), .A2(n16243), .A3(n16242), .ZN(P2_U2899) );
  AOI22_X1 U19478 ( .A1(n19166), .A2(n19314), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19190), .ZN(n16250) );
  AOI22_X1 U19479 ( .A1(n19168), .A2(BUF1_REG_18__SCAN_IN), .B1(n19167), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16249) );
  AOI22_X1 U19480 ( .A1(n16247), .A2(n19194), .B1(n16246), .B2(n16245), .ZN(
        n16248) );
  NAND3_X1 U19481 ( .A1(n16250), .A2(n16249), .A3(n16248), .ZN(P2_U2901) );
  AOI22_X1 U19482 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19275), .B1(n19274), 
        .B2(n16251), .ZN(n16256) );
  OAI22_X1 U19483 ( .A1(n16253), .A2(n16292), .B1(n19282), .B2(n16252), .ZN(
        n16254) );
  AOI21_X1 U19484 ( .B1(n19278), .B2(n9875), .A(n16254), .ZN(n16255) );
  OAI211_X1 U19485 ( .C1(n19288), .C2(n9925), .A(n16256), .B(n16255), .ZN(
        P2_U2991) );
  AOI22_X1 U19486 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19275), .ZN(n16264) );
  NAND3_X1 U19487 ( .A1(n16258), .A2(n16257), .A3(n16310), .ZN(n16259) );
  OAI21_X1 U19488 ( .B1(n16317), .B2(n16260), .A(n16259), .ZN(n16261) );
  AOI21_X1 U19489 ( .B1(n16262), .B2(n19276), .A(n16261), .ZN(n16263) );
  OAI211_X1 U19490 ( .C1(n16314), .C2(n16265), .A(n16264), .B(n16263), .ZN(
        P2_U2992) );
  AOI22_X1 U19491 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19275), .ZN(n16270) );
  INV_X1 U19492 ( .A(n16266), .ZN(n16267) );
  AOI222_X1 U19493 ( .A1(n16268), .A2(n19276), .B1(n19278), .B2(n19081), .C1(
        n16310), .C2(n16267), .ZN(n16269) );
  OAI211_X1 U19494 ( .C1(n16314), .C2(n16271), .A(n16270), .B(n16269), .ZN(
        P2_U3002) );
  AOI22_X1 U19495 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19275), .B1(n19274), 
        .B2(n16272), .ZN(n16277) );
  OAI22_X1 U19496 ( .A1(n16274), .A2(n19282), .B1(n16273), .B2(n16292), .ZN(
        n16275) );
  AOI21_X1 U19497 ( .B1(n19278), .B2(n19095), .A(n16275), .ZN(n16276) );
  OAI211_X1 U19498 ( .C1(n19288), .C2(n19085), .A(n16277), .B(n16276), .ZN(
        P2_U3003) );
  AOI22_X1 U19499 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19275), .ZN(n16289) );
  AOI21_X1 U19500 ( .B1(n16278), .B2(n15644), .A(n9843), .ZN(n16329) );
  NOR2_X1 U19501 ( .A1(n16280), .A2(n16279), .ZN(n16284) );
  NAND2_X1 U19502 ( .A1(n16282), .A2(n16281), .ZN(n16283) );
  XNOR2_X1 U19503 ( .A(n16284), .B(n16283), .ZN(n16332) );
  OAI22_X1 U19504 ( .A1(n16332), .A2(n16292), .B1(n16317), .B2(n16285), .ZN(
        n16286) );
  AOI21_X1 U19505 ( .B1(n16329), .B2(n16287), .A(n16286), .ZN(n16288) );
  OAI211_X1 U19506 ( .C1(n16314), .C2(n19108), .A(n16289), .B(n16288), .ZN(
        P2_U3004) );
  AOI22_X1 U19507 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19275), .B1(n19274), 
        .B2(n16290), .ZN(n16297) );
  INV_X1 U19508 ( .A(n19119), .ZN(n16295) );
  OAI22_X1 U19509 ( .A1(n16293), .A2(n19282), .B1(n16292), .B2(n16291), .ZN(
        n16294) );
  AOI21_X1 U19510 ( .B1(n19278), .B2(n16295), .A(n16294), .ZN(n16296) );
  OAI211_X1 U19511 ( .C1(n19288), .C2(n16298), .A(n16297), .B(n16296), .ZN(
        P2_U3005) );
  AOI22_X1 U19512 ( .A1(n16299), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19275), .ZN(n16312) );
  NAND2_X1 U19513 ( .A1(n16301), .A2(n16300), .ZN(n16305) );
  NAND2_X1 U19514 ( .A1(n16303), .A2(n16302), .ZN(n16304) );
  XNOR2_X1 U19515 ( .A(n16305), .B(n16304), .ZN(n16340) );
  OAI21_X1 U19516 ( .B1(n16308), .B2(n16307), .A(n16306), .ZN(n16309) );
  INV_X1 U19517 ( .A(n16309), .ZN(n16336) );
  AOI222_X1 U19518 ( .A1(n16340), .A2(n19276), .B1(n19278), .B2(n16338), .C1(
        n16310), .C2(n16336), .ZN(n16311) );
  OAI211_X1 U19519 ( .C1(n16314), .C2(n16313), .A(n16312), .B(n16311), .ZN(
        P2_U3006) );
  AOI22_X1 U19520 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19275), .B1(n19274), 
        .B2(n16315), .ZN(n16322) );
  OAI22_X1 U19521 ( .A1(n16318), .A2(n19282), .B1(n16317), .B2(n16316), .ZN(
        n16319) );
  AOI21_X1 U19522 ( .B1(n19276), .B2(n16320), .A(n16319), .ZN(n16321) );
  OAI211_X1 U19523 ( .C1(n19288), .C2(n16323), .A(n16322), .B(n16321), .ZN(
        P2_U3008) );
  NOR2_X1 U19524 ( .A1(n11445), .A2(n19131), .ZN(n16327) );
  XNOR2_X1 U19525 ( .A(n13157), .B(n16324), .ZN(n19186) );
  OAI22_X1 U19526 ( .A1(n19186), .A2(n16360), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16325), .ZN(n16326) );
  AOI211_X1 U19527 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16328), .A(
        n16327), .B(n16326), .ZN(n16331) );
  AOI22_X1 U19528 ( .A1(n16329), .A2(n16337), .B1(n16339), .B2(n19110), .ZN(
        n16330) );
  OAI211_X1 U19529 ( .C1(n16332), .C2(n16369), .A(n16331), .B(n16330), .ZN(
        P2_U3036) );
  OAI22_X1 U19530 ( .A1(n16334), .A2(n16333), .B1(n16360), .B2(n19189), .ZN(
        n16335) );
  INV_X1 U19531 ( .A(n16335), .ZN(n16346) );
  AOI222_X1 U19532 ( .A1(n16340), .A2(n19303), .B1(n16339), .B2(n16338), .C1(
        n16337), .C2(n16336), .ZN(n16345) );
  NAND2_X1 U19533 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19275), .ZN(n16344) );
  OAI211_X1 U19534 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16342), .B(n16341), .ZN(n16343) );
  NAND4_X1 U19535 ( .A1(n16346), .A2(n16345), .A3(n16344), .A4(n16343), .ZN(
        P2_U3038) );
  OAI21_X1 U19536 ( .B1(n13154), .B2(n19296), .A(n16347), .ZN(n16348) );
  AOI21_X1 U19537 ( .B1(n16349), .B2(n19301), .A(n16348), .ZN(n16350) );
  OAI21_X1 U19538 ( .B1(n16351), .B2(n19295), .A(n16350), .ZN(n16352) );
  AOI21_X1 U19539 ( .B1(n16353), .B2(n19303), .A(n16352), .ZN(n16354) );
  OAI221_X1 U19540 ( .B1(n16357), .B2(n16356), .C1(n16357), .C2(n16355), .A(
        n16354), .ZN(P2_U3043) );
  INV_X1 U19541 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16365) );
  OAI22_X1 U19542 ( .A1(n16365), .A2(n16358), .B1(n19296), .B2(n10073), .ZN(
        n16363) );
  OAI22_X1 U19543 ( .A1(n19295), .A2(n16361), .B1(n16360), .B2(n16359), .ZN(
        n16362) );
  AOI211_X1 U19544 ( .C1(n16365), .C2(n16364), .A(n16363), .B(n16362), .ZN(
        n16367) );
  OAI211_X1 U19545 ( .C1(n16369), .C2(n16368), .A(n16367), .B(n16366), .ZN(
        P2_U3046) );
  MUX2_X1 U19546 ( .A(n16371), .B(n16370), .S(n16404), .Z(n16407) );
  INV_X1 U19547 ( .A(n16404), .ZN(n16381) );
  INV_X1 U19548 ( .A(n16372), .ZN(n16374) );
  OAI211_X1 U19549 ( .C1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16374), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16373), .ZN(n16376) );
  NAND2_X1 U19550 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16374), .ZN(
        n16375) );
  AND2_X1 U19551 ( .A1(n16376), .A2(n16375), .ZN(n16377) );
  NAND2_X1 U19552 ( .A1(n16381), .A2(n16377), .ZN(n16378) );
  AOI21_X1 U19553 ( .B1(n16407), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16378), .ZN(n16385) );
  AND2_X1 U19554 ( .A1(n16404), .A2(n16379), .ZN(n16380) );
  AOI21_X1 U19555 ( .B1(n16382), .B2(n16381), .A(n16380), .ZN(n16384) );
  NOR2_X1 U19556 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16407), .ZN(
        n16383) );
  NOR3_X1 U19557 ( .A1(n16385), .A2(n16384), .A3(n16383), .ZN(n16387) );
  INV_X1 U19558 ( .A(n16384), .ZN(n16406) );
  INV_X1 U19559 ( .A(n16385), .ZN(n16386) );
  OAI22_X1 U19560 ( .A1(n16387), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n16406), .B2(n16386), .ZN(n16409) );
  INV_X1 U19561 ( .A(n11360), .ZN(n16390) );
  NOR4_X1 U19562 ( .A1(n16398), .A2(n16390), .A3(n16389), .A4(n16388), .ZN(
        n18966) );
  OAI21_X1 U19563 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18966), .ZN(n16396) );
  INV_X1 U19564 ( .A(n16391), .ZN(n16392) );
  NAND3_X1 U19565 ( .A1(n16394), .A2(n16393), .A3(n16392), .ZN(n16395) );
  OAI211_X1 U19566 ( .C1(n16397), .C2(n10538), .A(n16396), .B(n16395), .ZN(
        n16403) );
  AOI22_X1 U19567 ( .A1(n16402), .A2(n16399), .B1(n11360), .B2(n16398), .ZN(
        n16400) );
  OAI21_X1 U19568 ( .B1(n16402), .B2(n16401), .A(n16400), .ZN(n19960) );
  AOI211_X1 U19569 ( .C1(n16404), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16403), .B(n19960), .ZN(n16405) );
  OAI21_X1 U19570 ( .B1(n16407), .B2(n16406), .A(n16405), .ZN(n16408) );
  AOI21_X1 U19571 ( .B1(n16409), .B2(n15885), .A(n16408), .ZN(n16422) );
  NOR3_X1 U19572 ( .A1(n11337), .A2(n16410), .A3(n19969), .ZN(n16412) );
  INV_X1 U19573 ( .A(n19980), .ZN(n16411) );
  NOR3_X1 U19574 ( .A1(n16412), .A2(n16411), .A3(n19975), .ZN(n16418) );
  AOI22_X1 U19575 ( .A1(n19977), .A2(n16413), .B1(n19976), .B2(n16418), .ZN(
        n16416) );
  AOI211_X1 U19576 ( .C1(n16416), .C2(n20977), .A(n16415), .B(n16414), .ZN(
        n16421) );
  NOR3_X1 U19577 ( .A1(n16417), .A2(n19975), .A3(n16419), .ZN(n19953) );
  OAI221_X1 U19578 ( .B1(n16419), .B2(n20977), .C1(n16422), .C2(n20977), .A(
        n16418), .ZN(n16424) );
  INV_X1 U19579 ( .A(n16424), .ZN(n19842) );
  OAI21_X1 U19580 ( .B1(n19953), .B2(n19842), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16420) );
  OAI211_X1 U19581 ( .C1(n16422), .C2(n18965), .A(n16421), .B(n16420), .ZN(
        P2_U3176) );
  OAI221_X1 U19582 ( .B1(n19951), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19951), 
        .C2(n16424), .A(n16423), .ZN(P2_U3593) );
  NOR2_X1 U19583 ( .A1(n16427), .A2(n17720), .ZN(n17611) );
  INV_X1 U19584 ( .A(n17611), .ZN(n17630) );
  AOI21_X1 U19585 ( .B1(n16614), .B2(n16430), .A(n16429), .ZN(n16434) );
  OAI21_X1 U19586 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16445), .A(
        n16431), .ZN(n16613) );
  OAI21_X1 U19587 ( .B1(n17769), .B2(n16613), .A(n16432), .ZN(n16433) );
  AOI211_X1 U19588 ( .C1(n17573), .C2(n16435), .A(n16434), .B(n16433), .ZN(
        n16439) );
  NOR2_X1 U19589 ( .A1(n16436), .A2(n17920), .ZN(n16454) );
  NOR2_X1 U19590 ( .A1(n16437), .A2(n17753), .ZN(n16441) );
  OAI21_X1 U19591 ( .B1(n16454), .B2(n16441), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16438) );
  OAI211_X1 U19592 ( .C1(n16440), .C2(n17823), .A(n16439), .B(n16438), .ZN(
        P3_U2800) );
  OR2_X1 U19593 ( .A1(n17923), .A2(n16453), .ZN(n16475) );
  INV_X1 U19594 ( .A(n16441), .ZN(n16442) );
  AOI21_X1 U19595 ( .B1(n16443), .B2(n16475), .A(n16442), .ZN(n16451) );
  NAND2_X1 U19596 ( .A1(n18140), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16448) );
  AOI21_X1 U19597 ( .B1(n9948), .B2(n16605), .A(n16445), .ZN(n16622) );
  OAI21_X1 U19598 ( .B1(n16446), .B2(n17667), .A(n16622), .ZN(n16447) );
  OAI211_X1 U19599 ( .C1(n16449), .C2(n9949), .A(n16448), .B(n16447), .ZN(
        n16450) );
  AOI211_X1 U19600 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16452), .A(
        n16451), .B(n16450), .ZN(n16456) );
  NOR2_X1 U19601 ( .A1(n16453), .A2(n17924), .ZN(n16472) );
  OAI21_X1 U19602 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16472), .A(
        n16454), .ZN(n16455) );
  OAI211_X1 U19603 ( .C1(n16457), .C2(n17823), .A(n16456), .B(n16455), .ZN(
        P3_U2801) );
  NAND2_X1 U19604 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18900), .ZN(
        n16459) );
  NOR4_X1 U19605 ( .A1(n17948), .A2(n16459), .A3(n16458), .A4(n18245), .ZN(
        n16463) );
  NAND2_X1 U19606 ( .A1(n18224), .A2(n18149), .ZN(n18231) );
  AOI221_X1 U19607 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16460), 
        .C1(n18231), .C2(n16460), .A(n18900), .ZN(n16462) );
  AOI211_X1 U19608 ( .C1(n16464), .C2(n16463), .A(n16462), .B(n16461), .ZN(
        n16468) );
  INV_X1 U19609 ( .A(n18088), .ZN(n18159) );
  AOI22_X1 U19610 ( .A1(n16466), .A2(n18159), .B1(n16465), .B2(n18244), .ZN(
        n16467) );
  OAI211_X1 U19611 ( .C1(n16469), .C2(n18161), .A(n16468), .B(n16467), .ZN(
        P3_U2831) );
  AOI22_X1 U19612 ( .A1(n17820), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n17551), .B2(n11132), .ZN(n17562) );
  OAI21_X1 U19613 ( .B1(n16485), .B2(n11132), .A(n17568), .ZN(n17561) );
  NAND2_X1 U19614 ( .A1(n17562), .A2(n17561), .ZN(n17560) );
  NAND4_X1 U19615 ( .A1(n18727), .A2(n16471), .A3(n16470), .A4(n17560), .ZN(
        n16479) );
  OR2_X1 U19616 ( .A1(n16472), .A2(n18723), .ZN(n16477) );
  INV_X1 U19617 ( .A(n16473), .ZN(n16474) );
  AOI21_X1 U19618 ( .B1(n16475), .B2(n18111), .A(n16474), .ZN(n16476) );
  AND2_X1 U19619 ( .A1(n16477), .A2(n16476), .ZN(n16478) );
  INV_X1 U19620 ( .A(n16481), .ZN(n18006) );
  AND3_X1 U19621 ( .A1(n17996), .A2(n16482), .A3(n18006), .ZN(n17960) );
  NOR2_X1 U19622 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16483), .ZN(
        n17547) );
  AND3_X1 U19623 ( .A1(n16485), .A2(n18242), .A3(n16484), .ZN(n16487) );
  NAND2_X1 U19624 ( .A1(n18140), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17556) );
  INV_X1 U19625 ( .A(n17556), .ZN(n16486) );
  AOI211_X1 U19626 ( .C1(n17960), .C2(n17547), .A(n16487), .B(n16486), .ZN(
        n16489) );
  OR3_X1 U19627 ( .A1(n17568), .A2(n18161), .A3(n17562), .ZN(n16488) );
  OAI211_X1 U19628 ( .C1(n17551), .C2(n16490), .A(n16489), .B(n16488), .ZN(
        P3_U2834) );
  NOR3_X1 U19629 ( .A1(P3_BE_N_REG_0__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16492) );
  NOR4_X1 U19630 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16491) );
  INV_X2 U19631 ( .A(n16566), .ZN(U215) );
  NAND4_X1 U19632 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16492), .A3(n16491), .A4(
        U215), .ZN(U213) );
  INV_X1 U19633 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19207) );
  INV_X2 U19634 ( .A(U214), .ZN(n20885) );
  NOR2_X1 U19635 ( .A1(n20885), .A2(n16493), .ZN(n20887) );
  INV_X1 U19636 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16571) );
  OAI222_X1 U19637 ( .A1(U212), .A2(n19207), .B1(n16536), .B2(n19338), .C1(
        U214), .C2(n16571), .ZN(U216) );
  AOI22_X1 U19638 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20885), .ZN(n16494) );
  OAI21_X1 U19639 ( .B1(n21113), .B2(n16536), .A(n16494), .ZN(U217) );
  AOI222_X1 U19640 ( .A1(n20885), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n20887), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n20886), .C2(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n16495) );
  INV_X1 U19641 ( .A(n16495), .ZN(U218) );
  AOI22_X1 U19642 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n20885), .ZN(n16496) );
  OAI21_X1 U19643 ( .B1(n16497), .B2(n16536), .A(n16496), .ZN(U219) );
  INV_X1 U19644 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16499) );
  AOI22_X1 U19645 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n20885), .ZN(n16498) );
  OAI21_X1 U19646 ( .B1(n16499), .B2(n16536), .A(n16498), .ZN(U220) );
  INV_X1 U19647 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16501) );
  AOI22_X1 U19648 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n20885), .ZN(n16500) );
  OAI21_X1 U19649 ( .B1(n16501), .B2(n16536), .A(n16500), .ZN(U221) );
  AOI22_X1 U19650 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n20885), .ZN(n16502) );
  OAI21_X1 U19651 ( .B1(n16503), .B2(n16536), .A(n16502), .ZN(U222) );
  INV_X1 U19652 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n21129) );
  AOI22_X1 U19653 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20887), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n20885), .ZN(n16504) );
  OAI21_X1 U19654 ( .B1(n21129), .B2(U212), .A(n16504), .ZN(U223) );
  INV_X1 U19655 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16506) );
  AOI22_X1 U19656 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n20885), .ZN(n16505) );
  OAI21_X1 U19657 ( .B1(n16506), .B2(n16536), .A(n16505), .ZN(U224) );
  AOI222_X1 U19658 ( .A1(n20885), .A2(P1_DATAO_REG_22__SCAN_IN), .B1(n20887), 
        .B2(BUF1_REG_22__SCAN_IN), .C1(n20886), .C2(P2_DATAO_REG_22__SCAN_IN), 
        .ZN(n16507) );
  INV_X1 U19659 ( .A(n16507), .ZN(U225) );
  AOI22_X1 U19660 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n20885), .ZN(n16508) );
  OAI21_X1 U19661 ( .B1(n16509), .B2(n16536), .A(n16508), .ZN(U226) );
  INV_X1 U19662 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19327) );
  AOI22_X1 U19663 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n20885), .ZN(n16510) );
  OAI21_X1 U19664 ( .B1(n19327), .B2(n16536), .A(n16510), .ZN(U227) );
  INV_X1 U19665 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n19321) );
  AOI22_X1 U19666 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n20885), .ZN(n16511) );
  OAI21_X1 U19667 ( .B1(n19321), .B2(n16536), .A(n16511), .ZN(U228) );
  AOI22_X1 U19668 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n20885), .ZN(n16512) );
  OAI21_X1 U19669 ( .B1(n19315), .B2(n16536), .A(n16512), .ZN(U229) );
  INV_X1 U19670 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20237) );
  AOI22_X1 U19671 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n20885), .ZN(n16513) );
  OAI21_X1 U19672 ( .B1(n20237), .B2(n16536), .A(n16513), .ZN(U230) );
  AOI22_X1 U19673 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20885), .ZN(n16514) );
  OAI21_X1 U19674 ( .B1(n21083), .B2(n16536), .A(n16514), .ZN(U231) );
  INV_X1 U19675 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16516) );
  AOI22_X1 U19676 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n20887), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n20885), .ZN(n16515) );
  OAI21_X1 U19677 ( .B1(n16516), .B2(U212), .A(n16515), .ZN(U232) );
  INV_X1 U19678 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16518) );
  AOI22_X1 U19679 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n20887), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n20885), .ZN(n16517) );
  OAI21_X1 U19680 ( .B1(n16518), .B2(U212), .A(n16517), .ZN(U233) );
  INV_X1 U19681 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16552) );
  AOI22_X1 U19682 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n20887), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n20885), .ZN(n16519) );
  OAI21_X1 U19683 ( .B1(n16552), .B2(U212), .A(n16519), .ZN(U234) );
  INV_X1 U19684 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n21116) );
  INV_X1 U19685 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16551) );
  OAI222_X1 U19686 ( .A1(U214), .A2(n21116), .B1(n16536), .B2(n16520), .C1(
        U212), .C2(n16551), .ZN(U235) );
  AOI22_X1 U19687 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n20885), .ZN(n16521) );
  OAI21_X1 U19688 ( .B1(n12889), .B2(n16536), .A(n16521), .ZN(U236) );
  AOI22_X1 U19689 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n20885), .ZN(n16522) );
  OAI21_X1 U19690 ( .B1(n16523), .B2(n16536), .A(n16522), .ZN(U237) );
  AOI22_X1 U19691 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n20885), .ZN(n16524) );
  OAI21_X1 U19692 ( .B1(n16525), .B2(n16536), .A(n16524), .ZN(U238) );
  AOI22_X1 U19693 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n20885), .ZN(n16526) );
  OAI21_X1 U19694 ( .B1(n16527), .B2(n16536), .A(n16526), .ZN(U239) );
  INV_X1 U19695 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16529) );
  AOI22_X1 U19696 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n20885), .ZN(n16528) );
  OAI21_X1 U19697 ( .B1(n16529), .B2(n16536), .A(n16528), .ZN(U240) );
  AOI222_X1 U19698 ( .A1(n20885), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n20887), 
        .B2(BUF1_REG_6__SCAN_IN), .C1(n20886), .C2(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n16530) );
  INV_X1 U19699 ( .A(n16530), .ZN(U241) );
  INV_X1 U19700 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16543) );
  AOI22_X1 U19701 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n20887), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n20885), .ZN(n16531) );
  OAI21_X1 U19702 ( .B1(n16543), .B2(U212), .A(n16531), .ZN(U242) );
  INV_X1 U19703 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16533) );
  AOI22_X1 U19704 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n20885), .ZN(n16532) );
  OAI21_X1 U19705 ( .B1(n16533), .B2(n16536), .A(n16532), .ZN(U243) );
  INV_X1 U19706 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16541) );
  AOI22_X1 U19707 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n20887), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n20885), .ZN(n16534) );
  OAI21_X1 U19708 ( .B1(n16541), .B2(U212), .A(n16534), .ZN(U244) );
  INV_X1 U19709 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16537) );
  AOI22_X1 U19710 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n20886), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n20885), .ZN(n16535) );
  OAI21_X1 U19711 ( .B1(n16537), .B2(n16536), .A(n16535), .ZN(U245) );
  AOI222_X1 U19712 ( .A1(n20885), .A2(P1_DATAO_REG_0__SCAN_IN), .B1(n20887), 
        .B2(BUF1_REG_0__SCAN_IN), .C1(n20886), .C2(P2_DATAO_REG_0__SCAN_IN), 
        .ZN(n16538) );
  INV_X1 U19713 ( .A(n16538), .ZN(U247) );
  INV_X1 U19714 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n21161) );
  INV_X1 U19715 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18264) );
  AOI22_X1 U19716 ( .A1(n16566), .A2(n21161), .B1(n18264), .B2(U215), .ZN(U251) );
  OAI22_X1 U19717 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16566), .ZN(n16539) );
  INV_X1 U19718 ( .A(n16539), .ZN(U252) );
  OAI22_X1 U19719 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16566), .ZN(n16540) );
  INV_X1 U19720 ( .A(n16540), .ZN(U253) );
  INV_X1 U19721 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18277) );
  AOI22_X1 U19722 ( .A1(n16566), .A2(n16541), .B1(n18277), .B2(U215), .ZN(U254) );
  OAI22_X1 U19723 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16566), .ZN(n16542) );
  INV_X1 U19724 ( .A(n16542), .ZN(U255) );
  INV_X1 U19725 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18286) );
  AOI22_X1 U19726 ( .A1(n16566), .A2(n16543), .B1(n18286), .B2(U215), .ZN(U256) );
  INV_X1 U19727 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16544) );
  INV_X1 U19728 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18290) );
  AOI22_X1 U19729 ( .A1(n16566), .A2(n16544), .B1(n18290), .B2(U215), .ZN(U257) );
  OAI22_X1 U19730 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16566), .ZN(n16545) );
  INV_X1 U19731 ( .A(n16545), .ZN(U258) );
  INV_X1 U19732 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16547) );
  INV_X1 U19733 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n16546) );
  AOI22_X1 U19734 ( .A1(n16569), .A2(n16547), .B1(n16546), .B2(U215), .ZN(U259) );
  OAI22_X1 U19735 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16566), .ZN(n16548) );
  INV_X1 U19736 ( .A(n16548), .ZN(U260) );
  OAI22_X1 U19737 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16566), .ZN(n16549) );
  INV_X1 U19738 ( .A(n16549), .ZN(U261) );
  OAI22_X1 U19739 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16566), .ZN(n16550) );
  INV_X1 U19740 ( .A(n16550), .ZN(U262) );
  INV_X1 U19741 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U19742 ( .A1(n16566), .A2(n16551), .B1(n17388), .B2(U215), .ZN(U263) );
  INV_X1 U19743 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U19744 ( .A1(n16569), .A2(n16552), .B1(n17383), .B2(U215), .ZN(U264) );
  OAI22_X1 U19745 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16566), .ZN(n16553) );
  INV_X1 U19746 ( .A(n16553), .ZN(U265) );
  OAI22_X1 U19747 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16566), .ZN(n16554) );
  INV_X1 U19748 ( .A(n16554), .ZN(U266) );
  OAI22_X1 U19749 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16569), .ZN(n16555) );
  INV_X1 U19750 ( .A(n16555), .ZN(U267) );
  OAI22_X1 U19751 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16569), .ZN(n16556) );
  INV_X1 U19752 ( .A(n16556), .ZN(U268) );
  OAI22_X1 U19753 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16569), .ZN(n16557) );
  INV_X1 U19754 ( .A(n16557), .ZN(U269) );
  OAI22_X1 U19755 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16569), .ZN(n16558) );
  INV_X1 U19756 ( .A(n16558), .ZN(U270) );
  OAI22_X1 U19757 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16569), .ZN(n16559) );
  INV_X1 U19758 ( .A(n16559), .ZN(U271) );
  OAI22_X1 U19759 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16566), .ZN(n16560) );
  INV_X1 U19760 ( .A(n16560), .ZN(U272) );
  INV_X1 U19761 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n21115) );
  INV_X1 U19762 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n17331) );
  AOI22_X1 U19763 ( .A1(n16566), .A2(n21115), .B1(n17331), .B2(U215), .ZN(U273) );
  OAI22_X1 U19764 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16569), .ZN(n16561) );
  INV_X1 U19765 ( .A(n16561), .ZN(U274) );
  AOI22_X1 U19766 ( .A1(n16566), .A2(n21129), .B1(n15261), .B2(U215), .ZN(U275) );
  OAI22_X1 U19767 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16566), .ZN(n16562) );
  INV_X1 U19768 ( .A(n16562), .ZN(U276) );
  OAI22_X1 U19769 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16569), .ZN(n16563) );
  INV_X1 U19770 ( .A(n16563), .ZN(U277) );
  OAI22_X1 U19771 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16566), .ZN(n16564) );
  INV_X1 U19772 ( .A(n16564), .ZN(U278) );
  OAI22_X1 U19773 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16566), .ZN(n16565) );
  INV_X1 U19774 ( .A(n16565), .ZN(U279) );
  INV_X1 U19775 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n21208) );
  INV_X1 U19776 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n17298) );
  AOI22_X1 U19777 ( .A1(n16566), .A2(n21208), .B1(n17298), .B2(U215), .ZN(U280) );
  OAI22_X1 U19778 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16566), .ZN(n16567) );
  INV_X1 U19779 ( .A(n16567), .ZN(U281) );
  INV_X1 U19780 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19336) );
  AOI22_X1 U19781 ( .A1(n16569), .A2(n19207), .B1(n19336), .B2(U215), .ZN(U282) );
  INV_X1 U19782 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16570) );
  AOI222_X1 U19783 ( .A1(n19207), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16571), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16570), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16572) );
  INV_X2 U19784 ( .A(n16574), .ZN(n16573) );
  INV_X1 U19785 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18840) );
  INV_X1 U19786 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19875) );
  AOI22_X1 U19787 ( .A1(n16573), .A2(n18840), .B1(n19875), .B2(n16574), .ZN(
        U347) );
  INV_X1 U19788 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18838) );
  INV_X1 U19789 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U19790 ( .A1(n16572), .A2(n18838), .B1(n19874), .B2(n16574), .ZN(
        U348) );
  INV_X1 U19791 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n21077) );
  INV_X1 U19792 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n21175) );
  AOI22_X1 U19793 ( .A1(n16573), .A2(n21077), .B1(n21175), .B2(n16574), .ZN(
        U349) );
  INV_X1 U19794 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18835) );
  INV_X1 U19795 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20991) );
  AOI22_X1 U19796 ( .A1(n16573), .A2(n18835), .B1(n20991), .B2(n16574), .ZN(
        U350) );
  INV_X1 U19797 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18833) );
  INV_X1 U19798 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19871) );
  AOI22_X1 U19799 ( .A1(n16573), .A2(n18833), .B1(n19871), .B2(n16574), .ZN(
        U351) );
  INV_X1 U19800 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18831) );
  AOI22_X1 U19801 ( .A1(n16573), .A2(n18831), .B1(n21024), .B2(n16574), .ZN(
        U352) );
  INV_X1 U19802 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18828) );
  INV_X1 U19803 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19869) );
  AOI22_X1 U19804 ( .A1(n16573), .A2(n18828), .B1(n19869), .B2(n16574), .ZN(
        U353) );
  INV_X1 U19805 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18825) );
  INV_X1 U19806 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19867) );
  AOI22_X1 U19807 ( .A1(n16573), .A2(n18825), .B1(n19867), .B2(n16574), .ZN(
        U354) );
  INV_X1 U19808 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18879) );
  INV_X1 U19809 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19913) );
  AOI22_X1 U19810 ( .A1(n16573), .A2(n18879), .B1(n19913), .B2(n16574), .ZN(
        U355) );
  INV_X1 U19811 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18877) );
  INV_X1 U19812 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19910) );
  AOI22_X1 U19813 ( .A1(n16573), .A2(n18877), .B1(n19910), .B2(n16574), .ZN(
        U356) );
  INV_X1 U19814 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18875) );
  INV_X1 U19815 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19908) );
  AOI22_X1 U19816 ( .A1(n16573), .A2(n18875), .B1(n19908), .B2(n16574), .ZN(
        U357) );
  INV_X1 U19817 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18874) );
  INV_X1 U19818 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U19819 ( .A1(n16573), .A2(n18874), .B1(n19905), .B2(n16574), .ZN(
        U358) );
  INV_X1 U19820 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18872) );
  INV_X1 U19821 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19904) );
  AOI22_X1 U19822 ( .A1(n16573), .A2(n18872), .B1(n19904), .B2(n16574), .ZN(
        U359) );
  INV_X1 U19823 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18871) );
  INV_X1 U19824 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19902) );
  AOI22_X1 U19825 ( .A1(n16573), .A2(n18871), .B1(n19902), .B2(n16574), .ZN(
        U360) );
  INV_X1 U19826 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18868) );
  INV_X1 U19827 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19900) );
  AOI22_X1 U19828 ( .A1(n16573), .A2(n18868), .B1(n19900), .B2(n16574), .ZN(
        U361) );
  INV_X1 U19829 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18865) );
  INV_X1 U19830 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19898) );
  AOI22_X1 U19831 ( .A1(n16573), .A2(n18865), .B1(n19898), .B2(n16574), .ZN(
        U362) );
  INV_X1 U19832 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18864) );
  INV_X1 U19833 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19896) );
  AOI22_X1 U19834 ( .A1(n16573), .A2(n18864), .B1(n19896), .B2(n16574), .ZN(
        U363) );
  INV_X1 U19835 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18861) );
  INV_X1 U19836 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U19837 ( .A1(n16573), .A2(n18861), .B1(n19894), .B2(n16574), .ZN(
        U364) );
  INV_X1 U19838 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n21092) );
  INV_X1 U19839 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19865) );
  AOI22_X1 U19840 ( .A1(n16573), .A2(n21092), .B1(n19865), .B2(n16574), .ZN(
        U365) );
  INV_X1 U19841 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18860) );
  INV_X1 U19842 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19892) );
  AOI22_X1 U19843 ( .A1(n16573), .A2(n18860), .B1(n19892), .B2(n16574), .ZN(
        U366) );
  INV_X1 U19844 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18858) );
  INV_X1 U19845 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U19846 ( .A1(n16573), .A2(n18858), .B1(n19890), .B2(n16574), .ZN(
        U367) );
  INV_X1 U19847 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18856) );
  INV_X1 U19848 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19889) );
  AOI22_X1 U19849 ( .A1(n16573), .A2(n18856), .B1(n19889), .B2(n16574), .ZN(
        U368) );
  INV_X1 U19850 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18854) );
  INV_X1 U19851 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19888) );
  AOI22_X1 U19852 ( .A1(n16573), .A2(n18854), .B1(n19888), .B2(n16574), .ZN(
        U369) );
  INV_X1 U19853 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18852) );
  INV_X1 U19854 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19886) );
  AOI22_X1 U19855 ( .A1(n16573), .A2(n18852), .B1(n19886), .B2(n16574), .ZN(
        U370) );
  INV_X1 U19856 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18850) );
  INV_X1 U19857 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U19858 ( .A1(n16572), .A2(n18850), .B1(n19884), .B2(n16574), .ZN(
        U371) );
  INV_X1 U19859 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18847) );
  INV_X1 U19860 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19882) );
  AOI22_X1 U19861 ( .A1(n16573), .A2(n18847), .B1(n19882), .B2(n16574), .ZN(
        U372) );
  INV_X1 U19862 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18846) );
  INV_X1 U19863 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19880) );
  AOI22_X1 U19864 ( .A1(n16573), .A2(n18846), .B1(n19880), .B2(n16574), .ZN(
        U373) );
  INV_X1 U19865 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18844) );
  INV_X1 U19866 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U19867 ( .A1(n16573), .A2(n18844), .B1(n19879), .B2(n16574), .ZN(
        U374) );
  INV_X1 U19868 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18842) );
  INV_X1 U19869 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19877) );
  AOI22_X1 U19870 ( .A1(n16572), .A2(n18842), .B1(n19877), .B2(n16574), .ZN(
        U375) );
  INV_X1 U19871 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18823) );
  INV_X1 U19872 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19863) );
  AOI22_X1 U19873 ( .A1(n16572), .A2(n18823), .B1(n19863), .B2(n16574), .ZN(
        U376) );
  INV_X1 U19874 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18822) );
  NAND2_X1 U19875 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18822), .ZN(n18810) );
  AOI22_X1 U19876 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18810), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18820), .ZN(n18888) );
  AOI21_X1 U19877 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18888), .ZN(n16575) );
  INV_X1 U19878 ( .A(n16575), .ZN(P3_U2633) );
  INV_X1 U19879 ( .A(n18796), .ZN(n16577) );
  OAI21_X1 U19880 ( .B1(n16582), .B2(n17443), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16576) );
  OAI21_X1 U19881 ( .B1(n16578), .B2(n16577), .A(n16576), .ZN(P3_U2634) );
  AOI21_X1 U19882 ( .B1(n18820), .B2(n18822), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16579) );
  AOI22_X1 U19883 ( .A1(n18945), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16579), 
        .B2(n18946), .ZN(P3_U2635) );
  OAI21_X1 U19884 ( .B1(n18806), .B2(BS16), .A(n18888), .ZN(n18886) );
  OAI21_X1 U19885 ( .B1(n18888), .B2(n16580), .A(n18886), .ZN(P3_U2636) );
  NOR3_X1 U19886 ( .A1(n16582), .A2(n16581), .A3(n18725), .ZN(n18780) );
  NOR2_X1 U19887 ( .A1(n18780), .A2(n18784), .ZN(n18928) );
  OAI21_X1 U19888 ( .B1(n18928), .B2(n18250), .A(n16583), .ZN(P3_U2637) );
  NOR4_X1 U19889 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_18__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n16587) );
  NOR4_X1 U19890 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_14__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(n16586) );
  NOR4_X1 U19891 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16585) );
  NOR4_X1 U19892 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_23__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16584) );
  NAND4_X1 U19893 ( .A1(n16587), .A2(n16586), .A3(n16585), .A4(n16584), .ZN(
        n16593) );
  NOR4_X1 U19894 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n16591) );
  AOI211_X1 U19895 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_29__SCAN_IN), .B(
        P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(n16590) );
  NOR4_X1 U19896 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n16589) );
  NOR4_X1 U19897 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n16588) );
  NAND4_X1 U19898 ( .A1(n16591), .A2(n16590), .A3(n16589), .A4(n16588), .ZN(
        n16592) );
  NOR2_X1 U19899 ( .A1(n16593), .A2(n16592), .ZN(n18922) );
  INV_X1 U19900 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16595) );
  NOR3_X1 U19901 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16596) );
  OAI21_X1 U19902 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16596), .A(n18922), .ZN(
        n16594) );
  OAI21_X1 U19903 ( .B1(n18922), .B2(n16595), .A(n16594), .ZN(P3_U2638) );
  INV_X1 U19904 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18918) );
  INV_X1 U19905 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18887) );
  AOI21_X1 U19906 ( .B1(n18918), .B2(n18887), .A(n16596), .ZN(n16598) );
  INV_X1 U19907 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16597) );
  INV_X1 U19908 ( .A(n18922), .ZN(n18925) );
  AOI22_X1 U19909 ( .A1(n18922), .A2(n16598), .B1(n16597), .B2(n18925), .ZN(
        P3_U2639) );
  INV_X1 U19910 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17007) );
  NAND2_X1 U19911 ( .A1(n16647), .A2(n17007), .ZN(n16646) );
  NOR2_X1 U19912 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16646), .ZN(n16630) );
  INV_X1 U19913 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16995) );
  NAND2_X1 U19914 ( .A1(n16630), .A2(n16995), .ZN(n16612) );
  NOR2_X1 U19915 ( .A1(n16947), .A2(n16612), .ZN(n16618) );
  INV_X1 U19916 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16967) );
  INV_X1 U19917 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18880) );
  NAND4_X1 U19918 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16640), .ZN(n16603) );
  NOR3_X1 U19919 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18880), .A3(n16603), 
        .ZN(n16602) );
  AOI22_X1 U19920 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16939), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16955), .ZN(n16600) );
  INV_X1 U19921 ( .A(n16600), .ZN(n16601) );
  AOI211_X1 U19922 ( .C1(n16618), .C2(n16967), .A(n16602), .B(n16601), .ZN(
        n16611) );
  NOR2_X1 U19923 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16603), .ZN(n16617) );
  NAND3_X1 U19924 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16604) );
  AOI21_X1 U19925 ( .B1(n16935), .B2(n16604), .A(n16645), .ZN(n16615) );
  INV_X1 U19926 ( .A(n16615), .ZN(n16625) );
  OAI21_X1 U19927 ( .B1(n16617), .B2(n16625), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16610) );
  INV_X1 U19928 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17571) );
  NOR2_X1 U19929 ( .A1(n17571), .A2(n16607), .ZN(n16606) );
  OAI21_X1 U19930 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16606), .A(
        n16605), .ZN(n17557) );
  INV_X1 U19931 ( .A(n17557), .ZN(n16633) );
  AOI21_X1 U19932 ( .B1(n17571), .B2(n16607), .A(n16606), .ZN(n17566) );
  NOR2_X1 U19933 ( .A1(n16608), .A2(n16884), .ZN(n16642) );
  NOR2_X1 U19934 ( .A1(n16622), .A2(n16621), .ZN(n16620) );
  NAND4_X1 U19935 ( .A1(n16913), .A2(n16941), .A3(n16620), .A4(n16613), .ZN(
        n16609) );
  NAND3_X1 U19936 ( .A1(n16611), .A2(n16610), .A3(n16609), .ZN(P3_U2640) );
  NAND2_X1 U19937 ( .A1(n16954), .A2(n16612), .ZN(n16628) );
  OAI22_X1 U19938 ( .A1(n16615), .A2(n18880), .B1(n16614), .B2(n16938), .ZN(
        n16616) );
  OAI21_X1 U19939 ( .B1(n16955), .B2(n16618), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16619) );
  NOR2_X1 U19940 ( .A1(n16630), .A2(n16995), .ZN(n16629) );
  AOI211_X1 U19941 ( .C1(n16622), .C2(n16621), .A(n16620), .B(n18800), .ZN(
        n16624) );
  OAI22_X1 U19942 ( .A1(n9948), .A2(n16938), .B1(n16942), .B2(n16995), .ZN(
        n16623) );
  AOI211_X1 U19943 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16625), .A(n16624), 
        .B(n16623), .ZN(n16627) );
  INV_X1 U19944 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20979) );
  NAND4_X1 U19945 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16640), .A4(n20979), .ZN(n16626) );
  OAI211_X1 U19946 ( .C1(n16629), .C2(n16628), .A(n16627), .B(n16626), .ZN(
        P3_U2642) );
  INV_X1 U19947 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16639) );
  AOI22_X1 U19948 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16645), .B1(n16955), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16638) );
  INV_X1 U19949 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18873) );
  INV_X1 U19950 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18876) );
  AOI22_X1 U19951 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .B1(n18873), .B2(n18876), .ZN(n16636) );
  AOI211_X1 U19952 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16646), .A(n16630), .B(
        n16947), .ZN(n16635) );
  AOI211_X1 U19953 ( .C1(n16633), .C2(n16632), .A(n16631), .B(n18800), .ZN(
        n16634) );
  AOI211_X1 U19954 ( .C1(n16640), .C2(n16636), .A(n16635), .B(n16634), .ZN(
        n16637) );
  OAI211_X1 U19955 ( .C1(n16639), .C2(n16938), .A(n16638), .B(n16637), .ZN(
        P3_U2643) );
  INV_X1 U19956 ( .A(n16640), .ZN(n16650) );
  AOI211_X1 U19957 ( .C1(n17566), .C2(n16642), .A(n16641), .B(n18800), .ZN(
        n16644) );
  OAI22_X1 U19958 ( .A1(n17571), .A2(n16938), .B1(n16942), .B2(n17007), .ZN(
        n16643) );
  AOI211_X1 U19959 ( .C1(n16645), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16644), 
        .B(n16643), .ZN(n16649) );
  OAI211_X1 U19960 ( .C1(n16647), .C2(n17007), .A(n16954), .B(n16646), .ZN(
        n16648) );
  OAI211_X1 U19961 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16650), .A(n16649), 
        .B(n16648), .ZN(P3_U2644) );
  INV_X1 U19962 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18867) );
  OAI21_X1 U19963 ( .B1(n16673), .B2(n16943), .A(n16957), .ZN(n16670) );
  AOI21_X1 U19964 ( .B1(n16935), .B2(n18867), .A(n16670), .ZN(n16661) );
  INV_X1 U19965 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18870) );
  AOI211_X1 U19966 ( .C1(n17590), .C2(n16652), .A(n16651), .B(n18800), .ZN(
        n16655) );
  OAI22_X1 U19967 ( .A1(n16653), .A2(n16938), .B1(n16942), .B2(n16658), .ZN(
        n16654) );
  AOI211_X1 U19968 ( .C1(n16656), .C2(n18870), .A(n16655), .B(n16654), .ZN(
        n16660) );
  OAI211_X1 U19969 ( .C1(n16663), .C2(n16658), .A(n16954), .B(n16657), .ZN(
        n16659) );
  OAI211_X1 U19970 ( .C1(n16661), .C2(n18870), .A(n16660), .B(n16659), .ZN(
        P3_U2646) );
  NOR2_X1 U19971 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16943), .ZN(n16662) );
  AOI22_X1 U19972 ( .A1(n16955), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16673), 
        .B2(n16662), .ZN(n16669) );
  AOI211_X1 U19973 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16678), .A(n16663), .B(
        n16947), .ZN(n16667) );
  AOI211_X1 U19974 ( .C1(n17602), .C2(n16665), .A(n16664), .B(n18800), .ZN(
        n16666) );
  AOI211_X1 U19975 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16670), .A(n16667), 
        .B(n16666), .ZN(n16668) );
  OAI211_X1 U19976 ( .C1(n17604), .C2(n16938), .A(n16669), .B(n16668), .ZN(
        P3_U2647) );
  INV_X1 U19977 ( .A(n16670), .ZN(n16682) );
  AOI211_X1 U19978 ( .C1(n16672), .C2(n9856), .A(n16671), .B(n18800), .ZN(
        n16677) );
  INV_X1 U19979 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17619) );
  OR2_X1 U19980 ( .A1(n16943), .A2(n16673), .ZN(n16674) );
  OAI22_X1 U19981 ( .A1(n17619), .A2(n16938), .B1(n16675), .B2(n16674), .ZN(
        n16676) );
  AOI211_X1 U19982 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16955), .A(n16677), .B(
        n16676), .ZN(n16681) );
  OAI211_X1 U19983 ( .C1(n16685), .C2(n16679), .A(n16954), .B(n16678), .ZN(
        n16680) );
  OAI211_X1 U19984 ( .C1(n16682), .C2(n18866), .A(n16681), .B(n16680), .ZN(
        P3_U2648) );
  NOR2_X1 U19985 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16943), .ZN(n16683) );
  AOI22_X1 U19986 ( .A1(n16955), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n16684), 
        .B2(n16683), .ZN(n16692) );
  AOI21_X1 U19987 ( .B1(n16935), .B2(n16703), .A(n16950), .ZN(n16714) );
  OAI21_X1 U19988 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16943), .A(n16714), 
        .ZN(n16690) );
  AOI211_X1 U19989 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16700), .A(n16685), .B(
        n16947), .ZN(n16689) );
  AOI211_X1 U19990 ( .C1(n17638), .C2(n16687), .A(n16686), .B(n18800), .ZN(
        n16688) );
  AOI211_X1 U19991 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16690), .A(n16689), 
        .B(n16688), .ZN(n16691) );
  OAI211_X1 U19992 ( .C1(n16693), .C2(n16938), .A(n16692), .B(n16691), .ZN(
        P3_U2649) );
  NAND2_X1 U19993 ( .A1(n16935), .A2(n18862), .ZN(n16704) );
  INV_X1 U19994 ( .A(n16714), .ZN(n16699) );
  AOI211_X1 U19995 ( .C1(n16696), .C2(n16695), .A(n16694), .B(n18800), .ZN(
        n16698) );
  INV_X1 U19996 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17649) );
  OAI22_X1 U19997 ( .A1(n17649), .A2(n16938), .B1(n16942), .B2(n17051), .ZN(
        n16697) );
  AOI211_X1 U19998 ( .C1(n16699), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16698), 
        .B(n16697), .ZN(n16702) );
  OAI211_X1 U19999 ( .C1(n16705), .C2(n17051), .A(n16954), .B(n16700), .ZN(
        n16701) );
  OAI211_X1 U20000 ( .C1(n16704), .C2(n16703), .A(n16702), .B(n16701), .ZN(
        P3_U2650) );
  INV_X1 U20001 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18859) );
  AOI22_X1 U20002 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16939), .B1(
        n16955), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16713) );
  NOR2_X1 U20003 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16943), .ZN(n16710) );
  AOI211_X1 U20004 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16719), .A(n16705), .B(
        n16947), .ZN(n16709) );
  AOI211_X1 U20005 ( .C1(n17666), .C2(n16707), .A(n16706), .B(n18800), .ZN(
        n16708) );
  AOI211_X1 U20006 ( .C1(n16711), .C2(n16710), .A(n16709), .B(n16708), .ZN(
        n16712) );
  OAI211_X1 U20007 ( .C1(n18859), .C2(n16714), .A(n16713), .B(n16712), .ZN(
        P3_U2651) );
  INV_X1 U20008 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17692) );
  NOR2_X1 U20009 ( .A1(n17692), .A2(n16729), .ZN(n16716) );
  OAI21_X1 U20010 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16716), .A(
        n16715), .ZN(n17676) );
  NAND2_X1 U20011 ( .A1(n17672), .A2(n16752), .ZN(n16730) );
  OAI21_X1 U20012 ( .B1(n17692), .B2(n16730), .A(n16913), .ZN(n16717) );
  XNOR2_X1 U20013 ( .A(n17676), .B(n16717), .ZN(n16728) );
  OAI211_X1 U20014 ( .C1(n16733), .C2(n16721), .A(n16954), .B(n16719), .ZN(
        n16720) );
  OAI211_X1 U20015 ( .C1(n16942), .C2(n16721), .A(n16718), .B(n16720), .ZN(
        n16726) );
  INV_X1 U20016 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18851) );
  NOR2_X1 U20017 ( .A1(n16943), .A2(n16722), .ZN(n16765) );
  NAND2_X1 U20018 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16765), .ZN(n16762) );
  NOR2_X1 U20019 ( .A1(n18851), .A2(n16762), .ZN(n16740) );
  NAND2_X1 U20020 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16740), .ZN(n16739) );
  XOR2_X1 U20021 ( .A(P3_REIP_REG_19__SCAN_IN), .B(n18855), .Z(n16724) );
  NOR2_X1 U20022 ( .A1(n16950), .A2(n16722), .ZN(n16778) );
  NOR2_X1 U20023 ( .A1(n16902), .A2(n16778), .ZN(n16781) );
  AOI21_X1 U20024 ( .B1(n16723), .B2(n16956), .A(n16781), .ZN(n16744) );
  OAI22_X1 U20025 ( .A1(n16739), .A2(n16724), .B1(n18857), .B2(n16744), .ZN(
        n16725) );
  AOI211_X1 U20026 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n16939), .A(
        n16726), .B(n16725), .ZN(n16727) );
  OAI21_X1 U20027 ( .B1(n18800), .B2(n16728), .A(n16727), .ZN(P3_U2652) );
  AOI22_X1 U20028 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16729), .B1(
        n17672), .B2(n17692), .ZN(n17689) );
  NAND2_X1 U20029 ( .A1(n16913), .A2(n16730), .ZN(n16732) );
  OAI21_X1 U20030 ( .B1(n17689), .B2(n16732), .A(n16941), .ZN(n16731) );
  AOI21_X1 U20031 ( .B1(n17689), .B2(n16732), .A(n16731), .ZN(n16737) );
  AOI211_X1 U20032 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16746), .A(n16733), .B(
        n16947), .ZN(n16736) );
  AOI22_X1 U20033 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16939), .B1(
        n16955), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16734) );
  INV_X1 U20034 ( .A(n16734), .ZN(n16735) );
  NOR4_X1 U20035 ( .A1(n18140), .A2(n16737), .A3(n16736), .A4(n16735), .ZN(
        n16738) );
  OAI221_X1 U20036 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16739), .C1(n18855), 
        .C2(n16744), .A(n16738), .ZN(P3_U2653) );
  INV_X1 U20037 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16749) );
  NOR2_X1 U20038 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16740), .ZN(n16743) );
  NAND2_X1 U20039 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17705), .ZN(
        n16750) );
  AOI21_X1 U20040 ( .B1(n16749), .B2(n16750), .A(n17672), .ZN(n17700) );
  AOI21_X1 U20041 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16752), .A(
        n16884), .ZN(n16741) );
  XNOR2_X1 U20042 ( .A(n17700), .B(n16741), .ZN(n16742) );
  OAI22_X1 U20043 ( .A1(n16744), .A2(n16743), .B1(n18800), .B2(n16742), .ZN(
        n16745) );
  AOI211_X1 U20044 ( .C1(n16955), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18235), .B(
        n16745), .ZN(n16748) );
  OAI211_X1 U20045 ( .C1(n16755), .C2(n17094), .A(n16954), .B(n16746), .ZN(
        n16747) );
  OAI211_X1 U20046 ( .C1(n16938), .C2(n16749), .A(n16748), .B(n16747), .ZN(
        P3_U2654) );
  INV_X1 U20047 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18849) );
  AOI21_X1 U20048 ( .B1(n16765), .B2(n18849), .A(n16781), .ZN(n16761) );
  INV_X1 U20049 ( .A(n16764), .ZN(n16751) );
  OAI21_X1 U20050 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16751), .A(
        n16750), .ZN(n17716) );
  INV_X1 U20051 ( .A(n17716), .ZN(n16754) );
  NOR2_X1 U20052 ( .A1(n16752), .A2(n16884), .ZN(n16753) );
  INV_X1 U20053 ( .A(n16753), .ZN(n16763) );
  AOI221_X1 U20054 ( .B1(n16754), .B2(n16753), .C1(n17716), .C2(n16763), .A(
        n18800), .ZN(n16759) );
  AOI211_X1 U20055 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16767), .A(n16755), .B(
        n16947), .ZN(n16758) );
  AOI22_X1 U20056 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16939), .B1(
        n16955), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16756) );
  INV_X1 U20057 ( .A(n16756), .ZN(n16757) );
  NOR4_X1 U20058 ( .A1(n18235), .A2(n16759), .A3(n16758), .A4(n16757), .ZN(
        n16760) );
  OAI221_X1 U20059 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16762), .C1(n18851), 
        .C2(n16761), .A(n16760), .ZN(P3_U2655) );
  INV_X1 U20060 ( .A(n16781), .ZN(n16774) );
  NOR2_X1 U20061 ( .A1(n18800), .A2(n16763), .ZN(n16766) );
  OAI21_X1 U20062 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17711), .A(
        n16764), .ZN(n17722) );
  AOI22_X1 U20063 ( .A1(n16766), .A2(n17722), .B1(n16765), .B2(n18849), .ZN(
        n16773) );
  INV_X1 U20064 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16886) );
  NOR2_X1 U20065 ( .A1(n16884), .A2(n16886), .ZN(n16940) );
  OR2_X1 U20066 ( .A1(n18800), .A2(n16940), .ZN(n16953) );
  AOI211_X1 U20067 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16913), .A(
        n17722), .B(n16953), .ZN(n16771) );
  OAI211_X1 U20068 ( .C1(n16776), .C2(n16769), .A(n16954), .B(n16767), .ZN(
        n16768) );
  OAI211_X1 U20069 ( .C1(n16942), .C2(n16769), .A(n16718), .B(n16768), .ZN(
        n16770) );
  AOI211_X1 U20070 ( .C1(n16939), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16771), .B(n16770), .ZN(n16772) );
  OAI211_X1 U20071 ( .C1(n18849), .C2(n16774), .A(n16773), .B(n16772), .ZN(
        P3_U2656) );
  INV_X1 U20072 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16775) );
  NAND2_X1 U20073 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17731), .ZN(
        n16787) );
  AOI21_X1 U20074 ( .B1(n16775), .B2(n16787), .A(n17711), .ZN(n17732) );
  NOR2_X1 U20075 ( .A1(n17910), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16928) );
  AND2_X1 U20076 ( .A1(n17817), .A2(n16928), .ZN(n16873) );
  AOI21_X1 U20077 ( .B1(n16786), .B2(n16873), .A(n16884), .ZN(n16804) );
  AOI21_X1 U20078 ( .B1(n16913), .B2(n17748), .A(n16804), .ZN(n16785) );
  XOR2_X1 U20079 ( .A(n17732), .B(n16785), .Z(n16784) );
  AOI22_X1 U20080 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16939), .B1(
        n16955), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16783) );
  AOI211_X1 U20081 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16794), .A(n16776), .B(
        n16947), .ZN(n16780) );
  NAND3_X1 U20082 ( .A1(n16935), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n16790), 
        .ZN(n16777) );
  OAI21_X1 U20083 ( .B1(n16778), .B2(n16777), .A(n16718), .ZN(n16779) );
  AOI211_X1 U20084 ( .C1(n16781), .C2(P3_REIP_REG_14__SCAN_IN), .A(n16780), 
        .B(n16779), .ZN(n16782) );
  OAI211_X1 U20085 ( .C1(n18800), .C2(n16784), .A(n16783), .B(n16782), .ZN(
        P3_U2657) );
  NOR2_X1 U20086 ( .A1(n16785), .A2(n18800), .ZN(n16788) );
  INV_X1 U20087 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17764) );
  NOR2_X1 U20088 ( .A1(n17910), .A2(n17777), .ZN(n16883) );
  NAND2_X1 U20089 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16883), .ZN(
        n16860) );
  INV_X1 U20090 ( .A(n16860), .ZN(n16870) );
  NAND2_X1 U20091 ( .A1(n16786), .A2(n16870), .ZN(n17743) );
  NOR2_X1 U20092 ( .A1(n17764), .A2(n17743), .ZN(n16789) );
  OAI21_X1 U20093 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16789), .A(
        n16787), .ZN(n17751) );
  AOI22_X1 U20094 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16939), .B1(
        n16788), .B2(n17751), .ZN(n16799) );
  INV_X1 U20095 ( .A(n16789), .ZN(n16805) );
  AOI211_X1 U20096 ( .C1(n16913), .C2(n16805), .A(n17751), .B(n16953), .ZN(
        n16793) );
  NAND2_X1 U20097 ( .A1(n16935), .A2(n16790), .ZN(n16791) );
  OAI22_X1 U20098 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16791), .B1(n16942), 
        .B2(n16795), .ZN(n16792) );
  NOR3_X1 U20099 ( .A1(n18235), .A2(n16793), .A3(n16792), .ZN(n16798) );
  OAI21_X1 U20100 ( .B1(n16803), .B2(n16943), .A(n16957), .ZN(n16821) );
  NOR2_X1 U20101 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16943), .ZN(n16802) );
  OAI21_X1 U20102 ( .B1(n16821), .B2(n16802), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16797) );
  OAI211_X1 U20103 ( .C1(n16800), .C2(n16795), .A(n16954), .B(n16794), .ZN(
        n16796) );
  NAND4_X1 U20104 ( .A1(n16799), .A2(n16798), .A3(n16797), .A4(n16796), .ZN(
        P3_U2658) );
  AOI22_X1 U20105 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16939), .B1(
        n16955), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16810) );
  AOI211_X1 U20106 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16815), .A(n16800), .B(
        n16947), .ZN(n16801) );
  AOI211_X1 U20107 ( .C1(n16803), .C2(n16802), .A(n18235), .B(n16801), .ZN(
        n16809) );
  INV_X1 U20108 ( .A(n16804), .ZN(n16814) );
  INV_X1 U20109 ( .A(n17743), .ZN(n16806) );
  OAI21_X1 U20110 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16806), .A(
        n16805), .ZN(n17768) );
  XOR2_X1 U20111 ( .A(n16814), .B(n17768), .Z(n16807) );
  AOI22_X1 U20112 ( .A1(n16941), .A2(n16807), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16821), .ZN(n16808) );
  NAND3_X1 U20113 ( .A1(n16810), .A2(n16809), .A3(n16808), .ZN(P3_U2659) );
  NAND2_X1 U20114 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16812) );
  NAND2_X1 U20115 ( .A1(n16935), .A2(n16811), .ZN(n16836) );
  OAI21_X1 U20116 ( .B1(n16812), .B2(n16836), .A(n18841), .ZN(n16820) );
  INV_X1 U20117 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17792) );
  NOR2_X1 U20118 ( .A1(n17826), .A2(n16860), .ZN(n16847) );
  NAND2_X1 U20119 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16847), .ZN(
        n16835) );
  NOR2_X1 U20120 ( .A1(n17792), .A2(n16835), .ZN(n16826) );
  OAI21_X1 U20121 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16826), .A(
        n17743), .ZN(n17781) );
  NAND2_X1 U20122 ( .A1(n16941), .A2(n16884), .ZN(n16931) );
  OAI221_X1 U20123 ( .B1(n17781), .B2(n16826), .C1(n17781), .C2(n16886), .A(
        n16941), .ZN(n16813) );
  AOI22_X1 U20124 ( .A1(n17781), .A2(n16814), .B1(n16931), .B2(n16813), .ZN(
        n16819) );
  INV_X1 U20125 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16817) );
  OAI211_X1 U20126 ( .C1(n16829), .C2(n16823), .A(n16954), .B(n16815), .ZN(
        n16816) );
  OAI21_X1 U20127 ( .B1(n16938), .B2(n16817), .A(n16816), .ZN(n16818) );
  AOI211_X1 U20128 ( .C1(n16821), .C2(n16820), .A(n16819), .B(n16818), .ZN(
        n16822) );
  OAI211_X1 U20129 ( .C1(n16942), .C2(n16823), .A(n16822), .B(n16718), .ZN(
        P3_U2660) );
  AOI21_X1 U20130 ( .B1(n16935), .B2(n16824), .A(n16950), .ZN(n16854) );
  AOI221_X1 U20131 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .C1(n18839), .C2(n18837), .A(n16836), .ZN(n16825) );
  AOI211_X1 U20132 ( .C1(n16955), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18235), .B(
        n16825), .ZN(n16834) );
  AOI21_X1 U20133 ( .B1(n17792), .B2(n16835), .A(n16826), .ZN(n17795) );
  OAI21_X1 U20134 ( .B1(n16835), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16913), .ZN(n16827) );
  INV_X1 U20135 ( .A(n16827), .ZN(n16837) );
  OAI21_X1 U20136 ( .B1(n17795), .B2(n16837), .A(n16941), .ZN(n16828) );
  AOI21_X1 U20137 ( .B1(n17795), .B2(n16837), .A(n16828), .ZN(n16832) );
  AOI211_X1 U20138 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16830), .A(n16829), .B(
        n16947), .ZN(n16831) );
  AOI211_X1 U20139 ( .C1(n16939), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16832), .B(n16831), .ZN(n16833) );
  OAI211_X1 U20140 ( .C1(n18839), .C2(n16854), .A(n16834), .B(n16833), .ZN(
        P3_U2661) );
  AOI21_X1 U20141 ( .B1(n16954), .B2(n16839), .A(n16955), .ZN(n16845) );
  OAI21_X1 U20142 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16847), .A(
        n16835), .ZN(n17807) );
  OAI22_X1 U20143 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16836), .B1(n16931), 
        .B2(n17807), .ZN(n16843) );
  OAI221_X1 U20144 ( .B1(n17807), .B2(n17778), .C1(n17807), .C2(n16873), .A(
        n16837), .ZN(n16838) );
  OAI22_X1 U20145 ( .A1(n18800), .A2(n16838), .B1(n18837), .B2(n16854), .ZN(
        n16842) );
  OR2_X1 U20146 ( .A1(n16947), .A2(n16839), .ZN(n16851) );
  INV_X1 U20147 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16840) );
  OAI22_X1 U20148 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16851), .B1(n16840), .B2(
        n16938), .ZN(n16841) );
  NOR4_X1 U20149 ( .A1(n18140), .A2(n16843), .A3(n16842), .A4(n16841), .ZN(
        n16844) );
  OAI21_X1 U20150 ( .B1(n16846), .B2(n16845), .A(n16844), .ZN(P3_U2662) );
  NAND2_X1 U20151 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16870), .ZN(
        n16848) );
  AOI21_X1 U20152 ( .B1(n16849), .B2(n16848), .A(n16847), .ZN(n17818) );
  AND2_X1 U20153 ( .A1(n17817), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17827) );
  AOI21_X1 U20154 ( .B1(n17827), .B2(n16928), .A(n16884), .ZN(n16850) );
  XNOR2_X1 U20155 ( .A(n17818), .B(n16850), .ZN(n16859) );
  AOI21_X1 U20156 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16862), .A(n16851), .ZN(
        n16852) );
  AOI21_X1 U20157 ( .B1(n16939), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16852), .ZN(n16858) );
  INV_X1 U20158 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18826) );
  NAND3_X1 U20159 ( .A1(n16935), .A2(P3_REIP_REG_1__SCAN_IN), .A3(
        P3_REIP_REG_2__SCAN_IN), .ZN(n16910) );
  NOR2_X1 U20160 ( .A1(n18826), .A2(n16910), .ZN(n16907) );
  NOR2_X1 U20161 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16853), .ZN(n16856) );
  OAI22_X1 U20162 ( .A1(n16942), .A2(n17249), .B1(n18836), .B2(n16854), .ZN(
        n16855) );
  AOI211_X1 U20163 ( .C1(n16907), .C2(n16856), .A(n18235), .B(n16855), .ZN(
        n16857) );
  OAI211_X1 U20164 ( .C1(n18800), .C2(n16859), .A(n16858), .B(n16857), .ZN(
        P3_U2663) );
  AOI22_X1 U20165 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16870), .B1(
        n16860), .B2(n17834), .ZN(n17839) );
  NOR2_X1 U20166 ( .A1(n16873), .A2(n16884), .ZN(n16861) );
  XNOR2_X1 U20167 ( .A(n17839), .B(n16861), .ZN(n16869) );
  OAI211_X1 U20168 ( .C1(n16872), .C2(n16863), .A(n16954), .B(n16862), .ZN(
        n16864) );
  OAI211_X1 U20169 ( .C1(n17834), .C2(n16938), .A(n16718), .B(n16864), .ZN(
        n16865) );
  AOI21_X1 U20170 ( .B1(n16955), .B2(P3_EBX_REG_7__SCAN_IN), .A(n16865), .ZN(
        n16868) );
  INV_X1 U20171 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18830) );
  NAND2_X1 U20172 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16907), .ZN(n16888) );
  NOR2_X1 U20173 ( .A1(n18830), .A2(n16888), .ZN(n16879) );
  NAND2_X1 U20174 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n16866) );
  NOR3_X1 U20175 ( .A1(n16950), .A2(n16866), .A3(n16900), .ZN(n16887) );
  AOI21_X1 U20176 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16887), .A(n16902), .ZN(
        n16878) );
  INV_X1 U20177 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18834) );
  OAI222_X1 U20178 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16879), .C1(n16878), .C2(n18834), 
        .ZN(n16867) );
  OAI211_X1 U20179 ( .C1(n18800), .C2(n16869), .A(n16868), .B(n16867), .ZN(
        P3_U2664) );
  AOI22_X1 U20180 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16939), .B1(
        n16955), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n16882) );
  INV_X1 U20181 ( .A(n16883), .ZN(n16871) );
  AOI21_X1 U20182 ( .B1(n17847), .B2(n16871), .A(n16870), .ZN(n16874) );
  INV_X1 U20183 ( .A(n16874), .ZN(n17853) );
  AOI211_X1 U20184 ( .C1(n16913), .C2(n16871), .A(n17853), .B(n16953), .ZN(
        n16877) );
  AOI211_X1 U20185 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16889), .A(n16872), .B(
        n16947), .ZN(n16876) );
  NOR4_X1 U20186 ( .A1(n16874), .A2(n16873), .A3(n18800), .A4(n16884), .ZN(
        n16875) );
  NOR4_X1 U20187 ( .A1(n18235), .A2(n16877), .A3(n16876), .A4(n16875), .ZN(
        n16881) );
  OAI21_X1 U20188 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16879), .A(n16878), .ZN(
        n16880) );
  NAND3_X1 U20189 ( .A1(n16882), .A2(n16881), .A3(n16880), .ZN(P3_U2665) );
  INV_X1 U20190 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16891) );
  NAND2_X1 U20191 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17862), .ZN(
        n16903) );
  AOI21_X1 U20192 ( .B1(n16891), .B2(n16903), .A(n16883), .ZN(n17864) );
  INV_X1 U20193 ( .A(n16903), .ZN(n16885) );
  AOI21_X1 U20194 ( .B1(n16886), .B2(n16885), .A(n16884), .ZN(n16904) );
  XOR2_X1 U20195 ( .A(n17864), .B(n16904), .Z(n16894) );
  AOI211_X1 U20196 ( .C1(n18830), .C2(n16888), .A(n16887), .B(n16902), .ZN(
        n16893) );
  OAI211_X1 U20197 ( .C1(n16896), .C2(n17257), .A(n16954), .B(n16889), .ZN(
        n16890) );
  OAI21_X1 U20198 ( .B1(n16938), .B2(n16891), .A(n16890), .ZN(n16892) );
  AOI211_X1 U20199 ( .C1(n16941), .C2(n16894), .A(n16893), .B(n16892), .ZN(
        n16895) );
  OAI211_X1 U20200 ( .C1(n16942), .C2(n17257), .A(n16895), .B(n16718), .ZN(
        P3_U2666) );
  AOI211_X1 U20201 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16920), .A(n16896), .B(
        n16947), .ZN(n16899) );
  NAND2_X1 U20202 ( .A1(n18268), .A2(n18951), .ZN(n16946) );
  OAI221_X1 U20203 ( .B1(n16946), .B2(n11076), .C1(n16946), .C2(n16897), .A(
        n16718), .ZN(n16898) );
  AOI211_X1 U20204 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16955), .A(n16899), .B(
        n16898), .ZN(n16909) );
  NOR2_X1 U20205 ( .A1(n16950), .A2(n16900), .ZN(n16901) );
  NOR2_X1 U20206 ( .A1(n16902), .A2(n16901), .ZN(n16919) );
  INV_X1 U20207 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18827) );
  NOR2_X1 U20208 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17892), .ZN(
        n17873) );
  NOR2_X1 U20209 ( .A1(n17910), .A2(n17892), .ZN(n16911) );
  OAI21_X1 U20210 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16911), .A(
        n16903), .ZN(n17878) );
  AOI22_X1 U20211 ( .A1(n16928), .A2(n17873), .B1(n16904), .B2(n17878), .ZN(
        n16905) );
  AOI221_X1 U20212 ( .B1(n16913), .B2(n16905), .C1(n17878), .C2(n16905), .A(
        n18800), .ZN(n16906) );
  AOI221_X1 U20213 ( .B1(n16919), .B2(P3_REIP_REG_4__SCAN_IN), .C1(n16907), 
        .C2(n18827), .A(n16906), .ZN(n16908) );
  OAI211_X1 U20214 ( .C1(n17877), .C2(n16938), .A(n16909), .B(n16908), .ZN(
        P3_U2667) );
  INV_X1 U20215 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17888) );
  NAND2_X1 U20216 ( .A1(n18826), .A2(n16910), .ZN(n16918) );
  NAND2_X1 U20217 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16925) );
  AOI21_X1 U20218 ( .B1(n17888), .B2(n16925), .A(n16911), .ZN(n16912) );
  INV_X1 U20219 ( .A(n16912), .ZN(n17890) );
  OAI21_X1 U20220 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16925), .A(
        n16913), .ZN(n16926) );
  OAI21_X1 U20221 ( .B1(n17890), .B2(n16926), .A(n16941), .ZN(n16914) );
  AOI21_X1 U20222 ( .B1(n17890), .B2(n16926), .A(n16914), .ZN(n16917) );
  NOR2_X1 U20223 ( .A1(n18910), .A2(n9798), .ZN(n18748) );
  INV_X1 U20224 ( .A(n18748), .ZN(n18740) );
  NOR2_X1 U20225 ( .A1(n18916), .A2(n18740), .ZN(n18738) );
  OAI21_X1 U20226 ( .B1(n18897), .B2(n18738), .A(n17186), .ZN(n18895) );
  AOI22_X1 U20227 ( .A1(n18895), .A2(n18953), .B1(n16955), .B2(
        P3_EBX_REG_3__SCAN_IN), .ZN(n16915) );
  INV_X1 U20228 ( .A(n16915), .ZN(n16916) );
  AOI211_X1 U20229 ( .C1(n16919), .C2(n16918), .A(n16917), .B(n16916), .ZN(
        n16922) );
  OAI211_X1 U20230 ( .C1(n16923), .C2(n17263), .A(n16954), .B(n16920), .ZN(
        n16921) );
  OAI211_X1 U20231 ( .C1(n16938), .C2(n17888), .A(n16922), .B(n16921), .ZN(
        P3_U2668) );
  INV_X1 U20232 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21003) );
  NAND2_X1 U20233 ( .A1(n17283), .A2(n17277), .ZN(n16924) );
  AOI211_X1 U20234 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16924), .A(n16923), .B(
        n16947), .ZN(n16933) );
  OAI21_X1 U20235 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16925), .ZN(n17900) );
  NOR2_X1 U20236 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18744), .ZN(
        n18741) );
  NOR2_X1 U20237 ( .A1(n18738), .A2(n18741), .ZN(n18901) );
  AOI22_X1 U20238 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16950), .B1(n18901), 
        .B2(n18953), .ZN(n16930) );
  INV_X1 U20239 ( .A(n16926), .ZN(n16927) );
  OAI211_X1 U20240 ( .C1(n16928), .C2(n17900), .A(n16941), .B(n16927), .ZN(
        n16929) );
  OAI211_X1 U20241 ( .C1(n16931), .C2(n17900), .A(n16930), .B(n16929), .ZN(
        n16932) );
  AOI211_X1 U20242 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16955), .A(n16933), .B(
        n16932), .ZN(n16937) );
  NAND2_X1 U20243 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16934) );
  OAI211_X1 U20244 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16935), .B(n16934), .ZN(n16936) );
  OAI211_X1 U20245 ( .C1(n16938), .C2(n21003), .A(n16937), .B(n16936), .ZN(
        P3_U2669) );
  AOI21_X1 U20246 ( .B1(n16941), .B2(n16940), .A(n16939), .ZN(n16952) );
  OAI22_X1 U20247 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16943), .B1(n16942), 
        .B2(n17277), .ZN(n16949) );
  AOI21_X1 U20248 ( .B1(n17283), .B2(n17277), .A(n17271), .ZN(n16944) );
  INV_X1 U20249 ( .A(n16944), .ZN(n17279) );
  NOR2_X1 U20250 ( .A1(n16945), .A2(n18744), .ZN(n18907) );
  INV_X1 U20251 ( .A(n18907), .ZN(n18763) );
  OAI22_X1 U20252 ( .A1(n16947), .A2(n17279), .B1(n18763), .B2(n16946), .ZN(
        n16948) );
  AOI211_X1 U20253 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n16950), .A(n16949), .B(
        n16948), .ZN(n16951) );
  OAI221_X1 U20254 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16953), .C1(
        n17910), .C2(n16952), .A(n16951), .ZN(P3_U2670) );
  NOR2_X1 U20255 ( .A1(n16955), .A2(n16954), .ZN(n16960) );
  AOI22_X1 U20256 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16956), .B1(n18953), 
        .B2(n18916), .ZN(n16959) );
  NAND3_X1 U20257 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18892), .A3(
        n16957), .ZN(n16958) );
  OAI211_X1 U20258 ( .C1(n16960), .C2(n17283), .A(n16959), .B(n16958), .ZN(
        P3_U2671) );
  INV_X1 U20259 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16962) );
  NAND4_X1 U20260 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_20__SCAN_IN), .A4(n17083), .ZN(n16961) );
  NOR4_X1 U20261 ( .A1(n16995), .A2(n16962), .A3(n17051), .A4(n16961), .ZN(
        n16963) );
  NAND4_X1 U20262 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n16996), .A4(n16963), .ZN(n16966) );
  NAND2_X1 U20263 ( .A1(n17275), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16965) );
  NAND2_X1 U20264 ( .A1(n16994), .A2(n18297), .ZN(n16964) );
  OAI22_X1 U20265 ( .A1(n16994), .A2(n16965), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16964), .ZN(P3_U2672) );
  NAND2_X1 U20266 ( .A1(n16967), .A2(n16966), .ZN(n16968) );
  NAND2_X1 U20267 ( .A1(n16968), .A2(n17275), .ZN(n16993) );
  AOI22_X1 U20268 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16978) );
  AOI22_X1 U20269 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20270 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16976) );
  OAI22_X1 U20271 ( .A1(n11056), .A2(n17150), .B1(n11037), .B2(n18506), .ZN(
        n16974) );
  AOI22_X1 U20272 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20273 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20274 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16970) );
  NAND2_X1 U20275 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n16969) );
  NAND4_X1 U20276 ( .A1(n16972), .A2(n16971), .A3(n16970), .A4(n16969), .ZN(
        n16973) );
  AOI211_X1 U20277 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n16974), .B(n16973), .ZN(n16975) );
  NAND4_X1 U20278 ( .A1(n16978), .A2(n16977), .A3(n16976), .A4(n16975), .ZN(
        n16998) );
  NAND3_X1 U20279 ( .A1(n16997), .A2(n17003), .A3(n16998), .ZN(n16992) );
  AOI22_X1 U20280 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n11051), .ZN(n16979) );
  OAI21_X1 U20281 ( .B1(n17177), .B2(n17126), .A(n16979), .ZN(n16990) );
  AOI22_X1 U20282 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11065), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17195), .ZN(n16987) );
  AOI22_X1 U20283 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n9801), .ZN(n16980) );
  OAI21_X1 U20284 ( .B1(n16981), .B2(n11054), .A(n16980), .ZN(n16985) );
  AOI22_X1 U20285 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17105), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20286 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16982) );
  OAI211_X1 U20287 ( .C1(n18618), .C2(n17246), .A(n16983), .B(n16982), .ZN(
        n16984) );
  AOI211_X1 U20288 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n16985), .B(n16984), .ZN(n16986) );
  OAI211_X1 U20289 ( .C1(n16988), .C2(n11055), .A(n16987), .B(n16986), .ZN(
        n16989) );
  AOI211_X1 U20290 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16990), .B(n16989), .ZN(n16991) );
  XNOR2_X1 U20291 ( .A(n16992), .B(n16991), .ZN(n17289) );
  OAI22_X1 U20292 ( .A1(n16994), .A2(n16993), .B1(n17289), .B2(n17275), .ZN(
        P3_U2673) );
  NAND2_X1 U20293 ( .A1(n16996), .A2(n16995), .ZN(n17002) );
  NAND2_X1 U20294 ( .A1(n16997), .A2(n17003), .ZN(n16999) );
  XNOR2_X1 U20295 ( .A(n16999), .B(n16998), .ZN(n17293) );
  AOI22_X1 U20296 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17000), .B1(n17281), 
        .B2(n17293), .ZN(n17001) );
  OAI21_X1 U20297 ( .B1(n17008), .B2(n17002), .A(n17001), .ZN(P3_U2674) );
  AOI21_X1 U20298 ( .B1(n17004), .B2(n17009), .A(n17003), .ZN(n17303) );
  NAND2_X1 U20299 ( .A1(n17281), .A2(n17303), .ZN(n17005) );
  OAI221_X1 U20300 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17008), .C1(n17007), 
        .C2(n17006), .A(n17005), .ZN(P3_U2676) );
  AOI21_X1 U20301 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17275), .A(n17017), .ZN(
        n17012) );
  OAI21_X1 U20302 ( .B1(n17011), .B2(n17010), .A(n17009), .ZN(n17311) );
  OAI22_X1 U20303 ( .A1(n17013), .A2(n17012), .B1(n17275), .B2(n17311), .ZN(
        P3_U2677) );
  INV_X1 U20304 ( .A(n17014), .ZN(n17022) );
  AOI21_X1 U20305 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17275), .A(n17022), .ZN(
        n17016) );
  XNOR2_X1 U20306 ( .A(n17015), .B(n17018), .ZN(n17316) );
  OAI22_X1 U20307 ( .A1(n17017), .A2(n17016), .B1(n17275), .B2(n17316), .ZN(
        P3_U2678) );
  AOI21_X1 U20308 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17275), .A(n17027), .ZN(
        n17021) );
  OAI21_X1 U20309 ( .B1(n17020), .B2(n17019), .A(n17018), .ZN(n17322) );
  OAI22_X1 U20310 ( .A1(n17022), .A2(n17021), .B1(n17275), .B2(n17322), .ZN(
        P3_U2679) );
  INV_X1 U20311 ( .A(n17023), .ZN(n17039) );
  AOI21_X1 U20312 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17275), .A(n17039), .ZN(
        n17026) );
  XNOR2_X1 U20313 ( .A(n17025), .B(n17024), .ZN(n17328) );
  OAI22_X1 U20314 ( .A1(n17027), .A2(n17026), .B1(n17275), .B2(n17328), .ZN(
        P3_U2680) );
  AOI22_X1 U20315 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17275), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n17052), .ZN(n17038) );
  AOI22_X1 U20316 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17028) );
  OAI21_X1 U20317 ( .B1(n11076), .B2(n17150), .A(n17028), .ZN(n17037) );
  INV_X1 U20318 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20319 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17035) );
  INV_X1 U20320 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20321 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11065), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17029) );
  OAI21_X1 U20322 ( .B1(n17163), .B2(n17141), .A(n17029), .ZN(n17033) );
  AOI22_X1 U20323 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20324 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17030) );
  OAI211_X1 U20325 ( .C1(n11056), .C2(n17143), .A(n17031), .B(n17030), .ZN(
        n17032) );
  AOI211_X1 U20326 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17033), .B(n17032), .ZN(n17034) );
  OAI211_X1 U20327 ( .C1(n11054), .C2(n17254), .A(n17035), .B(n17034), .ZN(
        n17036) );
  AOI211_X1 U20328 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17037), .B(n17036), .ZN(n17330) );
  OAI22_X1 U20329 ( .A1(n17039), .A2(n17038), .B1(n17330), .B2(n17275), .ZN(
        P3_U2681) );
  AOI22_X1 U20330 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17040) );
  OAI21_X1 U20331 ( .B1(n17072), .B2(n17041), .A(n17040), .ZN(n17050) );
  AOI22_X1 U20332 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20333 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17042) );
  OAI21_X1 U20334 ( .B1(n11076), .B2(n21130), .A(n17042), .ZN(n17046) );
  AOI22_X1 U20335 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20336 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17043) );
  OAI211_X1 U20337 ( .C1(n17246), .C2(n21086), .A(n17044), .B(n17043), .ZN(
        n17045) );
  AOI211_X1 U20338 ( .C1(n17216), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n17046), .B(n17045), .ZN(n17047) );
  OAI211_X1 U20339 ( .C1(n11054), .C2(n17261), .A(n17048), .B(n17047), .ZN(
        n17049) );
  AOI211_X1 U20340 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n17050), .B(n17049), .ZN(n17341) );
  AOI21_X1 U20341 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17083), .A(n17281), .ZN(
        n17065) );
  AOI22_X1 U20342 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17065), .B1(n17052), 
        .B2(n17051), .ZN(n17053) );
  OAI21_X1 U20343 ( .B1(n17341), .B2(n17275), .A(n17053), .ZN(P3_U2682) );
  INV_X1 U20344 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20345 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17054) );
  OAI21_X1 U20346 ( .B1(n11055), .B2(n17055), .A(n17054), .ZN(n17064) );
  INV_X1 U20347 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18606) );
  AOI22_X1 U20348 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11065), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17062) );
  OAI22_X1 U20349 ( .A1(n11054), .A2(n17264), .B1(n9841), .B2(n17170), .ZN(
        n17060) );
  AOI22_X1 U20350 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20351 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20352 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17056) );
  NAND3_X1 U20353 ( .A1(n17058), .A2(n17057), .A3(n17056), .ZN(n17059) );
  AOI211_X1 U20354 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17060), .B(n17059), .ZN(n17061) );
  OAI211_X1 U20355 ( .C1(n10227), .C2(n18606), .A(n17062), .B(n17061), .ZN(
        n17063) );
  AOI211_X1 U20356 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17064), .B(n17063), .ZN(n17343) );
  OAI21_X1 U20357 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17066), .A(n17065), .ZN(
        n17067) );
  OAI21_X1 U20358 ( .B1(n17343), .B2(n17275), .A(n17067), .ZN(P3_U2683) );
  INV_X1 U20359 ( .A(n17068), .ZN(n17095) );
  OAI21_X1 U20360 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17095), .A(n17275), .ZN(
        n17082) );
  AOI22_X1 U20361 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17069) );
  OAI21_X1 U20362 ( .B1(n11076), .B2(n17070), .A(n17069), .ZN(n17081) );
  AOI22_X1 U20363 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17079) );
  OAI22_X1 U20364 ( .A1(n11054), .A2(n17268), .B1(n17072), .B2(n17071), .ZN(
        n17077) );
  AOI22_X1 U20365 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U20366 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20367 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17073) );
  NAND3_X1 U20368 ( .A1(n17075), .A2(n17074), .A3(n17073), .ZN(n17076) );
  AOI211_X1 U20369 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17077), .B(n17076), .ZN(n17078) );
  OAI211_X1 U20370 ( .C1(n11037), .C2(n17176), .A(n17079), .B(n17078), .ZN(
        n17080) );
  AOI211_X1 U20371 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17081), .B(n17080), .ZN(n17350) );
  OAI22_X1 U20372 ( .A1(n17083), .A2(n17082), .B1(n17350), .B2(n17275), .ZN(
        P3_U2684) );
  AOI22_X1 U20373 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17084) );
  OAI21_X1 U20374 ( .B1(n10227), .B2(n18598), .A(n17084), .ZN(n17093) );
  AOI22_X1 U20375 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17235), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17091) );
  OAI22_X1 U20376 ( .A1(n17177), .A2(n18494), .B1(n17163), .B2(n17201), .ZN(
        n17089) );
  AOI22_X1 U20377 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U20378 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20379 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17085) );
  NAND3_X1 U20380 ( .A1(n17087), .A2(n17086), .A3(n17085), .ZN(n17088) );
  AOI211_X1 U20381 ( .C1(n17237), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17089), .B(n17088), .ZN(n17090) );
  OAI211_X1 U20382 ( .C1(n11038), .C2(n17194), .A(n17091), .B(n17090), .ZN(
        n17092) );
  AOI211_X1 U20383 ( .C1(n17236), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n17093), .B(n17092), .ZN(n17355) );
  NAND3_X1 U20384 ( .A1(n18297), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17112), 
        .ZN(n17111) );
  NOR2_X1 U20385 ( .A1(n17094), .A2(n17111), .ZN(n17097) );
  NOR2_X1 U20386 ( .A1(n17281), .A2(n17095), .ZN(n17096) );
  OAI21_X1 U20387 ( .B1(n17097), .B2(P3_EBX_REG_18__SCAN_IN), .A(n17096), .ZN(
        n17098) );
  OAI21_X1 U20388 ( .B1(n17355), .B2(n17275), .A(n17098), .ZN(P3_U2685) );
  INV_X1 U20389 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U20390 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17099) );
  OAI21_X1 U20391 ( .B1(n17186), .B2(n17214), .A(n17099), .ZN(n17109) );
  AOI22_X1 U20392 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17107) );
  INV_X1 U20393 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17276) );
  OAI22_X1 U20394 ( .A1(n11054), .A2(n17276), .B1(n10227), .B2(n21111), .ZN(
        n17104) );
  AOI22_X1 U20395 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20396 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20397 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17100) );
  NAND3_X1 U20398 ( .A1(n17102), .A2(n17101), .A3(n17100), .ZN(n17103) );
  AOI211_X1 U20399 ( .C1(n17105), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n17104), .B(n17103), .ZN(n17106) );
  OAI211_X1 U20400 ( .C1(n17246), .C2(n17212), .A(n17107), .B(n17106), .ZN(
        n17108) );
  AOI211_X1 U20401 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n17109), .B(n17108), .ZN(n17361) );
  NAND3_X1 U20402 ( .A1(n17111), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17275), 
        .ZN(n17110) );
  OAI221_X1 U20403 ( .B1(n17111), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n17275), 
        .C2(n17361), .A(n17110), .ZN(P3_U2686) );
  NAND2_X1 U20404 ( .A1(n18297), .A2(n17112), .ZN(n17124) );
  NOR2_X1 U20405 ( .A1(n17281), .A2(n17112), .ZN(n17137) );
  AOI22_X1 U20406 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20407 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17121) );
  OAI22_X1 U20408 ( .A1(n10244), .A2(n18542), .B1(n11054), .B2(n17234), .ZN(
        n17119) );
  AOI22_X1 U20409 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11065), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20410 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20411 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17113) );
  OAI211_X1 U20412 ( .C1(n17163), .C2(n21045), .A(n17114), .B(n17113), .ZN(
        n17115) );
  AOI21_X1 U20413 ( .B1(n17215), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n17115), .ZN(n17116) );
  OAI211_X1 U20414 ( .C1(n11056), .C2(n18304), .A(n17117), .B(n17116), .ZN(
        n17118) );
  AOI211_X1 U20415 ( .C1(n17236), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n17119), .B(n17118), .ZN(n17120) );
  NAND3_X1 U20416 ( .A1(n17122), .A2(n17121), .A3(n17120), .ZN(n17362) );
  AOI22_X1 U20417 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17137), .B1(n17281), 
        .B2(n17362), .ZN(n17123) );
  OAI21_X1 U20418 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17124), .A(n17123), .ZN(
        P3_U2687) );
  AOI22_X1 U20419 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17125) );
  OAI21_X1 U20420 ( .B1(n10244), .B2(n17126), .A(n17125), .ZN(n17135) );
  AOI22_X1 U20421 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11065), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17105), .ZN(n17133) );
  INV_X1 U20422 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18562) );
  AOI22_X1 U20423 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17210), .ZN(n17127) );
  OAI21_X1 U20424 ( .B1(n18562), .B2(n17246), .A(n17127), .ZN(n17131) );
  AOI22_X1 U20425 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17229), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n9799), .ZN(n17129) );
  AOI22_X1 U20426 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n11051), .ZN(n17128) );
  OAI211_X1 U20427 ( .C1(n11056), .C2(n17252), .A(n17129), .B(n17128), .ZN(
        n17130) );
  AOI211_X1 U20428 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n17131), .B(n17130), .ZN(n17132) );
  OAI211_X1 U20429 ( .C1(n18618), .C2(n11038), .A(n17133), .B(n17132), .ZN(
        n17134) );
  AOI211_X1 U20430 ( .C1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .C2(n9806), .A(
        n17135), .B(n17134), .ZN(n17371) );
  INV_X1 U20431 ( .A(n17136), .ZN(n17138) );
  OAI21_X1 U20432 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17138), .A(n17137), .ZN(
        n17139) );
  OAI21_X1 U20433 ( .B1(n17371), .B2(n17275), .A(n17139), .ZN(P3_U2688) );
  AOI22_X1 U20434 ( .A1(n17236), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17140) );
  OAI21_X1 U20435 ( .B1(n11055), .B2(n17141), .A(n17140), .ZN(n17153) );
  AOI22_X1 U20436 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20437 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11145), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17142) );
  OAI21_X1 U20438 ( .B1(n11076), .B2(n17143), .A(n17142), .ZN(n17147) );
  AOI22_X1 U20439 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U20440 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17144) );
  OAI211_X1 U20441 ( .C1(n11056), .C2(n17254), .A(n17145), .B(n17144), .ZN(
        n17146) );
  AOI211_X1 U20442 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17147), .B(n17146), .ZN(n17148) );
  OAI211_X1 U20443 ( .C1(n17151), .C2(n17150), .A(n17149), .B(n17148), .ZN(
        n17152) );
  AOI211_X1 U20444 ( .C1(n17195), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17153), .B(n17152), .ZN(n17379) );
  OAI21_X1 U20445 ( .B1(n17155), .B2(n17154), .A(P3_EBX_REG_14__SCAN_IN), .ZN(
        n17159) );
  INV_X1 U20446 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17156) );
  NAND3_X1 U20447 ( .A1(n18297), .A2(n17157), .A3(n17156), .ZN(n17158) );
  OAI211_X1 U20448 ( .C1(n17379), .C2(n17275), .A(n17159), .B(n17158), .ZN(
        P3_U2689) );
  AOI22_X1 U20449 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17160) );
  OAI21_X1 U20450 ( .B1(n17186), .B2(n18500), .A(n17160), .ZN(n17172) );
  AOI22_X1 U20451 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17169) );
  INV_X1 U20452 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20453 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17161) );
  OAI21_X1 U20454 ( .B1(n17163), .B2(n17162), .A(n17161), .ZN(n17167) );
  AOI22_X1 U20455 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17210), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20456 ( .A1(n13905), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17164) );
  OAI211_X1 U20457 ( .C1(n11056), .C2(n17264), .A(n17165), .B(n17164), .ZN(
        n17166) );
  AOI211_X1 U20458 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17167), .B(n17166), .ZN(n17168) );
  OAI211_X1 U20459 ( .C1(n11037), .C2(n17170), .A(n17169), .B(n17168), .ZN(
        n17171) );
  AOI211_X1 U20460 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17172), .B(n17171), .ZN(n17385) );
  NOR2_X1 U20461 ( .A1(n17189), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n17174) );
  OAI22_X1 U20462 ( .A1(n17385), .A2(n17275), .B1(n17174), .B2(n17173), .ZN(
        P3_U2691) );
  AOI22_X1 U20463 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17175) );
  OAI21_X1 U20464 ( .B1(n17177), .B2(n17176), .A(n17175), .ZN(n17188) );
  AOI22_X1 U20465 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17185) );
  OAI22_X1 U20466 ( .A1(n9842), .A2(n17178), .B1(n11056), .B2(n17268), .ZN(
        n17183) );
  AOI22_X1 U20467 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20468 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17105), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20469 ( .A1(n11145), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17179) );
  NAND3_X1 U20470 ( .A1(n17181), .A2(n17180), .A3(n17179), .ZN(n17182) );
  AOI211_X1 U20471 ( .C1(n11065), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n17183), .B(n17182), .ZN(n17184) );
  OAI211_X1 U20472 ( .C1(n17186), .C2(n18497), .A(n17185), .B(n17184), .ZN(
        n17187) );
  AOI211_X1 U20473 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n17188), .B(n17187), .ZN(n17389) );
  OAI21_X1 U20474 ( .B1(n17208), .B2(n17227), .A(n17275), .ZN(n17209) );
  NAND2_X1 U20475 ( .A1(n18297), .A2(n17189), .ZN(n17190) );
  OAI21_X1 U20476 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17209), .A(n17190), .ZN(
        n17191) );
  AOI21_X1 U20477 ( .B1(n17281), .B2(n17389), .A(n17191), .ZN(P3_U2692) );
  AOI22_X1 U20478 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U20479 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17205) );
  OAI22_X1 U20480 ( .A1(n9842), .A2(n17194), .B1(n11037), .B2(n17193), .ZN(
        n17203) );
  AOI22_X1 U20481 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U20482 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20483 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9799), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17196) );
  OAI211_X1 U20484 ( .C1(n17246), .C2(n21093), .A(n17197), .B(n17196), .ZN(
        n17198) );
  AOI21_X1 U20485 ( .B1(n17216), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17198), .ZN(n17199) );
  OAI211_X1 U20486 ( .C1(n11055), .C2(n17201), .A(n17200), .B(n17199), .ZN(
        n17202) );
  AOI211_X1 U20487 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17203), .B(n17202), .ZN(n17204) );
  NAND3_X1 U20488 ( .A1(n17206), .A2(n17205), .A3(n17204), .ZN(n17396) );
  NAND2_X1 U20489 ( .A1(n17281), .A2(n17396), .ZN(n17207) );
  OAI221_X1 U20490 ( .B1(n17209), .B2(n17208), .C1(n17209), .C2(n17227), .A(
        n17207), .ZN(P3_U2693) );
  AOI22_X1 U20491 ( .A1(n17210), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17211) );
  OAI21_X1 U20492 ( .B1(n10227), .B2(n17212), .A(n17211), .ZN(n17226) );
  INV_X1 U20493 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20494 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17223) );
  OAI22_X1 U20495 ( .A1(n10244), .A2(n17214), .B1(n11054), .B2(n17213), .ZN(
        n17221) );
  AOI22_X1 U20496 ( .A1(n9806), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11226), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17219) );
  AOI22_X1 U20497 ( .A1(n17192), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20498 ( .A1(n17216), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17215), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17217) );
  NAND3_X1 U20499 ( .A1(n17219), .A2(n17218), .A3(n17217), .ZN(n17220) );
  AOI211_X1 U20500 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n17221), .B(n17220), .ZN(n17222) );
  OAI211_X1 U20501 ( .C1(n11037), .C2(n17224), .A(n17223), .B(n17222), .ZN(
        n17225) );
  AOI211_X1 U20502 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n17226), .B(n17225), .ZN(n17400) );
  OAI21_X1 U20503 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17247), .A(n17227), .ZN(
        n17228) );
  AOI22_X1 U20504 ( .A1(n17281), .A2(n17400), .B1(n17228), .B2(n17275), .ZN(
        P3_U2694) );
  AOI22_X1 U20505 ( .A1(n11065), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13905), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17245) );
  AOI22_X1 U20506 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11051), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20507 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9806), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17232) );
  OAI211_X1 U20508 ( .C1(n11056), .C2(n17234), .A(n17233), .B(n17232), .ZN(
        n17243) );
  AOI22_X1 U20509 ( .A1(n11226), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20510 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9801), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U20511 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17239) );
  NAND2_X1 U20512 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n17238) );
  NAND4_X1 U20513 ( .A1(n17241), .A2(n17240), .A3(n17239), .A4(n17238), .ZN(
        n17242) );
  AOI211_X1 U20514 ( .C1(n11145), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17243), .B(n17242), .ZN(n17244) );
  OAI211_X1 U20515 ( .C1(n17246), .C2(n18542), .A(n17245), .B(n17244), .ZN(
        n17406) );
  AOI21_X1 U20516 ( .B1(n17249), .B2(n17248), .A(n17247), .ZN(n17250) );
  MUX2_X1 U20517 ( .A(n17406), .B(n17250), .S(n17275), .Z(P3_U2695) );
  NAND4_X1 U20518 ( .A1(n18297), .A2(P3_EBX_REG_6__SCAN_IN), .A3(
        P3_EBX_REG_5__SCAN_IN), .A4(n17258), .ZN(n17253) );
  NAND3_X1 U20519 ( .A1(n17253), .A2(P3_EBX_REG_7__SCAN_IN), .A3(n17275), .ZN(
        n17251) );
  OAI221_X1 U20520 ( .B1(n17253), .B2(P3_EBX_REG_7__SCAN_IN), .C1(n17275), 
        .C2(n17252), .A(n17251), .ZN(P3_U2696) );
  INV_X1 U20521 ( .A(n17253), .ZN(n17256) );
  INV_X1 U20522 ( .A(n17258), .ZN(n17259) );
  NOR2_X1 U20523 ( .A1(n17333), .A2(n17259), .ZN(n17266) );
  AOI22_X1 U20524 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17275), .B1(
        P3_EBX_REG_5__SCAN_IN), .B2(n17266), .ZN(n17255) );
  OAI22_X1 U20525 ( .A1(n17256), .A2(n17255), .B1(n17254), .B2(n17275), .ZN(
        P3_U2697) );
  AOI22_X1 U20526 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17259), .B1(n17258), .B2(
        n17257), .ZN(n17260) );
  AOI22_X1 U20527 ( .A1(n17281), .A2(n17261), .B1(n17260), .B2(n17275), .ZN(
        P3_U2698) );
  INV_X1 U20528 ( .A(n17278), .ZN(n17280) );
  NAND2_X1 U20529 ( .A1(n17262), .A2(n17280), .ZN(n17267) );
  NOR2_X1 U20530 ( .A1(n17263), .A2(n17267), .ZN(n17270) );
  AOI21_X1 U20531 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17275), .A(n17270), .ZN(
        n17265) );
  OAI22_X1 U20532 ( .A1(n17266), .A2(n17265), .B1(n17264), .B2(n17275), .ZN(
        P3_U2699) );
  INV_X1 U20533 ( .A(n17267), .ZN(n17272) );
  AOI21_X1 U20534 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17275), .A(n17272), .ZN(
        n17269) );
  OAI22_X1 U20535 ( .A1(n17270), .A2(n17269), .B1(n17268), .B2(n17275), .ZN(
        P3_U2700) );
  INV_X1 U20536 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17274) );
  AOI221_X1 U20537 ( .B1(n17271), .B2(n17284), .C1(n17333), .C2(n17284), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17273) );
  AOI211_X1 U20538 ( .C1(n17281), .C2(n17274), .A(n17273), .B(n17272), .ZN(
        P3_U2701) );
  OAI222_X1 U20539 ( .A1(n17279), .A2(n17278), .B1(n17277), .B2(n17284), .C1(
        n17276), .C2(n17275), .ZN(P3_U2702) );
  AOI22_X1 U20540 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17281), .B1(
        n17280), .B2(n17283), .ZN(n17282) );
  OAI21_X1 U20541 ( .B1(n17284), .B2(n17283), .A(n17282), .ZN(P3_U2703) );
  INV_X1 U20542 ( .A(n17363), .ZN(n17342) );
  INV_X1 U20543 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17503) );
  INV_X1 U20544 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17499) );
  INV_X1 U20545 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17497) );
  INV_X1 U20546 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17486) );
  INV_X1 U20547 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17546) );
  NAND3_X1 U20548 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n17373) );
  INV_X1 U20549 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17519) );
  INV_X1 U20550 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17517) );
  NOR2_X1 U20551 ( .A1(n17519), .A2(n17517), .ZN(n17285) );
  NAND4_X1 U20552 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(n17285), .ZN(n17374) );
  NOR2_X1 U20553 ( .A1(n17373), .A2(n17374), .ZN(n17404) );
  INV_X1 U20554 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17529) );
  INV_X1 U20555 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17527) );
  NAND4_X1 U20556 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n17286)
         );
  NOR3_X1 U20557 ( .A1(n17529), .A2(n17527), .A3(n17286), .ZN(n17375) );
  NAND4_X1 U20558 ( .A1(n17429), .A2(P3_EAX_REG_14__SCAN_IN), .A3(n17404), 
        .A4(n17375), .ZN(n17376) );
  INV_X1 U20559 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17495) );
  NOR2_X1 U20560 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17294), .ZN(n17287) );
  OAI21_X1 U20561 ( .B1(n19336), .B2(n17342), .A(n17288), .ZN(P3_U2704) );
  INV_X1 U20562 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17509) );
  NAND2_X1 U20563 ( .A1(n18287), .A2(n17394), .ZN(n17367) );
  OAI22_X1 U20564 ( .A1(n17289), .A2(n17422), .B1(n14378), .B2(n17342), .ZN(
        n17290) );
  AOI21_X1 U20565 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17356), .A(n17290), .ZN(
        n17291) );
  OAI221_X1 U20566 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17294), .C1(n17509), 
        .C2(n17292), .A(n17291), .ZN(P3_U2705) );
  AOI22_X1 U20567 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17356), .B1(n17293), .B2(
        n17434), .ZN(n17297) );
  OAI211_X1 U20568 ( .C1(n17295), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17438), .B(
        n17294), .ZN(n17296) );
  OAI211_X1 U20569 ( .C1(n17342), .C2(n17298), .A(n17297), .B(n17296), .ZN(
        P3_U2706) );
  AOI22_X1 U20570 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17363), .B1(n17299), .B2(
        n17434), .ZN(n17302) );
  OAI211_X1 U20571 ( .C1(n17304), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17438), .B(
        n17300), .ZN(n17301) );
  OAI211_X1 U20572 ( .C1(n17367), .C2(n17388), .A(n17302), .B(n17301), .ZN(
        P3_U2707) );
  INV_X1 U20573 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20574 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n17363), .B1(n17303), .B2(
        n17434), .ZN(n17307) );
  AOI211_X1 U20575 ( .C1(n17503), .C2(n17308), .A(n17304), .B(n17394), .ZN(
        n17305) );
  INV_X1 U20576 ( .A(n17305), .ZN(n17306) );
  OAI211_X1 U20577 ( .C1(n17367), .C2(n17392), .A(n17307), .B(n17306), .ZN(
        P3_U2708) );
  AOI22_X1 U20578 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17356), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17363), .ZN(n17310) );
  OAI211_X1 U20579 ( .C1(n17312), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17438), .B(
        n17308), .ZN(n17309) );
  OAI211_X1 U20580 ( .C1(n17311), .C2(n17422), .A(n17310), .B(n17309), .ZN(
        P3_U2709) );
  AOI22_X1 U20581 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17356), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17363), .ZN(n17315) );
  AOI211_X1 U20582 ( .C1(n17499), .C2(n17318), .A(n17312), .B(n17394), .ZN(
        n17313) );
  INV_X1 U20583 ( .A(n17313), .ZN(n17314) );
  OAI211_X1 U20584 ( .C1(n17316), .C2(n17422), .A(n17315), .B(n17314), .ZN(
        P3_U2710) );
  AOI22_X1 U20585 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17356), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17363), .ZN(n17321) );
  OAI21_X1 U20586 ( .B1(n17497), .B2(n17394), .A(n17317), .ZN(n17319) );
  NAND2_X1 U20587 ( .A1(n17319), .A2(n17318), .ZN(n17320) );
  OAI211_X1 U20588 ( .C1(n17322), .C2(n17422), .A(n17321), .B(n17320), .ZN(
        P3_U2711) );
  AOI211_X1 U20589 ( .C1(n17495), .C2(n17324), .A(n17394), .B(n17323), .ZN(
        n17325) );
  AOI21_X1 U20590 ( .B1(n17363), .B2(BUF2_REG_23__SCAN_IN), .A(n17325), .ZN(
        n17327) );
  NAND2_X1 U20591 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17356), .ZN(n17326) );
  OAI211_X1 U20592 ( .C1(n17328), .C2(n17422), .A(n17327), .B(n17326), .ZN(
        P3_U2712) );
  NAND2_X1 U20593 ( .A1(n18297), .A2(n17329), .ZN(n17337) );
  OAI22_X1 U20594 ( .A1(n17331), .A2(n17342), .B1(n17422), .B2(n17330), .ZN(
        n17332) );
  INV_X1 U20595 ( .A(n17332), .ZN(n17336) );
  NOR2_X1 U20596 ( .A1(n17333), .A2(n17364), .ZN(n17358) );
  NAND2_X1 U20597 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17358), .ZN(n17357) );
  OR2_X1 U20598 ( .A1(n17394), .A2(n17338), .ZN(n17346) );
  OAI21_X1 U20599 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17372), .A(n17346), .ZN(
        n17334) );
  AOI22_X1 U20600 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17356), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17334), .ZN(n17335) );
  OAI211_X1 U20601 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17337), .A(n17336), .B(
        n17335), .ZN(P3_U2713) );
  AOI22_X1 U20602 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17356), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17363), .ZN(n17340) );
  OAI211_X1 U20603 ( .C1(n17338), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17438), .B(
        n17337), .ZN(n17339) );
  OAI211_X1 U20604 ( .C1(n17341), .C2(n17422), .A(n17340), .B(n17339), .ZN(
        P3_U2714) );
  NAND2_X1 U20605 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17351), .ZN(n17347) );
  INV_X1 U20606 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n21095) );
  INV_X1 U20607 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19328) );
  OAI22_X1 U20608 ( .A1(n17343), .A2(n17422), .B1(n19328), .B2(n17342), .ZN(
        n17344) );
  AOI21_X1 U20609 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n17356), .A(n17344), .ZN(
        n17345) );
  OAI221_X1 U20610 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n17347), .C1(n21095), 
        .C2(n17346), .A(n17345), .ZN(P3_U2715) );
  AOI22_X1 U20611 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17356), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17363), .ZN(n17349) );
  OAI211_X1 U20612 ( .C1(n17351), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17438), .B(
        n17347), .ZN(n17348) );
  OAI211_X1 U20613 ( .C1(n17350), .C2(n17422), .A(n17349), .B(n17348), .ZN(
        P3_U2716) );
  AOI22_X1 U20614 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17356), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17363), .ZN(n17354) );
  AOI211_X1 U20615 ( .C1(n17486), .C2(n17357), .A(n17351), .B(n17394), .ZN(
        n17352) );
  INV_X1 U20616 ( .A(n17352), .ZN(n17353) );
  OAI211_X1 U20617 ( .C1(n17355), .C2(n17422), .A(n17354), .B(n17353), .ZN(
        P3_U2717) );
  AOI22_X1 U20618 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17356), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17363), .ZN(n17360) );
  OAI211_X1 U20619 ( .C1(n17358), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17438), .B(
        n17357), .ZN(n17359) );
  OAI211_X1 U20620 ( .C1(n17361), .C2(n17422), .A(n17360), .B(n17359), .ZN(
        P3_U2718) );
  AOI22_X1 U20621 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17363), .B1(n17434), .B2(
        n17362), .ZN(n17366) );
  OAI211_X1 U20622 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17368), .A(n17438), .B(
        n17364), .ZN(n17365) );
  OAI211_X1 U20623 ( .C1(n17367), .C2(n18264), .A(n17366), .B(n17365), .ZN(
        P3_U2719) );
  AOI211_X1 U20624 ( .C1(n17546), .C2(n17376), .A(n17394), .B(n17368), .ZN(
        n17369) );
  AOI21_X1 U20625 ( .B1(n17435), .B2(BUF2_REG_15__SCAN_IN), .A(n17369), .ZN(
        n17370) );
  OAI21_X1 U20626 ( .B1(n17371), .B2(n17422), .A(n17370), .ZN(P3_U2720) );
  AND2_X1 U20627 ( .A1(n17375), .A2(n17412), .ZN(n17381) );
  INV_X1 U20628 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17541) );
  AOI22_X1 U20629 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17435), .B1(n17381), .B2(
        n17541), .ZN(n17378) );
  NAND3_X1 U20630 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17438), .A3(n17376), 
        .ZN(n17377) );
  OAI211_X1 U20631 ( .C1(n17379), .C2(n17422), .A(n17378), .B(n17377), .ZN(
        P3_U2721) );
  INV_X1 U20632 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17536) );
  INV_X1 U20633 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17531) );
  NAND3_X1 U20634 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n17412), .ZN(n17399) );
  NAND2_X1 U20635 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17393), .ZN(n17384) );
  NOR2_X1 U20636 ( .A1(n17536), .A2(n17384), .ZN(n17387) );
  AOI21_X1 U20637 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17438), .A(n17387), .ZN(
        n17382) );
  OAI222_X1 U20638 ( .A1(n17425), .A2(n17383), .B1(n17382), .B2(n17381), .C1(
        n17422), .C2(n17380), .ZN(P3_U2722) );
  INV_X1 U20639 ( .A(n17384), .ZN(n17391) );
  AOI21_X1 U20640 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17438), .A(n17391), .ZN(
        n17386) );
  OAI222_X1 U20641 ( .A1(n17425), .A2(n17388), .B1(n17387), .B2(n17386), .C1(
        n17422), .C2(n17385), .ZN(P3_U2723) );
  AOI21_X1 U20642 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17438), .A(n17393), .ZN(
        n17390) );
  OAI222_X1 U20643 ( .A1(n17425), .A2(n17392), .B1(n17391), .B2(n17390), .C1(
        n17422), .C2(n17389), .ZN(P3_U2724) );
  INV_X1 U20644 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17398) );
  AOI211_X1 U20645 ( .C1(n17531), .C2(n17399), .A(n17394), .B(n17393), .ZN(
        n17395) );
  AOI21_X1 U20646 ( .B1(n17434), .B2(n17396), .A(n17395), .ZN(n17397) );
  OAI21_X1 U20647 ( .B1(n17398), .B2(n17425), .A(n17397), .ZN(P3_U2725) );
  INV_X1 U20648 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17403) );
  INV_X1 U20649 ( .A(n17399), .ZN(n17402) );
  AOI22_X1 U20650 ( .A1(n17412), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17438), .ZN(n17401) );
  OAI222_X1 U20651 ( .A1(n17425), .A2(n17403), .B1(n17402), .B2(n17401), .C1(
        n17422), .C2(n17400), .ZN(P3_U2726) );
  INV_X1 U20652 ( .A(n17412), .ZN(n17409) );
  INV_X1 U20653 ( .A(n17404), .ZN(n17405) );
  AOI21_X1 U20654 ( .B1(n18297), .B2(n17405), .A(n17436), .ZN(n17408) );
  AOI22_X1 U20655 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17435), .B1(n17434), .B2(
        n17406), .ZN(n17407) );
  OAI221_X1 U20656 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17409), .C1(n17527), 
        .C2(n17408), .A(n17407), .ZN(P3_U2727) );
  INV_X1 U20657 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18294) );
  INV_X1 U20658 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17523) );
  NOR3_X1 U20659 ( .A1(n17519), .A2(n17517), .A3(n17428), .ZN(n17424) );
  NAND2_X1 U20660 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17424), .ZN(n17413) );
  NOR2_X1 U20661 ( .A1(n17523), .A2(n17413), .ZN(n17416) );
  AOI21_X1 U20662 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17438), .A(n17416), .ZN(
        n17411) );
  OAI222_X1 U20663 ( .A1(n17425), .A2(n18294), .B1(n17412), .B2(n17411), .C1(
        n17422), .C2(n17410), .ZN(P3_U2728) );
  INV_X1 U20664 ( .A(n17413), .ZN(n17419) );
  AOI21_X1 U20665 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17438), .A(n17419), .ZN(
        n17415) );
  OAI222_X1 U20666 ( .A1(n18290), .A2(n17425), .B1(n17416), .B2(n17415), .C1(
        n17422), .C2(n17414), .ZN(P3_U2729) );
  AOI21_X1 U20667 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17438), .A(n17424), .ZN(
        n17418) );
  OAI222_X1 U20668 ( .A1(n18286), .A2(n17425), .B1(n17419), .B2(n17418), .C1(
        n17422), .C2(n17417), .ZN(P3_U2730) );
  INV_X1 U20669 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18281) );
  NOR2_X1 U20670 ( .A1(n17517), .A2(n17428), .ZN(n17420) );
  AOI21_X1 U20671 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17438), .A(n17420), .ZN(
        n17423) );
  OAI222_X1 U20672 ( .A1(n18281), .A2(n17425), .B1(n17424), .B2(n17423), .C1(
        n17422), .C2(n17421), .ZN(P3_U2731) );
  NAND2_X1 U20673 ( .A1(n17438), .A2(n17428), .ZN(n17432) );
  AOI22_X1 U20674 ( .A1(n17435), .A2(BUF2_REG_3__SCAN_IN), .B1(n17434), .B2(
        n17426), .ZN(n17427) );
  OAI221_X1 U20675 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17428), .C1(n17517), 
        .C2(n17432), .A(n17427), .ZN(P3_U2732) );
  INV_X1 U20676 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17515) );
  NAND3_X1 U20677 ( .A1(n17429), .A2(P3_EAX_REG_1__SCAN_IN), .A3(
        P3_EAX_REG_0__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U20678 ( .A1(n17435), .A2(BUF2_REG_2__SCAN_IN), .B1(n17434), .B2(
        n17430), .ZN(n17431) );
  OAI221_X1 U20679 ( .B1(n17432), .B2(n17515), .C1(n17432), .C2(n17437), .A(
        n17431), .ZN(P3_U2733) );
  AOI22_X1 U20680 ( .A1(n17435), .A2(BUF2_REG_1__SCAN_IN), .B1(n17434), .B2(
        n17433), .ZN(n17441) );
  NOR2_X1 U20681 ( .A1(n17436), .A2(n17511), .ZN(n17439) );
  OAI211_X1 U20682 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17439), .A(n17438), .B(
        n17437), .ZN(n17440) );
  NAND2_X1 U20683 ( .A1(n17441), .A2(n17440), .ZN(P3_U2734) );
  INV_X2 U20684 ( .A(n18940), .ZN(n18793) );
  NOR2_X4 U20685 ( .A1(n18793), .A2(n17461), .ZN(n17471) );
  AND2_X1 U20686 ( .A1(n17471), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AOI22_X1 U20687 ( .A1(n18793), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17445) );
  OAI21_X1 U20688 ( .B1(n17509), .B2(n17460), .A(n17445), .ZN(P3_U2737) );
  INV_X1 U20689 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U20690 ( .A1(n18793), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17446) );
  OAI21_X1 U20691 ( .B1(n17507), .B2(n17460), .A(n17446), .ZN(P3_U2738) );
  INV_X1 U20692 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17505) );
  AOI22_X1 U20693 ( .A1(n18793), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20694 ( .B1(n17505), .B2(n17460), .A(n17447), .ZN(P3_U2739) );
  AOI22_X1 U20695 ( .A1(n18793), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17448) );
  OAI21_X1 U20696 ( .B1(n17503), .B2(n17460), .A(n17448), .ZN(P3_U2740) );
  INV_X1 U20697 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17501) );
  AOI22_X1 U20698 ( .A1(n18793), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20699 ( .B1(n17501), .B2(n17460), .A(n17449), .ZN(P3_U2741) );
  AOI22_X1 U20700 ( .A1(n18793), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17450) );
  OAI21_X1 U20701 ( .B1(n17499), .B2(n17460), .A(n17450), .ZN(P3_U2742) );
  AOI22_X1 U20702 ( .A1(n18793), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17451) );
  OAI21_X1 U20703 ( .B1(n17497), .B2(n17460), .A(n17451), .ZN(P3_U2743) );
  AOI22_X1 U20704 ( .A1(n18793), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U20705 ( .B1(n17495), .B2(n17460), .A(n17452), .ZN(P3_U2744) );
  INV_X1 U20706 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U20707 ( .A1(n18793), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17453) );
  OAI21_X1 U20708 ( .B1(n17493), .B2(n17460), .A(n17453), .ZN(P3_U2745) );
  INV_X1 U20709 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17491) );
  AOI22_X1 U20710 ( .A1(n18793), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17454) );
  OAI21_X1 U20711 ( .B1(n17491), .B2(n17460), .A(n17454), .ZN(P3_U2746) );
  AOI22_X1 U20712 ( .A1(n18793), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17455) );
  OAI21_X1 U20713 ( .B1(n21095), .B2(n17460), .A(n17455), .ZN(P3_U2747) );
  INV_X1 U20714 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U20715 ( .A1(n18793), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17456) );
  OAI21_X1 U20716 ( .B1(n17488), .B2(n17460), .A(n17456), .ZN(P3_U2748) );
  AOI22_X1 U20717 ( .A1(n18793), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17457) );
  OAI21_X1 U20718 ( .B1(n17486), .B2(n17460), .A(n17457), .ZN(P3_U2749) );
  INV_X1 U20719 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n21000) );
  AOI22_X1 U20720 ( .A1(n18793), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17458) );
  OAI21_X1 U20721 ( .B1(n21000), .B2(n17460), .A(n17458), .ZN(P3_U2750) );
  INV_X1 U20722 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17483) );
  AOI22_X1 U20723 ( .A1(n18793), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20724 ( .B1(n17483), .B2(n17460), .A(n17459), .ZN(P3_U2751) );
  AOI22_X1 U20725 ( .A1(n18793), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17462) );
  OAI21_X1 U20726 ( .B1(n17546), .B2(n17479), .A(n17462), .ZN(P3_U2752) );
  AOI22_X1 U20727 ( .A1(n18793), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17463) );
  OAI21_X1 U20728 ( .B1(n17541), .B2(n17479), .A(n17463), .ZN(P3_U2753) );
  INV_X1 U20729 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U20730 ( .A1(n18793), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17464) );
  OAI21_X1 U20731 ( .B1(n17538), .B2(n17479), .A(n17464), .ZN(P3_U2754) );
  AOI22_X1 U20732 ( .A1(n18793), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17465) );
  OAI21_X1 U20733 ( .B1(n17536), .B2(n17479), .A(n17465), .ZN(P3_U2755) );
  INV_X1 U20734 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17533) );
  AOI22_X1 U20735 ( .A1(n18793), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20736 ( .B1(n17533), .B2(n17479), .A(n17466), .ZN(P3_U2756) );
  AOI22_X1 U20737 ( .A1(n18793), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17467) );
  OAI21_X1 U20738 ( .B1(n17531), .B2(n17479), .A(n17467), .ZN(P3_U2757) );
  AOI22_X1 U20739 ( .A1(n18793), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17468) );
  OAI21_X1 U20740 ( .B1(n17529), .B2(n17479), .A(n17468), .ZN(P3_U2758) );
  AOI22_X1 U20741 ( .A1(n18793), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20742 ( .B1(n17527), .B2(n17479), .A(n17469), .ZN(P3_U2759) );
  INV_X1 U20743 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U20744 ( .A1(n18793), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17470) );
  OAI21_X1 U20745 ( .B1(n17525), .B2(n17479), .A(n17470), .ZN(P3_U2760) );
  AOI22_X1 U20746 ( .A1(n18793), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17472) );
  OAI21_X1 U20747 ( .B1(n17523), .B2(n17479), .A(n17472), .ZN(P3_U2761) );
  INV_X1 U20748 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17521) );
  AOI22_X1 U20749 ( .A1(n18793), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17473) );
  OAI21_X1 U20750 ( .B1(n17521), .B2(n17479), .A(n17473), .ZN(P3_U2762) );
  AOI22_X1 U20751 ( .A1(n18793), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17474) );
  OAI21_X1 U20752 ( .B1(n17519), .B2(n17479), .A(n17474), .ZN(P3_U2763) );
  AOI22_X1 U20753 ( .A1(n18793), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17475) );
  OAI21_X1 U20754 ( .B1(n17517), .B2(n17479), .A(n17475), .ZN(P3_U2764) );
  AOI22_X1 U20755 ( .A1(n18793), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17476) );
  OAI21_X1 U20756 ( .B1(n17515), .B2(n17479), .A(n17476), .ZN(P3_U2765) );
  INV_X1 U20757 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U20758 ( .A1(n18793), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17477) );
  OAI21_X1 U20759 ( .B1(n17513), .B2(n17479), .A(n17477), .ZN(P3_U2766) );
  AOI22_X1 U20760 ( .A1(n18793), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17471), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17478) );
  OAI21_X1 U20761 ( .B1(n17511), .B2(n17479), .A(n17478), .ZN(P3_U2767) );
  NAND2_X2 U20762 ( .A1(n17480), .A2(n18786), .ZN(n17545) );
  AOI22_X1 U20763 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17543), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17542), .ZN(n17482) );
  OAI21_X1 U20764 ( .B1(n17483), .B2(n17545), .A(n17482), .ZN(P3_U2768) );
  AOI22_X1 U20765 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17543), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17542), .ZN(n17484) );
  OAI21_X1 U20766 ( .B1(n21000), .B2(n17545), .A(n17484), .ZN(P3_U2769) );
  AOI22_X1 U20767 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17543), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17542), .ZN(n17485) );
  OAI21_X1 U20768 ( .B1(n17486), .B2(n17545), .A(n17485), .ZN(P3_U2770) );
  AOI22_X1 U20769 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17542), .ZN(n17487) );
  OAI21_X1 U20770 ( .B1(n17488), .B2(n17545), .A(n17487), .ZN(P3_U2771) );
  AOI22_X1 U20771 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17542), .ZN(n17489) );
  OAI21_X1 U20772 ( .B1(n21095), .B2(n17545), .A(n17489), .ZN(P3_U2772) );
  AOI22_X1 U20773 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17542), .ZN(n17490) );
  OAI21_X1 U20774 ( .B1(n17491), .B2(n17545), .A(n17490), .ZN(P3_U2773) );
  AOI22_X1 U20775 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17542), .ZN(n17492) );
  OAI21_X1 U20776 ( .B1(n17493), .B2(n17545), .A(n17492), .ZN(P3_U2774) );
  AOI22_X1 U20777 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17542), .ZN(n17494) );
  OAI21_X1 U20778 ( .B1(n17495), .B2(n17545), .A(n17494), .ZN(P3_U2775) );
  AOI22_X1 U20779 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17542), .ZN(n17496) );
  OAI21_X1 U20780 ( .B1(n17497), .B2(n17545), .A(n17496), .ZN(P3_U2776) );
  AOI22_X1 U20781 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17542), .ZN(n17498) );
  OAI21_X1 U20782 ( .B1(n17499), .B2(n17545), .A(n17498), .ZN(P3_U2777) );
  AOI22_X1 U20783 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17542), .ZN(n17500) );
  OAI21_X1 U20784 ( .B1(n17501), .B2(n17545), .A(n17500), .ZN(P3_U2778) );
  AOI22_X1 U20785 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17542), .ZN(n17502) );
  OAI21_X1 U20786 ( .B1(n17503), .B2(n17545), .A(n17502), .ZN(P3_U2779) );
  AOI22_X1 U20787 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17543), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17542), .ZN(n17504) );
  OAI21_X1 U20788 ( .B1(n17505), .B2(n17545), .A(n17504), .ZN(P3_U2780) );
  AOI22_X1 U20789 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17543), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17542), .ZN(n17506) );
  OAI21_X1 U20790 ( .B1(n17507), .B2(n17545), .A(n17506), .ZN(P3_U2781) );
  AOI22_X1 U20791 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17543), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17542), .ZN(n17508) );
  OAI21_X1 U20792 ( .B1(n17509), .B2(n17545), .A(n17508), .ZN(P3_U2782) );
  AOI22_X1 U20793 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17542), .ZN(n17510) );
  OAI21_X1 U20794 ( .B1(n17511), .B2(n17545), .A(n17510), .ZN(P3_U2783) );
  AOI22_X1 U20795 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17542), .ZN(n17512) );
  OAI21_X1 U20796 ( .B1(n17513), .B2(n17545), .A(n17512), .ZN(P3_U2784) );
  AOI22_X1 U20797 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17542), .ZN(n17514) );
  OAI21_X1 U20798 ( .B1(n17515), .B2(n17545), .A(n17514), .ZN(P3_U2785) );
  AOI22_X1 U20799 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17539), .ZN(n17516) );
  OAI21_X1 U20800 ( .B1(n17517), .B2(n17545), .A(n17516), .ZN(P3_U2786) );
  AOI22_X1 U20801 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17539), .ZN(n17518) );
  OAI21_X1 U20802 ( .B1(n17519), .B2(n17545), .A(n17518), .ZN(P3_U2787) );
  AOI22_X1 U20803 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17539), .ZN(n17520) );
  OAI21_X1 U20804 ( .B1(n17521), .B2(n17545), .A(n17520), .ZN(P3_U2788) );
  AOI22_X1 U20805 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17539), .ZN(n17522) );
  OAI21_X1 U20806 ( .B1(n17523), .B2(n17545), .A(n17522), .ZN(P3_U2789) );
  AOI22_X1 U20807 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17539), .ZN(n17524) );
  OAI21_X1 U20808 ( .B1(n17525), .B2(n17545), .A(n17524), .ZN(P3_U2790) );
  AOI22_X1 U20809 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17539), .ZN(n17526) );
  OAI21_X1 U20810 ( .B1(n17527), .B2(n17545), .A(n17526), .ZN(P3_U2791) );
  AOI22_X1 U20811 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17539), .ZN(n17528) );
  OAI21_X1 U20812 ( .B1(n17529), .B2(n17545), .A(n17528), .ZN(P3_U2792) );
  AOI22_X1 U20813 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17542), .ZN(n17530) );
  OAI21_X1 U20814 ( .B1(n17531), .B2(n17545), .A(n17530), .ZN(P3_U2793) );
  AOI22_X1 U20815 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17539), .ZN(n17532) );
  OAI21_X1 U20816 ( .B1(n17533), .B2(n17545), .A(n17532), .ZN(P3_U2794) );
  AOI22_X1 U20817 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17542), .ZN(n17535) );
  OAI21_X1 U20818 ( .B1(n17536), .B2(n17545), .A(n17535), .ZN(P3_U2795) );
  AOI22_X1 U20819 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17539), .ZN(n17537) );
  OAI21_X1 U20820 ( .B1(n17538), .B2(n17545), .A(n17537), .ZN(P3_U2796) );
  AOI22_X1 U20821 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17539), .ZN(n17540) );
  OAI21_X1 U20822 ( .B1(n17541), .B2(n17545), .A(n17540), .ZN(P3_U2797) );
  AOI22_X1 U20823 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17543), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17542), .ZN(n17544) );
  OAI21_X1 U20824 ( .B1(n17546), .B2(n17545), .A(n17544), .ZN(P3_U2798) );
  INV_X1 U20825 ( .A(n17547), .ZN(n17565) );
  OAI21_X1 U20826 ( .B1(n17548), .B2(n18803), .A(n17916), .ZN(n17549) );
  AOI21_X1 U20827 ( .B1(n18252), .B2(n17553), .A(n17549), .ZN(n17586) );
  OAI21_X1 U20828 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17661), .A(
        n17586), .ZN(n17567) );
  NOR2_X1 U20829 ( .A1(n17825), .A2(n17909), .ZN(n17669) );
  AOI22_X1 U20830 ( .A1(n17923), .A2(n17825), .B1(n17924), .B2(n17909), .ZN(
        n17550) );
  INV_X1 U20831 ( .A(n17550), .ZN(n17582) );
  NOR2_X1 U20832 ( .A1(n17928), .A2(n17582), .ZN(n17552) );
  NOR3_X1 U20833 ( .A1(n17669), .A2(n17552), .A3(n17551), .ZN(n17559) );
  NOR2_X1 U20834 ( .A1(n17747), .A2(n17553), .ZN(n17572) );
  OAI211_X1 U20835 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17572), .B(n17554), .ZN(n17555) );
  OAI211_X1 U20836 ( .C1(n17769), .C2(n17557), .A(n17556), .B(n17555), .ZN(
        n17558) );
  AOI211_X1 U20837 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17567), .A(
        n17559), .B(n17558), .ZN(n17564) );
  OAI211_X1 U20838 ( .C1(n17562), .C2(n17561), .A(n17812), .B(n17560), .ZN(
        n17563) );
  OAI211_X1 U20839 ( .C1(n17565), .C2(n17630), .A(n17564), .B(n17563), .ZN(
        P3_U2802) );
  AOI22_X1 U20840 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17567), .B1(
        n17667), .B2(n17566), .ZN(n17576) );
  NAND2_X1 U20841 ( .A1(n17569), .A2(n17568), .ZN(n17570) );
  XOR2_X1 U20842 ( .A(n17570), .B(n17820), .Z(n17929) );
  AOI22_X1 U20843 ( .A1(n17812), .A2(n17929), .B1(n17572), .B2(n17571), .ZN(
        n17575) );
  AOI22_X1 U20844 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17582), .B1(
        n17573), .B2(n17928), .ZN(n17574) );
  NAND2_X1 U20845 ( .A1(n18235), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17930) );
  NAND4_X1 U20846 ( .A1(n17576), .A2(n17575), .A3(n17574), .A4(n17930), .ZN(
        P3_U2803) );
  AOI21_X1 U20847 ( .B1(n17577), .B2(n18392), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17585) );
  NAND2_X1 U20848 ( .A1(n17769), .A2(n17661), .ZN(n17699) );
  AOI22_X1 U20849 ( .A1(n18235), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17578), 
        .B2(n17699), .ZN(n17584) );
  AOI21_X1 U20850 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17580), .A(
        n17579), .ZN(n17941) );
  INV_X1 U20851 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17936) );
  NAND3_X1 U20852 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17945), .A3(
        n17936), .ZN(n17935) );
  OAI22_X1 U20853 ( .A1(n17941), .A2(n17823), .B1(n17630), .B2(n17935), .ZN(
        n17581) );
  AOI21_X1 U20854 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17582), .A(
        n17581), .ZN(n17583) );
  OAI211_X1 U20855 ( .C1(n17586), .C2(n17585), .A(n17584), .B(n17583), .ZN(
        P3_U2804) );
  NAND3_X1 U20856 ( .A1(n17945), .A2(n18057), .A3(n17946), .ZN(n17587) );
  XOR2_X1 U20857 ( .A(n17587), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17952) );
  INV_X1 U20858 ( .A(n17588), .ZN(n17621) );
  INV_X1 U20859 ( .A(n17916), .ZN(n17903) );
  AND2_X1 U20860 ( .A1(n17591), .A2(n18392), .ZN(n17589) );
  AOI211_X1 U20861 ( .C1(n17744), .C2(n17621), .A(n17903), .B(n17589), .ZN(
        n17624) );
  OAI21_X1 U20862 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17661), .A(
        n17624), .ZN(n17603) );
  INV_X1 U20863 ( .A(n17590), .ZN(n17594) );
  NOR2_X1 U20864 ( .A1(n17747), .A2(n17591), .ZN(n17605) );
  OAI211_X1 U20865 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17605), .B(n17592), .ZN(n17593) );
  NAND2_X1 U20866 ( .A1(n18140), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17949) );
  OAI211_X1 U20867 ( .C1(n17769), .C2(n17594), .A(n17593), .B(n17949), .ZN(
        n17600) );
  NAND3_X1 U20868 ( .A1(n17946), .A2(n17945), .A3(n18058), .ZN(n17595) );
  XOR2_X1 U20869 ( .A(n17595), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17958) );
  OAI21_X1 U20870 ( .B1(n11132), .B2(n17597), .A(n17596), .ZN(n17598) );
  XOR2_X1 U20871 ( .A(n17598), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17951) );
  OAI22_X1 U20872 ( .A1(n17753), .A2(n17958), .B1(n17823), .B2(n17951), .ZN(
        n17599) );
  AOI211_X1 U20873 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17603), .A(
        n17600), .B(n17599), .ZN(n17601) );
  OAI21_X1 U20874 ( .B1(n17920), .B2(n17952), .A(n17601), .ZN(P3_U2805) );
  INV_X1 U20875 ( .A(n17602), .ZN(n17614) );
  NOR2_X1 U20876 ( .A1(n16718), .A2(n18867), .ZN(n17959) );
  AOI221_X1 U20877 ( .B1(n17605), .B2(n17604), .C1(n17603), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17959), .ZN(n17613) );
  NOR2_X1 U20878 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17973), .ZN(
        n17961) );
  NAND2_X1 U20879 ( .A1(n18058), .A2(n17606), .ZN(n17964) );
  NAND2_X1 U20880 ( .A1(n18057), .A2(n17606), .ZN(n17962) );
  AOI22_X1 U20881 ( .A1(n17825), .A2(n17964), .B1(n17909), .B2(n17962), .ZN(
        n17629) );
  INV_X1 U20882 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17609) );
  AOI21_X1 U20883 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17608), .A(
        n17607), .ZN(n17972) );
  OAI22_X1 U20884 ( .A1(n17629), .A2(n17609), .B1(n17972), .B2(n17823), .ZN(
        n17610) );
  AOI21_X1 U20885 ( .B1(n17611), .B2(n17961), .A(n17610), .ZN(n17612) );
  OAI211_X1 U20886 ( .C1(n17769), .C2(n17614), .A(n17613), .B(n17612), .ZN(
        P3_U2806) );
  AOI22_X1 U20887 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n11132), .B1(
        n17615), .B2(n17631), .ZN(n17616) );
  NAND2_X1 U20888 ( .A1(n17659), .A2(n17616), .ZN(n17617) );
  XOR2_X1 U20889 ( .A(n17617), .B(n17973), .Z(n17977) );
  AOI21_X1 U20890 ( .B1(n17618), .B2(n18392), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17623) );
  NAND2_X1 U20891 ( .A1(n17620), .A2(n17619), .ZN(n17622) );
  OAI22_X1 U20892 ( .A1(n17624), .A2(n17623), .B1(n17622), .B2(n17621), .ZN(
        n17627) );
  OAI22_X1 U20893 ( .A1(n16718), .A2(n18866), .B1(n17769), .B2(n17625), .ZN(
        n17626) );
  AOI211_X1 U20894 ( .C1(n17812), .C2(n17977), .A(n17627), .B(n17626), .ZN(
        n17628) );
  OAI221_X1 U20895 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17630), 
        .C1(n17973), .C2(n17629), .A(n17628), .ZN(P3_U2807) );
  INV_X1 U20896 ( .A(n17631), .ZN(n17633) );
  NOR2_X1 U20897 ( .A1(n17632), .A2(n17983), .ZN(n17988) );
  OAI221_X1 U20898 ( .B1(n17633), .B2(n17988), .C1(n17633), .C2(n17709), .A(
        n17659), .ZN(n17634) );
  XOR2_X1 U20899 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17634), .Z(
        n17995) );
  OAI22_X1 U20900 ( .A1(n17753), .A2(n18058), .B1(n17920), .B2(n18057), .ZN(
        n17635) );
  OAI21_X1 U20901 ( .B1(n17669), .B2(n17988), .A(n17719), .ZN(n17656) );
  INV_X1 U20902 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18863) );
  OAI21_X1 U20903 ( .B1(n17636), .B2(n18803), .A(n17916), .ZN(n17637) );
  AOI21_X1 U20904 ( .B1(n18252), .B2(n17639), .A(n17637), .ZN(n17664) );
  OAI21_X1 U20905 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17661), .A(
        n17664), .ZN(n17648) );
  AOI22_X1 U20906 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17648), .B1(
        n17667), .B2(n17638), .ZN(n17642) );
  NOR2_X1 U20907 ( .A1(n17747), .A2(n17639), .ZN(n17650) );
  OAI211_X1 U20908 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17650), .B(n17640), .ZN(n17641) );
  OAI211_X1 U20909 ( .C1(n18863), .C2(n16718), .A(n17642), .B(n17641), .ZN(
        n17643) );
  AOI21_X1 U20910 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17656), .A(
        n17643), .ZN(n17645) );
  NAND3_X1 U20911 ( .A1(n17702), .A2(n17988), .A3(n17990), .ZN(n17644) );
  OAI211_X1 U20912 ( .C1(n17823), .C2(n17995), .A(n17645), .B(n17644), .ZN(
        P3_U2808) );
  NAND2_X1 U20913 ( .A1(n18000), .A2(n17655), .ZN(n18004) );
  NAND2_X1 U20914 ( .A1(n17996), .A2(n17702), .ZN(n17685) );
  OAI22_X1 U20915 ( .A1(n16718), .A2(n18862), .B1(n17769), .B2(n17646), .ZN(
        n17647) );
  AOI221_X1 U20916 ( .B1(n17650), .B2(n17649), .C1(n17648), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17647), .ZN(n17658) );
  INV_X1 U20917 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17652) );
  NOR3_X1 U20918 ( .A1(n11132), .A2(n17652), .A3(n17651), .ZN(n17678) );
  INV_X1 U20919 ( .A(n17688), .ZN(n17679) );
  AOI22_X1 U20920 ( .A1(n18000), .A2(n17678), .B1(n17679), .B2(n17653), .ZN(
        n17654) );
  XOR2_X1 U20921 ( .A(n17655), .B(n17654), .Z(n17997) );
  AOI22_X1 U20922 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17656), .B1(
        n17812), .B2(n17997), .ZN(n17657) );
  OAI211_X1 U20923 ( .C1(n18004), .C2(n17685), .A(n17658), .B(n17657), .ZN(
        P3_U2809) );
  OAI221_X1 U20924 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17686), 
        .C1(n17681), .C2(n17678), .A(n17659), .ZN(n17660) );
  XOR2_X1 U20925 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17660), .Z(
        n18014) );
  AOI21_X1 U20926 ( .B1(n17662), .B2(n18392), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17663) );
  OAI22_X1 U20927 ( .A1(n17664), .A2(n17663), .B1(n16718), .B2(n18859), .ZN(
        n17665) );
  AOI221_X1 U20928 ( .B1(n17667), .B2(n17666), .C1(n17620), .C2(n17666), .A(
        n17665), .ZN(n17671) );
  NAND2_X1 U20929 ( .A1(n17996), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18008) );
  INV_X1 U20930 ( .A(n18008), .ZN(n17668) );
  OAI21_X1 U20931 ( .B1(n17669), .B2(n17668), .A(n17719), .ZN(n17682) );
  NOR2_X1 U20932 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18008), .ZN(
        n18005) );
  AOI22_X1 U20933 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17682), .B1(
        n17702), .B2(n18005), .ZN(n17670) );
  OAI211_X1 U20934 ( .C1(n17823), .C2(n18014), .A(n17671), .B(n17670), .ZN(
        P3_U2810) );
  AOI21_X1 U20935 ( .B1(n18252), .B2(n17673), .A(n17903), .ZN(n17703) );
  OAI21_X1 U20936 ( .B1(n17672), .B2(n18803), .A(n17703), .ZN(n17691) );
  NOR2_X1 U20937 ( .A1(n17747), .A2(n17673), .ZN(n17693) );
  OAI211_X1 U20938 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17693), .B(n17674), .ZN(n17675) );
  NAND2_X1 U20939 ( .A1(n18140), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18017) );
  OAI211_X1 U20940 ( .C1(n17769), .C2(n17676), .A(n17675), .B(n18017), .ZN(
        n17677) );
  AOI21_X1 U20941 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17691), .A(
        n17677), .ZN(n17684) );
  AOI21_X1 U20942 ( .B1(n17686), .B2(n17679), .A(n17678), .ZN(n17680) );
  XOR2_X1 U20943 ( .A(n17681), .B(n17680), .Z(n18015) );
  AOI22_X1 U20944 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17682), .B1(
        n17812), .B2(n18015), .ZN(n17683) );
  OAI211_X1 U20945 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17685), .A(
        n17684), .B(n17683), .ZN(P3_U2811) );
  AOI21_X1 U20946 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17820), .A(
        n17686), .ZN(n17687) );
  XOR2_X1 U20947 ( .A(n17688), .B(n17687), .Z(n18036) );
  OAI22_X1 U20948 ( .A1(n16718), .A2(n18855), .B1(n17769), .B2(n17689), .ZN(
        n17690) );
  AOI221_X1 U20949 ( .B1(n17693), .B2(n17692), .C1(n17691), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17690), .ZN(n17696) );
  OAI21_X1 U20950 ( .B1(n18025), .B2(n17720), .A(n17719), .ZN(n17701) );
  INV_X1 U20951 ( .A(n18025), .ZN(n17694) );
  NOR2_X1 U20952 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17694), .ZN(
        n18032) );
  AOI22_X1 U20953 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17701), .B1(
        n17702), .B2(n18032), .ZN(n17695) );
  OAI211_X1 U20954 ( .C1(n17823), .C2(n18036), .A(n17696), .B(n17695), .ZN(
        P3_U2812) );
  OAI21_X1 U20955 ( .B1(n17698), .B2(n18040), .A(n17697), .ZN(n18039) );
  AOI22_X1 U20956 ( .A1(n17812), .A2(n18039), .B1(n17700), .B2(n17699), .ZN(
        n17708) );
  OAI221_X1 U20957 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17702), .A(n17701), .ZN(
        n17707) );
  NAND2_X1 U20958 ( .A1(n18140), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18042) );
  INV_X1 U20959 ( .A(n17703), .ZN(n17704) );
  OAI221_X1 U20960 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17705), .C1(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n18392), .A(n17704), .ZN(
        n17706) );
  NAND4_X1 U20961 ( .A1(n17708), .A2(n17707), .A3(n18042), .A4(n17706), .ZN(
        P3_U2813) );
  NAND2_X1 U20962 ( .A1(n17820), .A2(n17819), .ZN(n17803) );
  OAI22_X1 U20963 ( .A1(n17820), .A2(n17709), .B1(n17803), .B2(n18031), .ZN(
        n17710) );
  XOR2_X1 U20964 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17710), .Z(
        n18052) );
  AOI21_X1 U20965 ( .B1(n18252), .B2(n17712), .A(n17903), .ZN(n17742) );
  OAI21_X1 U20966 ( .B1(n17711), .B2(n18803), .A(n17742), .ZN(n17724) );
  AOI22_X1 U20967 ( .A1(n18140), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17724), .ZN(n17715) );
  NOR2_X1 U20968 ( .A1(n17747), .A2(n17712), .ZN(n17726) );
  OAI211_X1 U20969 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17726), .B(n17713), .ZN(n17714) );
  OAI211_X1 U20970 ( .C1(n17769), .C2(n17716), .A(n17715), .B(n17714), .ZN(
        n17717) );
  AOI21_X1 U20971 ( .B1(n17812), .B2(n18052), .A(n17717), .ZN(n17718) );
  OAI221_X1 U20972 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17720), 
        .C1(n18050), .C2(n17719), .A(n17718), .ZN(P3_U2814) );
  NOR2_X1 U20973 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17761), .ZN(
        n17733) );
  INV_X1 U20974 ( .A(n18100), .ZN(n18071) );
  NOR2_X1 U20975 ( .A1(n18071), .A2(n17803), .ZN(n17755) );
  NAND2_X1 U20976 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17756), .ZN(
        n18099) );
  OAI221_X1 U20977 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17733), 
        .C1(n18080), .C2(n17755), .A(n18099), .ZN(n17721) );
  XNOR2_X1 U20978 ( .A(n11127), .B(n17721), .ZN(n18065) );
  INV_X1 U20979 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17725) );
  NAND2_X1 U20980 ( .A1(n18140), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18067) );
  OAI21_X1 U20981 ( .B1(n17769), .B2(n17722), .A(n18067), .ZN(n17723) );
  AOI221_X1 U20982 ( .B1(n17726), .B2(n17725), .C1(n17724), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17723), .ZN(n17730) );
  NOR2_X1 U20983 ( .A1(n18058), .A2(n17753), .ZN(n17728) );
  NOR3_X1 U20984 ( .A1(n18110), .A2(n18071), .A3(n17756), .ZN(n17736) );
  NAND2_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17736), .ZN(
        n17735) );
  NAND2_X1 U20986 ( .A1(n11127), .A2(n17735), .ZN(n18060) );
  NOR2_X1 U20987 ( .A1(n18057), .A2(n17920), .ZN(n17727) );
  NAND2_X1 U20988 ( .A1(n11127), .A2(n17737), .ZN(n18062) );
  AOI22_X1 U20989 ( .A1(n17728), .A2(n18060), .B1(n17727), .B2(n18062), .ZN(
        n17729) );
  OAI211_X1 U20990 ( .C1(n17823), .C2(n18065), .A(n17730), .B(n17729), .ZN(
        P3_U2815) );
  AOI21_X1 U20991 ( .B1(n17731), .B2(n18392), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17741) );
  AOI22_X1 U20992 ( .A1(n18235), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17732), 
        .B2(n17699), .ZN(n17740) );
  OAI21_X1 U20993 ( .B1(n17755), .B2(n17733), .A(n18099), .ZN(n17734) );
  XOR2_X1 U20994 ( .A(n17734), .B(n18080), .Z(n18081) );
  OAI21_X1 U20995 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17736), .A(
        n17735), .ZN(n18087) );
  NOR2_X1 U20996 ( .A1(n18112), .A2(n18071), .ZN(n18091) );
  OAI221_X1 U20997 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18091), .A(n17737), .ZN(
        n18083) );
  OAI22_X1 U20998 ( .A1(n17753), .A2(n18087), .B1(n17920), .B2(n18083), .ZN(
        n17738) );
  AOI21_X1 U20999 ( .B1(n17812), .B2(n18081), .A(n17738), .ZN(n17739) );
  OAI211_X1 U21000 ( .C1(n17742), .C2(n17741), .A(n17740), .B(n17739), .ZN(
        P3_U2816) );
  INV_X1 U21001 ( .A(n17786), .ZN(n17815) );
  NOR2_X1 U21002 ( .A1(n17762), .A2(n17815), .ZN(n17772) );
  INV_X1 U21003 ( .A(n17772), .ZN(n17760) );
  AOI22_X1 U21004 ( .A1(n17744), .A2(n17743), .B1(n18252), .B2(n17746), .ZN(
        n17745) );
  NAND2_X1 U21005 ( .A1(n17745), .A2(n17916), .ZN(n17766) );
  NOR2_X1 U21006 ( .A1(n17747), .A2(n17746), .ZN(n17765) );
  OAI211_X1 U21007 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17765), .B(n17748), .ZN(n17750) );
  NAND2_X1 U21008 ( .A1(n18235), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17749) );
  OAI211_X1 U21009 ( .C1(n17769), .C2(n17751), .A(n17750), .B(n17749), .ZN(
        n17752) );
  AOI21_X1 U21010 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17766), .A(
        n17752), .ZN(n17759) );
  NOR2_X1 U21011 ( .A1(n18110), .A2(n18071), .ZN(n18093) );
  OAI22_X1 U21012 ( .A1(n18093), .A2(n17753), .B1(n18091), .B2(n17920), .ZN(
        n17771) );
  NOR2_X1 U21013 ( .A1(n17755), .A2(n17754), .ZN(n17757) );
  XOR2_X1 U21014 ( .A(n17757), .B(n17756), .Z(n18089) );
  AOI22_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17771), .B1(
        n17812), .B2(n18089), .ZN(n17758) );
  OAI211_X1 U21016 ( .C1(n18099), .C2(n17760), .A(n17759), .B(n17758), .ZN(
        P3_U2817) );
  OAI21_X1 U21017 ( .B1(n17762), .B2(n17803), .A(n17761), .ZN(n17763) );
  XOR2_X1 U21018 ( .A(n17763), .B(n21108), .Z(n18108) );
  AOI22_X1 U21019 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17766), .B1(
        n17765), .B2(n17764), .ZN(n17767) );
  NAND2_X1 U21020 ( .A1(n18140), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18106) );
  OAI211_X1 U21021 ( .C1(n17769), .C2(n17768), .A(n17767), .B(n18106), .ZN(
        n17770) );
  AOI221_X1 U21022 ( .B1(n17772), .B2(n21108), .C1(n17771), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17770), .ZN(n17773) );
  OAI21_X1 U21023 ( .B1(n18108), .B2(n17823), .A(n17773), .ZN(P3_U2818) );
  INV_X1 U21024 ( .A(n17774), .ZN(n17775) );
  OAI21_X1 U21025 ( .B1(n17803), .B2(n18117), .A(n17775), .ZN(n17776) );
  XOR2_X1 U21026 ( .A(n17776), .B(n17787), .Z(n18122) );
  NOR2_X1 U21027 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18117), .ZN(
        n18109) );
  NOR2_X1 U21028 ( .A1(n16718), .A2(n18841), .ZN(n17785) );
  NOR2_X1 U21029 ( .A1(n17777), .A2(n18666), .ZN(n17848) );
  AND2_X1 U21030 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17848), .ZN(
        n17835) );
  NAND2_X1 U21031 ( .A1(n17778), .A2(n17835), .ZN(n17779) );
  INV_X1 U21032 ( .A(n17779), .ZN(n17806) );
  NAND2_X1 U21033 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17806), .ZN(
        n17805) );
  NOR2_X1 U21034 ( .A1(n17792), .A2(n17805), .ZN(n17791) );
  AOI21_X1 U21035 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17911), .A(
        n17791), .ZN(n17783) );
  NOR2_X1 U21036 ( .A1(n17780), .A2(n17779), .ZN(n17782) );
  OAI22_X1 U21037 ( .A1(n17783), .A2(n17782), .B1(n17901), .B2(n17781), .ZN(
        n17784) );
  AOI211_X1 U21038 ( .C1(n18109), .C2(n17786), .A(n17785), .B(n17784), .ZN(
        n17790) );
  NAND2_X1 U21039 ( .A1(n18117), .A2(n17786), .ZN(n17800) );
  AOI22_X1 U21040 ( .A1(n18110), .A2(n17825), .B1(n17909), .B2(n18112), .ZN(
        n17814) );
  AOI21_X1 U21041 ( .B1(n17800), .B2(n17814), .A(n17787), .ZN(n17788) );
  INV_X1 U21042 ( .A(n17788), .ZN(n17789) );
  OAI211_X1 U21043 ( .C1(n18122), .C2(n17823), .A(n17790), .B(n17789), .ZN(
        P3_U2819) );
  AOI211_X1 U21044 ( .C1(n17805), .C2(n17792), .A(n17849), .B(n17791), .ZN(
        n17794) );
  NOR2_X1 U21045 ( .A1(n16718), .A2(n18839), .ZN(n17793) );
  AOI211_X1 U21046 ( .C1(n17795), .C2(n17699), .A(n17794), .B(n17793), .ZN(
        n17799) );
  INV_X1 U21047 ( .A(n17814), .ZN(n17797) );
  INV_X1 U21048 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18143) );
  AOI22_X1 U21049 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17803), .B1(
        n17802), .B2(n18143), .ZN(n17796) );
  XOR2_X1 U21050 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17796), .Z(
        n18124) );
  AOI22_X1 U21051 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17797), .B1(
        n17812), .B2(n18124), .ZN(n17798) );
  OAI211_X1 U21052 ( .C1(n17801), .C2(n17800), .A(n17799), .B(n17798), .ZN(
        P3_U2820) );
  NAND2_X1 U21053 ( .A1(n17803), .A2(n17802), .ZN(n17804) );
  XOR2_X1 U21054 ( .A(n17804), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18138) );
  NOR2_X1 U21055 ( .A1(n16718), .A2(n18837), .ZN(n17811) );
  INV_X1 U21056 ( .A(n17805), .ZN(n17809) );
  AOI21_X1 U21057 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17911), .A(
        n17806), .ZN(n17808) );
  OAI22_X1 U21058 ( .A1(n17809), .A2(n17808), .B1(n17901), .B2(n17807), .ZN(
        n17810) );
  AOI211_X1 U21059 ( .C1(n17812), .C2(n18138), .A(n17811), .B(n17810), .ZN(
        n17813) );
  OAI221_X1 U21060 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17815), .C1(
        n18143), .C2(n17814), .A(n17813), .ZN(P3_U2821) );
  OAI21_X1 U21061 ( .B1(n17817), .B2(n17816), .A(n17916), .ZN(n17833) );
  AOI22_X1 U21062 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17833), .B1(
        n17818), .B2(n17699), .ZN(n17830) );
  AOI21_X1 U21063 ( .B1(n9849), .B2(n21098), .A(n17819), .ZN(n18158) );
  XOR2_X1 U21064 ( .A(n18158), .B(n17820), .Z(n18162) );
  OAI21_X1 U21065 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17822), .A(
        n17821), .ZN(n18156) );
  OAI22_X1 U21066 ( .A1(n18162), .A2(n17823), .B1(n17920), .B2(n18156), .ZN(
        n17824) );
  AOI21_X1 U21067 ( .B1(n17825), .B2(n18158), .A(n17824), .ZN(n17829) );
  NAND2_X1 U21068 ( .A1(n18140), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18154) );
  OAI211_X1 U21069 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17827), .A(
        n18392), .B(n17826), .ZN(n17828) );
  NAND4_X1 U21070 ( .A1(n17830), .A2(n17829), .A3(n18154), .A4(n17828), .ZN(
        P3_U2822) );
  OAI21_X1 U21071 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17832), .A(
        n17831), .ZN(n18171) );
  NOR2_X1 U21072 ( .A1(n16718), .A2(n18834), .ZN(n18163) );
  AOI221_X1 U21073 ( .B1(n17835), .B2(n17834), .C1(n17833), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18163), .ZN(n17841) );
  NOR2_X1 U21074 ( .A1(n17837), .A2(n17836), .ZN(n17838) );
  XOR2_X1 U21075 ( .A(n17838), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18167) );
  AOI22_X1 U21076 ( .A1(n17909), .A2(n18167), .B1(n17839), .B2(n17699), .ZN(
        n17840) );
  OAI211_X1 U21077 ( .C1(n17919), .C2(n18171), .A(n17841), .B(n17840), .ZN(
        P3_U2823) );
  AOI22_X1 U21078 ( .A1(n17844), .A2(n17859), .B1(n17843), .B2(n17842), .ZN(
        n17846) );
  XNOR2_X1 U21079 ( .A(n17846), .B(n17845), .ZN(n18176) );
  AOI22_X1 U21080 ( .A1(n18140), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17848), 
        .B2(n17847), .ZN(n17856) );
  NOR2_X1 U21081 ( .A1(n17849), .A2(n17848), .ZN(n17866) );
  OAI21_X1 U21082 ( .B1(n17852), .B2(n17851), .A(n17850), .ZN(n18174) );
  OAI22_X1 U21083 ( .A1(n17901), .A2(n17853), .B1(n17919), .B2(n18174), .ZN(
        n17854) );
  AOI21_X1 U21084 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17866), .A(
        n17854), .ZN(n17855) );
  OAI211_X1 U21085 ( .C1(n18176), .C2(n17920), .A(n17856), .B(n17855), .ZN(
        P3_U2824) );
  OAI21_X1 U21086 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17858), .A(
        n17857), .ZN(n18190) );
  AOI21_X1 U21087 ( .B1(n17861), .B2(n17860), .A(n17859), .ZN(n18188) );
  AOI22_X1 U21088 ( .A1(n17909), .A2(n18188), .B1(n18140), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17868) );
  AOI21_X1 U21089 ( .B1(n17916), .B2(n17862), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17863) );
  INV_X1 U21090 ( .A(n17863), .ZN(n17865) );
  AOI22_X1 U21091 ( .A1(n17866), .A2(n17865), .B1(n17864), .B2(n17699), .ZN(
        n17867) );
  OAI211_X1 U21092 ( .C1(n17919), .C2(n18190), .A(n17868), .B(n17867), .ZN(
        P3_U2825) );
  OAI21_X1 U21093 ( .B1(n17871), .B2(n17870), .A(n17869), .ZN(n17872) );
  XOR2_X1 U21094 ( .A(n17872), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18201) );
  AOI22_X1 U21095 ( .A1(n18140), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18392), 
        .B2(n17873), .ZN(n17881) );
  AOI21_X1 U21096 ( .B1(n17876), .B2(n17875), .A(n17874), .ZN(n18198) );
  AOI21_X1 U21097 ( .B1(n18252), .B2(n17892), .A(n17903), .ZN(n17889) );
  OAI22_X1 U21098 ( .A1(n17901), .A2(n17878), .B1(n17889), .B2(n17877), .ZN(
        n17879) );
  AOI21_X1 U21099 ( .B1(n17909), .B2(n18198), .A(n17879), .ZN(n17880) );
  OAI211_X1 U21100 ( .C1(n17919), .C2(n18201), .A(n17881), .B(n17880), .ZN(
        P3_U2826) );
  OAI21_X1 U21101 ( .B1(n17884), .B2(n17883), .A(n17882), .ZN(n18202) );
  AOI21_X1 U21102 ( .B1(n17887), .B2(n17886), .A(n17885), .ZN(n18205) );
  NOR2_X1 U21103 ( .A1(n16718), .A2(n18826), .ZN(n18203) );
  OAI22_X1 U21104 ( .A1(n17901), .A2(n17890), .B1(n17889), .B2(n17888), .ZN(
        n17891) );
  AOI211_X1 U21105 ( .C1(n17909), .C2(n18205), .A(n18203), .B(n17891), .ZN(
        n17894) );
  NAND4_X1 U21106 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18252), .A3(
        n17916), .A4(n17892), .ZN(n17893) );
  OAI211_X1 U21107 ( .C1(n18202), .C2(n17919), .A(n17894), .B(n17893), .ZN(
        P3_U2827) );
  OAI21_X1 U21108 ( .B1(n17897), .B2(n17896), .A(n17895), .ZN(n18228) );
  XNOR2_X1 U21109 ( .A(n17899), .B(n17898), .ZN(n18222) );
  OAI22_X1 U21110 ( .A1(n17901), .A2(n17900), .B1(n17920), .B2(n18222), .ZN(
        n17902) );
  AOI221_X1 U21111 ( .B1(n17903), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18392), .C2(n21003), .A(n17902), .ZN(n17904) );
  NAND2_X1 U21112 ( .A1(n18235), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18226) );
  OAI211_X1 U21113 ( .C1(n17919), .C2(n18228), .A(n17904), .B(n18226), .ZN(
        P3_U2828) );
  OAI21_X1 U21114 ( .B1(n17915), .B2(n17906), .A(n17905), .ZN(n18239) );
  OAI21_X1 U21115 ( .B1(n17908), .B2(n17914), .A(n17907), .ZN(n18234) );
  AOI22_X1 U21116 ( .A1(n17909), .A2(n18234), .B1(n18140), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17913) );
  AOI22_X1 U21117 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17911), .B1(
        n17699), .B2(n17910), .ZN(n17912) );
  OAI211_X1 U21118 ( .C1(n17919), .C2(n18239), .A(n17913), .B(n17912), .ZN(
        P3_U2829) );
  NOR2_X1 U21119 ( .A1(n17915), .A2(n17914), .ZN(n18241) );
  INV_X1 U21120 ( .A(n18241), .ZN(n18243) );
  NAND3_X1 U21121 ( .A1(n21022), .A2(n18803), .A3(n17916), .ZN(n17917) );
  AOI22_X1 U21122 ( .A1(n18235), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17917), .ZN(n17918) );
  OAI221_X1 U21123 ( .B1(n18241), .B2(n17920), .C1(n18243), .C2(n17919), .A(
        n17918), .ZN(P3_U2830) );
  AOI21_X1 U21124 ( .B1(n18224), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17921), .ZN(n17933) );
  AOI22_X1 U21125 ( .A1(n18739), .A2(n17950), .B1(n18759), .B2(n17922), .ZN(
        n17927) );
  AOI22_X1 U21126 ( .A1(n18113), .A2(n17924), .B1(n18111), .B2(n17923), .ZN(
        n17926) );
  NAND2_X1 U21127 ( .A1(n18759), .A2(n18913), .ZN(n18214) );
  NAND3_X1 U21128 ( .A1(n18020), .A2(n17946), .A3(n18214), .ZN(n17963) );
  INV_X1 U21129 ( .A(n18213), .ZN(n18146) );
  OAI21_X1 U21130 ( .B1(n17942), .B2(n17963), .A(n18146), .ZN(n17943) );
  NAND4_X1 U21131 ( .A1(n17927), .A2(n17926), .A3(n17925), .A4(n17943), .ZN(
        n17934) );
  AOI211_X1 U21132 ( .C1(n18739), .C2(n17936), .A(n17928), .B(n17934), .ZN(
        n17932) );
  AOI22_X1 U21133 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18225), .B1(
        n18139), .B2(n17929), .ZN(n17931) );
  OAI211_X1 U21134 ( .C1(n17933), .C2(n17932), .A(n17931), .B(n17930), .ZN(
        P3_U2835) );
  INV_X1 U21135 ( .A(n17934), .ZN(n17937) );
  NAND3_X1 U21136 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17988), .A3(
        n17987), .ZN(n17974) );
  OAI22_X1 U21137 ( .A1(n17937), .A2(n17936), .B1(n17935), .B2(n17974), .ZN(
        n17938) );
  AOI22_X1 U21138 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18225), .B1(
        n18224), .B2(n17938), .ZN(n17940) );
  NAND2_X1 U21139 ( .A1(n18140), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17939) );
  OAI211_X1 U21140 ( .C1(n17941), .C2(n18161), .A(n17940), .B(n17939), .ZN(
        P3_U2836) );
  AOI221_X1 U21141 ( .B1(n17942), .B2(n18220), .C1(n17967), .C2(n18220), .A(
        n17950), .ZN(n17944) );
  AOI21_X1 U21142 ( .B1(n17944), .B2(n17943), .A(n18245), .ZN(n17956) );
  NAND2_X1 U21143 ( .A1(n17946), .A2(n17945), .ZN(n17947) );
  OAI21_X1 U21144 ( .B1(n17948), .B2(n17947), .A(n17950), .ZN(n17955) );
  OAI21_X1 U21145 ( .B1(n18230), .B2(n17950), .A(n17949), .ZN(n17954) );
  OAI22_X1 U21146 ( .A1(n18175), .A2(n17952), .B1(n18161), .B2(n17951), .ZN(
        n17953) );
  AOI211_X1 U21147 ( .C1(n17956), .C2(n17955), .A(n17954), .B(n17953), .ZN(
        n17957) );
  OAI21_X1 U21148 ( .B1(n18088), .B2(n17958), .A(n17957), .ZN(P3_U2837) );
  AOI21_X1 U21149 ( .B1(n17961), .B2(n17960), .A(n17959), .ZN(n17971) );
  INV_X1 U21150 ( .A(n17962), .ZN(n17966) );
  AOI22_X1 U21151 ( .A1(n18111), .A2(n17964), .B1(n18146), .B2(n17963), .ZN(
        n17965) );
  OAI211_X1 U21152 ( .C1(n17966), .C2(n18723), .A(n17965), .B(n18230), .ZN(
        n17969) );
  AOI211_X1 U21153 ( .C1(n18220), .C2(n17967), .A(n17973), .B(n17969), .ZN(
        n17968) );
  NOR2_X1 U21154 ( .A1(n18235), .A2(n17968), .ZN(n17976) );
  OAI211_X1 U21155 ( .C1(n18149), .C2(n17969), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17976), .ZN(n17970) );
  OAI211_X1 U21156 ( .C1(n17972), .C2(n18161), .A(n17971), .B(n17970), .ZN(
        P3_U2838) );
  OAI21_X1 U21157 ( .B1(n18225), .B2(n17974), .A(n17973), .ZN(n17975) );
  AOI22_X1 U21158 ( .A1(n18139), .A2(n17977), .B1(n17976), .B2(n17975), .ZN(
        n17978) );
  OAI21_X1 U21159 ( .B1(n16718), .B2(n18866), .A(n17978), .ZN(P3_U2839) );
  OAI21_X1 U21160 ( .B1(n17990), .B2(n18759), .A(n17979), .ZN(n17980) );
  INV_X1 U21161 ( .A(n17980), .ZN(n17981) );
  OAI22_X1 U21162 ( .A1(n18723), .A2(n18057), .B1(n18092), .B2(n18058), .ZN(
        n18027) );
  AOI211_X1 U21163 ( .C1(n17983), .C2(n17982), .A(n17981), .B(n18027), .ZN(
        n17991) );
  OAI21_X1 U21164 ( .B1(n17984), .B2(n18008), .A(n18739), .ZN(n17985) );
  OAI221_X1 U21165 ( .B1(n18752), .B2(n17996), .C1(n18752), .C2(n18021), .A(
        n17985), .ZN(n18007) );
  NAND2_X1 U21166 ( .A1(n18723), .A2(n18092), .ZN(n18116) );
  INV_X1 U21167 ( .A(n18116), .ZN(n18024) );
  OAI22_X1 U21168 ( .A1(n18761), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17988), .B2(n18024), .ZN(n17986) );
  NOR2_X1 U21169 ( .A1(n18007), .A2(n17986), .ZN(n17999) );
  NAND2_X1 U21170 ( .A1(n17988), .A2(n17987), .ZN(n17989) );
  AOI22_X1 U21171 ( .A1(n17991), .A2(n17999), .B1(n17990), .B2(n17989), .ZN(
        n17992) );
  AOI22_X1 U21172 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18225), .B1(
        n18224), .B2(n17992), .ZN(n17994) );
  NAND2_X1 U21173 ( .A1(n18140), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17993) );
  OAI211_X1 U21174 ( .C1(n17995), .C2(n18161), .A(n17994), .B(n17993), .ZN(
        P3_U2840) );
  NAND2_X1 U21175 ( .A1(n17996), .A2(n18006), .ZN(n18019) );
  AOI22_X1 U21176 ( .A1(n18140), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18139), 
        .B2(n17997), .ZN(n18003) );
  OR2_X1 U21177 ( .A1(n18245), .A2(n18027), .ZN(n18049) );
  NOR2_X1 U21178 ( .A1(n18220), .A2(n18759), .ZN(n18229) );
  OR2_X1 U21179 ( .A1(n18749), .A2(n17998), .ZN(n18009) );
  OAI211_X1 U21180 ( .C1(n18229), .C2(n18000), .A(n18009), .B(n17999), .ZN(
        n18001) );
  OAI211_X1 U21181 ( .C1(n18049), .C2(n18001), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n16718), .ZN(n18002) );
  OAI211_X1 U21182 ( .C1(n18004), .C2(n18019), .A(n18003), .B(n18002), .ZN(
        P3_U2841) );
  AOI22_X1 U21183 ( .A1(n18235), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18006), 
        .B2(n18005), .ZN(n18013) );
  AOI211_X1 U21184 ( .C1(n18008), .C2(n18116), .A(n18049), .B(n18007), .ZN(
        n18010) );
  AOI21_X1 U21185 ( .B1(n18010), .B2(n18009), .A(n18235), .ZN(n18016) );
  NOR3_X1 U21186 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18229), .A3(
        n18948), .ZN(n18011) );
  OAI21_X1 U21187 ( .B1(n18016), .B2(n18011), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18012) );
  OAI211_X1 U21188 ( .C1(n18014), .C2(n18161), .A(n18013), .B(n18012), .ZN(
        P3_U2842) );
  AOI22_X1 U21189 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18016), .B1(
        n18139), .B2(n18015), .ZN(n18018) );
  OAI211_X1 U21190 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18019), .A(
        n18018), .B(n18017), .ZN(P3_U2843) );
  NAND3_X1 U21191 ( .A1(n18020), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18214), .ZN(n18028) );
  AOI21_X1 U21192 ( .B1(n18025), .B2(n18021), .A(n18752), .ZN(n18022) );
  INV_X1 U21193 ( .A(n18022), .ZN(n18023) );
  OAI211_X1 U21194 ( .C1(n18025), .C2(n18024), .A(n18023), .B(n18230), .ZN(
        n18026) );
  AOI211_X1 U21195 ( .C1(n18146), .C2(n18028), .A(n18027), .B(n18026), .ZN(
        n18037) );
  AOI221_X1 U21196 ( .B1(n18213), .B2(n18037), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18037), .A(n18235), .ZN(
        n18033) );
  INV_X1 U21197 ( .A(n18193), .ZN(n18211) );
  AOI22_X1 U21198 ( .A1(n18211), .A2(n18220), .B1(n18191), .B2(n18215), .ZN(
        n18150) );
  NOR2_X1 U21199 ( .A1(n18173), .A2(n18150), .ZN(n18164) );
  NAND2_X1 U21200 ( .A1(n18029), .A2(n18164), .ZN(n18076) );
  AOI21_X1 U21201 ( .B1(n18076), .B2(n18030), .A(n18245), .ZN(n18123) );
  INV_X1 U21202 ( .A(n18123), .ZN(n18144) );
  NOR2_X1 U21203 ( .A1(n18031), .A2(n18144), .ZN(n18051) );
  AOI22_X1 U21204 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18033), .B1(
        n18032), .B2(n18051), .ZN(n18035) );
  NAND2_X1 U21205 ( .A1(n18235), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18034) );
  OAI211_X1 U21206 ( .C1(n18036), .C2(n18161), .A(n18035), .B(n18034), .ZN(
        P3_U2844) );
  NOR3_X1 U21207 ( .A1(n18235), .A2(n18037), .A3(n18040), .ZN(n18038) );
  AOI21_X1 U21208 ( .B1(n18139), .B2(n18039), .A(n18038), .ZN(n18043) );
  NAND3_X1 U21209 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18051), .A3(
        n18040), .ZN(n18041) );
  NAND3_X1 U21210 ( .A1(n18043), .A2(n18042), .A3(n18041), .ZN(P3_U2845) );
  INV_X1 U21211 ( .A(n18070), .ZN(n18046) );
  INV_X1 U21212 ( .A(n18044), .ZN(n18145) );
  OAI21_X1 U21213 ( .B1(n18151), .B2(n18145), .A(n18739), .ZN(n18045) );
  OAI21_X1 U21214 ( .B1(n18046), .B2(n18752), .A(n18045), .ZN(n18137) );
  AOI21_X1 U21215 ( .B1(n18739), .B2(n21098), .A(n18137), .ZN(n18126) );
  OAI21_X1 U21216 ( .B1(n11127), .B2(n18759), .A(n18047), .ZN(n18048) );
  OAI211_X1 U21217 ( .C1(n18127), .C2(n18055), .A(n18126), .B(n18048), .ZN(
        n18063) );
  OAI221_X1 U21218 ( .B1(n18049), .B2(n18149), .C1(n18049), .C2(n18063), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18054) );
  AOI22_X1 U21219 ( .A1(n18139), .A2(n18052), .B1(n18051), .B2(n18050), .ZN(
        n18053) );
  OAI221_X1 U21220 ( .B1(n18140), .B2(n18054), .C1(n16718), .C2(n18851), .A(
        n18053), .ZN(P3_U2846) );
  INV_X1 U21221 ( .A(n18055), .ZN(n18056) );
  OAI21_X1 U21222 ( .B1(n18056), .B2(n18076), .A(n11127), .ZN(n18064) );
  NOR2_X1 U21223 ( .A1(n18057), .A2(n18723), .ZN(n18061) );
  NOR2_X1 U21224 ( .A1(n18058), .A2(n18092), .ZN(n18059) );
  AOI222_X1 U21225 ( .A1(n18064), .A2(n18063), .B1(n18062), .B2(n18061), .C1(
        n18060), .C2(n18059), .ZN(n18069) );
  INV_X1 U21226 ( .A(n18065), .ZN(n18066) );
  AOI22_X1 U21227 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18225), .B1(
        n18139), .B2(n18066), .ZN(n18068) );
  OAI211_X1 U21228 ( .C1(n18069), .C2(n18245), .A(n18068), .B(n18067), .ZN(
        P3_U2847) );
  AOI21_X1 U21229 ( .B1(n18100), .B2(n18135), .A(n18749), .ZN(n18096) );
  AOI221_X1 U21230 ( .B1(n18071), .B2(n18220), .C1(n18070), .C2(n18220), .A(
        n18080), .ZN(n18074) );
  OAI21_X1 U21231 ( .B1(n18077), .B2(n18072), .A(n18739), .ZN(n18073) );
  OAI211_X1 U21232 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18229), .A(
        n18074), .B(n18073), .ZN(n18075) );
  OAI21_X1 U21233 ( .B1(n18096), .B2(n18075), .A(n18224), .ZN(n18079) );
  OR2_X1 U21234 ( .A1(n18077), .A2(n18076), .ZN(n18078) );
  AOI222_X1 U21235 ( .A1(n18080), .A2(n18079), .B1(n18080), .B2(n18078), .C1(
        n18079), .C2(n18230), .ZN(n18085) );
  INV_X1 U21236 ( .A(n18081), .ZN(n18082) );
  OAI22_X1 U21237 ( .A1(n18175), .A2(n18083), .B1(n18161), .B2(n18082), .ZN(
        n18084) );
  AOI211_X1 U21238 ( .C1(n18235), .C2(P3_REIP_REG_14__SCAN_IN), .A(n18085), 
        .B(n18084), .ZN(n18086) );
  OAI21_X1 U21239 ( .B1(n18088), .B2(n18087), .A(n18086), .ZN(P3_U2848) );
  NAND2_X1 U21240 ( .A1(n18090), .A2(n18123), .ZN(n18103) );
  AOI22_X1 U21241 ( .A1(n18235), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18139), 
        .B2(n18089), .ZN(n18098) );
  OAI21_X1 U21242 ( .B1(n18090), .B2(n18127), .A(n18126), .ZN(n18119) );
  OAI22_X1 U21243 ( .A1(n18093), .A2(n18092), .B1(n18091), .B2(n18723), .ZN(
        n18094) );
  NOR2_X1 U21244 ( .A1(n18119), .A2(n18094), .ZN(n18101) );
  OAI211_X1 U21245 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18127), .A(
        n18224), .B(n18101), .ZN(n18095) );
  OAI211_X1 U21246 ( .C1(n18096), .C2(n18095), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n16718), .ZN(n18097) );
  OAI211_X1 U21247 ( .C1(n18099), .C2(n18103), .A(n18098), .B(n18097), .ZN(
        P3_U2849) );
  AND2_X1 U21248 ( .A1(n18100), .A2(n18135), .ZN(n18102) );
  OAI211_X1 U21249 ( .C1(n18102), .C2(n18749), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18101), .ZN(n18105) );
  OAI21_X1 U21250 ( .B1(n18245), .B2(n21108), .A(n18103), .ZN(n18104) );
  AOI22_X1 U21251 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18225), .B1(
        n18105), .B2(n18104), .ZN(n18107) );
  OAI211_X1 U21252 ( .C1(n18108), .C2(n18161), .A(n18107), .B(n18106), .ZN(
        P3_U2850) );
  AOI22_X1 U21253 ( .A1(n18140), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18123), 
        .B2(n18109), .ZN(n18121) );
  AOI21_X1 U21254 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18135), .A(
        n18749), .ZN(n18115) );
  AOI22_X1 U21255 ( .A1(n18113), .A2(n18112), .B1(n18111), .B2(n18110), .ZN(
        n18114) );
  NAND2_X1 U21256 ( .A1(n18114), .A2(n18230), .ZN(n18132) );
  AOI211_X1 U21257 ( .C1(n18117), .C2(n18116), .A(n18115), .B(n18132), .ZN(
        n18125) );
  OAI21_X1 U21258 ( .B1(n18749), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18125), .ZN(n18118) );
  OAI211_X1 U21259 ( .C1(n18119), .C2(n18118), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16718), .ZN(n18120) );
  OAI211_X1 U21260 ( .C1(n18122), .C2(n18161), .A(n18121), .B(n18120), .ZN(
        P3_U2851) );
  NAND2_X1 U21261 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18123), .ZN(
        n18131) );
  AOI22_X1 U21262 ( .A1(n18235), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18139), 
        .B2(n18124), .ZN(n18130) );
  OAI211_X1 U21263 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18127), .A(
        n18126), .B(n18125), .ZN(n18128) );
  NAND3_X1 U21264 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16718), .A3(
        n18128), .ZN(n18129) );
  OAI211_X1 U21265 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n18131), .A(
        n18130), .B(n18129), .ZN(P3_U2852) );
  NAND2_X1 U21266 ( .A1(n18739), .A2(n21098), .ZN(n18134) );
  INV_X1 U21267 ( .A(n18132), .ZN(n18133) );
  OAI211_X1 U21268 ( .C1(n18135), .C2(n18749), .A(n18134), .B(n18133), .ZN(
        n18136) );
  OAI21_X1 U21269 ( .B1(n18137), .B2(n18136), .A(n16718), .ZN(n18142) );
  AOI22_X1 U21270 ( .A1(n18140), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18139), 
        .B2(n18138), .ZN(n18141) );
  OAI221_X1 U21271 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18144), .C1(
        n18143), .C2(n18142), .A(n18141), .ZN(P3_U2853) );
  NAND2_X1 U21272 ( .A1(n18146), .A2(n18145), .ZN(n18147) );
  OAI211_X1 U21273 ( .C1(n18148), .C2(n18752), .A(n18214), .B(n18147), .ZN(
        n18172) );
  AOI21_X1 U21274 ( .B1(n18149), .B2(n18151), .A(n18172), .ZN(n18165) );
  OAI21_X1 U21275 ( .B1(n18165), .B2(n18231), .A(n18230), .ZN(n18153) );
  OR2_X1 U21276 ( .A1(n18245), .A2(n18150), .ZN(n18209) );
  NOR3_X1 U21277 ( .A1(n18173), .A2(n18151), .A3(n18209), .ZN(n18152) );
  AOI22_X1 U21278 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18153), .B1(
        n18152), .B2(n21098), .ZN(n18155) );
  OAI211_X1 U21279 ( .C1(n18156), .C2(n18175), .A(n18155), .B(n18154), .ZN(
        n18157) );
  AOI21_X1 U21280 ( .B1(n18159), .B2(n18158), .A(n18157), .ZN(n18160) );
  OAI21_X1 U21281 ( .B1(n18162), .B2(n18161), .A(n18160), .ZN(P3_U2854) );
  AOI21_X1 U21282 ( .B1(n18225), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18163), .ZN(n18170) );
  INV_X1 U21283 ( .A(n18164), .ZN(n18166) );
  AOI221_X1 U21284 ( .B1(n18181), .B2(n21142), .C1(n18166), .C2(n21142), .A(
        n18165), .ZN(n18168) );
  AOI22_X1 U21285 ( .A1(n18224), .A2(n18168), .B1(n18244), .B2(n18167), .ZN(
        n18169) );
  OAI211_X1 U21286 ( .C1(n18238), .C2(n18171), .A(n18170), .B(n18169), .ZN(
        P3_U2855) );
  AOI21_X1 U21287 ( .B1(n18224), .B2(n18172), .A(n18225), .ZN(n18183) );
  NOR2_X1 U21288 ( .A1(n18173), .A2(n18209), .ZN(n18178) );
  OAI22_X1 U21289 ( .A1(n18176), .A2(n18175), .B1(n18238), .B2(n18174), .ZN(
        n18177) );
  AOI21_X1 U21290 ( .B1(n18178), .B2(n18181), .A(n18177), .ZN(n18180) );
  NAND2_X1 U21291 ( .A1(n18235), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18179) );
  OAI211_X1 U21292 ( .C1(n18183), .C2(n18181), .A(n18180), .B(n18179), .ZN(
        P3_U2856) );
  NOR2_X1 U21293 ( .A1(n16718), .A2(n18830), .ZN(n18187) );
  NAND2_X1 U21294 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18182) );
  NOR2_X1 U21295 ( .A1(n18182), .A2(n18209), .ZN(n18185) );
  INV_X1 U21296 ( .A(n18183), .ZN(n18184) );
  MUX2_X1 U21297 ( .A(n18185), .B(n18184), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18186) );
  AOI211_X1 U21298 ( .C1(n18244), .C2(n18188), .A(n18187), .B(n18186), .ZN(
        n18189) );
  OAI21_X1 U21299 ( .B1(n18238), .B2(n18190), .A(n18189), .ZN(P3_U2857) );
  OAI211_X1 U21300 ( .C1(n18213), .C2(n18191), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18214), .ZN(n18192) );
  AOI21_X1 U21301 ( .B1(n18220), .B2(n18193), .A(n18192), .ZN(n18210) );
  AOI221_X1 U21302 ( .B1(n18210), .B2(n18230), .C1(n18231), .C2(n18230), .A(
        n18194), .ZN(n18197) );
  NOR3_X1 U21303 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18195), .A3(
        n18209), .ZN(n18196) );
  AOI211_X1 U21304 ( .C1(n18198), .C2(n18244), .A(n18197), .B(n18196), .ZN(
        n18200) );
  NAND2_X1 U21305 ( .A1(n18235), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18199) );
  OAI211_X1 U21306 ( .C1(n18238), .C2(n18201), .A(n18200), .B(n18199), .ZN(
        P3_U2858) );
  INV_X1 U21307 ( .A(n18202), .ZN(n18204) );
  AOI21_X1 U21308 ( .B1(n18242), .B2(n18204), .A(n18203), .ZN(n18208) );
  OAI21_X1 U21309 ( .B1(n18210), .B2(n18245), .A(n18230), .ZN(n18206) );
  AOI22_X1 U21310 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18206), .B1(
        n18244), .B2(n18205), .ZN(n18207) );
  OAI211_X1 U21311 ( .C1(n18210), .C2(n18209), .A(n18208), .B(n18207), .ZN(
        P3_U2859) );
  OAI21_X1 U21312 ( .B1(n18913), .B2(n18212), .A(n18211), .ZN(n18219) );
  AOI211_X1 U21313 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18214), .A(
        n18213), .B(n18216), .ZN(n18218) );
  AND3_X1 U21314 ( .A1(n18216), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n18215), .ZN(n18217) );
  AOI211_X1 U21315 ( .C1(n18220), .C2(n18219), .A(n18218), .B(n18217), .ZN(
        n18221) );
  OAI21_X1 U21316 ( .B1(n18723), .B2(n18222), .A(n18221), .ZN(n18223) );
  AOI22_X1 U21317 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18225), .B1(
        n18224), .B2(n18223), .ZN(n18227) );
  OAI211_X1 U21318 ( .C1(n18238), .C2(n18228), .A(n18227), .B(n18226), .ZN(
        P3_U2860) );
  OR3_X1 U21319 ( .A1(n18245), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18229), .ZN(n18247) );
  AOI21_X1 U21320 ( .B1(n18230), .B2(n18247), .A(n20976), .ZN(n18233) );
  AOI211_X1 U21321 ( .C1(n18761), .C2(n18913), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18231), .ZN(n18232) );
  AOI211_X1 U21322 ( .C1(n18244), .C2(n18234), .A(n18233), .B(n18232), .ZN(
        n18237) );
  NAND2_X1 U21323 ( .A1(n18235), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18236) );
  OAI211_X1 U21324 ( .C1(n18239), .C2(n18238), .A(n18237), .B(n18236), .ZN(
        P3_U2861) );
  INV_X1 U21325 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18924) );
  NOR2_X1 U21326 ( .A1(n16718), .A2(n18924), .ZN(n18240) );
  AOI221_X1 U21327 ( .B1(n18244), .B2(n18243), .C1(n18242), .C2(n18241), .A(
        n18240), .ZN(n18248) );
  OAI211_X1 U21328 ( .C1(n18739), .C2(n18245), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n16718), .ZN(n18246) );
  NAND3_X1 U21329 ( .A1(n18248), .A2(n18247), .A3(n18246), .ZN(P3_U2862) );
  AOI211_X1 U21330 ( .C1(n18250), .C2(n18249), .A(n18948), .B(n21022), .ZN(
        n18787) );
  OAI21_X1 U21331 ( .B1(n18787), .B2(n18301), .A(n18260), .ZN(n18251) );
  OAI221_X1 U21332 ( .B1(n18765), .B2(n18938), .C1(n18765), .C2(n18260), .A(
        n18251), .ZN(P3_U2863) );
  NOR2_X1 U21333 ( .A1(n18938), .A2(n18252), .ZN(n18253) );
  OAI21_X1 U21334 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18253), .A(n18767), 
        .ZN(n18254) );
  AND2_X1 U21335 ( .A1(n18255), .A2(n18254), .ZN(n18259) );
  OAI221_X1 U21336 ( .B1(n18564), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18564), .C2(n18256), .A(n18260), .ZN(n18257) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18259), .B1(
        n18257), .B2(n18772), .ZN(P3_U2865) );
  INV_X1 U21338 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18262) );
  NAND2_X1 U21339 ( .A1(n18772), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18514) );
  INV_X1 U21340 ( .A(n18514), .ZN(n18563) );
  NAND2_X1 U21341 ( .A1(n18262), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18389) );
  INV_X1 U21342 ( .A(n18389), .ZN(n18437) );
  NOR2_X1 U21343 ( .A1(n18563), .A2(n18437), .ZN(n18258) );
  OAI22_X1 U21344 ( .A1(n18259), .A2(n18262), .B1(n18258), .B2(n18257), .ZN(
        P3_U2866) );
  NOR2_X1 U21345 ( .A1(n18261), .A2(n18260), .ZN(P3_U2867) );
  NOR2_X1 U21346 ( .A1(n18772), .A2(n18262), .ZN(n18265) );
  NAND2_X1 U21347 ( .A1(n18767), .A2(n18265), .ZN(n18665) );
  NOR2_X2 U21348 ( .A1(n18765), .A2(n18665), .ZN(n18714) );
  INV_X1 U21349 ( .A(n18714), .ZN(n18698) );
  NAND2_X1 U21350 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18392), .ZN(n18671) );
  NOR2_X2 U21351 ( .A1(n18666), .A2(n18263), .ZN(n18662) );
  NOR2_X1 U21352 ( .A1(n18767), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18413) );
  NAND2_X1 U21353 ( .A1(n18265), .A2(n18413), .ZN(n18629) );
  INV_X1 U21354 ( .A(n18629), .ZN(n18655) );
  NOR2_X2 U21355 ( .A1(n18459), .A2(n18264), .ZN(n18661) );
  NAND2_X1 U21356 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18265), .ZN(
        n18664) );
  NOR2_X2 U21357 ( .A1(n18765), .A2(n18664), .ZN(n18716) );
  INV_X1 U21358 ( .A(n18716), .ZN(n18678) );
  NOR2_X1 U21359 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18364) );
  NOR2_X1 U21360 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18343) );
  NAND2_X1 U21361 ( .A1(n18364), .A2(n18343), .ZN(n18354) );
  NAND2_X1 U21362 ( .A1(n18678), .A2(n18354), .ZN(n18323) );
  AND2_X1 U21363 ( .A1(n18794), .A2(n18323), .ZN(n18295) );
  AOI22_X1 U21364 ( .A1(n18662), .A2(n18655), .B1(n18661), .B2(n18295), .ZN(
        n18270) );
  NAND2_X1 U21365 ( .A1(n18767), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18388) );
  INV_X1 U21366 ( .A(n18388), .ZN(n18486) );
  NOR2_X1 U21367 ( .A1(n18413), .A2(n18486), .ZN(n18566) );
  INV_X1 U21368 ( .A(n18265), .ZN(n18589) );
  NOR2_X1 U21369 ( .A1(n18566), .A2(n18589), .ZN(n18619) );
  AOI21_X1 U21370 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18459), .ZN(n18414) );
  AOI22_X1 U21371 ( .A1(n18392), .A2(n18619), .B1(n18414), .B2(n18323), .ZN(
        n18298) );
  NAND2_X1 U21372 ( .A1(n18267), .A2(n18266), .ZN(n18296) );
  NOR2_X1 U21373 ( .A1(n18268), .A2(n18296), .ZN(n18668) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18298), .B1(
        n18361), .B2(n18668), .ZN(n18269) );
  OAI211_X1 U21375 ( .C1(n18698), .C2(n18671), .A(n18270), .B(n18269), .ZN(
        P3_U2868) );
  NOR2_X2 U21376 ( .A1(n18271), .A2(n18666), .ZN(n18673) );
  INV_X1 U21377 ( .A(n18673), .ZN(n18634) );
  AND2_X1 U21378 ( .A1(n18392), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18674) );
  AND2_X1 U21379 ( .A1(n18625), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18672) );
  AOI22_X1 U21380 ( .A1(n18655), .A2(n18674), .B1(n18295), .B2(n18672), .ZN(
        n18274) );
  NOR2_X1 U21381 ( .A1(n18272), .A2(n18296), .ZN(n18631) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18298), .B1(
        n18361), .B2(n18631), .ZN(n18273) );
  OAI211_X1 U21383 ( .C1(n18698), .C2(n18634), .A(n18274), .B(n18273), .ZN(
        P3_U2869) );
  INV_X1 U21384 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19316) );
  INV_X1 U21385 ( .A(n18680), .ZN(n18638) );
  NAND2_X1 U21386 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18392), .ZN(n18684) );
  INV_X1 U21387 ( .A(n18684), .ZN(n18635) );
  INV_X1 U21388 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n21025) );
  NOR2_X2 U21389 ( .A1(n18459), .A2(n21025), .ZN(n18679) );
  AOI22_X1 U21390 ( .A1(n18714), .A2(n18635), .B1(n18295), .B2(n18679), .ZN(
        n18276) );
  NOR2_X2 U21391 ( .A1(n9815), .A2(n18296), .ZN(n18681) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18298), .B1(
        n18361), .B2(n18681), .ZN(n18275) );
  OAI211_X1 U21393 ( .C1(n18629), .C2(n18638), .A(n18276), .B(n18275), .ZN(
        P3_U2870) );
  INV_X1 U21394 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19322) );
  NOR2_X1 U21395 ( .A1(n18666), .A2(n19322), .ZN(n18599) );
  INV_X1 U21396 ( .A(n18599), .ZN(n18690) );
  NAND2_X1 U21397 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18392), .ZN(n18603) );
  INV_X1 U21398 ( .A(n18603), .ZN(n18686) );
  NOR2_X2 U21399 ( .A1(n18459), .A2(n18277), .ZN(n18685) );
  AOI22_X1 U21400 ( .A1(n18714), .A2(n18686), .B1(n18295), .B2(n18685), .ZN(
        n18280) );
  NOR2_X2 U21401 ( .A1(n18278), .A2(n18296), .ZN(n18687) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18298), .B1(
        n18361), .B2(n18687), .ZN(n18279) );
  OAI211_X1 U21403 ( .C1(n18629), .C2(n18690), .A(n18280), .B(n18279), .ZN(
        P3_U2871) );
  NOR2_X1 U21404 ( .A1(n18666), .A2(n19328), .ZN(n18641) );
  INV_X1 U21405 ( .A(n18641), .ZN(n18697) );
  NAND2_X1 U21406 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18392), .ZN(n18644) );
  INV_X1 U21407 ( .A(n18644), .ZN(n18692) );
  NOR2_X2 U21408 ( .A1(n18459), .A2(n18281), .ZN(n18693) );
  AOI22_X1 U21409 ( .A1(n18714), .A2(n18692), .B1(n18295), .B2(n18693), .ZN(
        n18284) );
  NOR2_X2 U21410 ( .A1(n18282), .A2(n18296), .ZN(n18694) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18298), .B1(
        n18361), .B2(n18694), .ZN(n18283) );
  OAI211_X1 U21412 ( .C1(n18629), .C2(n18697), .A(n18284), .B(n18283), .ZN(
        P3_U2872) );
  NOR2_X1 U21413 ( .A1(n18666), .A2(n18285), .ZN(n18700) );
  NAND2_X1 U21414 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18392), .ZN(n18704) );
  INV_X1 U21415 ( .A(n18704), .ZN(n18645) );
  NOR2_X2 U21416 ( .A1(n18459), .A2(n18286), .ZN(n18699) );
  AOI22_X1 U21417 ( .A1(n18714), .A2(n18645), .B1(n18295), .B2(n18699), .ZN(
        n18289) );
  NOR2_X2 U21418 ( .A1(n18287), .A2(n18296), .ZN(n18701) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18298), .B1(
        n18361), .B2(n18701), .ZN(n18288) );
  OAI211_X1 U21420 ( .C1(n18629), .C2(n18648), .A(n18289), .B(n18288), .ZN(
        P3_U2873) );
  NOR2_X1 U21421 ( .A1(n14378), .A2(n18666), .ZN(n18650) );
  INV_X1 U21422 ( .A(n18650), .ZN(n18710) );
  NAND2_X1 U21423 ( .A1(n18392), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18653) );
  INV_X1 U21424 ( .A(n18653), .ZN(n18706) );
  NOR2_X2 U21425 ( .A1(n18459), .A2(n18290), .ZN(n18705) );
  AOI22_X1 U21426 ( .A1(n18655), .A2(n18706), .B1(n18295), .B2(n18705), .ZN(
        n18293) );
  NOR2_X2 U21427 ( .A1(n18291), .A2(n18296), .ZN(n18707) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18298), .B1(
        n18361), .B2(n18707), .ZN(n18292) );
  OAI211_X1 U21429 ( .C1(n18698), .C2(n18710), .A(n18293), .B(n18292), .ZN(
        P3_U2874) );
  NOR2_X1 U21430 ( .A1(n18666), .A2(n19336), .ZN(n18614) );
  INV_X1 U21431 ( .A(n18614), .ZN(n18721) );
  NAND2_X1 U21432 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18392), .ZN(n18538) );
  INV_X1 U21433 ( .A(n18538), .ZN(n18713) );
  NOR2_X2 U21434 ( .A1(n18294), .A2(n18459), .ZN(n18712) );
  AOI22_X1 U21435 ( .A1(n18655), .A2(n18713), .B1(n18295), .B2(n18712), .ZN(
        n18300) );
  NOR2_X2 U21436 ( .A1(n18297), .A2(n18296), .ZN(n18715) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18298), .B1(
        n18361), .B2(n18715), .ZN(n18299) );
  OAI211_X1 U21438 ( .C1(n18698), .C2(n18721), .A(n18300), .B(n18299), .ZN(
        P3_U2875) );
  OR2_X1 U21439 ( .A1(n18301), .A2(n18459), .ZN(n18663) );
  NOR2_X1 U21440 ( .A1(n18663), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18390) );
  INV_X1 U21441 ( .A(n18390), .ZN(n18588) );
  OAI22_X1 U21442 ( .A1(n18666), .A2(n18664), .B1(n18342), .B2(n18588), .ZN(
        n18308) );
  NAND2_X1 U21443 ( .A1(n18767), .A2(n18794), .ZN(n18485) );
  NOR2_X1 U21444 ( .A1(n18342), .A2(n18485), .ZN(n18319) );
  AOI22_X1 U21445 ( .A1(n18620), .A2(n18655), .B1(n18661), .B2(n18319), .ZN(
        n18303) );
  NAND2_X1 U21446 ( .A1(n18343), .A2(n18486), .ZN(n18382) );
  AOI22_X1 U21447 ( .A1(n18716), .A2(n18662), .B1(n18668), .B2(n18384), .ZN(
        n18302) );
  OAI211_X1 U21448 ( .C1(n18304), .C2(n18308), .A(n18303), .B(n18302), .ZN(
        P3_U2876) );
  INV_X1 U21449 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18307) );
  AOI22_X1 U21450 ( .A1(n18655), .A2(n18673), .B1(n18672), .B2(n18319), .ZN(
        n18306) );
  AOI22_X1 U21451 ( .A1(n18716), .A2(n18674), .B1(n18631), .B2(n18384), .ZN(
        n18305) );
  OAI211_X1 U21452 ( .C1(n18307), .C2(n18308), .A(n18306), .B(n18305), .ZN(
        P3_U2877) );
  AOI22_X1 U21453 ( .A1(n18655), .A2(n18635), .B1(n18679), .B2(n18319), .ZN(
        n18310) );
  INV_X1 U21454 ( .A(n18308), .ZN(n18320) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18320), .B1(
        n18681), .B2(n18384), .ZN(n18309) );
  OAI211_X1 U21456 ( .C1(n18678), .C2(n18638), .A(n18310), .B(n18309), .ZN(
        P3_U2878) );
  AOI22_X1 U21457 ( .A1(n18716), .A2(n18599), .B1(n18685), .B2(n18319), .ZN(
        n18312) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18320), .B1(
        n18687), .B2(n18384), .ZN(n18311) );
  OAI211_X1 U21459 ( .C1(n18629), .C2(n18603), .A(n18312), .B(n18311), .ZN(
        P3_U2879) );
  AOI22_X1 U21460 ( .A1(n18716), .A2(n18641), .B1(n18693), .B2(n18319), .ZN(
        n18314) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18320), .B1(
        n18694), .B2(n18384), .ZN(n18313) );
  OAI211_X1 U21462 ( .C1(n18629), .C2(n18644), .A(n18314), .B(n18313), .ZN(
        P3_U2880) );
  AOI22_X1 U21463 ( .A1(n18655), .A2(n18645), .B1(n18699), .B2(n18319), .ZN(
        n18316) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18320), .B1(
        n18701), .B2(n18384), .ZN(n18315) );
  OAI211_X1 U21465 ( .C1(n18678), .C2(n18648), .A(n18316), .B(n18315), .ZN(
        P3_U2881) );
  AOI22_X1 U21466 ( .A1(n18716), .A2(n18706), .B1(n18705), .B2(n18319), .ZN(
        n18318) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18320), .B1(
        n18707), .B2(n18384), .ZN(n18317) );
  OAI211_X1 U21468 ( .C1(n18629), .C2(n18710), .A(n18318), .B(n18317), .ZN(
        P3_U2882) );
  AOI22_X1 U21469 ( .A1(n18716), .A2(n18713), .B1(n18712), .B2(n18319), .ZN(
        n18322) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18320), .B1(
        n18715), .B2(n18384), .ZN(n18321) );
  OAI211_X1 U21471 ( .C1(n18629), .C2(n18721), .A(n18322), .B(n18321), .ZN(
        P3_U2883) );
  INV_X1 U21472 ( .A(n18668), .ZN(n18630) );
  INV_X1 U21473 ( .A(n18413), .ZN(n18513) );
  NOR2_X2 U21474 ( .A1(n18342), .A2(n18513), .ZN(n18409) );
  NAND2_X1 U21475 ( .A1(n18382), .A2(n18407), .ZN(n18365) );
  AND2_X1 U21476 ( .A1(n18794), .A2(n18365), .ZN(n18338) );
  AOI22_X1 U21477 ( .A1(n18620), .A2(n18716), .B1(n18661), .B2(n18338), .ZN(
        n18325) );
  OAI221_X1 U21478 ( .B1(n18365), .B2(n18564), .C1(n18365), .C2(n18323), .A(
        n18414), .ZN(n18339) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18339), .B1(
        n18361), .B2(n18662), .ZN(n18324) );
  OAI211_X1 U21480 ( .C1(n18630), .C2(n18407), .A(n18325), .B(n18324), .ZN(
        P3_U2884) );
  AOI22_X1 U21481 ( .A1(n18361), .A2(n18674), .B1(n18672), .B2(n18338), .ZN(
        n18327) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18339), .B1(
        n18631), .B2(n18409), .ZN(n18326) );
  OAI211_X1 U21483 ( .C1(n18678), .C2(n18634), .A(n18327), .B(n18326), .ZN(
        P3_U2885) );
  AOI22_X1 U21484 ( .A1(n18716), .A2(n18635), .B1(n18679), .B2(n18338), .ZN(
        n18329) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18339), .B1(
        n18681), .B2(n18409), .ZN(n18328) );
  OAI211_X1 U21486 ( .C1(n18354), .C2(n18638), .A(n18329), .B(n18328), .ZN(
        P3_U2886) );
  AOI22_X1 U21487 ( .A1(n18361), .A2(n18599), .B1(n18685), .B2(n18338), .ZN(
        n18331) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18339), .B1(
        n18687), .B2(n18409), .ZN(n18330) );
  OAI211_X1 U21489 ( .C1(n18678), .C2(n18603), .A(n18331), .B(n18330), .ZN(
        P3_U2887) );
  AOI22_X1 U21490 ( .A1(n18716), .A2(n18692), .B1(n18693), .B2(n18338), .ZN(
        n18333) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18339), .B1(
        n18694), .B2(n18409), .ZN(n18332) );
  OAI211_X1 U21492 ( .C1(n18354), .C2(n18697), .A(n18333), .B(n18332), .ZN(
        P3_U2888) );
  AOI22_X1 U21493 ( .A1(n18716), .A2(n18645), .B1(n18699), .B2(n18338), .ZN(
        n18335) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18339), .B1(
        n18701), .B2(n18409), .ZN(n18334) );
  OAI211_X1 U21495 ( .C1(n18354), .C2(n18648), .A(n18335), .B(n18334), .ZN(
        P3_U2889) );
  AOI22_X1 U21496 ( .A1(n18716), .A2(n18650), .B1(n18705), .B2(n18338), .ZN(
        n18337) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18339), .B1(
        n18707), .B2(n18409), .ZN(n18336) );
  OAI211_X1 U21498 ( .C1(n18354), .C2(n18653), .A(n18337), .B(n18336), .ZN(
        P3_U2890) );
  AOI22_X1 U21499 ( .A1(n18716), .A2(n18614), .B1(n18712), .B2(n18338), .ZN(
        n18341) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18339), .B1(
        n18715), .B2(n18409), .ZN(n18340) );
  OAI211_X1 U21501 ( .C1(n18354), .C2(n18538), .A(n18341), .B(n18340), .ZN(
        P3_U2891) );
  NOR2_X1 U21502 ( .A1(n18767), .A2(n18342), .ZN(n18391) );
  NAND2_X1 U21503 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18391), .ZN(
        n18435) );
  AND2_X1 U21504 ( .A1(n18794), .A2(n18391), .ZN(n18359) );
  AOI22_X1 U21505 ( .A1(n18620), .A2(n18361), .B1(n18661), .B2(n18359), .ZN(
        n18345) );
  AOI21_X1 U21506 ( .B1(n18767), .B2(n18622), .A(n18459), .ZN(n18436) );
  OAI211_X1 U21507 ( .C1(n18420), .C2(n18626), .A(n18343), .B(n18436), .ZN(
        n18360) );
  AOI22_X1 U21508 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18360), .B1(
        n18662), .B2(n18384), .ZN(n18344) );
  OAI211_X1 U21509 ( .C1(n18630), .C2(n18435), .A(n18345), .B(n18344), .ZN(
        P3_U2892) );
  AOI22_X1 U21510 ( .A1(n18361), .A2(n18673), .B1(n18672), .B2(n18359), .ZN(
        n18347) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18360), .B1(
        n18674), .B2(n18384), .ZN(n18346) );
  OAI211_X1 U21512 ( .C1(n18677), .C2(n18435), .A(n18347), .B(n18346), .ZN(
        P3_U2893) );
  AOI22_X1 U21513 ( .A1(n18680), .A2(n18384), .B1(n18679), .B2(n18359), .ZN(
        n18349) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18360), .B1(
        n18681), .B2(n18420), .ZN(n18348) );
  OAI211_X1 U21515 ( .C1(n18354), .C2(n18684), .A(n18349), .B(n18348), .ZN(
        P3_U2894) );
  AOI22_X1 U21516 ( .A1(n18599), .A2(n18384), .B1(n18685), .B2(n18359), .ZN(
        n18351) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18360), .B1(
        n18687), .B2(n18420), .ZN(n18350) );
  OAI211_X1 U21518 ( .C1(n18354), .C2(n18603), .A(n18351), .B(n18350), .ZN(
        P3_U2895) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18360), .B1(
        n18693), .B2(n18359), .ZN(n18353) );
  AOI22_X1 U21520 ( .A1(n18641), .A2(n18384), .B1(n18694), .B2(n18420), .ZN(
        n18352) );
  OAI211_X1 U21521 ( .C1(n18354), .C2(n18644), .A(n18353), .B(n18352), .ZN(
        P3_U2896) );
  AOI22_X1 U21522 ( .A1(n18361), .A2(n18645), .B1(n18699), .B2(n18359), .ZN(
        n18356) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18360), .B1(
        n18701), .B2(n18420), .ZN(n18355) );
  OAI211_X1 U21524 ( .C1(n18648), .C2(n18382), .A(n18356), .B(n18355), .ZN(
        P3_U2897) );
  AOI22_X1 U21525 ( .A1(n18361), .A2(n18650), .B1(n18705), .B2(n18359), .ZN(
        n18358) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18360), .B1(
        n18707), .B2(n18420), .ZN(n18357) );
  OAI211_X1 U21527 ( .C1(n18653), .C2(n18382), .A(n18358), .B(n18357), .ZN(
        P3_U2898) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18360), .B1(
        n18712), .B2(n18359), .ZN(n18363) );
  AOI22_X1 U21529 ( .A1(n18361), .A2(n18614), .B1(n18715), .B2(n18420), .ZN(
        n18362) );
  OAI211_X1 U21530 ( .C1(n18538), .C2(n18382), .A(n18363), .B(n18362), .ZN(
        P3_U2899) );
  INV_X1 U21531 ( .A(n18364), .ZN(n18768) );
  NOR2_X2 U21532 ( .A1(n18768), .A2(n18389), .ZN(n18450) );
  OAI221_X1 U21533 ( .B1(n18420), .B2(n18564), .C1(n18420), .C2(n18365), .A(
        n18626), .ZN(n18366) );
  AOI21_X1 U21534 ( .B1(n18457), .B2(n18366), .A(n18459), .ZN(n18369) );
  AOI21_X1 U21535 ( .B1(n18435), .B2(n18457), .A(n18660), .ZN(n18383) );
  AOI22_X1 U21536 ( .A1(n18620), .A2(n18384), .B1(n18661), .B2(n18383), .ZN(
        n18368) );
  AOI22_X1 U21537 ( .A1(n18668), .A2(n18450), .B1(n18662), .B2(n18409), .ZN(
        n18367) );
  OAI211_X1 U21538 ( .C1(n18369), .C2(n21045), .A(n18368), .B(n18367), .ZN(
        P3_U2900) );
  AOI22_X1 U21539 ( .A1(n18673), .A2(n18384), .B1(n18672), .B2(n18383), .ZN(
        n18371) );
  INV_X1 U21540 ( .A(n18369), .ZN(n18385) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18385), .B1(
        n18674), .B2(n18409), .ZN(n18370) );
  OAI211_X1 U21542 ( .C1(n18677), .C2(n18457), .A(n18371), .B(n18370), .ZN(
        P3_U2901) );
  AOI22_X1 U21543 ( .A1(n18680), .A2(n18409), .B1(n18679), .B2(n18383), .ZN(
        n18373) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18385), .B1(
        n18681), .B2(n18450), .ZN(n18372) );
  OAI211_X1 U21545 ( .C1(n18684), .C2(n18382), .A(n18373), .B(n18372), .ZN(
        P3_U2902) );
  AOI22_X1 U21546 ( .A1(n18686), .A2(n18384), .B1(n18685), .B2(n18383), .ZN(
        n18375) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18385), .B1(
        n18687), .B2(n18450), .ZN(n18374) );
  OAI211_X1 U21548 ( .C1(n18690), .C2(n18407), .A(n18375), .B(n18374), .ZN(
        P3_U2903) );
  AOI22_X1 U21549 ( .A1(n18693), .A2(n18383), .B1(n18692), .B2(n18384), .ZN(
        n18377) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18385), .B1(
        n18694), .B2(n18450), .ZN(n18376) );
  OAI211_X1 U21551 ( .C1(n18697), .C2(n18407), .A(n18377), .B(n18376), .ZN(
        P3_U2904) );
  AOI22_X1 U21552 ( .A1(n18700), .A2(n18409), .B1(n18699), .B2(n18383), .ZN(
        n18379) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18385), .B1(
        n18701), .B2(n18450), .ZN(n18378) );
  OAI211_X1 U21554 ( .C1(n18704), .C2(n18382), .A(n18379), .B(n18378), .ZN(
        P3_U2905) );
  AOI22_X1 U21555 ( .A1(n18705), .A2(n18383), .B1(n18706), .B2(n18409), .ZN(
        n18381) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18385), .B1(
        n18707), .B2(n18450), .ZN(n18380) );
  OAI211_X1 U21557 ( .C1(n18710), .C2(n18382), .A(n18381), .B(n18380), .ZN(
        P3_U2906) );
  AOI22_X1 U21558 ( .A1(n18614), .A2(n18384), .B1(n18712), .B2(n18383), .ZN(
        n18387) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18385), .B1(
        n18715), .B2(n18450), .ZN(n18386) );
  OAI211_X1 U21560 ( .C1(n18538), .C2(n18407), .A(n18387), .B(n18386), .ZN(
        P3_U2907) );
  NOR2_X2 U21561 ( .A1(n18389), .A2(n18388), .ZN(n18479) );
  INV_X1 U21562 ( .A(n18479), .ZN(n18475) );
  NOR2_X1 U21563 ( .A1(n18389), .A2(n18485), .ZN(n18408) );
  AOI22_X1 U21564 ( .A1(n18662), .A2(n18420), .B1(n18661), .B2(n18408), .ZN(
        n18394) );
  AOI22_X1 U21565 ( .A1(n18392), .A2(n18391), .B1(n18437), .B2(n18390), .ZN(
        n18410) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18410), .B1(
        n18620), .B2(n18409), .ZN(n18393) );
  OAI211_X1 U21567 ( .C1(n18630), .C2(n18475), .A(n18394), .B(n18393), .ZN(
        P3_U2908) );
  AOI22_X1 U21568 ( .A1(n18673), .A2(n18409), .B1(n18672), .B2(n18408), .ZN(
        n18396) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18410), .B1(
        n18674), .B2(n18420), .ZN(n18395) );
  OAI211_X1 U21570 ( .C1(n18677), .C2(n18475), .A(n18396), .B(n18395), .ZN(
        P3_U2909) );
  AOI22_X1 U21571 ( .A1(n18680), .A2(n18420), .B1(n18679), .B2(n18408), .ZN(
        n18398) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18410), .B1(
        n18681), .B2(n18479), .ZN(n18397) );
  OAI211_X1 U21573 ( .C1(n18684), .C2(n18407), .A(n18398), .B(n18397), .ZN(
        P3_U2910) );
  AOI22_X1 U21574 ( .A1(n18686), .A2(n18409), .B1(n18685), .B2(n18408), .ZN(
        n18400) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18410), .B1(
        n18687), .B2(n18479), .ZN(n18399) );
  OAI211_X1 U21576 ( .C1(n18690), .C2(n18435), .A(n18400), .B(n18399), .ZN(
        P3_U2911) );
  AOI22_X1 U21577 ( .A1(n18641), .A2(n18420), .B1(n18693), .B2(n18408), .ZN(
        n18402) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18410), .B1(
        n18694), .B2(n18479), .ZN(n18401) );
  OAI211_X1 U21579 ( .C1(n18644), .C2(n18407), .A(n18402), .B(n18401), .ZN(
        P3_U2912) );
  AOI22_X1 U21580 ( .A1(n18645), .A2(n18409), .B1(n18699), .B2(n18408), .ZN(
        n18404) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18410), .B1(
        n18701), .B2(n18479), .ZN(n18403) );
  OAI211_X1 U21582 ( .C1(n18648), .C2(n18435), .A(n18404), .B(n18403), .ZN(
        P3_U2913) );
  AOI22_X1 U21583 ( .A1(n18705), .A2(n18408), .B1(n18706), .B2(n18420), .ZN(
        n18406) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18410), .B1(
        n18707), .B2(n18479), .ZN(n18405) );
  OAI211_X1 U21585 ( .C1(n18710), .C2(n18407), .A(n18406), .B(n18405), .ZN(
        P3_U2914) );
  AOI22_X1 U21586 ( .A1(n18614), .A2(n18409), .B1(n18712), .B2(n18408), .ZN(
        n18412) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18410), .B1(
        n18715), .B2(n18479), .ZN(n18411) );
  OAI211_X1 U21588 ( .C1(n18538), .C2(n18435), .A(n18412), .B(n18411), .ZN(
        P3_U2915) );
  NAND2_X1 U21589 ( .A1(n18437), .A2(n18413), .ZN(n18483) );
  NAND2_X1 U21590 ( .A1(n18475), .A2(n18483), .ZN(n18458) );
  AND2_X1 U21591 ( .A1(n18794), .A2(n18458), .ZN(n18431) );
  AOI22_X1 U21592 ( .A1(n18662), .A2(n18450), .B1(n18661), .B2(n18431), .ZN(
        n18417) );
  NAND2_X1 U21593 ( .A1(n18435), .A2(n18457), .ZN(n18415) );
  OAI221_X1 U21594 ( .B1(n18458), .B2(n18564), .C1(n18458), .C2(n18415), .A(
        n18414), .ZN(n18432) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18432), .B1(
        n18668), .B2(n18508), .ZN(n18416) );
  OAI211_X1 U21596 ( .C1(n18671), .C2(n18435), .A(n18417), .B(n18416), .ZN(
        P3_U2916) );
  AOI22_X1 U21597 ( .A1(n18673), .A2(n18420), .B1(n18672), .B2(n18431), .ZN(
        n18419) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18432), .B1(
        n18674), .B2(n18450), .ZN(n18418) );
  OAI211_X1 U21599 ( .C1(n18677), .C2(n18483), .A(n18419), .B(n18418), .ZN(
        P3_U2917) );
  AOI22_X1 U21600 ( .A1(n18679), .A2(n18431), .B1(n18635), .B2(n18420), .ZN(
        n18422) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18432), .B1(
        n18681), .B2(n18508), .ZN(n18421) );
  OAI211_X1 U21602 ( .C1(n18638), .C2(n18457), .A(n18422), .B(n18421), .ZN(
        P3_U2918) );
  AOI22_X1 U21603 ( .A1(n18599), .A2(n18450), .B1(n18685), .B2(n18431), .ZN(
        n18424) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18432), .B1(
        n18687), .B2(n18508), .ZN(n18423) );
  OAI211_X1 U21605 ( .C1(n18603), .C2(n18435), .A(n18424), .B(n18423), .ZN(
        P3_U2919) );
  AOI22_X1 U21606 ( .A1(n18641), .A2(n18450), .B1(n18693), .B2(n18431), .ZN(
        n18426) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18432), .B1(
        n18694), .B2(n18508), .ZN(n18425) );
  OAI211_X1 U21608 ( .C1(n18644), .C2(n18435), .A(n18426), .B(n18425), .ZN(
        P3_U2920) );
  AOI22_X1 U21609 ( .A1(n18700), .A2(n18450), .B1(n18699), .B2(n18431), .ZN(
        n18428) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18432), .B1(
        n18701), .B2(n18508), .ZN(n18427) );
  OAI211_X1 U21611 ( .C1(n18704), .C2(n18435), .A(n18428), .B(n18427), .ZN(
        P3_U2921) );
  AOI22_X1 U21612 ( .A1(n18705), .A2(n18431), .B1(n18706), .B2(n18450), .ZN(
        n18430) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18432), .B1(
        n18707), .B2(n18508), .ZN(n18429) );
  OAI211_X1 U21614 ( .C1(n18710), .C2(n18435), .A(n18430), .B(n18429), .ZN(
        P3_U2922) );
  AOI22_X1 U21615 ( .A1(n18713), .A2(n18450), .B1(n18712), .B2(n18431), .ZN(
        n18434) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18432), .B1(
        n18715), .B2(n18508), .ZN(n18433) );
  OAI211_X1 U21617 ( .C1(n18721), .C2(n18435), .A(n18434), .B(n18433), .ZN(
        P3_U2923) );
  NAND2_X1 U21618 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18437), .ZN(
        n18484) );
  INV_X1 U21619 ( .A(n18527), .ZN(n18530) );
  OAI211_X1 U21620 ( .C1(n18530), .C2(n18626), .A(n18437), .B(n18436), .ZN(
        n18454) );
  NOR2_X1 U21621 ( .A1(n18660), .A2(n18484), .ZN(n18453) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18454), .B1(
        n18661), .B2(n18453), .ZN(n18439) );
  AOI22_X1 U21623 ( .A1(n18668), .A2(n18530), .B1(n18662), .B2(n18479), .ZN(
        n18438) );
  OAI211_X1 U21624 ( .C1(n18671), .C2(n18457), .A(n18439), .B(n18438), .ZN(
        P3_U2924) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18454), .B1(
        n18672), .B2(n18453), .ZN(n18441) );
  AOI22_X1 U21626 ( .A1(n18631), .A2(n18530), .B1(n18674), .B2(n18479), .ZN(
        n18440) );
  OAI211_X1 U21627 ( .C1(n18634), .C2(n18457), .A(n18441), .B(n18440), .ZN(
        P3_U2925) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18454), .B1(
        n18679), .B2(n18453), .ZN(n18443) );
  AOI22_X1 U21629 ( .A1(n18680), .A2(n18479), .B1(n18681), .B2(n18530), .ZN(
        n18442) );
  OAI211_X1 U21630 ( .C1(n18684), .C2(n18457), .A(n18443), .B(n18442), .ZN(
        P3_U2926) );
  AOI22_X1 U21631 ( .A1(n18686), .A2(n18450), .B1(n18685), .B2(n18453), .ZN(
        n18445) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18454), .B1(
        n18687), .B2(n18530), .ZN(n18444) );
  OAI211_X1 U21633 ( .C1(n18690), .C2(n18475), .A(n18445), .B(n18444), .ZN(
        P3_U2927) );
  AOI22_X1 U21634 ( .A1(n18693), .A2(n18453), .B1(n18692), .B2(n18450), .ZN(
        n18447) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18454), .B1(
        n18694), .B2(n18530), .ZN(n18446) );
  OAI211_X1 U21636 ( .C1(n18697), .C2(n18475), .A(n18447), .B(n18446), .ZN(
        P3_U2928) );
  AOI22_X1 U21637 ( .A1(n18645), .A2(n18450), .B1(n18699), .B2(n18453), .ZN(
        n18449) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18454), .B1(
        n18701), .B2(n18530), .ZN(n18448) );
  OAI211_X1 U21639 ( .C1(n18648), .C2(n18475), .A(n18449), .B(n18448), .ZN(
        P3_U2929) );
  AOI22_X1 U21640 ( .A1(n18650), .A2(n18450), .B1(n18705), .B2(n18453), .ZN(
        n18452) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18454), .B1(
        n18707), .B2(n18530), .ZN(n18451) );
  OAI211_X1 U21642 ( .C1(n18653), .C2(n18475), .A(n18452), .B(n18451), .ZN(
        P3_U2930) );
  AOI22_X1 U21643 ( .A1(n18713), .A2(n18479), .B1(n18712), .B2(n18453), .ZN(
        n18456) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18454), .B1(
        n18715), .B2(n18530), .ZN(n18455) );
  OAI211_X1 U21645 ( .C1(n18721), .C2(n18457), .A(n18456), .B(n18455), .ZN(
        P3_U2931) );
  NOR2_X2 U21646 ( .A1(n18768), .A2(n18514), .ZN(n18558) );
  OAI221_X1 U21647 ( .B1(n18530), .B2(n18564), .C1(n18534), .C2(n18458), .A(
        n18626), .ZN(n18460) );
  AOI21_X1 U21648 ( .B1(n18553), .B2(n18460), .A(n18459), .ZN(n18464) );
  AOI21_X1 U21649 ( .B1(n18527), .B2(n18553), .A(n18660), .ZN(n18478) );
  AOI22_X1 U21650 ( .A1(n18620), .A2(n18479), .B1(n18661), .B2(n18478), .ZN(
        n18462) );
  AOI22_X1 U21651 ( .A1(n18668), .A2(n18558), .B1(n18662), .B2(n18508), .ZN(
        n18461) );
  OAI211_X1 U21652 ( .C1(n18464), .C2(n18463), .A(n18462), .B(n18461), .ZN(
        P3_U2932) );
  AOI22_X1 U21653 ( .A1(n18674), .A2(n18508), .B1(n18672), .B2(n18478), .ZN(
        n18466) );
  INV_X1 U21654 ( .A(n18464), .ZN(n18480) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18480), .B1(
        n18631), .B2(n18558), .ZN(n18465) );
  OAI211_X1 U21656 ( .C1(n18634), .C2(n18475), .A(n18466), .B(n18465), .ZN(
        P3_U2933) );
  AOI22_X1 U21657 ( .A1(n18680), .A2(n18508), .B1(n18679), .B2(n18478), .ZN(
        n18468) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18480), .B1(
        n18681), .B2(n18558), .ZN(n18467) );
  OAI211_X1 U21659 ( .C1(n18684), .C2(n18475), .A(n18468), .B(n18467), .ZN(
        P3_U2934) );
  AOI22_X1 U21660 ( .A1(n18599), .A2(n18508), .B1(n18685), .B2(n18478), .ZN(
        n18470) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18480), .B1(
        n18687), .B2(n18558), .ZN(n18469) );
  OAI211_X1 U21662 ( .C1(n18603), .C2(n18475), .A(n18470), .B(n18469), .ZN(
        P3_U2935) );
  AOI22_X1 U21663 ( .A1(n18641), .A2(n18508), .B1(n18693), .B2(n18478), .ZN(
        n18472) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18480), .B1(
        n18694), .B2(n18558), .ZN(n18471) );
  OAI211_X1 U21665 ( .C1(n18644), .C2(n18475), .A(n18472), .B(n18471), .ZN(
        P3_U2936) );
  AOI22_X1 U21666 ( .A1(n18700), .A2(n18508), .B1(n18699), .B2(n18478), .ZN(
        n18474) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18480), .B1(
        n18701), .B2(n18558), .ZN(n18473) );
  OAI211_X1 U21668 ( .C1(n18704), .C2(n18475), .A(n18474), .B(n18473), .ZN(
        P3_U2937) );
  AOI22_X1 U21669 ( .A1(n18650), .A2(n18479), .B1(n18705), .B2(n18478), .ZN(
        n18477) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18480), .B1(
        n18707), .B2(n18558), .ZN(n18476) );
  OAI211_X1 U21671 ( .C1(n18653), .C2(n18483), .A(n18477), .B(n18476), .ZN(
        P3_U2938) );
  AOI22_X1 U21672 ( .A1(n18614), .A2(n18479), .B1(n18712), .B2(n18478), .ZN(
        n18482) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18480), .B1(
        n18715), .B2(n18558), .ZN(n18481) );
  OAI211_X1 U21674 ( .C1(n18538), .C2(n18483), .A(n18482), .B(n18481), .ZN(
        P3_U2939) );
  NAND2_X1 U21675 ( .A1(n18563), .A2(n18767), .ZN(n18539) );
  OAI22_X1 U21676 ( .A1(n18666), .A2(n18484), .B1(n18663), .B2(n18539), .ZN(
        n18509) );
  NOR2_X1 U21677 ( .A1(n18514), .A2(n18485), .ZN(n18507) );
  AOI22_X1 U21678 ( .A1(n18662), .A2(n18534), .B1(n18661), .B2(n18507), .ZN(
        n18488) );
  NAND2_X1 U21679 ( .A1(n18563), .A2(n18486), .ZN(n18587) );
  AOI22_X1 U21680 ( .A1(n18620), .A2(n18508), .B1(n18668), .B2(n18576), .ZN(
        n18487) );
  OAI211_X1 U21681 ( .C1(n18489), .C2(n18509), .A(n18488), .B(n18487), .ZN(
        P3_U2940) );
  AOI22_X1 U21682 ( .A1(n18673), .A2(n18508), .B1(n18672), .B2(n18507), .ZN(
        n18491) );
  AOI22_X1 U21683 ( .A1(n18631), .A2(n18576), .B1(n18674), .B2(n18530), .ZN(
        n18490) );
  OAI211_X1 U21684 ( .C1(n20981), .C2(n18509), .A(n18491), .B(n18490), .ZN(
        P3_U2941) );
  AOI22_X1 U21685 ( .A1(n18680), .A2(n18534), .B1(n18679), .B2(n18507), .ZN(
        n18493) );
  AOI22_X1 U21686 ( .A1(n18681), .A2(n18576), .B1(n18635), .B2(n18508), .ZN(
        n18492) );
  OAI211_X1 U21687 ( .C1(n18494), .C2(n18509), .A(n18493), .B(n18492), .ZN(
        P3_U2942) );
  AOI22_X1 U21688 ( .A1(n18599), .A2(n18534), .B1(n18685), .B2(n18507), .ZN(
        n18496) );
  AOI22_X1 U21689 ( .A1(n18687), .A2(n18576), .B1(n18686), .B2(n18508), .ZN(
        n18495) );
  OAI211_X1 U21690 ( .C1(n18497), .C2(n18509), .A(n18496), .B(n18495), .ZN(
        P3_U2943) );
  AOI22_X1 U21691 ( .A1(n18641), .A2(n18534), .B1(n18693), .B2(n18507), .ZN(
        n18499) );
  AOI22_X1 U21692 ( .A1(n18694), .A2(n18576), .B1(n18692), .B2(n18508), .ZN(
        n18498) );
  OAI211_X1 U21693 ( .C1(n18500), .C2(n18509), .A(n18499), .B(n18498), .ZN(
        P3_U2944) );
  AOI22_X1 U21694 ( .A1(n18645), .A2(n18508), .B1(n18699), .B2(n18507), .ZN(
        n18502) );
  AOI22_X1 U21695 ( .A1(n18700), .A2(n18530), .B1(n18701), .B2(n18576), .ZN(
        n18501) );
  OAI211_X1 U21696 ( .C1(n18503), .C2(n18509), .A(n18502), .B(n18501), .ZN(
        P3_U2945) );
  AOI22_X1 U21697 ( .A1(n18705), .A2(n18507), .B1(n18706), .B2(n18530), .ZN(
        n18505) );
  AOI22_X1 U21698 ( .A1(n18650), .A2(n18508), .B1(n18707), .B2(n18576), .ZN(
        n18504) );
  OAI211_X1 U21699 ( .C1(n18506), .C2(n18509), .A(n18505), .B(n18504), .ZN(
        P3_U2946) );
  AOI22_X1 U21700 ( .A1(n18614), .A2(n18508), .B1(n18712), .B2(n18507), .ZN(
        n18512) );
  INV_X1 U21701 ( .A(n18509), .ZN(n18510) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18510), .B1(
        n18715), .B2(n18576), .ZN(n18511) );
  OAI211_X1 U21703 ( .C1(n18538), .C2(n18527), .A(n18512), .B(n18511), .ZN(
        P3_U2947) );
  INV_X1 U21704 ( .A(n18613), .ZN(n18602) );
  AOI21_X1 U21705 ( .B1(n18587), .B2(n18602), .A(n18660), .ZN(n18533) );
  AOI22_X1 U21706 ( .A1(n18620), .A2(n18534), .B1(n18661), .B2(n18533), .ZN(
        n18518) );
  NOR2_X1 U21707 ( .A1(n18530), .A2(n18558), .ZN(n18515) );
  OAI211_X1 U21708 ( .C1(n18515), .C2(n18622), .A(n18587), .B(n18602), .ZN(
        n18516) );
  OAI211_X1 U21709 ( .C1(n18613), .C2(n18626), .A(n18625), .B(n18516), .ZN(
        n18535) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18535), .B1(
        n18662), .B2(n18558), .ZN(n18517) );
  OAI211_X1 U21711 ( .C1(n18630), .C2(n18602), .A(n18518), .B(n18517), .ZN(
        P3_U2948) );
  AOI22_X1 U21712 ( .A1(n18673), .A2(n18534), .B1(n18672), .B2(n18533), .ZN(
        n18520) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18535), .B1(
        n18674), .B2(n18558), .ZN(n18519) );
  OAI211_X1 U21714 ( .C1(n18677), .C2(n18602), .A(n18520), .B(n18519), .ZN(
        P3_U2949) );
  AOI22_X1 U21715 ( .A1(n18680), .A2(n18558), .B1(n18679), .B2(n18533), .ZN(
        n18522) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18535), .B1(
        n18681), .B2(n18613), .ZN(n18521) );
  OAI211_X1 U21717 ( .C1(n18684), .C2(n18527), .A(n18522), .B(n18521), .ZN(
        P3_U2950) );
  AOI22_X1 U21718 ( .A1(n18686), .A2(n18534), .B1(n18685), .B2(n18533), .ZN(
        n18524) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18535), .B1(
        n18687), .B2(n18613), .ZN(n18523) );
  OAI211_X1 U21720 ( .C1(n18690), .C2(n18553), .A(n18524), .B(n18523), .ZN(
        P3_U2951) );
  AOI22_X1 U21721 ( .A1(n18641), .A2(n18558), .B1(n18693), .B2(n18533), .ZN(
        n18526) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18535), .B1(
        n18694), .B2(n18613), .ZN(n18525) );
  OAI211_X1 U21723 ( .C1(n18644), .C2(n18527), .A(n18526), .B(n18525), .ZN(
        P3_U2952) );
  AOI22_X1 U21724 ( .A1(n18645), .A2(n18534), .B1(n18699), .B2(n18533), .ZN(
        n18529) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18535), .B1(
        n18701), .B2(n18613), .ZN(n18528) );
  OAI211_X1 U21726 ( .C1(n18648), .C2(n18553), .A(n18529), .B(n18528), .ZN(
        P3_U2953) );
  AOI22_X1 U21727 ( .A1(n18650), .A2(n18530), .B1(n18705), .B2(n18533), .ZN(
        n18532) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18535), .B1(
        n18707), .B2(n18613), .ZN(n18531) );
  OAI211_X1 U21729 ( .C1(n18653), .C2(n18553), .A(n18532), .B(n18531), .ZN(
        P3_U2954) );
  AOI22_X1 U21730 ( .A1(n18614), .A2(n18534), .B1(n18712), .B2(n18533), .ZN(
        n18537) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18535), .B1(
        n18715), .B2(n18613), .ZN(n18536) );
  OAI211_X1 U21732 ( .C1(n18538), .C2(n18553), .A(n18537), .B(n18536), .ZN(
        P3_U2955) );
  NAND2_X1 U21733 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18563), .ZN(
        n18590) );
  OAI22_X1 U21734 ( .A1(n18666), .A2(n18539), .B1(n18663), .B2(n18590), .ZN(
        n18561) );
  NOR2_X1 U21735 ( .A1(n18660), .A2(n18590), .ZN(n18557) );
  AOI22_X1 U21736 ( .A1(n18620), .A2(n18558), .B1(n18661), .B2(n18557), .ZN(
        n18541) );
  NOR2_X2 U21737 ( .A1(n18765), .A2(n18590), .ZN(n18649) );
  AOI22_X1 U21738 ( .A1(n18668), .A2(n18649), .B1(n18662), .B2(n18576), .ZN(
        n18540) );
  OAI211_X1 U21739 ( .C1(n18542), .C2(n18561), .A(n18541), .B(n18540), .ZN(
        P3_U2956) );
  INV_X1 U21740 ( .A(n18649), .ZN(n18659) );
  AOI22_X1 U21741 ( .A1(n18673), .A2(n18558), .B1(n18672), .B2(n18557), .ZN(
        n18544) );
  INV_X1 U21742 ( .A(n18561), .ZN(n18554) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18554), .B1(
        n18674), .B2(n18576), .ZN(n18543) );
  OAI211_X1 U21744 ( .C1(n18677), .C2(n18659), .A(n18544), .B(n18543), .ZN(
        P3_U2957) );
  AOI22_X1 U21745 ( .A1(n18680), .A2(n18576), .B1(n18679), .B2(n18557), .ZN(
        n18546) );
  AOI22_X1 U21746 ( .A1(n18681), .A2(n18649), .B1(n18635), .B2(n18558), .ZN(
        n18545) );
  OAI211_X1 U21747 ( .C1(n21093), .C2(n18561), .A(n18546), .B(n18545), .ZN(
        P3_U2958) );
  AOI22_X1 U21748 ( .A1(n18599), .A2(n18576), .B1(n18685), .B2(n18557), .ZN(
        n18548) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18554), .B1(
        n18687), .B2(n18649), .ZN(n18547) );
  OAI211_X1 U21750 ( .C1(n18603), .C2(n18553), .A(n18548), .B(n18547), .ZN(
        P3_U2959) );
  AOI22_X1 U21751 ( .A1(n18641), .A2(n18576), .B1(n18693), .B2(n18557), .ZN(
        n18550) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18554), .B1(
        n18694), .B2(n18649), .ZN(n18549) );
  OAI211_X1 U21753 ( .C1(n18644), .C2(n18553), .A(n18550), .B(n18549), .ZN(
        P3_U2960) );
  AOI22_X1 U21754 ( .A1(n18700), .A2(n18576), .B1(n18699), .B2(n18557), .ZN(
        n18552) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18554), .B1(
        n18701), .B2(n18649), .ZN(n18551) );
  OAI211_X1 U21756 ( .C1(n18704), .C2(n18553), .A(n18552), .B(n18551), .ZN(
        P3_U2961) );
  AOI22_X1 U21757 ( .A1(n18650), .A2(n18558), .B1(n18705), .B2(n18557), .ZN(
        n18556) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18554), .B1(
        n18707), .B2(n18649), .ZN(n18555) );
  OAI211_X1 U21759 ( .C1(n18653), .C2(n18587), .A(n18556), .B(n18555), .ZN(
        P3_U2962) );
  AOI22_X1 U21760 ( .A1(n18614), .A2(n18558), .B1(n18712), .B2(n18557), .ZN(
        n18560) );
  AOI22_X1 U21761 ( .A1(n18715), .A2(n18649), .B1(n18713), .B2(n18576), .ZN(
        n18559) );
  OAI211_X1 U21762 ( .C1(n18562), .C2(n18561), .A(n18560), .B(n18559), .ZN(
        P3_U2963) );
  NOR2_X2 U21763 ( .A1(n18665), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18691) );
  NOR2_X1 U21764 ( .A1(n18649), .A2(n18691), .ZN(n18623) );
  NOR2_X1 U21765 ( .A1(n18660), .A2(n18623), .ZN(n18583) );
  AOI22_X1 U21766 ( .A1(n18662), .A2(n18613), .B1(n18661), .B2(n18583), .ZN(
        n18569) );
  NAND2_X1 U21767 ( .A1(n18564), .A2(n18563), .ZN(n18565) );
  OAI21_X1 U21768 ( .B1(n18566), .B2(n18565), .A(n18623), .ZN(n18567) );
  OAI211_X1 U21769 ( .C1(n18691), .C2(n18626), .A(n18625), .B(n18567), .ZN(
        n18584) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18584), .B1(
        n18620), .B2(n18576), .ZN(n18568) );
  OAI211_X1 U21771 ( .C1(n18630), .C2(n18720), .A(n18569), .B(n18568), .ZN(
        P3_U2964) );
  AOI22_X1 U21772 ( .A1(n18673), .A2(n18576), .B1(n18672), .B2(n18583), .ZN(
        n18571) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18584), .B1(
        n18674), .B2(n18613), .ZN(n18570) );
  OAI211_X1 U21774 ( .C1(n18677), .C2(n18720), .A(n18571), .B(n18570), .ZN(
        P3_U2965) );
  AOI22_X1 U21775 ( .A1(n18680), .A2(n18613), .B1(n18679), .B2(n18583), .ZN(
        n18573) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18584), .B1(
        n18681), .B2(n18691), .ZN(n18572) );
  OAI211_X1 U21777 ( .C1(n18684), .C2(n18587), .A(n18573), .B(n18572), .ZN(
        P3_U2966) );
  AOI22_X1 U21778 ( .A1(n18599), .A2(n18613), .B1(n18685), .B2(n18583), .ZN(
        n18575) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18584), .B1(
        n18687), .B2(n18691), .ZN(n18574) );
  OAI211_X1 U21780 ( .C1(n18603), .C2(n18587), .A(n18575), .B(n18574), .ZN(
        P3_U2967) );
  AOI22_X1 U21781 ( .A1(n18693), .A2(n18583), .B1(n18692), .B2(n18576), .ZN(
        n18578) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18584), .B1(
        n18694), .B2(n18691), .ZN(n18577) );
  OAI211_X1 U21783 ( .C1(n18697), .C2(n18602), .A(n18578), .B(n18577), .ZN(
        P3_U2968) );
  AOI22_X1 U21784 ( .A1(n18700), .A2(n18613), .B1(n18699), .B2(n18583), .ZN(
        n18580) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18584), .B1(
        n18701), .B2(n18691), .ZN(n18579) );
  OAI211_X1 U21786 ( .C1(n18704), .C2(n18587), .A(n18580), .B(n18579), .ZN(
        P3_U2969) );
  AOI22_X1 U21787 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18584), .B1(
        n18705), .B2(n18583), .ZN(n18582) );
  AOI22_X1 U21788 ( .A1(n18707), .A2(n18691), .B1(n18706), .B2(n18613), .ZN(
        n18581) );
  OAI211_X1 U21789 ( .C1(n18710), .C2(n18587), .A(n18582), .B(n18581), .ZN(
        P3_U2970) );
  AOI22_X1 U21790 ( .A1(n18713), .A2(n18613), .B1(n18712), .B2(n18583), .ZN(
        n18586) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18584), .B1(
        n18715), .B2(n18691), .ZN(n18585) );
  OAI211_X1 U21792 ( .C1(n18721), .C2(n18587), .A(n18586), .B(n18585), .ZN(
        P3_U2971) );
  OAI22_X1 U21793 ( .A1(n18666), .A2(n18590), .B1(n18589), .B2(n18588), .ZN(
        n18617) );
  NOR2_X1 U21794 ( .A1(n18660), .A2(n18665), .ZN(n18612) );
  AOI22_X1 U21795 ( .A1(n18620), .A2(n18613), .B1(n18661), .B2(n18612), .ZN(
        n18592) );
  AOI22_X1 U21796 ( .A1(n18714), .A2(n18668), .B1(n18662), .B2(n18649), .ZN(
        n18591) );
  OAI211_X1 U21797 ( .C1(n18593), .C2(n18617), .A(n18592), .B(n18591), .ZN(
        P3_U2972) );
  AOI22_X1 U21798 ( .A1(n18673), .A2(n18613), .B1(n18672), .B2(n18612), .ZN(
        n18595) );
  AOI22_X1 U21799 ( .A1(n18714), .A2(n18631), .B1(n18674), .B2(n18649), .ZN(
        n18594) );
  OAI211_X1 U21800 ( .C1(n21111), .C2(n18617), .A(n18595), .B(n18594), .ZN(
        P3_U2973) );
  AOI22_X1 U21801 ( .A1(n18679), .A2(n18612), .B1(n18635), .B2(n18613), .ZN(
        n18597) );
  AOI22_X1 U21802 ( .A1(n18714), .A2(n18681), .B1(n18680), .B2(n18649), .ZN(
        n18596) );
  OAI211_X1 U21803 ( .C1(n18598), .C2(n18617), .A(n18597), .B(n18596), .ZN(
        P3_U2974) );
  AOI22_X1 U21804 ( .A1(n18599), .A2(n18649), .B1(n18685), .B2(n18612), .ZN(
        n18601) );
  INV_X1 U21805 ( .A(n18617), .ZN(n18609) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18609), .B1(
        n18714), .B2(n18687), .ZN(n18600) );
  OAI211_X1 U21807 ( .C1(n18603), .C2(n18602), .A(n18601), .B(n18600), .ZN(
        P3_U2975) );
  AOI22_X1 U21808 ( .A1(n18641), .A2(n18649), .B1(n18693), .B2(n18612), .ZN(
        n18605) );
  AOI22_X1 U21809 ( .A1(n18714), .A2(n18694), .B1(n18692), .B2(n18613), .ZN(
        n18604) );
  OAI211_X1 U21810 ( .C1(n18606), .C2(n18617), .A(n18605), .B(n18604), .ZN(
        P3_U2976) );
  AOI22_X1 U21811 ( .A1(n18645), .A2(n18613), .B1(n18699), .B2(n18612), .ZN(
        n18608) );
  AOI22_X1 U21812 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18609), .B1(
        n18714), .B2(n18701), .ZN(n18607) );
  OAI211_X1 U21813 ( .C1(n18648), .C2(n18659), .A(n18608), .B(n18607), .ZN(
        P3_U2977) );
  AOI22_X1 U21814 ( .A1(n18650), .A2(n18613), .B1(n18705), .B2(n18612), .ZN(
        n18611) );
  AOI22_X1 U21815 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18609), .B1(
        n18714), .B2(n18707), .ZN(n18610) );
  OAI211_X1 U21816 ( .C1(n18653), .C2(n18659), .A(n18611), .B(n18610), .ZN(
        P3_U2978) );
  AOI22_X1 U21817 ( .A1(n18614), .A2(n18613), .B1(n18712), .B2(n18612), .ZN(
        n18616) );
  AOI22_X1 U21818 ( .A1(n18714), .A2(n18715), .B1(n18713), .B2(n18649), .ZN(
        n18615) );
  OAI211_X1 U21819 ( .C1(n18618), .C2(n18617), .A(n18616), .B(n18615), .ZN(
        P3_U2979) );
  INV_X1 U21820 ( .A(n18619), .ZN(n18621) );
  NOR2_X1 U21821 ( .A1(n18660), .A2(n18621), .ZN(n18654) );
  AOI22_X1 U21822 ( .A1(n18620), .A2(n18649), .B1(n18661), .B2(n18654), .ZN(
        n18628) );
  OAI21_X1 U21823 ( .B1(n18623), .B2(n18622), .A(n18621), .ZN(n18624) );
  OAI211_X1 U21824 ( .C1(n18655), .C2(n18626), .A(n18625), .B(n18624), .ZN(
        n18656) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18656), .B1(
        n18662), .B2(n18691), .ZN(n18627) );
  OAI211_X1 U21826 ( .C1(n18630), .C2(n18629), .A(n18628), .B(n18627), .ZN(
        P3_U2980) );
  AOI22_X1 U21827 ( .A1(n18674), .A2(n18691), .B1(n18672), .B2(n18654), .ZN(
        n18633) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18656), .B1(
        n18655), .B2(n18631), .ZN(n18632) );
  OAI211_X1 U21829 ( .C1(n18634), .C2(n18659), .A(n18633), .B(n18632), .ZN(
        P3_U2981) );
  AOI22_X1 U21830 ( .A1(n18679), .A2(n18654), .B1(n18635), .B2(n18649), .ZN(
        n18637) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18656), .B1(
        n18655), .B2(n18681), .ZN(n18636) );
  OAI211_X1 U21832 ( .C1(n18638), .C2(n18720), .A(n18637), .B(n18636), .ZN(
        P3_U2982) );
  AOI22_X1 U21833 ( .A1(n18686), .A2(n18649), .B1(n18685), .B2(n18654), .ZN(
        n18640) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18656), .B1(
        n18655), .B2(n18687), .ZN(n18639) );
  OAI211_X1 U21835 ( .C1(n18690), .C2(n18720), .A(n18640), .B(n18639), .ZN(
        P3_U2983) );
  AOI22_X1 U21836 ( .A1(n18641), .A2(n18691), .B1(n18693), .B2(n18654), .ZN(
        n18643) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18656), .B1(
        n18655), .B2(n18694), .ZN(n18642) );
  OAI211_X1 U21838 ( .C1(n18644), .C2(n18659), .A(n18643), .B(n18642), .ZN(
        P3_U2984) );
  AOI22_X1 U21839 ( .A1(n18645), .A2(n18649), .B1(n18699), .B2(n18654), .ZN(
        n18647) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18656), .B1(
        n18655), .B2(n18701), .ZN(n18646) );
  OAI211_X1 U21841 ( .C1(n18648), .C2(n18720), .A(n18647), .B(n18646), .ZN(
        P3_U2985) );
  AOI22_X1 U21842 ( .A1(n18650), .A2(n18649), .B1(n18705), .B2(n18654), .ZN(
        n18652) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18656), .B1(
        n18655), .B2(n18707), .ZN(n18651) );
  OAI211_X1 U21844 ( .C1(n18653), .C2(n18720), .A(n18652), .B(n18651), .ZN(
        P3_U2986) );
  AOI22_X1 U21845 ( .A1(n18713), .A2(n18691), .B1(n18712), .B2(n18654), .ZN(
        n18658) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18656), .B1(
        n18655), .B2(n18715), .ZN(n18657) );
  OAI211_X1 U21847 ( .C1(n18721), .C2(n18659), .A(n18658), .B(n18657), .ZN(
        P3_U2987) );
  NOR2_X1 U21848 ( .A1(n18660), .A2(n18664), .ZN(n18711) );
  AOI22_X1 U21849 ( .A1(n18714), .A2(n18662), .B1(n18661), .B2(n18711), .ZN(
        n18670) );
  OAI22_X1 U21850 ( .A1(n18666), .A2(n18665), .B1(n18664), .B2(n18663), .ZN(
        n18667) );
  INV_X1 U21851 ( .A(n18667), .ZN(n18717) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18717), .B1(
        n18716), .B2(n18668), .ZN(n18669) );
  OAI211_X1 U21853 ( .C1(n18671), .C2(n18720), .A(n18670), .B(n18669), .ZN(
        P3_U2988) );
  AOI22_X1 U21854 ( .A1(n18673), .A2(n18691), .B1(n18672), .B2(n18711), .ZN(
        n18676) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18717), .B1(
        n18714), .B2(n18674), .ZN(n18675) );
  OAI211_X1 U21856 ( .C1(n18678), .C2(n18677), .A(n18676), .B(n18675), .ZN(
        P3_U2989) );
  AOI22_X1 U21857 ( .A1(n18714), .A2(n18680), .B1(n18679), .B2(n18711), .ZN(
        n18683) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18717), .B1(
        n18716), .B2(n18681), .ZN(n18682) );
  OAI211_X1 U21859 ( .C1(n18684), .C2(n18720), .A(n18683), .B(n18682), .ZN(
        P3_U2990) );
  AOI22_X1 U21860 ( .A1(n18686), .A2(n18691), .B1(n18685), .B2(n18711), .ZN(
        n18689) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18717), .B1(
        n18716), .B2(n18687), .ZN(n18688) );
  OAI211_X1 U21862 ( .C1(n18698), .C2(n18690), .A(n18689), .B(n18688), .ZN(
        P3_U2991) );
  AOI22_X1 U21863 ( .A1(n18693), .A2(n18711), .B1(n18692), .B2(n18691), .ZN(
        n18696) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18717), .B1(
        n18716), .B2(n18694), .ZN(n18695) );
  OAI211_X1 U21865 ( .C1(n18698), .C2(n18697), .A(n18696), .B(n18695), .ZN(
        P3_U2992) );
  AOI22_X1 U21866 ( .A1(n18714), .A2(n18700), .B1(n18699), .B2(n18711), .ZN(
        n18703) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18717), .B1(
        n18716), .B2(n18701), .ZN(n18702) );
  OAI211_X1 U21868 ( .C1(n18704), .C2(n18720), .A(n18703), .B(n18702), .ZN(
        P3_U2993) );
  AOI22_X1 U21869 ( .A1(n18714), .A2(n18706), .B1(n18705), .B2(n18711), .ZN(
        n18709) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18717), .B1(
        n18716), .B2(n18707), .ZN(n18708) );
  OAI211_X1 U21871 ( .C1(n18710), .C2(n18720), .A(n18709), .B(n18708), .ZN(
        P3_U2994) );
  AOI22_X1 U21872 ( .A1(n18714), .A2(n18713), .B1(n18712), .B2(n18711), .ZN(
        n18719) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18717), .B1(
        n18716), .B2(n18715), .ZN(n18718) );
  OAI211_X1 U21874 ( .C1(n18721), .C2(n18720), .A(n18719), .B(n18718), .ZN(
        P3_U2995) );
  NAND2_X1 U21875 ( .A1(n21022), .A2(n18948), .ZN(n18935) );
  OAI22_X1 U21876 ( .A1(n18722), .A2(n18935), .B1(n18809), .B2(n18940), .ZN(
        n18792) );
  NAND2_X1 U21877 ( .A1(n18752), .A2(n18723), .ZN(n18729) );
  NAND2_X1 U21878 ( .A1(n18724), .A2(n18747), .ZN(n18726) );
  AOI222_X1 U21879 ( .A1(n18730), .A2(n18729), .B1(n18728), .B2(n18727), .C1(
        n18726), .C2(n18725), .ZN(n18930) );
  AOI211_X1 U21880 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18770), .A(
        n18732), .B(n18731), .ZN(n18783) );
  OAI21_X1 U21881 ( .B1(n18735), .B2(n18734), .A(n18733), .ZN(n18745) );
  AOI21_X1 U21882 ( .B1(n18739), .B2(n18740), .A(n18745), .ZN(n18737) );
  INV_X1 U21883 ( .A(n18741), .ZN(n18736) );
  OAI21_X1 U21884 ( .B1(n18738), .B2(n18737), .A(n18736), .ZN(n18896) );
  NOR2_X1 U21885 ( .A1(n18770), .A2(n18896), .ZN(n18743) );
  NOR2_X1 U21886 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18739), .ZN(
        n18762) );
  OAI22_X1 U21887 ( .A1(n18741), .A2(n18752), .B1(n18762), .B2(n18740), .ZN(
        n18893) );
  NAND2_X1 U21888 ( .A1(n18897), .A2(n18893), .ZN(n18742) );
  OAI22_X1 U21889 ( .A1(n18743), .A2(n18897), .B1(n18770), .B2(n18742), .ZN(
        n18779) );
  NOR2_X1 U21890 ( .A1(n18744), .A2(n21179), .ZN(n18756) );
  AOI21_X1 U21891 ( .B1(n18910), .B2(n12833), .A(n18745), .ZN(n18746) );
  INV_X1 U21892 ( .A(n18746), .ZN(n18755) );
  AOI211_X1 U21893 ( .C1(n18910), .C2(n9798), .A(n18748), .B(n18747), .ZN(
        n18754) );
  NOR2_X1 U21894 ( .A1(n18749), .A2(n18916), .ZN(n18750) );
  OAI211_X1 U21895 ( .C1(n18750), .C2(n12833), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n21179), .ZN(n18751) );
  OAI21_X1 U21896 ( .B1(n18901), .B2(n18752), .A(n18751), .ZN(n18753) );
  AOI211_X1 U21897 ( .C1(n18756), .C2(n18755), .A(n18754), .B(n18753), .ZN(
        n18757) );
  INV_X1 U21898 ( .A(n18757), .ZN(n18903) );
  OAI22_X1 U21899 ( .A1(n18758), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18903), .B2(n18770), .ZN(n18775) );
  INV_X1 U21900 ( .A(n18775), .ZN(n18773) );
  NOR2_X1 U21901 ( .A1(n18760), .A2(n18759), .ZN(n18764) );
  AOI22_X1 U21902 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18761), .B1(
        n18764), .B2(n18916), .ZN(n18912) );
  OAI22_X1 U21903 ( .A1(n18764), .A2(n18763), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18762), .ZN(n18908) );
  OR3_X1 U21904 ( .A1(n18912), .A2(n18767), .A3(n18765), .ZN(n18766) );
  AOI22_X1 U21905 ( .A1(n18912), .A2(n18767), .B1(n18908), .B2(n18766), .ZN(
        n18769) );
  OAI21_X1 U21906 ( .B1(n18770), .B2(n18769), .A(n18768), .ZN(n18771) );
  OAI21_X1 U21907 ( .B1(n18773), .B2(n18772), .A(n18771), .ZN(n18774) );
  OAI221_X1 U21908 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n18774), .A(n18775), .ZN(
        n18778) );
  NOR2_X1 U21909 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18777) );
  OAI21_X1 U21910 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18775), .A(
        n18774), .ZN(n18776) );
  AOI22_X1 U21911 ( .A1(n18779), .A2(n18778), .B1(n18777), .B2(n18776), .ZN(
        n18782) );
  OAI21_X1 U21912 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18780), .ZN(n18781) );
  NAND4_X1 U21913 ( .A1(n18930), .A2(n18783), .A3(n18782), .A4(n18781), .ZN(
        n18789) );
  AOI211_X1 U21914 ( .C1(n18786), .C2(n18785), .A(n18784), .B(n18789), .ZN(
        n18889) );
  AOI21_X1 U21915 ( .B1(n18941), .B2(n18948), .A(n18889), .ZN(n18795) );
  INV_X1 U21916 ( .A(n18787), .ZN(n18788) );
  OAI211_X1 U21917 ( .C1(P3_STATE2_REG_1__SCAN_IN), .C2(n18794), .A(n18795), 
        .B(n18788), .ZN(n18790) );
  AOI22_X1 U21918 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18790), .B1(n18939), 
        .B2(n18789), .ZN(n18791) );
  OAI21_X1 U21919 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18792), .A(n18791), 
        .ZN(P3_U2996) );
  NAND2_X1 U21920 ( .A1(n18941), .A2(n18793), .ZN(n18799) );
  NOR4_X1 U21921 ( .A1(n18936), .A2(n21022), .A3(n18809), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18801) );
  INV_X1 U21922 ( .A(n18801), .ZN(n18798) );
  NAND3_X1 U21923 ( .A1(n18796), .A2(n18795), .A3(n18794), .ZN(n18797) );
  NAND4_X1 U21924 ( .A1(n18800), .A2(n18799), .A3(n18798), .A4(n18797), .ZN(
        P3_U2997) );
  NOR2_X1 U21925 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATEBS16_REG_SCAN_IN), .ZN(n18804) );
  AOI221_X1 U21926 ( .B1(n18804), .B2(n18803), .C1(n18802), .C2(n18803), .A(
        n18801), .ZN(P3_U2998) );
  AND2_X1 U21927 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18805), .ZN(
        P3_U2999) );
  AND2_X1 U21928 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18805), .ZN(
        P3_U3000) );
  AND2_X1 U21929 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18805), .ZN(
        P3_U3001) );
  AND2_X1 U21930 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18805), .ZN(
        P3_U3002) );
  AND2_X1 U21931 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18805), .ZN(
        P3_U3003) );
  AND2_X1 U21932 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18805), .ZN(
        P3_U3004) );
  AND2_X1 U21933 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18805), .ZN(
        P3_U3005) );
  INV_X1 U21934 ( .A(P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(n20974) );
  NOR2_X1 U21935 ( .A1(n20974), .A2(n18888), .ZN(P3_U3006) );
  AND2_X1 U21936 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18805), .ZN(
        P3_U3007) );
  AND2_X1 U21937 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18805), .ZN(
        P3_U3008) );
  AND2_X1 U21938 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18805), .ZN(
        P3_U3009) );
  AND2_X1 U21939 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18805), .ZN(
        P3_U3010) );
  AND2_X1 U21940 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18805), .ZN(
        P3_U3011) );
  AND2_X1 U21941 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18805), .ZN(
        P3_U3012) );
  AND2_X1 U21942 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18805), .ZN(
        P3_U3013) );
  AND2_X1 U21943 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18805), .ZN(
        P3_U3014) );
  AND2_X1 U21944 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18805), .ZN(
        P3_U3015) );
  AND2_X1 U21945 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18805), .ZN(
        P3_U3016) );
  AND2_X1 U21946 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18805), .ZN(
        P3_U3017) );
  AND2_X1 U21947 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18805), .ZN(
        P3_U3018) );
  AND2_X1 U21948 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18805), .ZN(
        P3_U3019) );
  AND2_X1 U21949 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18805), .ZN(
        P3_U3020) );
  AND2_X1 U21950 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18805), .ZN(P3_U3021) );
  AND2_X1 U21951 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18805), .ZN(P3_U3022) );
  AND2_X1 U21952 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18805), .ZN(P3_U3023) );
  AND2_X1 U21953 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18805), .ZN(P3_U3024) );
  AND2_X1 U21954 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18805), .ZN(P3_U3025) );
  AND2_X1 U21955 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18805), .ZN(P3_U3026) );
  AND2_X1 U21956 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18805), .ZN(P3_U3027) );
  AND2_X1 U21957 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18805), .ZN(P3_U3028) );
  INV_X1 U21958 ( .A(HOLD), .ZN(n20782) );
  OAI21_X1 U21959 ( .B1(n18806), .B2(n20782), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18807) );
  AOI22_X1 U21960 ( .A1(n18820), .A2(n18822), .B1(n18946), .B2(n18807), .ZN(
        n18808) );
  INV_X1 U21961 ( .A(NA), .ZN(n20786) );
  OR3_X1 U21962 ( .A1(n20786), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18815) );
  OAI211_X1 U21963 ( .C1(n18809), .C2(n18810), .A(n18808), .B(n18815), .ZN(
        P3_U3029) );
  INV_X1 U21964 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18811) );
  NOR2_X1 U21965 ( .A1(n18822), .A2(n20782), .ZN(n18818) );
  OAI22_X1 U21966 ( .A1(n18811), .A2(n18818), .B1(n20782), .B2(n18810), .ZN(
        n18812) );
  INV_X1 U21967 ( .A(n18812), .ZN(n18814) );
  NAND2_X1 U21968 ( .A1(n18941), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18816) );
  INV_X1 U21969 ( .A(n18932), .ZN(n18813) );
  OAI211_X1 U21970 ( .C1(n18814), .C2(n18820), .A(n18816), .B(n18813), .ZN(
        P3_U3030) );
  AOI22_X1 U21971 ( .A1(n18941), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18820), 
        .B2(n18815), .ZN(n18821) );
  OAI22_X1 U21972 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18816), .ZN(n18817) );
  OAI22_X1 U21973 ( .A1(n18818), .A2(n18817), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18819) );
  OAI22_X1 U21974 ( .A1(n18821), .A2(n18822), .B1(n18820), .B2(n18819), .ZN(
        P3_U3031) );
  INV_X2 U21975 ( .A(n18829), .ZN(n18881) );
  INV_X1 U21976 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18824) );
  OAI222_X1 U21977 ( .A1(n18918), .A2(n18881), .B1(n18823), .B2(n18945), .C1(
        n18824), .C2(n18869), .ZN(P3_U3032) );
  OAI222_X1 U21978 ( .A1(n18869), .A2(n18826), .B1(n21092), .B2(n18945), .C1(
        n18824), .C2(n18881), .ZN(P3_U3033) );
  OAI222_X1 U21979 ( .A1(n18826), .A2(n18881), .B1(n18825), .B2(n18945), .C1(
        n18827), .C2(n18869), .ZN(P3_U3034) );
  OAI222_X1 U21980 ( .A1(n18869), .A2(n18830), .B1(n18828), .B2(n18945), .C1(
        n18827), .C2(n18881), .ZN(P3_U3035) );
  INV_X1 U21981 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18832) );
  OAI222_X1 U21982 ( .A1(n18869), .A2(n18832), .B1(n18831), .B2(n18945), .C1(
        n18830), .C2(n18881), .ZN(P3_U3036) );
  OAI222_X1 U21983 ( .A1(n18869), .A2(n18834), .B1(n18833), .B2(n18945), .C1(
        n18832), .C2(n18881), .ZN(P3_U3037) );
  OAI222_X1 U21984 ( .A1(n18869), .A2(n18836), .B1(n18835), .B2(n18945), .C1(
        n18834), .C2(n18881), .ZN(P3_U3038) );
  OAI222_X1 U21985 ( .A1(n18836), .A2(n18881), .B1(n21077), .B2(n18945), .C1(
        n18837), .C2(n18869), .ZN(P3_U3039) );
  OAI222_X1 U21986 ( .A1(n18869), .A2(n18839), .B1(n18838), .B2(n18945), .C1(
        n18837), .C2(n18881), .ZN(P3_U3040) );
  OAI222_X1 U21987 ( .A1(n18869), .A2(n18841), .B1(n18840), .B2(n18945), .C1(
        n18839), .C2(n18881), .ZN(P3_U3041) );
  INV_X1 U21988 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18843) );
  OAI222_X1 U21989 ( .A1(n18869), .A2(n18843), .B1(n18842), .B2(n18945), .C1(
        n18841), .C2(n18881), .ZN(P3_U3042) );
  INV_X1 U21990 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18845) );
  OAI222_X1 U21991 ( .A1(n18869), .A2(n18845), .B1(n18844), .B2(n18945), .C1(
        n18843), .C2(n18881), .ZN(P3_U3043) );
  INV_X1 U21992 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18848) );
  OAI222_X1 U21993 ( .A1(n18869), .A2(n18848), .B1(n18846), .B2(n18945), .C1(
        n18845), .C2(n18881), .ZN(P3_U3044) );
  OAI222_X1 U21994 ( .A1(n18848), .A2(n18881), .B1(n18847), .B2(n18945), .C1(
        n18849), .C2(n18869), .ZN(P3_U3045) );
  OAI222_X1 U21995 ( .A1(n18869), .A2(n18851), .B1(n18850), .B2(n18945), .C1(
        n18849), .C2(n18881), .ZN(P3_U3046) );
  INV_X1 U21996 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18853) );
  OAI222_X1 U21997 ( .A1(n18869), .A2(n18853), .B1(n18852), .B2(n18945), .C1(
        n18851), .C2(n18881), .ZN(P3_U3047) );
  OAI222_X1 U21998 ( .A1(n18869), .A2(n18855), .B1(n18854), .B2(n18945), .C1(
        n18853), .C2(n18881), .ZN(P3_U3048) );
  OAI222_X1 U21999 ( .A1(n18869), .A2(n18857), .B1(n18856), .B2(n18945), .C1(
        n18855), .C2(n18881), .ZN(P3_U3049) );
  OAI222_X1 U22000 ( .A1(n18869), .A2(n18859), .B1(n18858), .B2(n18945), .C1(
        n18857), .C2(n18881), .ZN(P3_U3050) );
  OAI222_X1 U22001 ( .A1(n18869), .A2(n18862), .B1(n18860), .B2(n18945), .C1(
        n18859), .C2(n18881), .ZN(P3_U3051) );
  OAI222_X1 U22002 ( .A1(n18862), .A2(n18881), .B1(n18861), .B2(n18945), .C1(
        n18863), .C2(n18869), .ZN(P3_U3052) );
  OAI222_X1 U22003 ( .A1(n18869), .A2(n18866), .B1(n18864), .B2(n18945), .C1(
        n18863), .C2(n18881), .ZN(P3_U3053) );
  OAI222_X1 U22004 ( .A1(n18866), .A2(n18881), .B1(n18865), .B2(n18945), .C1(
        n18867), .C2(n18869), .ZN(P3_U3054) );
  OAI222_X1 U22005 ( .A1(n18869), .A2(n18870), .B1(n18868), .B2(n18945), .C1(
        n18867), .C2(n18881), .ZN(P3_U3055) );
  OAI222_X1 U22006 ( .A1(n18869), .A2(n21158), .B1(n18871), .B2(n18945), .C1(
        n18870), .C2(n18881), .ZN(P3_U3056) );
  OAI222_X1 U22007 ( .A1(n18869), .A2(n18873), .B1(n18872), .B2(n18945), .C1(
        n21158), .C2(n18881), .ZN(P3_U3057) );
  OAI222_X1 U22008 ( .A1(n18869), .A2(n18876), .B1(n18874), .B2(n18945), .C1(
        n18873), .C2(n18881), .ZN(P3_U3058) );
  OAI222_X1 U22009 ( .A1(n18876), .A2(n18881), .B1(n18875), .B2(n18945), .C1(
        n20979), .C2(n18869), .ZN(P3_U3059) );
  OAI222_X1 U22010 ( .A1(n18869), .A2(n18880), .B1(n18877), .B2(n18945), .C1(
        n20979), .C2(n18881), .ZN(P3_U3060) );
  OAI222_X1 U22011 ( .A1(n18881), .A2(n18880), .B1(n18879), .B2(n18945), .C1(
        n18878), .C2(n18869), .ZN(P3_U3061) );
  OAI22_X1 U22012 ( .A1(n18946), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18945), .ZN(n18882) );
  INV_X1 U22013 ( .A(n18882), .ZN(P3_U3274) );
  OAI22_X1 U22014 ( .A1(n18946), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18945), .ZN(n18883) );
  INV_X1 U22015 ( .A(n18883), .ZN(P3_U3275) );
  OAI22_X1 U22016 ( .A1(n18946), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18945), .ZN(n18884) );
  INV_X1 U22017 ( .A(n18884), .ZN(P3_U3276) );
  INV_X1 U22018 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18926) );
  INV_X1 U22019 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n21150) );
  AOI22_X1 U22020 ( .A1(n18945), .A2(n18926), .B1(n21150), .B2(n18946), .ZN(
        P3_U3277) );
  OAI21_X1 U22021 ( .B1(n18888), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18886), 
        .ZN(n18885) );
  INV_X1 U22022 ( .A(n18885), .ZN(P3_U3280) );
  OAI21_X1 U22023 ( .B1(n18888), .B2(n18887), .A(n18886), .ZN(P3_U3281) );
  OAI21_X1 U22024 ( .B1(n18936), .B2(n18889), .A(P3_STATE2_REG_3__SCAN_IN), 
        .ZN(n18891) );
  NAND2_X1 U22025 ( .A1(n18891), .A2(n18890), .ZN(P3_U3282) );
  NOR2_X1 U22026 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18892), .ZN(
        n18894) );
  AOI22_X1 U22027 ( .A1(n18911), .A2(n18895), .B1(n18894), .B2(n18893), .ZN(
        n18899) );
  AOI21_X1 U22028 ( .B1(n18949), .B2(n18896), .A(n18917), .ZN(n18898) );
  OAI22_X1 U22029 ( .A1(n18917), .A2(n18899), .B1(n18898), .B2(n18897), .ZN(
        P3_U3285) );
  NOR2_X1 U22030 ( .A1(n21022), .A2(n18913), .ZN(n18905) );
  OAI22_X1 U22031 ( .A1(n18900), .A2(n20976), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18906) );
  INV_X1 U22032 ( .A(n18906), .ZN(n18902) );
  AOI222_X1 U22033 ( .A1(n18903), .A2(n18949), .B1(n18905), .B2(n18902), .C1(
        n18911), .C2(n18901), .ZN(n18904) );
  AOI22_X1 U22034 ( .A1(n18917), .A2(n9798), .B1(n18904), .B2(n18914), .ZN(
        P3_U3288) );
  AOI222_X1 U22035 ( .A1(n18908), .A2(n18949), .B1(n18911), .B2(n18907), .C1(
        n18906), .C2(n18905), .ZN(n18909) );
  AOI22_X1 U22036 ( .A1(n18917), .A2(n18910), .B1(n18909), .B2(n18914), .ZN(
        P3_U3289) );
  AOI222_X1 U22037 ( .A1(n18913), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18949), 
        .B2(n18912), .C1(n18916), .C2(n18911), .ZN(n18915) );
  AOI22_X1 U22038 ( .A1(n18917), .A2(n18916), .B1(n18915), .B2(n18914), .ZN(
        P3_U3290) );
  AOI21_X1 U22039 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18919) );
  AOI22_X1 U22040 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18919), .B2(n18918), .ZN(n18921) );
  INV_X1 U22041 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18920) );
  AOI22_X1 U22042 ( .A1(n18922), .A2(n18921), .B1(n18920), .B2(n18925), .ZN(
        P3_U3292) );
  NOR2_X1 U22043 ( .A1(n18925), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18923) );
  AOI22_X1 U22044 ( .A1(n18926), .A2(n18925), .B1(n18924), .B2(n18923), .ZN(
        P3_U3293) );
  INV_X1 U22045 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18952) );
  OAI22_X1 U22046 ( .A1(n18946), .A2(n18952), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18945), .ZN(n18927) );
  INV_X1 U22047 ( .A(n18927), .ZN(P3_U3294) );
  INV_X1 U22048 ( .A(n18928), .ZN(n18931) );
  NAND2_X1 U22049 ( .A1(n18931), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18929) );
  OAI21_X1 U22050 ( .B1(n18931), .B2(n18930), .A(n18929), .ZN(P3_U3295) );
  OAI21_X1 U22051 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18933), .A(n18932), 
        .ZN(n18934) );
  AOI211_X1 U22052 ( .C1(n18950), .C2(n18934), .A(n18941), .B(n18948), .ZN(
        n18937) );
  OAI21_X1 U22053 ( .B1(n18937), .B2(n18936), .A(n18935), .ZN(n18944) );
  OAI22_X1 U22054 ( .A1(n18941), .A2(n18940), .B1(n18939), .B2(n18938), .ZN(
        n18942) );
  NOR2_X1 U22055 ( .A1(n18951), .A2(n18942), .ZN(n18943) );
  MUX2_X1 U22056 ( .A(n18944), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18943), 
        .Z(P3_U3296) );
  OAI22_X1 U22057 ( .A1(n18946), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18945), .ZN(n18947) );
  INV_X1 U22058 ( .A(n18947), .ZN(P3_U3297) );
  AOI21_X1 U22059 ( .B1(n18949), .B2(n18948), .A(n18951), .ZN(n18955) );
  AOI22_X1 U22060 ( .A1(n18955), .A2(n18952), .B1(n18951), .B2(n18950), .ZN(
        P3_U3298) );
  INV_X1 U22061 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18954) );
  AOI21_X1 U22062 ( .B1(n18955), .B2(n18954), .A(n18953), .ZN(P3_U3299) );
  AOI211_X1 U22063 ( .C1(n18958), .C2(P2_MEMORYFETCH_REG_SCAN_IN), .A(n18957), 
        .B(n18956), .ZN(n18959) );
  INV_X1 U22064 ( .A(n18959), .ZN(P2_U2814) );
  AND2_X1 U22065 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19861), .ZN(n19851) );
  NOR2_X1 U22066 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n18962) );
  AOI21_X1 U22067 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19851), .A(n18962), 
        .ZN(n19844) );
  INV_X1 U22068 ( .A(n19844), .ZN(n19922) );
  AOI21_X1 U22069 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19922), .ZN(n18960) );
  INV_X1 U22070 ( .A(n18960), .ZN(P2_U2815) );
  INV_X1 U22071 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18963) );
  OAI22_X1 U22072 ( .A1(n18961), .A2(n19722), .B1(n19981), .B2(n18963), .ZN(
        P2_U2816) );
  INV_X1 U22073 ( .A(n18962), .ZN(n19850) );
  AOI22_X1 U22074 ( .A1(n19988), .A2(n18963), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19986), .ZN(n18964) );
  OAI21_X1 U22075 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n19850), .A(n18964), 
        .ZN(P2_U2817) );
  OAI21_X1 U22076 ( .B1(n19845), .B2(BS16), .A(n19922), .ZN(n19920) );
  OAI21_X1 U22077 ( .B1(n19922), .B2(n10593), .A(n19920), .ZN(P2_U2818) );
  NOR2_X1 U22078 ( .A1(n18966), .A2(n18965), .ZN(n19967) );
  OAI21_X1 U22079 ( .B1(n19967), .B2(n18968), .A(n18967), .ZN(P2_U2819) );
  NOR4_X1 U22080 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18978) );
  NOR4_X1 U22081 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18977) );
  NOR4_X1 U22082 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18969) );
  INV_X1 U22083 ( .A(P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n21146) );
  INV_X1 U22084 ( .A(P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20992) );
  NAND3_X1 U22085 ( .A1(n18969), .A2(n21146), .A3(n20992), .ZN(n18975) );
  NOR4_X1 U22086 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18973) );
  NOR4_X1 U22087 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18972) );
  NOR4_X1 U22088 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18971) );
  NOR4_X1 U22089 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18970) );
  NAND4_X1 U22090 ( .A1(n18973), .A2(n18972), .A3(n18971), .A4(n18970), .ZN(
        n18974) );
  AOI211_X1 U22091 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n18975), .B(n18974), .ZN(n18976) );
  NAND3_X1 U22092 ( .A1(n18978), .A2(n18977), .A3(n18976), .ZN(n18987) );
  NOR2_X1 U22093 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18987), .ZN(n18981) );
  INV_X1 U22094 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18979) );
  AOI22_X1 U22095 ( .A1(n18981), .A2(n18982), .B1(n18987), .B2(n18979), .ZN(
        P2_U2820) );
  OR3_X1 U22096 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18986) );
  INV_X1 U22097 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18980) );
  AOI22_X1 U22098 ( .A1(n18981), .A2(n18986), .B1(n18987), .B2(n18980), .ZN(
        P2_U2821) );
  INV_X1 U22099 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19921) );
  NAND2_X1 U22100 ( .A1(n18981), .A2(n19921), .ZN(n18985) );
  INV_X1 U22101 ( .A(n18987), .ZN(n18988) );
  OAI21_X1 U22102 ( .B1(n19862), .B2(n18982), .A(n18988), .ZN(n18983) );
  OAI21_X1 U22103 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18988), .A(n18983), 
        .ZN(n18984) );
  OAI221_X1 U22104 ( .B1(n18985), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18985), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18984), .ZN(P2_U2822) );
  INV_X1 U22105 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21126) );
  OAI221_X1 U22106 ( .B1(n18988), .B2(n21126), .C1(n18987), .C2(n18986), .A(
        n18985), .ZN(P2_U2823) );
  INV_X1 U22107 ( .A(n18989), .ZN(n18994) );
  AOI22_X1 U22108 ( .A1(n19128), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19145), .ZN(n18991) );
  NAND2_X1 U22109 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n19138), .ZN(
        n18990) );
  OAI211_X1 U22110 ( .C1(n18992), .C2(n19142), .A(n18991), .B(n18990), .ZN(
        n18993) );
  AOI21_X1 U22111 ( .B1(n18994), .B2(n19109), .A(n18993), .ZN(n18998) );
  OAI211_X1 U22112 ( .C1(n18996), .C2(n19000), .A(n19154), .B(n18995), .ZN(
        n18997) );
  OAI211_X1 U22113 ( .C1(n19150), .C2(n18999), .A(n18998), .B(n18997), .ZN(
        P2_U2834) );
  AOI21_X1 U22114 ( .B1(n19004), .B2(n19001), .A(n19000), .ZN(n19003) );
  AOI22_X1 U22115 ( .A1(n19003), .A2(n19154), .B1(n19129), .B2(n19002), .ZN(
        n19010) );
  AOI22_X1 U22116 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19145), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n19128), .ZN(n19009) );
  AOI22_X1 U22117 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19138), .B1(
        n19004), .B2(n19028), .ZN(n19008) );
  AOI22_X1 U22118 ( .A1(n19006), .A2(n19109), .B1(n19005), .B2(n19089), .ZN(
        n19007) );
  NAND4_X1 U22119 ( .A1(n19010), .A2(n19009), .A3(n19008), .A4(n19007), .ZN(
        P2_U2835) );
  NOR2_X1 U22120 ( .A1(n19147), .A2(n19011), .ZN(n19012) );
  XOR2_X1 U22121 ( .A(n19013), .B(n19012), .Z(n19025) );
  OAI21_X1 U22122 ( .B1(n21177), .B2(n19133), .A(n19131), .ZN(n19018) );
  INV_X1 U22123 ( .A(n19014), .ZN(n19016) );
  INV_X1 U22124 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19015) );
  OAI22_X1 U22125 ( .A1(n19016), .A2(n19142), .B1(n19158), .B2(n19015), .ZN(
        n19017) );
  AOI211_X1 U22126 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19128), .A(n19018), .B(
        n19017), .ZN(n19024) );
  INV_X1 U22127 ( .A(n19019), .ZN(n19020) );
  OAI22_X1 U22128 ( .A1(n19021), .A2(n19151), .B1(n19020), .B2(n19150), .ZN(
        n19022) );
  INV_X1 U22129 ( .A(n19022), .ZN(n19023) );
  OAI211_X1 U22130 ( .C1(n19840), .C2(n19025), .A(n19024), .B(n19023), .ZN(
        P2_U2836) );
  INV_X1 U22131 ( .A(n19035), .ZN(n19029) );
  INV_X1 U22132 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U22133 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19138), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19128), .ZN(n19026) );
  OAI211_X1 U22134 ( .C1(n19133), .C2(n19887), .A(n19026), .B(n19131), .ZN(
        n19027) );
  AOI21_X1 U22135 ( .B1(n19029), .B2(n19028), .A(n19027), .ZN(n19030) );
  OAI21_X1 U22136 ( .B1(n19031), .B2(n19142), .A(n19030), .ZN(n19032) );
  AOI21_X1 U22137 ( .B1(n19033), .B2(n19109), .A(n19032), .ZN(n19038) );
  OAI21_X1 U22138 ( .B1(n19036), .B2(n19035), .A(n19034), .ZN(n19037) );
  OAI211_X1 U22139 ( .C1(n19150), .C2(n19039), .A(n19038), .B(n19037), .ZN(
        P2_U2838) );
  NOR2_X1 U22140 ( .A1(n19147), .A2(n19040), .ZN(n19042) );
  XOR2_X1 U22141 ( .A(n19042), .B(n19041), .Z(n19051) );
  INV_X1 U22142 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U22143 ( .A1(n19043), .A2(n19129), .B1(P2_EBX_REG_15__SCAN_IN), 
        .B2(n19128), .ZN(n19044) );
  OAI211_X1 U22144 ( .C1(n19883), .C2(n19133), .A(n19044), .B(n19131), .ZN(
        n19049) );
  INV_X1 U22145 ( .A(n19045), .ZN(n19047) );
  OAI22_X1 U22146 ( .A1(n19047), .A2(n19151), .B1(n19046), .B2(n19150), .ZN(
        n19048) );
  AOI211_X1 U22147 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19138), .A(
        n19049), .B(n19048), .ZN(n19050) );
  OAI21_X1 U22148 ( .B1(n19840), .B2(n19051), .A(n19050), .ZN(P2_U2840) );
  NAND2_X1 U22149 ( .A1(n19075), .A2(n19052), .ZN(n19061) );
  XOR2_X1 U22150 ( .A(n19053), .B(n19061), .Z(n19060) );
  AOI22_X1 U22151 ( .A1(n19054), .A2(n19129), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19138), .ZN(n19055) );
  OAI211_X1 U22152 ( .C1(n19881), .C2(n19133), .A(n19055), .B(n19131), .ZN(
        n19056) );
  AOI21_X1 U22153 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19128), .A(n19056), .ZN(
        n19059) );
  AOI22_X1 U22154 ( .A1(n19057), .A2(n19109), .B1(n19177), .B2(n19089), .ZN(
        n19058) );
  OAI211_X1 U22155 ( .C1(n19840), .C2(n19060), .A(n19059), .B(n19058), .ZN(
        P2_U2841) );
  INV_X1 U22156 ( .A(n19061), .ZN(n19062) );
  OAI211_X1 U22157 ( .C1(n19063), .C2(n19068), .A(n19154), .B(n19062), .ZN(
        n19065) );
  AOI22_X1 U22158 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19138), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19128), .ZN(n19064) );
  OAI211_X1 U22159 ( .C1(n19066), .C2(n19142), .A(n19065), .B(n19064), .ZN(
        n19067) );
  AOI211_X1 U22160 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19145), .A(n19088), 
        .B(n19067), .ZN(n19072) );
  OAI22_X1 U22161 ( .A1(n19069), .A2(n19151), .B1(n19102), .B2(n19068), .ZN(
        n19070) );
  INV_X1 U22162 ( .A(n19070), .ZN(n19071) );
  OAI211_X1 U22163 ( .C1(n19073), .C2(n19150), .A(n19072), .B(n19071), .ZN(
        P2_U2842) );
  NAND2_X1 U22164 ( .A1(n19075), .A2(n19074), .ZN(n19096) );
  XOR2_X1 U22165 ( .A(n19076), .B(n19096), .Z(n19084) );
  AOI22_X1 U22166 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19138), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19128), .ZN(n19077) );
  OAI21_X1 U22167 ( .B1(n19078), .B2(n19142), .A(n19077), .ZN(n19079) );
  AOI211_X1 U22168 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19145), .A(n19275), 
        .B(n19079), .ZN(n19083) );
  AOI22_X1 U22169 ( .A1(n19081), .A2(n19109), .B1(n19080), .B2(n19089), .ZN(
        n19082) );
  OAI211_X1 U22170 ( .C1(n19840), .C2(n19084), .A(n19083), .B(n19082), .ZN(
        P2_U2843) );
  OAI22_X1 U22171 ( .A1(n19143), .A2(n10449), .B1(n19085), .B2(n19158), .ZN(
        n19094) );
  INV_X1 U22172 ( .A(n19086), .ZN(n19092) );
  NOR2_X1 U22173 ( .A1(n19133), .A2(n19876), .ZN(n19087) );
  AOI211_X1 U22174 ( .C1(n19090), .C2(n19089), .A(n19088), .B(n19087), .ZN(
        n19091) );
  OAI21_X1 U22175 ( .B1(n19092), .B2(n19142), .A(n19091), .ZN(n19093) );
  AOI211_X1 U22176 ( .C1(n19095), .C2(n19109), .A(n19094), .B(n19093), .ZN(
        n19100) );
  INV_X1 U22177 ( .A(n19096), .ZN(n19097) );
  OAI211_X1 U22178 ( .C1(n19098), .C2(n19101), .A(n19154), .B(n19097), .ZN(
        n19099) );
  OAI211_X1 U22179 ( .C1(n19102), .C2(n19101), .A(n19100), .B(n19099), .ZN(
        P2_U2844) );
  OAI21_X1 U22180 ( .B1(n11445), .B2(n19133), .A(n19131), .ZN(n19105) );
  OAI22_X1 U22181 ( .A1(n19103), .A2(n19142), .B1(n19143), .B2(n10009), .ZN(
        n19104) );
  AOI211_X1 U22182 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19138), .A(
        n19105), .B(n19104), .ZN(n19113) );
  NAND2_X1 U22183 ( .A1(n19075), .A2(n19106), .ZN(n19107) );
  XOR2_X1 U22184 ( .A(n19108), .B(n19107), .Z(n19111) );
  AOI22_X1 U22185 ( .A1(n19111), .A2(n19154), .B1(n19110), .B2(n19109), .ZN(
        n19112) );
  OAI211_X1 U22186 ( .C1(n19186), .C2(n19150), .A(n19113), .B(n19112), .ZN(
        P2_U2845) );
  NOR2_X1 U22187 ( .A1(n19147), .A2(n19114), .ZN(n19116) );
  XOR2_X1 U22188 ( .A(n19116), .B(n19115), .Z(n19124) );
  AOI22_X1 U22189 ( .A1(n19117), .A2(n19129), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19128), .ZN(n19118) );
  OAI211_X1 U22190 ( .C1(n19873), .C2(n19133), .A(n19118), .B(n19131), .ZN(
        n19122) );
  OAI22_X1 U22191 ( .A1(n19120), .A2(n19150), .B1(n19151), .B2(n19119), .ZN(
        n19121) );
  AOI211_X1 U22192 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19138), .A(
        n19122), .B(n19121), .ZN(n19123) );
  OAI21_X1 U22193 ( .B1(n19840), .B2(n19124), .A(n19123), .ZN(P2_U2846) );
  NOR2_X1 U22194 ( .A1(n19147), .A2(n19125), .ZN(n19126) );
  XOR2_X1 U22195 ( .A(n19127), .B(n19126), .Z(n19140) );
  AOI22_X1 U22196 ( .A1(n19130), .A2(n19129), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19128), .ZN(n19132) );
  OAI211_X1 U22197 ( .C1(n19872), .C2(n19133), .A(n19132), .B(n19131), .ZN(
        n19137) );
  OAI22_X1 U22198 ( .A1(n19135), .A2(n19151), .B1(n19150), .B2(n19134), .ZN(
        n19136) );
  AOI211_X1 U22199 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19138), .A(
        n19137), .B(n19136), .ZN(n19139) );
  OAI21_X1 U22200 ( .B1(n19840), .B2(n19140), .A(n19139), .ZN(P2_U2848) );
  OAI22_X1 U22201 ( .A1(n19143), .A2(n10429), .B1(n19142), .B2(n19141), .ZN(
        n19144) );
  AOI211_X1 U22202 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19145), .A(n19275), .B(
        n19144), .ZN(n19157) );
  NOR2_X1 U22203 ( .A1(n19147), .A2(n19146), .ZN(n19148) );
  XNOR2_X1 U22204 ( .A(n19149), .B(n19148), .ZN(n19155) );
  OAI22_X1 U22205 ( .A1(n19152), .A2(n19151), .B1(n19199), .B2(n19150), .ZN(
        n19153) );
  AOI21_X1 U22206 ( .B1(n19155), .B2(n19154), .A(n19153), .ZN(n19156) );
  OAI211_X1 U22207 ( .C1(n19159), .C2(n19158), .A(n19157), .B(n19156), .ZN(
        P2_U2850) );
  OAI22_X1 U22208 ( .A1(n19161), .A2(n19170), .B1(n19160), .B2(n19338), .ZN(
        n19162) );
  INV_X1 U22209 ( .A(n19162), .ZN(n19164) );
  AOI22_X1 U22210 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19190), .B1(n19167), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19163) );
  NAND2_X1 U22211 ( .A1(n19164), .A2(n19163), .ZN(P2_U2888) );
  AOI22_X1 U22212 ( .A1(n19166), .A2(n19165), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19190), .ZN(n19176) );
  AOI22_X1 U22213 ( .A1(n19168), .A2(BUF1_REG_16__SCAN_IN), .B1(n19167), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19175) );
  OAI22_X1 U22214 ( .A1(n19172), .A2(n19171), .B1(n19170), .B2(n19169), .ZN(
        n19173) );
  INV_X1 U22215 ( .A(n19173), .ZN(n19174) );
  NAND3_X1 U22216 ( .A1(n19176), .A2(n19175), .A3(n19174), .ZN(P2_U2903) );
  INV_X1 U22217 ( .A(n19177), .ZN(n19180) );
  AOI22_X1 U22218 ( .A1(n19192), .A2(n19178), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19190), .ZN(n19179) );
  OAI21_X1 U22219 ( .B1(n19200), .B2(n19180), .A(n19179), .ZN(P2_U2905) );
  AOI22_X1 U22220 ( .A1(n19192), .A2(n19181), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19190), .ZN(n19182) );
  OAI21_X1 U22221 ( .B1(n19200), .B2(n19183), .A(n19182), .ZN(P2_U2907) );
  AOI22_X1 U22222 ( .A1(n19192), .A2(n19184), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19190), .ZN(n19185) );
  OAI21_X1 U22223 ( .B1(n19200), .B2(n19186), .A(n19185), .ZN(P2_U2909) );
  AOI22_X1 U22224 ( .A1(n19192), .A2(n19187), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19190), .ZN(n19188) );
  OAI21_X1 U22225 ( .B1(n19200), .B2(n19189), .A(n19188), .ZN(P2_U2911) );
  AOI22_X1 U22226 ( .A1(n19192), .A2(n19191), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19190), .ZN(n19198) );
  INV_X1 U22227 ( .A(n19193), .ZN(n19195) );
  NAND3_X1 U22228 ( .A1(n19196), .A2(n19195), .A3(n19194), .ZN(n19197) );
  OAI211_X1 U22229 ( .C1(n19200), .C2(n19199), .A(n19198), .B(n19197), .ZN(
        P2_U2914) );
  OAI21_X1 U22230 ( .B1(n19203), .B2(n19202), .A(n19201), .ZN(n19205) );
  INV_X1 U22231 ( .A(n19204), .ZN(n19972) );
  NOR2_X1 U22232 ( .A1(n19272), .A2(n19207), .ZN(P2_U2920) );
  INV_X2 U22233 ( .A(n19272), .ZN(n19265) );
  AOI22_X1 U22234 ( .A1(n19269), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U22235 ( .B1(n19210), .B2(n19237), .A(n19209), .ZN(P2_U2921) );
  AOI22_X1 U22236 ( .A1(n19269), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19211) );
  OAI21_X1 U22237 ( .B1(n19212), .B2(n19237), .A(n19211), .ZN(P2_U2922) );
  AOI22_X1 U22238 ( .A1(n19269), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U22239 ( .B1(n19214), .B2(n19237), .A(n19213), .ZN(P2_U2923) );
  AOI22_X1 U22240 ( .A1(n19269), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19215) );
  OAI21_X1 U22241 ( .B1(n19216), .B2(n19237), .A(n19215), .ZN(P2_U2924) );
  AOI22_X1 U22242 ( .A1(n19269), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19217) );
  OAI21_X1 U22243 ( .B1(n19218), .B2(n19237), .A(n19217), .ZN(P2_U2925) );
  AOI22_X1 U22244 ( .A1(n19269), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19219) );
  OAI21_X1 U22245 ( .B1(n19220), .B2(n19237), .A(n19219), .ZN(P2_U2926) );
  AOI22_X1 U22246 ( .A1(n19269), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19221) );
  OAI21_X1 U22247 ( .B1(n19222), .B2(n19237), .A(n19221), .ZN(P2_U2927) );
  AOI22_X1 U22248 ( .A1(n19269), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19223) );
  OAI21_X1 U22249 ( .B1(n19224), .B2(n19237), .A(n19223), .ZN(P2_U2928) );
  INV_X1 U22250 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19226) );
  AOI22_X1 U22251 ( .A1(n19269), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19225) );
  OAI21_X1 U22252 ( .B1(n19226), .B2(n19237), .A(n19225), .ZN(P2_U2929) );
  AOI22_X1 U22253 ( .A1(n19269), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19227) );
  OAI21_X1 U22254 ( .B1(n19228), .B2(n19237), .A(n19227), .ZN(P2_U2930) );
  INV_X1 U22255 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19230) );
  AOI22_X1 U22256 ( .A1(n19269), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19229) );
  OAI21_X1 U22257 ( .B1(n19230), .B2(n19237), .A(n19229), .ZN(P2_U2931) );
  AOI22_X1 U22258 ( .A1(n19269), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19231) );
  OAI21_X1 U22259 ( .B1(n19232), .B2(n19237), .A(n19231), .ZN(P2_U2932) );
  INV_X1 U22260 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19234) );
  AOI22_X1 U22261 ( .A1(n19269), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19233) );
  OAI21_X1 U22262 ( .B1(n19234), .B2(n19237), .A(n19233), .ZN(P2_U2933) );
  AOI22_X1 U22263 ( .A1(n19269), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19235) );
  OAI21_X1 U22264 ( .B1(n21133), .B2(n19237), .A(n19235), .ZN(P2_U2934) );
  AOI22_X1 U22265 ( .A1(n19269), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19236) );
  OAI21_X1 U22266 ( .B1(n19238), .B2(n19237), .A(n19236), .ZN(P2_U2935) );
  AOI22_X1 U22267 ( .A1(n19269), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19239) );
  OAI21_X1 U22268 ( .B1(n12991), .B2(n19267), .A(n19239), .ZN(P2_U2936) );
  AOI22_X1 U22269 ( .A1(n19269), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19240) );
  OAI21_X1 U22270 ( .B1(n19241), .B2(n19267), .A(n19240), .ZN(P2_U2937) );
  AOI22_X1 U22271 ( .A1(n19269), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19242) );
  OAI21_X1 U22272 ( .B1(n19243), .B2(n19267), .A(n19242), .ZN(P2_U2938) );
  AOI22_X1 U22273 ( .A1(n19269), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19244) );
  OAI21_X1 U22274 ( .B1(n19245), .B2(n19267), .A(n19244), .ZN(P2_U2939) );
  AOI22_X1 U22275 ( .A1(n19269), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19246) );
  OAI21_X1 U22276 ( .B1(n19247), .B2(n19267), .A(n19246), .ZN(P2_U2940) );
  AOI22_X1 U22277 ( .A1(n19269), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19248) );
  OAI21_X1 U22278 ( .B1(n19249), .B2(n19267), .A(n19248), .ZN(P2_U2941) );
  AOI22_X1 U22279 ( .A1(n19269), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19250) );
  OAI21_X1 U22280 ( .B1(n21085), .B2(n19267), .A(n19250), .ZN(P2_U2942) );
  AOI22_X1 U22281 ( .A1(n19269), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19251) );
  OAI21_X1 U22282 ( .B1(n19252), .B2(n19267), .A(n19251), .ZN(P2_U2943) );
  AOI22_X1 U22283 ( .A1(n19269), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19253) );
  OAI21_X1 U22284 ( .B1(n19254), .B2(n19267), .A(n19253), .ZN(P2_U2944) );
  AOI22_X1 U22285 ( .A1(n19269), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19255) );
  OAI21_X1 U22286 ( .B1(n19256), .B2(n19267), .A(n19255), .ZN(P2_U2945) );
  INV_X1 U22287 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19258) );
  AOI22_X1 U22288 ( .A1(n19269), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19257) );
  OAI21_X1 U22289 ( .B1(n19258), .B2(n19267), .A(n19257), .ZN(P2_U2946) );
  INV_X1 U22290 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19260) );
  AOI22_X1 U22291 ( .A1(n19269), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19259) );
  OAI21_X1 U22292 ( .B1(n19260), .B2(n19267), .A(n19259), .ZN(P2_U2947) );
  INV_X1 U22293 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19262) );
  AOI22_X1 U22294 ( .A1(n19269), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19261) );
  OAI21_X1 U22295 ( .B1(n19262), .B2(n19267), .A(n19261), .ZN(P2_U2948) );
  INV_X1 U22296 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19264) );
  AOI22_X1 U22297 ( .A1(n19269), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19263) );
  OAI21_X1 U22298 ( .B1(n19264), .B2(n19267), .A(n19263), .ZN(P2_U2949) );
  INV_X1 U22299 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19268) );
  AOI22_X1 U22300 ( .A1(n19269), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19265), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19266) );
  OAI21_X1 U22301 ( .B1(n19268), .B2(n19267), .A(n19266), .ZN(P2_U2950) );
  AOI22_X1 U22302 ( .A1(P2_EAX_REG_0__SCAN_IN), .A2(n19270), .B1(n19269), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n19271) );
  OAI21_X1 U22303 ( .B1(n19272), .B2(n21161), .A(n19271), .ZN(P2_U2951) );
  AOI22_X1 U22304 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19275), .B1(n19274), 
        .B2(n19273), .ZN(n19286) );
  NAND2_X1 U22305 ( .A1(n19277), .A2(n19276), .ZN(n19281) );
  NAND2_X1 U22306 ( .A1(n19279), .A2(n19278), .ZN(n19280) );
  OAI211_X1 U22307 ( .C1(n19283), .C2(n19282), .A(n19281), .B(n19280), .ZN(
        n19284) );
  INV_X1 U22308 ( .A(n19284), .ZN(n19285) );
  OAI211_X1 U22309 ( .C1(n19288), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P2_U3010) );
  OAI21_X1 U22310 ( .B1(n19291), .B2(n19290), .A(n19289), .ZN(n19292) );
  OAI211_X1 U22311 ( .C1(n19295), .C2(n19294), .A(n19293), .B(n19292), .ZN(
        n19300) );
  OAI22_X1 U22312 ( .A1(n19298), .A2(n19297), .B1(n10626), .B2(n19296), .ZN(
        n19299) );
  AOI211_X1 U22313 ( .C1(n19301), .C2(n19940), .A(n19300), .B(n19299), .ZN(
        n19305) );
  NAND2_X1 U22314 ( .A1(n19303), .A2(n19302), .ZN(n19304) );
  OAI211_X1 U22315 ( .C1(n19307), .C2(n19306), .A(n19305), .B(n19304), .ZN(
        P2_U3044) );
  AOI22_X1 U22316 ( .A1(n19727), .A2(n19814), .B1(n19774), .B2(n19341), .ZN(
        n19309) );
  AOI22_X1 U22317 ( .A1(n19775), .A2(n19345), .B1(n19378), .B2(n19783), .ZN(
        n19308) );
  OAI211_X1 U22318 ( .C1(n19349), .C2(n19310), .A(n19309), .B(n19308), .ZN(
        P2_U3048) );
  AOI22_X1 U22319 ( .A1(n19789), .A2(n19814), .B1(n19341), .B2(n19787), .ZN(
        n19312) );
  AOI22_X1 U22320 ( .A1(n19788), .A2(n19345), .B1(n19378), .B2(n19737), .ZN(
        n19311) );
  OAI211_X1 U22321 ( .C1(n19349), .C2(n19313), .A(n19312), .B(n19311), .ZN(
        P2_U3049) );
  AOI22_X1 U22322 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19344), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19343), .ZN(n19798) );
  INV_X1 U22323 ( .A(n19798), .ZN(n19741) );
  NOR2_X2 U22324 ( .A1(n10364), .A2(n19339), .ZN(n19793) );
  AOI22_X1 U22325 ( .A1(n19741), .A2(n19814), .B1(n19341), .B2(n19793), .ZN(
        n19318) );
  NAND2_X1 U22326 ( .A1(n19314), .A2(n19777), .ZN(n19744) );
  OAI22_X2 U22327 ( .A1(n19316), .A2(n19335), .B1(n19315), .B2(n19337), .ZN(
        n19795) );
  AOI22_X1 U22328 ( .A1(n19794), .A2(n19345), .B1(n19378), .B2(n19795), .ZN(
        n19317) );
  OAI211_X1 U22329 ( .C1(n19349), .C2(n14211), .A(n19318), .B(n19317), .ZN(
        P2_U3050) );
  INV_X1 U22330 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19325) );
  AOI22_X1 U22331 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19344), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19343), .ZN(n19804) );
  INV_X1 U22332 ( .A(n19804), .ZN(n19745) );
  AOI22_X1 U22333 ( .A1(n19745), .A2(n19814), .B1(n19341), .B2(n19799), .ZN(
        n19324) );
  NOR2_X2 U22334 ( .A1(n19320), .A2(n9793), .ZN(n19800) );
  OAI22_X2 U22335 ( .A1(n19322), .A2(n19335), .B1(n19321), .B2(n19337), .ZN(
        n19801) );
  AOI22_X1 U22336 ( .A1(n19800), .A2(n19345), .B1(n19378), .B2(n19801), .ZN(
        n19323) );
  OAI211_X1 U22337 ( .C1(n19349), .C2(n19325), .A(n19324), .B(n19323), .ZN(
        P2_U3051) );
  AOI22_X1 U22338 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19344), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19343), .ZN(n19810) );
  INV_X1 U22339 ( .A(n19810), .ZN(n19749) );
  NOR2_X2 U22340 ( .A1(n10354), .A2(n19339), .ZN(n19805) );
  AOI22_X1 U22341 ( .A1(n19749), .A2(n19814), .B1(n19341), .B2(n19805), .ZN(
        n19330) );
  NAND2_X1 U22342 ( .A1(n19326), .A2(n19777), .ZN(n19752) );
  OAI22_X2 U22343 ( .A1(n19328), .A2(n19335), .B1(n19327), .B2(n19337), .ZN(
        n19807) );
  AOI22_X1 U22344 ( .A1(n19806), .A2(n19345), .B1(n19378), .B2(n19807), .ZN(
        n19329) );
  OAI211_X1 U22345 ( .C1(n19349), .C2(n19331), .A(n19330), .B(n19329), .ZN(
        P2_U3052) );
  INV_X1 U22346 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19334) );
  AOI22_X1 U22347 ( .A1(n19821), .A2(n19814), .B1(n19341), .B2(n19819), .ZN(
        n19333) );
  AOI22_X1 U22348 ( .A1(n19820), .A2(n19345), .B1(n19378), .B2(n19757), .ZN(
        n19332) );
  OAI211_X1 U22349 ( .C1(n19349), .C2(n19334), .A(n19333), .B(n19332), .ZN(
        P2_U3054) );
  OAI22_X2 U22350 ( .A1(n19338), .A2(n19337), .B1(n19336), .B2(n19335), .ZN(
        n19829) );
  NOR2_X2 U22351 ( .A1(n19340), .A2(n19339), .ZN(n19825) );
  AOI22_X1 U22352 ( .A1(n19829), .A2(n19814), .B1(n19341), .B2(n19825), .ZN(
        n19347) );
  NOR2_X2 U22353 ( .A1(n19342), .A2(n9793), .ZN(n19827) );
  INV_X1 U22354 ( .A(n19835), .ZN(n19762) );
  AOI22_X1 U22355 ( .A1(n19827), .A2(n19345), .B1(n19378), .B2(n19762), .ZN(
        n19346) );
  OAI211_X1 U22356 ( .C1(n19349), .C2(n19348), .A(n19347), .B(n19346), .ZN(
        P2_U3055) );
  NAND2_X1 U22357 ( .A1(n19950), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19572) );
  NOR2_X1 U22358 ( .A1(n19572), .A2(n19406), .ZN(n19376) );
  OR2_X1 U22359 ( .A1(n19376), .A2(n19975), .ZN(n19350) );
  NOR2_X1 U22360 ( .A1(n19351), .A2(n19350), .ZN(n19356) );
  INV_X1 U22361 ( .A(n19357), .ZN(n19352) );
  NOR2_X1 U22362 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19352), .ZN(n19353) );
  NOR3_X2 U22363 ( .A1(n19356), .A2(n19510), .A3(n19353), .ZN(n19377) );
  AOI22_X1 U22364 ( .A1(n19775), .A2(n19377), .B1(n19774), .B2(n19376), .ZN(
        n19361) );
  AND2_X1 U22365 ( .A1(n19354), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19512) );
  NAND2_X1 U22366 ( .A1(n19512), .A2(n19355), .ZN(n19358) );
  AOI21_X1 U22367 ( .B1(n19358), .B2(n19357), .A(n19356), .ZN(n19359) );
  OAI211_X1 U22368 ( .C1(n19376), .C2(n19951), .A(n19359), .B(n19777), .ZN(
        n19379) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19379), .B1(
        n19401), .B2(n19783), .ZN(n19360) );
  OAI211_X1 U22370 ( .C1(n19786), .C2(n19373), .A(n19361), .B(n19360), .ZN(
        P2_U3056) );
  INV_X1 U22371 ( .A(n19401), .ZN(n19382) );
  AOI22_X1 U22372 ( .A1(n19377), .A2(n19788), .B1(n19787), .B2(n19376), .ZN(
        n19363) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19379), .B1(
        n19378), .B2(n19789), .ZN(n19362) );
  OAI211_X1 U22374 ( .C1(n19792), .C2(n19382), .A(n19363), .B(n19362), .ZN(
        P2_U3057) );
  AOI22_X1 U22375 ( .A1(n19794), .A2(n19377), .B1(n19793), .B2(n19376), .ZN(
        n19365) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19379), .B1(
        n19401), .B2(n19795), .ZN(n19364) );
  OAI211_X1 U22377 ( .C1(n19798), .C2(n19373), .A(n19365), .B(n19364), .ZN(
        P2_U3058) );
  AOI22_X1 U22378 ( .A1(n19377), .A2(n19800), .B1(n19799), .B2(n19376), .ZN(
        n19367) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19379), .B1(
        n19401), .B2(n19801), .ZN(n19366) );
  OAI211_X1 U22380 ( .C1(n19804), .C2(n19373), .A(n19367), .B(n19366), .ZN(
        P2_U3059) );
  AOI22_X1 U22381 ( .A1(n19806), .A2(n19377), .B1(n19805), .B2(n19376), .ZN(
        n19369) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19379), .B1(
        n19401), .B2(n19807), .ZN(n19368) );
  OAI211_X1 U22383 ( .C1(n19810), .C2(n19373), .A(n19369), .B(n19368), .ZN(
        P2_U3060) );
  AOI22_X1 U22384 ( .A1(n19377), .A2(n19812), .B1(n19811), .B2(n19376), .ZN(
        n19372) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19379), .B1(
        n19401), .B2(n19813), .ZN(n19371) );
  OAI211_X1 U22386 ( .C1(n19818), .C2(n19373), .A(n19372), .B(n19371), .ZN(
        P2_U3061) );
  AOI22_X1 U22387 ( .A1(n19820), .A2(n19377), .B1(n19819), .B2(n19376), .ZN(
        n19375) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19379), .B1(
        n19378), .B2(n19821), .ZN(n19374) );
  OAI211_X1 U22389 ( .C1(n19824), .C2(n19382), .A(n19375), .B(n19374), .ZN(
        P2_U3062) );
  AOI22_X1 U22390 ( .A1(n19377), .A2(n19827), .B1(n19825), .B2(n19376), .ZN(
        n19381) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19379), .B1(
        n19378), .B2(n19829), .ZN(n19380) );
  OAI211_X1 U22392 ( .C1(n19835), .C2(n19382), .A(n19381), .B(n19380), .ZN(
        P2_U3063) );
  INV_X1 U22393 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n19385) );
  AOI22_X1 U22394 ( .A1(n19400), .A2(n19788), .B1(n19399), .B2(n19787), .ZN(
        n19384) );
  AOI22_X1 U22395 ( .A1(n19401), .A2(n19789), .B1(n19430), .B2(n19737), .ZN(
        n19383) );
  OAI211_X1 U22396 ( .C1(n19405), .C2(n19385), .A(n19384), .B(n19383), .ZN(
        P2_U3065) );
  AOI22_X1 U22397 ( .A1(n19794), .A2(n19400), .B1(n19399), .B2(n19793), .ZN(
        n19387) );
  AOI22_X1 U22398 ( .A1(n19430), .A2(n19795), .B1(n19401), .B2(n19741), .ZN(
        n19386) );
  OAI211_X1 U22399 ( .C1(n19405), .C2(n14210), .A(n19387), .B(n19386), .ZN(
        P2_U3066) );
  INV_X1 U22400 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n19390) );
  AOI22_X1 U22401 ( .A1(n19400), .A2(n19800), .B1(n19399), .B2(n19799), .ZN(
        n19389) );
  AOI22_X1 U22402 ( .A1(n19430), .A2(n19801), .B1(n19401), .B2(n19745), .ZN(
        n19388) );
  OAI211_X1 U22403 ( .C1(n19405), .C2(n19390), .A(n19389), .B(n19388), .ZN(
        P2_U3067) );
  AOI22_X1 U22404 ( .A1(n19806), .A2(n19400), .B1(n19399), .B2(n19805), .ZN(
        n19392) );
  AOI22_X1 U22405 ( .A1(n19430), .A2(n19807), .B1(n19401), .B2(n19749), .ZN(
        n19391) );
  OAI211_X1 U22406 ( .C1(n19405), .C2(n14261), .A(n19392), .B(n19391), .ZN(
        P2_U3068) );
  INV_X1 U22407 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n19395) );
  AOI22_X1 U22408 ( .A1(n19400), .A2(n19812), .B1(n19399), .B2(n19811), .ZN(
        n19394) );
  AOI22_X1 U22409 ( .A1(n19430), .A2(n19813), .B1(n19401), .B2(n19753), .ZN(
        n19393) );
  OAI211_X1 U22410 ( .C1(n19405), .C2(n19395), .A(n19394), .B(n19393), .ZN(
        P2_U3069) );
  INV_X1 U22411 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n19398) );
  AOI22_X1 U22412 ( .A1(n19820), .A2(n19400), .B1(n19399), .B2(n19819), .ZN(
        n19397) );
  AOI22_X1 U22413 ( .A1(n19401), .A2(n19821), .B1(n19430), .B2(n19757), .ZN(
        n19396) );
  OAI211_X1 U22414 ( .C1(n19405), .C2(n19398), .A(n19397), .B(n19396), .ZN(
        P2_U3070) );
  INV_X1 U22415 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19404) );
  AOI22_X1 U22416 ( .A1(n19400), .A2(n19827), .B1(n19399), .B2(n19825), .ZN(
        n19403) );
  AOI22_X1 U22417 ( .A1(n19401), .A2(n19829), .B1(n19430), .B2(n19762), .ZN(
        n19402) );
  OAI211_X1 U22418 ( .C1(n19405), .C2(n19404), .A(n19403), .B(n19402), .ZN(
        P2_U3071) );
  AOI21_X1 U22419 ( .B1(n19512), .B2(n19925), .A(n19722), .ZN(n19412) );
  NOR2_X1 U22420 ( .A1(n19950), .A2(n19406), .ZN(n19410) );
  NOR2_X1 U22421 ( .A1(n19407), .A2(n19406), .ZN(n19429) );
  INV_X1 U22422 ( .A(n19429), .ZN(n19408) );
  AOI21_X1 U22423 ( .B1(n10713), .B2(n19408), .A(n19975), .ZN(n19409) );
  AOI22_X1 U22424 ( .A1(n19727), .A2(n19430), .B1(n19774), .B2(n19429), .ZN(
        n19416) );
  AOI21_X1 U22425 ( .B1(n10713), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19414) );
  INV_X1 U22426 ( .A(n19410), .ZN(n19411) );
  NAND2_X1 U22427 ( .A1(n19412), .A2(n19411), .ZN(n19413) );
  OAI211_X1 U22428 ( .C1(n19429), .C2(n19414), .A(n19413), .B(n19777), .ZN(
        n19431) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19431), .B1(
        n19449), .B2(n19783), .ZN(n19415) );
  OAI211_X1 U22430 ( .C1(n19434), .C2(n19736), .A(n19416), .B(n19415), .ZN(
        P2_U3072) );
  INV_X1 U22431 ( .A(n19788), .ZN(n19740) );
  AOI22_X1 U22432 ( .A1(n19737), .A2(n19449), .B1(n19787), .B2(n19429), .ZN(
        n19418) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19431), .B1(
        n19430), .B2(n19789), .ZN(n19417) );
  OAI211_X1 U22434 ( .C1(n19434), .C2(n19740), .A(n19418), .B(n19417), .ZN(
        P2_U3073) );
  AOI22_X1 U22435 ( .A1(n19795), .A2(n19449), .B1(n19429), .B2(n19793), .ZN(
        n19420) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19431), .B1(
        n19430), .B2(n19741), .ZN(n19419) );
  OAI211_X1 U22437 ( .C1(n19434), .C2(n19744), .A(n19420), .B(n19419), .ZN(
        P2_U3074) );
  INV_X1 U22438 ( .A(n19800), .ZN(n19748) );
  AOI22_X1 U22439 ( .A1(n19801), .A2(n19449), .B1(n19429), .B2(n19799), .ZN(
        n19422) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19431), .B1(
        n19430), .B2(n19745), .ZN(n19421) );
  OAI211_X1 U22441 ( .C1(n19434), .C2(n19748), .A(n19422), .B(n19421), .ZN(
        P2_U3075) );
  AOI22_X1 U22442 ( .A1(n19807), .A2(n19449), .B1(n19429), .B2(n19805), .ZN(
        n19424) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19431), .B1(
        n19430), .B2(n19749), .ZN(n19423) );
  OAI211_X1 U22444 ( .C1(n19434), .C2(n19752), .A(n19424), .B(n19423), .ZN(
        P2_U3076) );
  INV_X1 U22445 ( .A(n19812), .ZN(n19756) );
  AOI22_X1 U22446 ( .A1(n19813), .A2(n19449), .B1(n19811), .B2(n19429), .ZN(
        n19426) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19431), .B1(
        n19430), .B2(n19753), .ZN(n19425) );
  OAI211_X1 U22448 ( .C1(n19434), .C2(n19756), .A(n19426), .B(n19425), .ZN(
        P2_U3077) );
  AOI22_X1 U22449 ( .A1(n19821), .A2(n19430), .B1(n19819), .B2(n19429), .ZN(
        n19428) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19431), .B1(
        n19449), .B2(n19757), .ZN(n19427) );
  OAI211_X1 U22451 ( .C1(n19434), .C2(n19760), .A(n19428), .B(n19427), .ZN(
        P2_U3078) );
  INV_X1 U22452 ( .A(n19827), .ZN(n19767) );
  AOI22_X1 U22453 ( .A1(n19829), .A2(n19430), .B1(n19429), .B2(n19825), .ZN(
        n19433) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19431), .B1(
        n19449), .B2(n19762), .ZN(n19432) );
  OAI211_X1 U22455 ( .C1(n19434), .C2(n19767), .A(n19433), .B(n19432), .ZN(
        P2_U3079) );
  AOI22_X1 U22456 ( .A1(n19448), .A2(n19788), .B1(n19787), .B2(n19447), .ZN(
        n19436) );
  AOI22_X1 U22457 ( .A1(n19449), .A2(n19789), .B1(n19475), .B2(n19737), .ZN(
        n19435) );
  OAI211_X1 U22458 ( .C1(n19452), .C2(n14181), .A(n19436), .B(n19435), .ZN(
        P2_U3081) );
  INV_X1 U22459 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19439) );
  AOI22_X1 U22460 ( .A1(n19794), .A2(n19448), .B1(n19793), .B2(n19447), .ZN(
        n19438) );
  AOI22_X1 U22461 ( .A1(n19475), .A2(n19795), .B1(n19449), .B2(n19741), .ZN(
        n19437) );
  OAI211_X1 U22462 ( .C1(n19452), .C2(n19439), .A(n19438), .B(n19437), .ZN(
        P2_U3082) );
  AOI22_X1 U22463 ( .A1(n19448), .A2(n19800), .B1(n19799), .B2(n19447), .ZN(
        n19441) );
  AOI22_X1 U22464 ( .A1(n19475), .A2(n19801), .B1(n19449), .B2(n19745), .ZN(
        n19440) );
  OAI211_X1 U22465 ( .C1(n19452), .C2(n14239), .A(n19441), .B(n19440), .ZN(
        P2_U3083) );
  INV_X1 U22466 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n19444) );
  AOI22_X1 U22467 ( .A1(n19806), .A2(n19448), .B1(n19805), .B2(n19447), .ZN(
        n19443) );
  AOI22_X1 U22468 ( .A1(n19475), .A2(n19807), .B1(n19449), .B2(n19749), .ZN(
        n19442) );
  OAI211_X1 U22469 ( .C1(n19452), .C2(n19444), .A(n19443), .B(n19442), .ZN(
        P2_U3084) );
  AOI22_X1 U22470 ( .A1(n19820), .A2(n19448), .B1(n19819), .B2(n19447), .ZN(
        n19446) );
  AOI22_X1 U22471 ( .A1(n19449), .A2(n19821), .B1(n19475), .B2(n19757), .ZN(
        n19445) );
  OAI211_X1 U22472 ( .C1(n19452), .C2(n14319), .A(n19446), .B(n19445), .ZN(
        P2_U3086) );
  AOI22_X1 U22473 ( .A1(n19448), .A2(n19827), .B1(n19825), .B2(n19447), .ZN(
        n19451) );
  AOI22_X1 U22474 ( .A1(n19449), .A2(n19829), .B1(n19475), .B2(n19762), .ZN(
        n19450) );
  OAI211_X1 U22475 ( .C1(n19452), .C2(n14149), .A(n19451), .B(n19450), .ZN(
        P2_U3087) );
  INV_X1 U22476 ( .A(n19696), .ZN(n19694) );
  AOI21_X1 U22477 ( .B1(n19512), .B2(n19694), .A(n19722), .ZN(n19459) );
  INV_X1 U22478 ( .A(n19458), .ZN(n19454) );
  NOR2_X1 U22479 ( .A1(n19958), .A2(n19458), .ZN(n19480) );
  INV_X1 U22480 ( .A(n19480), .ZN(n19455) );
  AOI21_X1 U22481 ( .B1(n19456), .B2(n19455), .A(n19975), .ZN(n19453) );
  AOI22_X1 U22482 ( .A1(n19783), .A2(n19505), .B1(n19774), .B2(n19480), .ZN(
        n19462) );
  AND2_X1 U22483 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19455), .ZN(n19457) );
  AOI22_X1 U22484 ( .A1(n19459), .A2(n19458), .B1(n19457), .B2(n19456), .ZN(
        n19460) );
  OAI211_X1 U22485 ( .C1(n19480), .C2(n19951), .A(n19460), .B(n19777), .ZN(
        n19476) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19476), .B1(
        n19475), .B2(n19727), .ZN(n19461) );
  OAI211_X1 U22487 ( .C1(n19479), .C2(n19736), .A(n19462), .B(n19461), .ZN(
        P2_U3088) );
  AOI22_X1 U22488 ( .A1(n19789), .A2(n19475), .B1(n19787), .B2(n19480), .ZN(
        n19464) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19476), .B1(
        n19505), .B2(n19737), .ZN(n19463) );
  OAI211_X1 U22490 ( .C1(n19479), .C2(n19740), .A(n19464), .B(n19463), .ZN(
        P2_U3089) );
  AOI22_X1 U22491 ( .A1(n19795), .A2(n19505), .B1(n19480), .B2(n19793), .ZN(
        n19466) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19476), .B1(
        n19475), .B2(n19741), .ZN(n19465) );
  OAI211_X1 U22493 ( .C1(n19479), .C2(n19744), .A(n19466), .B(n19465), .ZN(
        P2_U3090) );
  AOI22_X1 U22494 ( .A1(n19745), .A2(n19475), .B1(n19480), .B2(n19799), .ZN(
        n19468) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19476), .B1(
        n19505), .B2(n19801), .ZN(n19467) );
  OAI211_X1 U22496 ( .C1(n19479), .C2(n19748), .A(n19468), .B(n19467), .ZN(
        P2_U3091) );
  AOI22_X1 U22497 ( .A1(n19749), .A2(n19475), .B1(n19480), .B2(n19805), .ZN(
        n19470) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19476), .B1(
        n19505), .B2(n19807), .ZN(n19469) );
  OAI211_X1 U22499 ( .C1(n19479), .C2(n19752), .A(n19470), .B(n19469), .ZN(
        P2_U3092) );
  AOI22_X1 U22500 ( .A1(n19753), .A2(n19475), .B1(n19811), .B2(n19480), .ZN(
        n19472) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19476), .B1(
        n19505), .B2(n19813), .ZN(n19471) );
  OAI211_X1 U22502 ( .C1(n19479), .C2(n19756), .A(n19472), .B(n19471), .ZN(
        P2_U3093) );
  AOI22_X1 U22503 ( .A1(n19757), .A2(n19505), .B1(n19819), .B2(n19480), .ZN(
        n19474) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19476), .B1(
        n19475), .B2(n19821), .ZN(n19473) );
  OAI211_X1 U22505 ( .C1(n19479), .C2(n19760), .A(n19474), .B(n19473), .ZN(
        P2_U3094) );
  AOI22_X1 U22506 ( .A1(n19829), .A2(n19475), .B1(n19480), .B2(n19825), .ZN(
        n19478) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19476), .B1(
        n19505), .B2(n19762), .ZN(n19477) );
  OAI211_X1 U22508 ( .C1(n19479), .C2(n19767), .A(n19478), .B(n19477), .ZN(
        P2_U3095) );
  NOR2_X1 U22509 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19724), .ZN(
        n19517) );
  INV_X1 U22510 ( .A(n19517), .ZN(n19511) );
  NOR2_X1 U22511 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19511), .ZN(
        n19503) );
  NOR2_X1 U22512 ( .A1(n19480), .A2(n19503), .ZN(n19485) );
  OAI21_X1 U22513 ( .B1(n19481), .B2(n19503), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19482) );
  OAI21_X1 U22514 ( .B1(n19485), .B2(n19722), .A(n19482), .ZN(n19504) );
  AOI22_X1 U22515 ( .A1(n19775), .A2(n19504), .B1(n19774), .B2(n19503), .ZN(
        n19489) );
  OAI21_X1 U22516 ( .B1(n19505), .B2(n19535), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19486) );
  AOI211_X1 U22517 ( .C1(n19481), .C2(n19951), .A(n19503), .B(n19924), .ZN(
        n19484) );
  AOI211_X1 U22518 ( .C1(n19486), .C2(n19485), .A(n9793), .B(n19484), .ZN(
        n19487) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19506), .B1(
        n19535), .B2(n19783), .ZN(n19488) );
  OAI211_X1 U22520 ( .C1(n19786), .C2(n19500), .A(n19489), .B(n19488), .ZN(
        P2_U3096) );
  AOI22_X1 U22521 ( .A1(n19504), .A2(n19788), .B1(n19787), .B2(n19503), .ZN(
        n19491) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19789), .ZN(n19490) );
  OAI211_X1 U22523 ( .C1(n19792), .C2(n19531), .A(n19491), .B(n19490), .ZN(
        P2_U3097) );
  AOI22_X1 U22524 ( .A1(n19794), .A2(n19504), .B1(n19793), .B2(n19503), .ZN(
        n19493) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19506), .B1(
        n19535), .B2(n19795), .ZN(n19492) );
  OAI211_X1 U22526 ( .C1(n19798), .C2(n19500), .A(n19493), .B(n19492), .ZN(
        P2_U3098) );
  AOI22_X1 U22527 ( .A1(n19504), .A2(n19800), .B1(n19799), .B2(n19503), .ZN(
        n19495) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19506), .B1(
        n19535), .B2(n19801), .ZN(n19494) );
  OAI211_X1 U22529 ( .C1(n19804), .C2(n19500), .A(n19495), .B(n19494), .ZN(
        P2_U3099) );
  AOI22_X1 U22530 ( .A1(n19806), .A2(n19504), .B1(n19805), .B2(n19503), .ZN(
        n19497) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19506), .B1(
        n19535), .B2(n19807), .ZN(n19496) );
  OAI211_X1 U22532 ( .C1(n19810), .C2(n19500), .A(n19497), .B(n19496), .ZN(
        P2_U3100) );
  AOI22_X1 U22533 ( .A1(n19504), .A2(n19812), .B1(n19811), .B2(n19503), .ZN(
        n19499) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19506), .B1(
        n19535), .B2(n19813), .ZN(n19498) );
  OAI211_X1 U22535 ( .C1(n19818), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        P2_U3101) );
  AOI22_X1 U22536 ( .A1(n19820), .A2(n19504), .B1(n19819), .B2(n19503), .ZN(
        n19502) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19821), .ZN(n19501) );
  OAI211_X1 U22538 ( .C1(n19824), .C2(n19531), .A(n19502), .B(n19501), .ZN(
        P2_U3102) );
  AOI22_X1 U22539 ( .A1(n19504), .A2(n19827), .B1(n19825), .B2(n19503), .ZN(
        n19508) );
  AOI22_X1 U22540 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19829), .ZN(n19507) );
  OAI211_X1 U22541 ( .C1(n19835), .C2(n19531), .A(n19508), .B(n19507), .ZN(
        P2_U3103) );
  NOR2_X1 U22542 ( .A1(n19958), .A2(n19511), .ZN(n19545) );
  INV_X1 U22543 ( .A(n19545), .ZN(n19542) );
  NAND2_X1 U22544 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19542), .ZN(n19509) );
  NOR2_X1 U22545 ( .A1(n10717), .A2(n19509), .ZN(n19515) );
  AOI211_X2 U22546 ( .C1(n19511), .C2(n19975), .A(n19510), .B(n19515), .ZN(
        n19534) );
  AOI22_X1 U22547 ( .A1(n19534), .A2(n19775), .B1(n19774), .B2(n19545), .ZN(
        n19520) );
  AND2_X1 U22548 ( .A1(n19512), .A2(n19781), .ZN(n19923) );
  AND2_X1 U22549 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19542), .ZN(n19513) );
  OR2_X1 U22550 ( .A1(n9793), .A2(n19513), .ZN(n19514) );
  NOR2_X1 U22551 ( .A1(n19515), .A2(n19514), .ZN(n19516) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19536), .B1(
        n19565), .B2(n19783), .ZN(n19519) );
  OAI211_X1 U22553 ( .C1(n19786), .C2(n19531), .A(n19520), .B(n19519), .ZN(
        P2_U3104) );
  AOI22_X1 U22554 ( .A1(n19534), .A2(n19788), .B1(n19787), .B2(n19545), .ZN(
        n19522) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19536), .B1(
        n19535), .B2(n19789), .ZN(n19521) );
  OAI211_X1 U22556 ( .C1(n19792), .C2(n19561), .A(n19522), .B(n19521), .ZN(
        P2_U3105) );
  AOI22_X1 U22557 ( .A1(n19534), .A2(n19794), .B1(n19793), .B2(n19545), .ZN(
        n19524) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19536), .B1(
        n19565), .B2(n19795), .ZN(n19523) );
  OAI211_X1 U22559 ( .C1(n19798), .C2(n19531), .A(n19524), .B(n19523), .ZN(
        P2_U3106) );
  AOI22_X1 U22560 ( .A1(n19534), .A2(n19800), .B1(n19799), .B2(n19545), .ZN(
        n19526) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19536), .B1(
        n19565), .B2(n19801), .ZN(n19525) );
  OAI211_X1 U22562 ( .C1(n19804), .C2(n19531), .A(n19526), .B(n19525), .ZN(
        P2_U3107) );
  AOI22_X1 U22563 ( .A1(n19534), .A2(n19806), .B1(n19805), .B2(n19545), .ZN(
        n19528) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19536), .B1(
        n19565), .B2(n19807), .ZN(n19527) );
  OAI211_X1 U22565 ( .C1(n19810), .C2(n19531), .A(n19528), .B(n19527), .ZN(
        P2_U3108) );
  AOI22_X1 U22566 ( .A1(n19534), .A2(n19812), .B1(n19811), .B2(n19545), .ZN(
        n19530) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19536), .B1(
        n19565), .B2(n19813), .ZN(n19529) );
  OAI211_X1 U22568 ( .C1(n19818), .C2(n19531), .A(n19530), .B(n19529), .ZN(
        P2_U3109) );
  AOI22_X1 U22569 ( .A1(n19534), .A2(n19820), .B1(n19819), .B2(n19545), .ZN(
        n19533) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19536), .B1(
        n19535), .B2(n19821), .ZN(n19532) );
  OAI211_X1 U22571 ( .C1(n19824), .C2(n19561), .A(n19533), .B(n19532), .ZN(
        P2_U3110) );
  AOI22_X1 U22572 ( .A1(n19534), .A2(n19827), .B1(n19825), .B2(n19545), .ZN(
        n19538) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19536), .B1(
        n19535), .B2(n19829), .ZN(n19537) );
  OAI211_X1 U22574 ( .C1(n19835), .C2(n19561), .A(n19538), .B(n19537), .ZN(
        P2_U3111) );
  NAND2_X1 U22575 ( .A1(n19539), .A2(n19950), .ZN(n19580) );
  NOR2_X1 U22576 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19580), .ZN(
        n19564) );
  AOI22_X1 U22577 ( .A1(n19783), .A2(n19598), .B1(n19774), .B2(n19564), .ZN(
        n19550) );
  AOI21_X1 U22578 ( .B1(n19540), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19722), 
        .ZN(n19544) );
  OAI21_X1 U22579 ( .B1(n19546), .B2(n19975), .A(n19951), .ZN(n19541) );
  AOI21_X1 U22580 ( .B1(n19544), .B2(n19542), .A(n19541), .ZN(n19543) );
  OAI21_X1 U22581 ( .B1(n19564), .B2(n19545), .A(n19544), .ZN(n19548) );
  OAI21_X1 U22582 ( .B1(n19546), .B2(n19564), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19547) );
  NAND2_X1 U22583 ( .A1(n19548), .A2(n19547), .ZN(n19566) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19567), .B1(
        n19775), .B2(n19566), .ZN(n19549) );
  OAI211_X1 U22585 ( .C1(n19786), .C2(n19561), .A(n19550), .B(n19549), .ZN(
        P2_U3112) );
  INV_X1 U22586 ( .A(n19598), .ZN(n19570) );
  AOI22_X1 U22587 ( .A1(n19789), .A2(n19565), .B1(n19787), .B2(n19564), .ZN(
        n19552) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19788), .ZN(n19551) );
  OAI211_X1 U22589 ( .C1(n19792), .C2(n19570), .A(n19552), .B(n19551), .ZN(
        P2_U3113) );
  AOI22_X1 U22590 ( .A1(n19795), .A2(n19598), .B1(n19793), .B2(n19564), .ZN(
        n19554) );
  AOI22_X1 U22591 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19794), .ZN(n19553) );
  OAI211_X1 U22592 ( .C1(n19798), .C2(n19561), .A(n19554), .B(n19553), .ZN(
        P2_U3114) );
  AOI22_X1 U22593 ( .A1(n19801), .A2(n19598), .B1(n19799), .B2(n19564), .ZN(
        n19556) );
  AOI22_X1 U22594 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19800), .ZN(n19555) );
  OAI211_X1 U22595 ( .C1(n19804), .C2(n19561), .A(n19556), .B(n19555), .ZN(
        P2_U3115) );
  AOI22_X1 U22596 ( .A1(n19807), .A2(n19598), .B1(n19805), .B2(n19564), .ZN(
        n19558) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19806), .ZN(n19557) );
  OAI211_X1 U22598 ( .C1(n19810), .C2(n19561), .A(n19558), .B(n19557), .ZN(
        P2_U3116) );
  AOI22_X1 U22599 ( .A1(n19813), .A2(n19598), .B1(n19811), .B2(n19564), .ZN(
        n19560) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19812), .ZN(n19559) );
  OAI211_X1 U22601 ( .C1(n19818), .C2(n19561), .A(n19560), .B(n19559), .ZN(
        P2_U3117) );
  AOI22_X1 U22602 ( .A1(n19821), .A2(n19565), .B1(n19819), .B2(n19564), .ZN(
        n19563) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19820), .ZN(n19562) );
  OAI211_X1 U22604 ( .C1(n19824), .C2(n19570), .A(n19563), .B(n19562), .ZN(
        P2_U3118) );
  AOI22_X1 U22605 ( .A1(n19829), .A2(n19565), .B1(n19564), .B2(n19825), .ZN(
        n19569) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19567), .B1(
        n19566), .B2(n19827), .ZN(n19568) );
  OAI211_X1 U22607 ( .C1(n19835), .C2(n19570), .A(n19569), .B(n19568), .ZN(
        P2_U3119) );
  OAI21_X1 U22608 ( .B1(n19689), .B2(n19577), .A(n19924), .ZN(n19581) );
  INV_X1 U22609 ( .A(n19580), .ZN(n19571) );
  OR2_X1 U22610 ( .A1(n19581), .A2(n19571), .ZN(n19576) );
  NAND2_X1 U22611 ( .A1(n10701), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19573) );
  NOR2_X1 U22612 ( .A1(n19572), .A2(n19607), .ZN(n19608) );
  AOI21_X1 U22613 ( .B1(n19573), .B2(n19951), .A(n19608), .ZN(n19574) );
  NOR2_X1 U22614 ( .A1(n9793), .A2(n19574), .ZN(n19575) );
  AOI22_X1 U22615 ( .A1(n19783), .A2(n19633), .B1(n19774), .B2(n19608), .ZN(
        n19583) );
  INV_X1 U22616 ( .A(n10701), .ZN(n19578) );
  OAI21_X1 U22617 ( .B1(n19578), .B2(n19608), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19579) );
  OAI21_X1 U22618 ( .B1(n19581), .B2(n19580), .A(n19579), .ZN(n19600) );
  AOI22_X1 U22619 ( .A1(n19775), .A2(n19600), .B1(n19598), .B2(n19727), .ZN(
        n19582) );
  OAI211_X1 U22620 ( .C1(n19599), .C2(n19584), .A(n19583), .B(n19582), .ZN(
        P2_U3120) );
  AOI22_X1 U22621 ( .A1(n19737), .A2(n19633), .B1(n19787), .B2(n19608), .ZN(
        n19586) );
  AOI22_X1 U22622 ( .A1(n19598), .A2(n19789), .B1(n19788), .B2(n19600), .ZN(
        n19585) );
  OAI211_X1 U22623 ( .C1(n19599), .C2(n14191), .A(n19586), .B(n19585), .ZN(
        P2_U3121) );
  INV_X1 U22624 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n21162) );
  AOI22_X1 U22625 ( .A1(n19741), .A2(n19598), .B1(n19793), .B2(n19608), .ZN(
        n19588) );
  AOI22_X1 U22626 ( .A1(n19794), .A2(n19600), .B1(n19633), .B2(n19795), .ZN(
        n19587) );
  OAI211_X1 U22627 ( .C1(n19599), .C2(n21162), .A(n19588), .B(n19587), .ZN(
        P2_U3122) );
  AOI22_X1 U22628 ( .A1(n19745), .A2(n19598), .B1(n19799), .B2(n19608), .ZN(
        n19590) );
  AOI22_X1 U22629 ( .A1(n19800), .A2(n19600), .B1(n19633), .B2(n19801), .ZN(
        n19589) );
  OAI211_X1 U22630 ( .C1(n19599), .C2(n14249), .A(n19590), .B(n19589), .ZN(
        P2_U3123) );
  INV_X1 U22631 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n19593) );
  AOI22_X1 U22632 ( .A1(n19807), .A2(n19633), .B1(n19805), .B2(n19608), .ZN(
        n19592) );
  AOI22_X1 U22633 ( .A1(n19598), .A2(n19749), .B1(n19806), .B2(n19600), .ZN(
        n19591) );
  OAI211_X1 U22634 ( .C1(n19599), .C2(n19593), .A(n19592), .B(n19591), .ZN(
        P2_U3124) );
  AOI22_X1 U22635 ( .A1(n19813), .A2(n19633), .B1(n19811), .B2(n19608), .ZN(
        n19595) );
  AOI22_X1 U22636 ( .A1(n19598), .A2(n19753), .B1(n19812), .B2(n19600), .ZN(
        n19594) );
  OAI211_X1 U22637 ( .C1(n19599), .C2(n14306), .A(n19595), .B(n19594), .ZN(
        P2_U3125) );
  AOI22_X1 U22638 ( .A1(n19757), .A2(n19633), .B1(n19819), .B2(n19608), .ZN(
        n19597) );
  AOI22_X1 U22639 ( .A1(n19598), .A2(n19821), .B1(n19820), .B2(n19600), .ZN(
        n19596) );
  OAI211_X1 U22640 ( .C1(n19599), .C2(n14327), .A(n19597), .B(n19596), .ZN(
        P2_U3126) );
  AOI22_X1 U22641 ( .A1(n19829), .A2(n19598), .B1(n19825), .B2(n19608), .ZN(
        n19603) );
  INV_X1 U22642 ( .A(n19599), .ZN(n19601) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19601), .B1(
        n19827), .B2(n19600), .ZN(n19602) );
  OAI211_X1 U22644 ( .C1(n19835), .C2(n19628), .A(n19603), .B(n19602), .ZN(
        P2_U3127) );
  INV_X1 U22645 ( .A(n10726), .ZN(n19611) );
  NOR2_X1 U22646 ( .A1(n19604), .A2(n19607), .ZN(n19631) );
  OAI21_X1 U22647 ( .B1(n19611), .B2(n19631), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19605) );
  OAI21_X1 U22648 ( .B1(n19607), .B2(n19606), .A(n19605), .ZN(n19632) );
  AOI22_X1 U22649 ( .A1(n19775), .A2(n19632), .B1(n19774), .B2(n19631), .ZN(
        n19617) );
  OAI21_X1 U22650 ( .B1(n19653), .B2(n19633), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19610) );
  INV_X1 U22651 ( .A(n19608), .ZN(n19609) );
  AOI21_X1 U22652 ( .B1(n19610), .B2(n19609), .A(n19722), .ZN(n19615) );
  NAND3_X1 U22653 ( .A1(n19611), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19951), 
        .ZN(n19613) );
  INV_X1 U22654 ( .A(n19631), .ZN(n19612) );
  NAND2_X1 U22655 ( .A1(n19613), .A2(n19612), .ZN(n19614) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19634), .B1(
        n19653), .B2(n19783), .ZN(n19616) );
  OAI211_X1 U22657 ( .C1(n19786), .C2(n19628), .A(n19617), .B(n19616), .ZN(
        P2_U3128) );
  AOI22_X1 U22658 ( .A1(n19632), .A2(n19788), .B1(n19787), .B2(n19631), .ZN(
        n19619) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19634), .B1(
        n19633), .B2(n19789), .ZN(n19618) );
  OAI211_X1 U22660 ( .C1(n19792), .C2(n19650), .A(n19619), .B(n19618), .ZN(
        P2_U3129) );
  AOI22_X1 U22661 ( .A1(n19794), .A2(n19632), .B1(n19793), .B2(n19631), .ZN(
        n19621) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19634), .B1(
        n19653), .B2(n19795), .ZN(n19620) );
  OAI211_X1 U22663 ( .C1(n19798), .C2(n19628), .A(n19621), .B(n19620), .ZN(
        P2_U3130) );
  AOI22_X1 U22664 ( .A1(n19632), .A2(n19800), .B1(n19799), .B2(n19631), .ZN(
        n19623) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19634), .B1(
        n19653), .B2(n19801), .ZN(n19622) );
  OAI211_X1 U22666 ( .C1(n19804), .C2(n19628), .A(n19623), .B(n19622), .ZN(
        P2_U3131) );
  AOI22_X1 U22667 ( .A1(n19806), .A2(n19632), .B1(n19805), .B2(n19631), .ZN(
        n19625) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19634), .B1(
        n19653), .B2(n19807), .ZN(n19624) );
  OAI211_X1 U22669 ( .C1(n19810), .C2(n19628), .A(n19625), .B(n19624), .ZN(
        P2_U3132) );
  AOI22_X1 U22670 ( .A1(n19632), .A2(n19812), .B1(n19811), .B2(n19631), .ZN(
        n19627) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19634), .B1(
        n19653), .B2(n19813), .ZN(n19626) );
  OAI211_X1 U22672 ( .C1(n19818), .C2(n19628), .A(n19627), .B(n19626), .ZN(
        P2_U3133) );
  AOI22_X1 U22673 ( .A1(n19820), .A2(n19632), .B1(n19819), .B2(n19631), .ZN(
        n19630) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19634), .B1(
        n19633), .B2(n19821), .ZN(n19629) );
  OAI211_X1 U22675 ( .C1(n19824), .C2(n19650), .A(n19630), .B(n19629), .ZN(
        P2_U3134) );
  AOI22_X1 U22676 ( .A1(n19632), .A2(n19827), .B1(n19825), .B2(n19631), .ZN(
        n19636) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19634), .B1(
        n19633), .B2(n19829), .ZN(n19635) );
  OAI211_X1 U22678 ( .C1(n19835), .C2(n19650), .A(n19636), .B(n19635), .ZN(
        P2_U3135) );
  INV_X1 U22679 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n19640) );
  INV_X1 U22680 ( .A(n19637), .ZN(n19651) );
  AOI22_X1 U22681 ( .A1(n19775), .A2(n19652), .B1(n19774), .B2(n19651), .ZN(
        n19639) );
  AOI22_X1 U22682 ( .A1(n19681), .A2(n19783), .B1(n19653), .B2(n19727), .ZN(
        n19638) );
  OAI211_X1 U22683 ( .C1(n19641), .C2(n19640), .A(n19639), .B(n19638), .ZN(
        P2_U3136) );
  AOI22_X1 U22684 ( .A1(n19794), .A2(n19652), .B1(n19651), .B2(n19793), .ZN(
        n19643) );
  AOI22_X1 U22685 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19654), .B1(
        n19681), .B2(n19795), .ZN(n19642) );
  OAI211_X1 U22686 ( .C1(n19798), .C2(n19650), .A(n19643), .B(n19642), .ZN(
        P2_U3138) );
  AOI22_X1 U22687 ( .A1(n19652), .A2(n19800), .B1(n19651), .B2(n19799), .ZN(
        n19645) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19654), .B1(
        n19681), .B2(n19801), .ZN(n19644) );
  OAI211_X1 U22689 ( .C1(n19804), .C2(n19650), .A(n19645), .B(n19644), .ZN(
        P2_U3139) );
  AOI22_X1 U22690 ( .A1(n19806), .A2(n19652), .B1(n19651), .B2(n19805), .ZN(
        n19647) );
  AOI22_X1 U22691 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19654), .B1(
        n19681), .B2(n19807), .ZN(n19646) );
  OAI211_X1 U22692 ( .C1(n19810), .C2(n19650), .A(n19647), .B(n19646), .ZN(
        P2_U3140) );
  AOI22_X1 U22693 ( .A1(n19652), .A2(n19812), .B1(n19811), .B2(n19651), .ZN(
        n19649) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19654), .B1(
        n19681), .B2(n19813), .ZN(n19648) );
  OAI211_X1 U22695 ( .C1(n19818), .C2(n19650), .A(n19649), .B(n19648), .ZN(
        P2_U3141) );
  AOI22_X1 U22696 ( .A1(n19652), .A2(n19827), .B1(n19651), .B2(n19825), .ZN(
        n19656) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19654), .B1(
        n19653), .B2(n19829), .ZN(n19655) );
  OAI211_X1 U22698 ( .C1(n19835), .C2(n19676), .A(n19656), .B(n19655), .ZN(
        P2_U3143) );
  NAND2_X1 U22699 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19657), .ZN(
        n19661) );
  NAND3_X1 U22700 ( .A1(n19950), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19688) );
  NOR2_X1 U22701 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19688), .ZN(
        n19679) );
  OAI21_X1 U22702 ( .B1(n19659), .B2(n19679), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19658) );
  OAI21_X1 U22703 ( .B1(n19661), .B2(n19722), .A(n19658), .ZN(n19680) );
  AOI22_X1 U22704 ( .A1(n19775), .A2(n19680), .B1(n19774), .B2(n19679), .ZN(
        n19665) );
  OAI21_X1 U22705 ( .B1(n19681), .B2(n19715), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19662) );
  AOI211_X1 U22706 ( .C1(n19659), .C2(n19951), .A(n19679), .B(n19924), .ZN(
        n19660) );
  AOI211_X1 U22707 ( .C1(n19662), .C2(n19661), .A(n9793), .B(n19660), .ZN(
        n19663) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19682), .B1(
        n19715), .B2(n19783), .ZN(n19664) );
  OAI211_X1 U22709 ( .C1(n19786), .C2(n19676), .A(n19665), .B(n19664), .ZN(
        P2_U3144) );
  AOI22_X1 U22710 ( .A1(n19680), .A2(n19788), .B1(n19787), .B2(n19679), .ZN(
        n19667) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19682), .B1(
        n19681), .B2(n19789), .ZN(n19666) );
  OAI211_X1 U22712 ( .C1(n19792), .C2(n19710), .A(n19667), .B(n19666), .ZN(
        P2_U3145) );
  AOI22_X1 U22713 ( .A1(n19794), .A2(n19680), .B1(n19793), .B2(n19679), .ZN(
        n19669) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19682), .B1(
        n19715), .B2(n19795), .ZN(n19668) );
  OAI211_X1 U22715 ( .C1(n19798), .C2(n19676), .A(n19669), .B(n19668), .ZN(
        P2_U3146) );
  AOI22_X1 U22716 ( .A1(n19680), .A2(n19800), .B1(n19799), .B2(n19679), .ZN(
        n19671) );
  AOI22_X1 U22717 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19682), .B1(
        n19715), .B2(n19801), .ZN(n19670) );
  OAI211_X1 U22718 ( .C1(n19804), .C2(n19676), .A(n19671), .B(n19670), .ZN(
        P2_U3147) );
  AOI22_X1 U22719 ( .A1(n19806), .A2(n19680), .B1(n19805), .B2(n19679), .ZN(
        n19673) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19682), .B1(
        n19715), .B2(n19807), .ZN(n19672) );
  OAI211_X1 U22721 ( .C1(n19810), .C2(n19676), .A(n19673), .B(n19672), .ZN(
        P2_U3148) );
  AOI22_X1 U22722 ( .A1(n19680), .A2(n19812), .B1(n19811), .B2(n19679), .ZN(
        n19675) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19682), .B1(
        n19715), .B2(n19813), .ZN(n19674) );
  OAI211_X1 U22724 ( .C1(n19818), .C2(n19676), .A(n19675), .B(n19674), .ZN(
        P2_U3149) );
  AOI22_X1 U22725 ( .A1(n19820), .A2(n19680), .B1(n19819), .B2(n19679), .ZN(
        n19678) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19682), .B1(
        n19681), .B2(n19821), .ZN(n19677) );
  OAI211_X1 U22727 ( .C1(n19824), .C2(n19710), .A(n19678), .B(n19677), .ZN(
        P2_U3150) );
  AOI22_X1 U22728 ( .A1(n19680), .A2(n19827), .B1(n19825), .B2(n19679), .ZN(
        n19684) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19682), .B1(
        n19681), .B2(n19829), .ZN(n19683) );
  OAI211_X1 U22730 ( .C1(n19835), .C2(n19710), .A(n19684), .B(n19683), .ZN(
        P2_U3151) );
  NOR2_X1 U22731 ( .A1(n19958), .A2(n19688), .ZN(n19713) );
  INV_X1 U22732 ( .A(n19713), .ZN(n19728) );
  AND2_X1 U22733 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19728), .ZN(n19685) );
  NAND2_X1 U22734 ( .A1(n19686), .A2(n19685), .ZN(n19690) );
  OAI21_X1 U22735 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19688), .A(n19975), 
        .ZN(n19687) );
  AND2_X1 U22736 ( .A1(n19690), .A2(n19687), .ZN(n19714) );
  AOI22_X1 U22737 ( .A1(n19775), .A2(n19714), .B1(n19774), .B2(n19713), .ZN(
        n19699) );
  INV_X1 U22738 ( .A(n19688), .ZN(n19695) );
  INV_X1 U22739 ( .A(n19689), .ZN(n19780) );
  INV_X1 U22740 ( .A(n19690), .ZN(n19692) );
  AOI211_X1 U22741 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19728), .A(n19692), 
        .B(n9793), .ZN(n19693) );
  OAI221_X1 U22742 ( .B1(n19695), .B2(n19694), .C1(n19695), .C2(n19780), .A(
        n19693), .ZN(n19716) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19716), .B1(
        n19763), .B2(n19783), .ZN(n19698) );
  OAI211_X1 U22744 ( .C1(n19786), .C2(n19710), .A(n19699), .B(n19698), .ZN(
        P2_U3152) );
  AOI22_X1 U22745 ( .A1(n19714), .A2(n19788), .B1(n19787), .B2(n19713), .ZN(
        n19701) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19789), .ZN(n19700) );
  OAI211_X1 U22747 ( .C1(n19792), .C2(n19721), .A(n19701), .B(n19700), .ZN(
        P2_U3153) );
  AOI22_X1 U22748 ( .A1(n19794), .A2(n19714), .B1(n19793), .B2(n19713), .ZN(
        n19703) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19716), .B1(
        n19763), .B2(n19795), .ZN(n19702) );
  OAI211_X1 U22750 ( .C1(n19798), .C2(n19710), .A(n19703), .B(n19702), .ZN(
        P2_U3154) );
  AOI22_X1 U22751 ( .A1(n19714), .A2(n19800), .B1(n19799), .B2(n19713), .ZN(
        n19705) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19716), .B1(
        n19763), .B2(n19801), .ZN(n19704) );
  OAI211_X1 U22753 ( .C1(n19804), .C2(n19710), .A(n19705), .B(n19704), .ZN(
        P2_U3155) );
  AOI22_X1 U22754 ( .A1(n19806), .A2(n19714), .B1(n19805), .B2(n19713), .ZN(
        n19707) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19716), .B1(
        n19763), .B2(n19807), .ZN(n19706) );
  OAI211_X1 U22756 ( .C1(n19810), .C2(n19710), .A(n19707), .B(n19706), .ZN(
        P2_U3156) );
  AOI22_X1 U22757 ( .A1(n19714), .A2(n19812), .B1(n19811), .B2(n19713), .ZN(
        n19709) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19716), .B1(
        n19763), .B2(n19813), .ZN(n19708) );
  OAI211_X1 U22759 ( .C1(n19818), .C2(n19710), .A(n19709), .B(n19708), .ZN(
        P2_U3157) );
  AOI22_X1 U22760 ( .A1(n19820), .A2(n19714), .B1(n19819), .B2(n19713), .ZN(
        n19712) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19821), .ZN(n19711) );
  OAI211_X1 U22762 ( .C1(n19824), .C2(n19721), .A(n19712), .B(n19711), .ZN(
        P2_U3158) );
  AOI22_X1 U22763 ( .A1(n19714), .A2(n19827), .B1(n19825), .B2(n19713), .ZN(
        n19718) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19829), .ZN(n19717) );
  OAI211_X1 U22765 ( .C1(n19835), .C2(n19721), .A(n19718), .B(n19717), .ZN(
        P2_U3159) );
  NAND2_X1 U22766 ( .A1(n19817), .A2(n19721), .ZN(n19723) );
  AOI21_X1 U22767 ( .B1(n19723), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19722), 
        .ZN(n19729) );
  NOR2_X1 U22768 ( .A1(n19935), .A2(n19724), .ZN(n19782) );
  INV_X1 U22769 ( .A(n19782), .ZN(n19771) );
  NOR2_X1 U22770 ( .A1(n19771), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19761) );
  INV_X1 U22771 ( .A(n19761), .ZN(n19730) );
  NAND2_X1 U22772 ( .A1(n19730), .A2(n19728), .ZN(n19726) );
  AOI21_X1 U22773 ( .B1(n19731), .B2(n19730), .A(n19975), .ZN(n19725) );
  AOI22_X1 U22774 ( .A1(n19727), .A2(n19763), .B1(n19774), .B2(n19761), .ZN(
        n19735) );
  OAI221_X1 U22775 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19729), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19728), .A(n19730), .ZN(n19733) );
  NAND3_X1 U22776 ( .A1(n19731), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19730), 
        .ZN(n19732) );
  NAND3_X1 U22777 ( .A1(n19733), .A2(n19777), .A3(n19732), .ZN(n19764) );
  AOI22_X1 U22778 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19764), .B1(
        n19830), .B2(n19783), .ZN(n19734) );
  OAI211_X1 U22779 ( .C1(n19768), .C2(n19736), .A(n19735), .B(n19734), .ZN(
        P2_U3160) );
  AOI22_X1 U22780 ( .A1(n19737), .A2(n19830), .B1(n19787), .B2(n19761), .ZN(
        n19739) );
  AOI22_X1 U22781 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19789), .ZN(n19738) );
  OAI211_X1 U22782 ( .C1(n19768), .C2(n19740), .A(n19739), .B(n19738), .ZN(
        P2_U3161) );
  AOI22_X1 U22783 ( .A1(n19795), .A2(n19830), .B1(n19793), .B2(n19761), .ZN(
        n19743) );
  AOI22_X1 U22784 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19741), .ZN(n19742) );
  OAI211_X1 U22785 ( .C1(n19768), .C2(n19744), .A(n19743), .B(n19742), .ZN(
        P2_U3162) );
  AOI22_X1 U22786 ( .A1(n19745), .A2(n19763), .B1(n19799), .B2(n19761), .ZN(
        n19747) );
  AOI22_X1 U22787 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19764), .B1(
        n19830), .B2(n19801), .ZN(n19746) );
  OAI211_X1 U22788 ( .C1(n19768), .C2(n19748), .A(n19747), .B(n19746), .ZN(
        P2_U3163) );
  AOI22_X1 U22789 ( .A1(n19807), .A2(n19830), .B1(n19805), .B2(n19761), .ZN(
        n19751) );
  AOI22_X1 U22790 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19749), .ZN(n19750) );
  OAI211_X1 U22791 ( .C1(n19768), .C2(n19752), .A(n19751), .B(n19750), .ZN(
        P2_U3164) );
  AOI22_X1 U22792 ( .A1(n19753), .A2(n19763), .B1(n19811), .B2(n19761), .ZN(
        n19755) );
  AOI22_X1 U22793 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19764), .B1(
        n19830), .B2(n19813), .ZN(n19754) );
  OAI211_X1 U22794 ( .C1(n19768), .C2(n19756), .A(n19755), .B(n19754), .ZN(
        P2_U3165) );
  AOI22_X1 U22795 ( .A1(n19757), .A2(n19830), .B1(n19819), .B2(n19761), .ZN(
        n19759) );
  AOI22_X1 U22796 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19821), .ZN(n19758) );
  OAI211_X1 U22797 ( .C1(n19768), .C2(n19760), .A(n19759), .B(n19758), .ZN(
        P2_U3166) );
  AOI22_X1 U22798 ( .A1(n19762), .A2(n19830), .B1(n19825), .B2(n19761), .ZN(
        n19766) );
  AOI22_X1 U22799 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19829), .ZN(n19765) );
  OAI211_X1 U22800 ( .C1(n19768), .C2(n19767), .A(n19766), .B(n19765), .ZN(
        P2_U3167) );
  AND2_X1 U22801 ( .A1(n19773), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19769) );
  NAND2_X1 U22802 ( .A1(n19770), .A2(n19769), .ZN(n19776) );
  OAI21_X1 U22803 ( .B1(n19771), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19975), 
        .ZN(n19772) );
  AND2_X1 U22804 ( .A1(n19776), .A2(n19772), .ZN(n19828) );
  INV_X1 U22805 ( .A(n19773), .ZN(n19826) );
  AOI22_X1 U22806 ( .A1(n19775), .A2(n19828), .B1(n19826), .B2(n19774), .ZN(
        n19785) );
  OAI211_X1 U22807 ( .C1(n19826), .C2(n19951), .A(n19777), .B(n19776), .ZN(
        n19778) );
  INV_X1 U22808 ( .A(n19778), .ZN(n19779) );
  OAI221_X1 U22809 ( .B1(n19782), .B2(n19781), .C1(n19782), .C2(n19780), .A(
        n19779), .ZN(n19831) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19831), .B1(
        n19814), .B2(n19783), .ZN(n19784) );
  OAI211_X1 U22811 ( .C1(n19786), .C2(n19817), .A(n19785), .B(n19784), .ZN(
        P2_U3168) );
  AOI22_X1 U22812 ( .A1(n19828), .A2(n19788), .B1(n19826), .B2(n19787), .ZN(
        n19791) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19831), .B1(
        n19830), .B2(n19789), .ZN(n19790) );
  OAI211_X1 U22814 ( .C1(n19792), .C2(n19834), .A(n19791), .B(n19790), .ZN(
        P2_U3169) );
  AOI22_X1 U22815 ( .A1(n19794), .A2(n19828), .B1(n19826), .B2(n19793), .ZN(
        n19797) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19831), .B1(
        n19814), .B2(n19795), .ZN(n19796) );
  OAI211_X1 U22817 ( .C1(n19798), .C2(n19817), .A(n19797), .B(n19796), .ZN(
        P2_U3170) );
  AOI22_X1 U22818 ( .A1(n19828), .A2(n19800), .B1(n19826), .B2(n19799), .ZN(
        n19803) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19831), .B1(
        n19814), .B2(n19801), .ZN(n19802) );
  OAI211_X1 U22820 ( .C1(n19804), .C2(n19817), .A(n19803), .B(n19802), .ZN(
        P2_U3171) );
  AOI22_X1 U22821 ( .A1(n19806), .A2(n19828), .B1(n19826), .B2(n19805), .ZN(
        n19809) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19831), .B1(
        n19814), .B2(n19807), .ZN(n19808) );
  OAI211_X1 U22823 ( .C1(n19810), .C2(n19817), .A(n19809), .B(n19808), .ZN(
        P2_U3172) );
  AOI22_X1 U22824 ( .A1(n19828), .A2(n19812), .B1(n19826), .B2(n19811), .ZN(
        n19816) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19831), .B1(
        n19814), .B2(n19813), .ZN(n19815) );
  OAI211_X1 U22826 ( .C1(n19818), .C2(n19817), .A(n19816), .B(n19815), .ZN(
        P2_U3173) );
  AOI22_X1 U22827 ( .A1(n19820), .A2(n19828), .B1(n19826), .B2(n19819), .ZN(
        n19823) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19831), .B1(
        n19830), .B2(n19821), .ZN(n19822) );
  OAI211_X1 U22829 ( .C1(n19824), .C2(n19834), .A(n19823), .B(n19822), .ZN(
        P2_U3174) );
  AOI22_X1 U22830 ( .A1(n19828), .A2(n19827), .B1(n19826), .B2(n19825), .ZN(
        n19833) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19831), .B1(
        n19830), .B2(n19829), .ZN(n19832) );
  OAI211_X1 U22832 ( .C1(n19835), .C2(n19834), .A(n19833), .B(n19832), .ZN(
        P2_U3175) );
  OAI211_X1 U22833 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19983), .A(n19837), 
        .B(n19836), .ZN(n19841) );
  NOR2_X1 U22834 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20977), .ZN(n19838) );
  OAI211_X1 U22835 ( .C1(n19842), .C2(n19838), .A(n19976), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19839) );
  OAI211_X1 U22836 ( .C1(n19842), .C2(n19841), .A(n19840), .B(n19839), .ZN(
        P2_U3177) );
  AND2_X1 U22837 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19844), .ZN(
        P2_U3179) );
  AND2_X1 U22838 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19844), .ZN(
        P2_U3180) );
  AND2_X1 U22839 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19844), .ZN(
        P2_U3181) );
  AND2_X1 U22840 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19844), .ZN(
        P2_U3182) );
  AND2_X1 U22841 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19844), .ZN(
        P2_U3183) );
  NOR2_X1 U22842 ( .A1(n21146), .A2(n19922), .ZN(P2_U3184) );
  AND2_X1 U22843 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19844), .ZN(
        P2_U3185) );
  AND2_X1 U22844 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19844), .ZN(
        P2_U3186) );
  AND2_X1 U22845 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19844), .ZN(
        P2_U3187) );
  AND2_X1 U22846 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19844), .ZN(
        P2_U3188) );
  AND2_X1 U22847 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19844), .ZN(
        P2_U3189) );
  AND2_X1 U22848 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19843), .ZN(
        P2_U3190) );
  AND2_X1 U22849 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19843), .ZN(
        P2_U3191) );
  AND2_X1 U22850 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19843), .ZN(
        P2_U3192) );
  AND2_X1 U22851 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19843), .ZN(
        P2_U3193) );
  AND2_X1 U22852 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19843), .ZN(
        P2_U3194) );
  AND2_X1 U22853 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19843), .ZN(
        P2_U3195) );
  AND2_X1 U22854 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19843), .ZN(
        P2_U3196) );
  AND2_X1 U22855 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19843), .ZN(
        P2_U3197) );
  AND2_X1 U22856 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19843), .ZN(
        P2_U3198) );
  AND2_X1 U22857 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19843), .ZN(
        P2_U3199) );
  AND2_X1 U22858 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19843), .ZN(
        P2_U3200) );
  AND2_X1 U22859 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19843), .ZN(P2_U3201) );
  NOR2_X1 U22860 ( .A1(n20992), .A2(n19922), .ZN(P2_U3202) );
  AND2_X1 U22861 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19844), .ZN(P2_U3203) );
  AND2_X1 U22862 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19844), .ZN(P2_U3204) );
  AND2_X1 U22863 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19844), .ZN(P2_U3205) );
  AND2_X1 U22864 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19843), .ZN(P2_U3206) );
  AND2_X1 U22865 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19843), .ZN(P2_U3207) );
  AND2_X1 U22866 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19844), .ZN(P2_U3208) );
  OAI21_X1 U22867 ( .B1(n20786), .B2(n19850), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19860) );
  NAND2_X1 U22868 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19976), .ZN(n19858) );
  NAND3_X1 U22869 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19858), .ZN(n19847) );
  AOI211_X1 U22870 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20782), .A(
        n19988), .B(n19845), .ZN(n19846) );
  AOI21_X1 U22871 ( .B1(n19860), .B2(n19847), .A(n19846), .ZN(n19848) );
  INV_X1 U22872 ( .A(n19848), .ZN(P2_U3209) );
  NOR2_X1 U22873 ( .A1(HOLD), .A2(n19849), .ZN(n19859) );
  AOI21_X1 U22874 ( .B1(n19861), .B2(n19850), .A(n19859), .ZN(n19854) );
  INV_X1 U22875 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19853) );
  AOI21_X1 U22876 ( .B1(HOLD), .B2(n19851), .A(n19972), .ZN(n19852) );
  OAI211_X1 U22877 ( .C1(n19854), .C2(n19853), .A(n19852), .B(n19858), .ZN(
        P2_U3210) );
  OAI22_X1 U22878 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19855), .B1(NA), 
        .B2(n19858), .ZN(n19856) );
  OAI211_X1 U22879 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19856), .ZN(n19857) );
  OAI221_X1 U22880 ( .B1(n19860), .B2(n19859), .C1(n19860), .C2(n19858), .A(
        n19857), .ZN(P2_U3211) );
  OAI222_X1 U22881 ( .A1(n19915), .A2(n19864), .B1(n19863), .B2(n19988), .C1(
        n19862), .C2(n19911), .ZN(P2_U3212) );
  OAI222_X1 U22882 ( .A1(n19915), .A2(n19866), .B1(n19865), .B2(n19988), .C1(
        n19864), .C2(n19911), .ZN(P2_U3213) );
  OAI222_X1 U22883 ( .A1(n19915), .A2(n19868), .B1(n19867), .B2(n19988), .C1(
        n19866), .C2(n19911), .ZN(P2_U3214) );
  OAI222_X1 U22884 ( .A1(n19915), .A2(n13589), .B1(n19869), .B2(n19988), .C1(
        n19868), .C2(n19911), .ZN(P2_U3215) );
  OAI222_X1 U22885 ( .A1(n19915), .A2(n19870), .B1(n21024), .B2(n19988), .C1(
        n13589), .C2(n19911), .ZN(P2_U3216) );
  OAI222_X1 U22886 ( .A1(n19915), .A2(n19872), .B1(n19871), .B2(n19988), .C1(
        n19870), .C2(n19911), .ZN(P2_U3217) );
  OAI222_X1 U22887 ( .A1(n19915), .A2(n13650), .B1(n20991), .B2(n19988), .C1(
        n19872), .C2(n19911), .ZN(P2_U3218) );
  OAI222_X1 U22888 ( .A1(n19915), .A2(n19873), .B1(n21175), .B2(n19988), .C1(
        n13650), .C2(n19911), .ZN(P2_U3219) );
  OAI222_X1 U22889 ( .A1(n19915), .A2(n11445), .B1(n19874), .B2(n19988), .C1(
        n19873), .C2(n19911), .ZN(P2_U3220) );
  OAI222_X1 U22890 ( .A1(n19915), .A2(n19876), .B1(n19875), .B2(n19988), .C1(
        n11445), .C2(n19911), .ZN(P2_U3221) );
  INV_X1 U22891 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19878) );
  OAI222_X1 U22892 ( .A1(n19915), .A2(n19878), .B1(n19877), .B2(n19988), .C1(
        n19876), .C2(n19911), .ZN(P2_U3222) );
  OAI222_X1 U22893 ( .A1(n19915), .A2(n21209), .B1(n19879), .B2(n19988), .C1(
        n19878), .C2(n19911), .ZN(P2_U3223) );
  OAI222_X1 U22894 ( .A1(n19915), .A2(n19881), .B1(n19880), .B2(n19988), .C1(
        n21209), .C2(n19911), .ZN(P2_U3224) );
  OAI222_X1 U22895 ( .A1(n19915), .A2(n19883), .B1(n19882), .B2(n19988), .C1(
        n19881), .C2(n19911), .ZN(P2_U3225) );
  INV_X1 U22896 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19885) );
  OAI222_X1 U22897 ( .A1(n19915), .A2(n19885), .B1(n19884), .B2(n19988), .C1(
        n19883), .C2(n19911), .ZN(P2_U3226) );
  OAI222_X1 U22898 ( .A1(n19915), .A2(n19887), .B1(n19886), .B2(n19988), .C1(
        n19885), .C2(n19911), .ZN(P2_U3227) );
  OAI222_X1 U22899 ( .A1(n19915), .A2(n15378), .B1(n19888), .B2(n19988), .C1(
        n19887), .C2(n19911), .ZN(P2_U3228) );
  OAI222_X1 U22900 ( .A1(n19915), .A2(n21177), .B1(n19889), .B2(n19988), .C1(
        n15378), .C2(n19911), .ZN(P2_U3229) );
  INV_X1 U22901 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19891) );
  OAI222_X1 U22902 ( .A1(n19915), .A2(n19891), .B1(n19890), .B2(n19988), .C1(
        n21177), .C2(n19911), .ZN(P2_U3230) );
  OAI222_X1 U22903 ( .A1(n19915), .A2(n19893), .B1(n19892), .B2(n19988), .C1(
        n19891), .C2(n19911), .ZN(P2_U3231) );
  INV_X1 U22904 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19895) );
  OAI222_X1 U22905 ( .A1(n19915), .A2(n19895), .B1(n19894), .B2(n19988), .C1(
        n19893), .C2(n19911), .ZN(P2_U3232) );
  OAI222_X1 U22906 ( .A1(n19915), .A2(n19897), .B1(n19896), .B2(n19988), .C1(
        n19895), .C2(n19911), .ZN(P2_U3233) );
  OAI222_X1 U22907 ( .A1(n19915), .A2(n19899), .B1(n19898), .B2(n19988), .C1(
        n19897), .C2(n19911), .ZN(P2_U3234) );
  OAI222_X1 U22908 ( .A1(n19915), .A2(n19901), .B1(n19900), .B2(n19988), .C1(
        n19899), .C2(n19911), .ZN(P2_U3235) );
  INV_X1 U22909 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19903) );
  OAI222_X1 U22910 ( .A1(n19915), .A2(n19903), .B1(n19902), .B2(n19988), .C1(
        n19901), .C2(n19911), .ZN(P2_U3236) );
  OAI222_X1 U22911 ( .A1(n19915), .A2(n19906), .B1(n19904), .B2(n19988), .C1(
        n19903), .C2(n19911), .ZN(P2_U3237) );
  OAI222_X1 U22912 ( .A1(n19911), .A2(n19906), .B1(n19905), .B2(n19988), .C1(
        n19907), .C2(n19915), .ZN(P2_U3238) );
  INV_X1 U22913 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19909) );
  OAI222_X1 U22914 ( .A1(n19915), .A2(n19909), .B1(n19908), .B2(n19988), .C1(
        n19907), .C2(n19911), .ZN(P2_U3239) );
  INV_X1 U22915 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19912) );
  OAI222_X1 U22916 ( .A1(n19915), .A2(n19912), .B1(n19910), .B2(n19988), .C1(
        n19909), .C2(n19911), .ZN(P2_U3240) );
  OAI222_X1 U22917 ( .A1(n19915), .A2(n19914), .B1(n19913), .B2(n19988), .C1(
        n19912), .C2(n19911), .ZN(P2_U3241) );
  OAI22_X1 U22918 ( .A1(n19986), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19988), .ZN(n19916) );
  INV_X1 U22919 ( .A(n19916), .ZN(P2_U3585) );
  MUX2_X1 U22920 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19986), .Z(P2_U3586) );
  OAI22_X1 U22921 ( .A1(n19986), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19988), .ZN(n19917) );
  INV_X1 U22922 ( .A(n19917), .ZN(P2_U3587) );
  OAI22_X1 U22923 ( .A1(n19986), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19988), .ZN(n19918) );
  INV_X1 U22924 ( .A(n19918), .ZN(P2_U3588) );
  OAI21_X1 U22925 ( .B1(n19922), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19920), 
        .ZN(n19919) );
  INV_X1 U22926 ( .A(n19919), .ZN(P2_U3591) );
  OAI21_X1 U22927 ( .B1(n19922), .B2(n19921), .A(n19920), .ZN(P2_U3592) );
  INV_X1 U22928 ( .A(n19956), .ZN(n19959) );
  NAND2_X1 U22929 ( .A1(n19923), .A2(n19924), .ZN(n19931) );
  AND2_X1 U22930 ( .A1(n19924), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19946) );
  NAND2_X1 U22931 ( .A1(n19925), .A2(n19946), .ZN(n19936) );
  NAND3_X1 U22932 ( .A1(n19944), .A2(n19926), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19927) );
  NAND2_X1 U22933 ( .A1(n19927), .A2(n19954), .ZN(n19937) );
  NAND2_X1 U22934 ( .A1(n19936), .A2(n19937), .ZN(n19929) );
  NAND2_X1 U22935 ( .A1(n19929), .A2(n19928), .ZN(n19930) );
  OAI211_X1 U22936 ( .C1(n19932), .C2(n19951), .A(n19931), .B(n19930), .ZN(
        n19933) );
  INV_X1 U22937 ( .A(n19933), .ZN(n19934) );
  AOI22_X1 U22938 ( .A1(n19959), .A2(n19935), .B1(n19934), .B2(n19956), .ZN(
        P2_U3602) );
  OAI21_X1 U22939 ( .B1(n19938), .B2(n19937), .A(n19936), .ZN(n19939) );
  AOI21_X1 U22940 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19940), .A(n19939), 
        .ZN(n19941) );
  AOI22_X1 U22941 ( .A1(n19959), .A2(n13038), .B1(n19941), .B2(n19956), .ZN(
        P2_U3603) );
  INV_X1 U22942 ( .A(n19954), .ZN(n19943) );
  NOR2_X1 U22943 ( .A1(n19943), .A2(n19942), .ZN(n19945) );
  MUX2_X1 U22944 ( .A(n19946), .B(n19945), .S(n19944), .Z(n19947) );
  AOI21_X1 U22945 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19948), .A(n19947), 
        .ZN(n19949) );
  AOI22_X1 U22946 ( .A1(n19959), .A2(n19950), .B1(n19949), .B2(n19956), .ZN(
        P2_U3604) );
  NOR2_X1 U22947 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19951), .ZN(
        n19952) );
  AOI211_X1 U22948 ( .C1(n19955), .C2(n19954), .A(n19953), .B(n19952), .ZN(
        n19957) );
  AOI22_X1 U22949 ( .A1(n19959), .A2(n19958), .B1(n19957), .B2(n19956), .ZN(
        P2_U3605) );
  INV_X1 U22950 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n21066) );
  AOI22_X1 U22951 ( .A1(n19988), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n21066), 
        .B2(n19986), .ZN(P2_U3608) );
  INV_X1 U22952 ( .A(n19960), .ZN(n19966) );
  AOI22_X1 U22953 ( .A1(n19964), .A2(n19963), .B1(n19962), .B2(n19961), .ZN(
        n19965) );
  NAND2_X1 U22954 ( .A1(n19966), .A2(n19965), .ZN(n19968) );
  MUX2_X1 U22955 ( .A(P2_MORE_REG_SCAN_IN), .B(n19968), .S(n19967), .Z(
        P2_U3609) );
  AOI21_X1 U22956 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19972), .A(n19969), 
        .ZN(n19974) );
  NOR3_X1 U22957 ( .A1(n19972), .A2(n19971), .A3(n19970), .ZN(n19973) );
  OAI21_X1 U22958 ( .B1(n19974), .B2(n19973), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19979) );
  OAI22_X1 U22959 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19977), .B1(n19976), 
        .B2(n19975), .ZN(n19978) );
  NAND2_X1 U22960 ( .A1(n19979), .A2(n19978), .ZN(n19985) );
  AOI21_X1 U22961 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19980), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19982) );
  AOI211_X1 U22962 ( .C1(n19269), .C2(n19983), .A(n19982), .B(n19981), .ZN(
        n19984) );
  MUX2_X1 U22963 ( .A(n19985), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19984), 
        .Z(P2_U3610) );
  INV_X1 U22964 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19987) );
  INV_X1 U22965 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n21171) );
  AOI22_X1 U22966 ( .A1(n19988), .A2(n19987), .B1(n21171), .B2(n19986), .ZN(
        P2_U3611) );
  INV_X1 U22967 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20795) );
  AOI21_X1 U22968 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20795), .A(n21063), 
        .ZN(n19997) );
  INV_X1 U22969 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19989) );
  AOI21_X1 U22970 ( .B1(n19997), .B2(n19989), .A(n20873), .ZN(P1_U2802) );
  NAND2_X1 U22971 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n19990), .ZN(n19995) );
  INV_X1 U22972 ( .A(n19991), .ZN(n19993) );
  OAI21_X1 U22973 ( .B1(n19993), .B2(n19992), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19994) );
  OAI21_X1 U22974 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19995), .A(n19994), 
        .ZN(P1_U2803) );
  INV_X2 U22975 ( .A(n20873), .ZN(n20884) );
  NOR2_X1 U22976 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19998) );
  OAI21_X1 U22977 ( .B1(n19998), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20884), .ZN(
        n19996) );
  OAI21_X1 U22978 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20884), .A(n19996), 
        .ZN(P1_U2804) );
  NOR2_X1 U22979 ( .A1(n19997), .A2(n20873), .ZN(n20844) );
  OAI21_X1 U22980 ( .B1(BS16), .B2(n19998), .A(n20844), .ZN(n20843) );
  OAI21_X1 U22981 ( .B1(n20844), .B2(n20847), .A(n20843), .ZN(P1_U2805) );
  OAI21_X1 U22982 ( .B1(n20001), .B2(n20000), .A(n19999), .ZN(P1_U2806) );
  NOR4_X1 U22983 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20005) );
  NOR4_X1 U22984 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20004) );
  NOR4_X1 U22985 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20003) );
  NOR4_X1 U22986 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20002) );
  NAND4_X1 U22987 ( .A1(n20005), .A2(n20004), .A3(n20003), .A4(n20002), .ZN(
        n20011) );
  NOR4_X1 U22988 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20009) );
  AOI211_X1 U22989 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_26__SCAN_IN), .B(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20008) );
  NOR4_X1 U22990 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20007) );
  NOR4_X1 U22991 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20006) );
  NAND4_X1 U22992 ( .A1(n20009), .A2(n20008), .A3(n20007), .A4(n20006), .ZN(
        n20010) );
  NOR2_X1 U22993 ( .A1(n20011), .A2(n20010), .ZN(n20871) );
  INV_X1 U22994 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20013) );
  NOR3_X1 U22995 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20014) );
  OAI21_X1 U22996 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20014), .A(n20871), .ZN(
        n20012) );
  OAI21_X1 U22997 ( .B1(n20871), .B2(n20013), .A(n20012), .ZN(P1_U2807) );
  INV_X1 U22998 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21065) );
  AOI21_X1 U22999 ( .B1(n20796), .B2(n21065), .A(n20014), .ZN(n20016) );
  INV_X1 U23000 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20015) );
  INV_X1 U23001 ( .A(n20871), .ZN(n20868) );
  AOI22_X1 U23002 ( .A1(n20871), .A2(n20016), .B1(n20015), .B2(n20868), .ZN(
        P1_U2808) );
  INV_X1 U23003 ( .A(n20017), .ZN(n20019) );
  AOI22_X1 U23004 ( .A1(n20019), .A2(n20050), .B1(n20086), .B2(n20018), .ZN(
        n20030) );
  INV_X1 U23005 ( .A(n20020), .ZN(n20021) );
  AOI22_X1 U23006 ( .A1(n20056), .A2(n20021), .B1(n20081), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n20023) );
  OAI211_X1 U23007 ( .C1(n20025), .C2(n20024), .A(n20023), .B(n20022), .ZN(
        n20026) );
  AOI221_X1 U23008 ( .B1(n20028), .B2(P1_REIP_REG_9__SCAN_IN), .C1(n20027), 
        .C2(n20806), .A(n20026), .ZN(n20029) );
  NAND2_X1 U23009 ( .A1(n20030), .A2(n20029), .ZN(P1_U2831) );
  INV_X1 U23010 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20804) );
  NAND2_X1 U23011 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20032) );
  OAI21_X1 U23012 ( .B1(n20032), .B2(n20060), .A(n20031), .ZN(n20047) );
  OAI22_X1 U23013 ( .A1(n20034), .A2(n20098), .B1(n20043), .B2(n20033), .ZN(
        n20035) );
  AOI211_X1 U23014 ( .C1(n20087), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20069), .B(n20035), .ZN(n20036) );
  OAI221_X1 U23015 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n20037), .C1(n20804), 
        .C2(n20047), .A(n20036), .ZN(n20038) );
  AOI21_X1 U23016 ( .B1(n20039), .B2(n20050), .A(n20038), .ZN(n20040) );
  OAI21_X1 U23017 ( .B1(n20041), .B2(n20078), .A(n20040), .ZN(P1_U2833) );
  NAND3_X1 U23018 ( .A1(n20084), .A2(n20054), .A3(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20048) );
  OAI22_X1 U23019 ( .A1(n20044), .A2(n20098), .B1(n20043), .B2(n20042), .ZN(
        n20045) );
  AOI211_X1 U23020 ( .C1(n20087), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20069), .B(n20045), .ZN(n20046) );
  OAI221_X1 U23021 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n20048), .C1(n16132), 
        .C2(n20047), .A(n20046), .ZN(n20049) );
  AOI21_X1 U23022 ( .B1(n20051), .B2(n20050), .A(n20049), .ZN(n20052) );
  OAI21_X1 U23023 ( .B1(n20053), .B2(n20078), .A(n20052), .ZN(P1_U2834) );
  NAND2_X1 U23024 ( .A1(n20084), .A2(n20054), .ZN(n20058) );
  AOI22_X1 U23025 ( .A1(n20056), .A2(n20055), .B1(n20081), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n20057) );
  OAI21_X1 U23026 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20058), .A(n20057), .ZN(
        n20059) );
  AOI211_X1 U23027 ( .C1(n20087), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20069), .B(n20059), .ZN(n20065) );
  INV_X1 U23028 ( .A(n20060), .ZN(n20061) );
  NOR2_X1 U23029 ( .A1(n20062), .A2(n20061), .ZN(n20070) );
  AOI22_X1 U23030 ( .A1(n20063), .A2(n20091), .B1(n20070), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20064) );
  OAI211_X1 U23031 ( .C1(n20066), .C2(n20078), .A(n20065), .B(n20064), .ZN(
        P1_U2835) );
  AOI22_X1 U23032 ( .A1(n20081), .A2(P1_EBX_REG_4__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20087), .ZN(n20067) );
  INV_X1 U23033 ( .A(n20067), .ZN(n20068) );
  AOI211_X1 U23034 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n20070), .A(n20069), .B(
        n20068), .ZN(n20077) );
  OAI22_X1 U23035 ( .A1(n20098), .A2(n20178), .B1(n20072), .B2(n20071), .ZN(
        n20075) );
  NOR3_X1 U23036 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n13687), .A3(n20073), .ZN(
        n20074) );
  AOI211_X1 U23037 ( .C1(n20158), .C2(n20091), .A(n20075), .B(n20074), .ZN(
        n20076) );
  OAI211_X1 U23038 ( .C1(n20162), .C2(n20078), .A(n20077), .B(n20076), .ZN(
        P1_U2836) );
  OAI21_X1 U23039 ( .B1(n20080), .B2(P1_REIP_REG_1__SCAN_IN), .A(n20079), .ZN(
        n20082) );
  AOI22_X1 U23040 ( .A1(n20082), .A2(P1_REIP_REG_2__SCAN_IN), .B1(n20081), 
        .B2(P1_EBX_REG_2__SCAN_IN), .ZN(n20097) );
  NAND3_X1 U23041 ( .A1(n20084), .A2(P1_REIP_REG_1__SCAN_IN), .A3(n20083), 
        .ZN(n20095) );
  AOI22_X1 U23042 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20087), .B1(
        n20086), .B2(n20085), .ZN(n20094) );
  NAND2_X1 U23043 ( .A1(n20089), .A2(n20088), .ZN(n20093) );
  NAND2_X1 U23044 ( .A1(n20091), .A2(n20090), .ZN(n20092) );
  OAI211_X1 U23045 ( .C1(n20098), .C2(n20196), .A(n20097), .B(n20096), .ZN(
        P1_U2838) );
  AOI22_X1 U23046 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20104), .B1(n20112), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20099) );
  OAI21_X1 U23047 ( .B1(n20100), .B2(n20106), .A(n20099), .ZN(P1_U2921) );
  AOI22_X1 U23048 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20101) );
  OAI21_X1 U23049 ( .B1(n14700), .B2(n20123), .A(n20101), .ZN(P1_U2922) );
  AOI22_X1 U23050 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20102) );
  OAI21_X1 U23051 ( .B1(n14702), .B2(n20123), .A(n20102), .ZN(P1_U2923) );
  AOI22_X1 U23052 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20103) );
  OAI21_X1 U23053 ( .B1(n14705), .B2(n20123), .A(n20103), .ZN(P1_U2924) );
  INV_X1 U23054 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n20107) );
  AOI22_X1 U23055 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n20104), .B1(n20112), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20105) );
  OAI21_X1 U23056 ( .B1(n20107), .B2(n20106), .A(n20105), .ZN(P1_U2925) );
  AOI22_X1 U23057 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20108) );
  OAI21_X1 U23058 ( .B1(n13761), .B2(n20123), .A(n20108), .ZN(P1_U2926) );
  AOI22_X1 U23059 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20109) );
  OAI21_X1 U23060 ( .B1(n13701), .B2(n20123), .A(n20109), .ZN(P1_U2927) );
  AOI22_X1 U23061 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20110) );
  OAI21_X1 U23062 ( .B1(n13491), .B2(n20123), .A(n20110), .ZN(P1_U2928) );
  AOI22_X1 U23063 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20111) );
  OAI21_X1 U23064 ( .B1(n12024), .B2(n20123), .A(n20111), .ZN(P1_U2929) );
  AOI22_X1 U23065 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20113) );
  OAI21_X1 U23066 ( .B1(n20114), .B2(n20123), .A(n20113), .ZN(P1_U2930) );
  AOI22_X1 U23067 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20115) );
  OAI21_X1 U23068 ( .B1(n11989), .B2(n20123), .A(n20115), .ZN(P1_U2931) );
  AOI22_X1 U23069 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20116) );
  OAI21_X1 U23070 ( .B1(n20117), .B2(n20123), .A(n20116), .ZN(P1_U2932) );
  AOI22_X1 U23071 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20118) );
  OAI21_X1 U23072 ( .B1(n11920), .B2(n20123), .A(n20118), .ZN(P1_U2933) );
  AOI22_X1 U23073 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20119) );
  OAI21_X1 U23074 ( .B1(n11927), .B2(n20123), .A(n20119), .ZN(P1_U2934) );
  AOI22_X1 U23075 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20120) );
  OAI21_X1 U23076 ( .B1(n11931), .B2(n20123), .A(n20120), .ZN(P1_U2935) );
  AOI22_X1 U23077 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20121), .B1(n20112), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20122) );
  OAI21_X1 U23078 ( .B1(n20124), .B2(n20123), .A(n20122), .ZN(P1_U2936) );
  AOI22_X1 U23079 ( .A1(n20151), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20150), .ZN(n20127) );
  INV_X1 U23080 ( .A(n20125), .ZN(n20126) );
  NAND2_X1 U23081 ( .A1(n20136), .A2(n20126), .ZN(n20138) );
  NAND2_X1 U23082 ( .A1(n20127), .A2(n20138), .ZN(P1_U2945) );
  AOI22_X1 U23083 ( .A1(n20151), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20130) );
  INV_X1 U23084 ( .A(n20128), .ZN(n20129) );
  NAND2_X1 U23085 ( .A1(n20136), .A2(n20129), .ZN(n20140) );
  NAND2_X1 U23086 ( .A1(n20130), .A2(n20140), .ZN(P1_U2946) );
  AOI22_X1 U23087 ( .A1(n20151), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20133) );
  INV_X1 U23088 ( .A(n20131), .ZN(n20132) );
  NAND2_X1 U23089 ( .A1(n20136), .A2(n20132), .ZN(n20142) );
  NAND2_X1 U23090 ( .A1(n20133), .A2(n20142), .ZN(P1_U2947) );
  AOI22_X1 U23091 ( .A1(n20151), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20150), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20137) );
  INV_X1 U23092 ( .A(n20134), .ZN(n20135) );
  NAND2_X1 U23093 ( .A1(n20136), .A2(n20135), .ZN(n20152) );
  NAND2_X1 U23094 ( .A1(n20137), .A2(n20152), .ZN(P1_U2951) );
  AOI22_X1 U23095 ( .A1(n20151), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20139) );
  NAND2_X1 U23096 ( .A1(n20139), .A2(n20138), .ZN(P1_U2960) );
  AOI22_X1 U23097 ( .A1(n20151), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20150), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20141) );
  NAND2_X1 U23098 ( .A1(n20141), .A2(n20140), .ZN(P1_U2961) );
  AOI22_X1 U23099 ( .A1(n20151), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20150), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20143) );
  NAND2_X1 U23100 ( .A1(n20143), .A2(n20142), .ZN(P1_U2962) );
  AOI22_X1 U23101 ( .A1(n20151), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20150), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20145) );
  NAND2_X1 U23102 ( .A1(n20145), .A2(n20144), .ZN(P1_U2963) );
  AOI22_X1 U23103 ( .A1(n20151), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20150), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20147) );
  NAND2_X1 U23104 ( .A1(n20147), .A2(n20146), .ZN(P1_U2964) );
  AOI22_X1 U23105 ( .A1(n20151), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20150), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20149) );
  NAND2_X1 U23106 ( .A1(n20149), .A2(n20148), .ZN(P1_U2965) );
  AOI22_X1 U23107 ( .A1(n20151), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20150), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20153) );
  NAND2_X1 U23108 ( .A1(n20153), .A2(n20152), .ZN(P1_U2966) );
  AOI22_X1 U23109 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20161) );
  OAI21_X1 U23110 ( .B1(n20156), .B2(n20155), .A(n20154), .ZN(n20157) );
  INV_X1 U23111 ( .A(n20157), .ZN(n20180) );
  AOI22_X1 U23112 ( .A1(n20180), .A2(n20169), .B1(n20159), .B2(n20158), .ZN(
        n20160) );
  OAI211_X1 U23113 ( .C1(n20163), .C2(n20162), .A(n20161), .B(n20160), .ZN(
        P1_U2995) );
  AOI22_X1 U23114 ( .A1(n20165), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20164), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20173) );
  OR2_X1 U23115 ( .A1(n20166), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20167) );
  AND2_X1 U23116 ( .A1(n20168), .A2(n20167), .ZN(n20211) );
  AOI22_X1 U23117 ( .A1(n20171), .A2(n20170), .B1(n20169), .B2(n20211), .ZN(
        n20172) );
  OAI211_X1 U23118 ( .C1(n20175), .C2(n20174), .A(n20173), .B(n20172), .ZN(
        P1_U2998) );
  OAI21_X1 U23119 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20176), .ZN(n20183) );
  INV_X1 U23120 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20177) );
  OAI22_X1 U23121 ( .A1(n20224), .A2(n20178), .B1(n20208), .B2(n20177), .ZN(
        n20179) );
  INV_X1 U23122 ( .A(n20179), .ZN(n20182) );
  AOI22_X1 U23123 ( .A1(n20189), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20180), .B2(n20228), .ZN(n20181) );
  OAI211_X1 U23124 ( .C1(n20192), .C2(n20183), .A(n20182), .B(n20181), .ZN(
        P1_U3027) );
  AOI21_X1 U23125 ( .B1(n20186), .B2(n20185), .A(n20184), .ZN(n20191) );
  INV_X1 U23126 ( .A(n20187), .ZN(n20188) );
  AOI22_X1 U23127 ( .A1(n20189), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20228), .B2(n20188), .ZN(n20190) );
  OAI211_X1 U23128 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20192), .A(
        n20191), .B(n20190), .ZN(P1_U3028) );
  OR2_X1 U23129 ( .A1(n20219), .A2(n20193), .ZN(n20205) );
  NAND2_X1 U23130 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20195) );
  OAI21_X1 U23131 ( .B1(n20204), .B2(n20195), .A(n20194), .ZN(n20201) );
  OAI22_X1 U23132 ( .A1(n20224), .A2(n20196), .B1(n20083), .B2(n20208), .ZN(
        n20200) );
  AND3_X1 U23133 ( .A1(n20198), .A2(n20197), .A3(n20228), .ZN(n20199) );
  AOI211_X1 U23134 ( .C1(n20206), .C2(n20201), .A(n20200), .B(n20199), .ZN(
        n20202) );
  OAI221_X1 U23135 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20205), .C1(
        n20204), .C2(n20203), .A(n20202), .ZN(P1_U3029) );
  NAND2_X1 U23136 ( .A1(n20206), .A2(n20233), .ZN(n20223) );
  NAND2_X1 U23137 ( .A1(n20219), .A2(n20207), .ZN(n20214) );
  OAI22_X1 U23138 ( .A1(n20224), .A2(n20209), .B1(n20208), .B2(n20796), .ZN(
        n20210) );
  INV_X1 U23139 ( .A(n20210), .ZN(n20213) );
  NAND2_X1 U23140 ( .A1(n20228), .A2(n20211), .ZN(n20212) );
  OAI211_X1 U23141 ( .C1(n20215), .C2(n20214), .A(n20213), .B(n20212), .ZN(
        n20216) );
  INV_X1 U23142 ( .A(n20216), .ZN(n20217) );
  OAI221_X1 U23143 ( .B1(n20219), .B2(n20218), .C1(n20219), .C2(n20223), .A(
        n20217), .ZN(P1_U3030) );
  INV_X1 U23144 ( .A(n20220), .ZN(n20232) );
  INV_X1 U23145 ( .A(n20221), .ZN(n20229) );
  OAI211_X1 U23146 ( .C1(n20225), .C2(n20224), .A(n20223), .B(n20222), .ZN(
        n20226) );
  AOI211_X1 U23147 ( .C1(n20229), .C2(n20228), .A(n20227), .B(n20226), .ZN(
        n20230) );
  OAI221_X1 U23148 ( .B1(n20233), .B2(n20232), .C1(n20233), .C2(n20231), .A(
        n20230), .ZN(P1_U3031) );
  NOR2_X1 U23149 ( .A1(n20234), .A2(n20864), .ZN(P1_U3032) );
  INV_X1 U23150 ( .A(DATAI_17_), .ZN(n20963) );
  OAI22_X1 U23151 ( .A1(n20237), .A2(n20236), .B1(n20963), .B2(n20235), .ZN(
        n20685) );
  INV_X1 U23152 ( .A(n20685), .ZN(n20733) );
  NOR2_X2 U23153 ( .A1(n20265), .A2(n20238), .ZN(n20729) );
  AOI22_X1 U23154 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20267), .B1(DATAI_25_), 
        .B2(n20266), .ZN(n20688) );
  INV_X1 U23155 ( .A(n20688), .ZN(n20730) );
  AOI22_X1 U23156 ( .A1(n20729), .A2(n20268), .B1(n20761), .B2(n20730), .ZN(
        n20241) );
  INV_X1 U23157 ( .A(n20263), .ZN(n20272) );
  NAND2_X1 U23158 ( .A1(n20239), .A2(n20269), .ZN(n20551) );
  AOI22_X1 U23159 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20272), .B1(
        n20728), .B2(n20271), .ZN(n20240) );
  OAI211_X1 U23160 ( .C1(n20733), .C2(n20292), .A(n20241), .B(n20240), .ZN(
        P1_U3034) );
  AOI22_X1 U23161 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20267), .B1(DATAI_18_), 
        .B2(n20266), .ZN(n20739) );
  NOR2_X2 U23162 ( .A1(n20265), .A2(n13784), .ZN(n20735) );
  AOI22_X1 U23163 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20267), .B1(DATAI_26_), 
        .B2(n20266), .ZN(n20692) );
  INV_X1 U23164 ( .A(n20692), .ZN(n20736) );
  AOI22_X1 U23165 ( .A1(n20735), .A2(n20268), .B1(n20761), .B2(n20736), .ZN(
        n20244) );
  NAND2_X1 U23166 ( .A1(n20242), .A2(n20269), .ZN(n20554) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20272), .B1(
        n20734), .B2(n20271), .ZN(n20243) );
  OAI211_X1 U23168 ( .C1(n20739), .C2(n20292), .A(n20244), .B(n20243), .ZN(
        P1_U3035) );
  AOI22_X1 U23169 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20267), .B1(DATAI_19_), 
        .B2(n20266), .ZN(n20745) );
  NOR2_X2 U23170 ( .A1(n20265), .A2(n20245), .ZN(n20741) );
  AOI22_X1 U23171 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20267), .B1(DATAI_27_), 
        .B2(n20266), .ZN(n20696) );
  INV_X1 U23172 ( .A(n20696), .ZN(n20742) );
  AOI22_X1 U23173 ( .A1(n20741), .A2(n20268), .B1(n20761), .B2(n20742), .ZN(
        n20248) );
  NAND2_X1 U23174 ( .A1(n20246), .A2(n20269), .ZN(n20557) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20272), .B1(
        n20740), .B2(n20271), .ZN(n20247) );
  OAI211_X1 U23176 ( .C1(n20745), .C2(n20292), .A(n20248), .B(n20247), .ZN(
        P1_U3036) );
  NOR2_X2 U23177 ( .A1(n20265), .A2(n20249), .ZN(n20747) );
  INV_X1 U23178 ( .A(n20751), .ZN(n20656) );
  AOI22_X1 U23179 ( .A1(n20747), .A2(n20268), .B1(n20761), .B2(n20656), .ZN(
        n20252) );
  NAND2_X1 U23180 ( .A1(n20250), .A2(n20269), .ZN(n20560) );
  INV_X1 U23181 ( .A(n20292), .ZN(n20299) );
  AOI22_X1 U23182 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20267), .B1(DATAI_20_), 
        .B2(n20266), .ZN(n20659) );
  INV_X1 U23183 ( .A(n20659), .ZN(n20748) );
  AOI22_X1 U23184 ( .A1(n20746), .A2(n20271), .B1(n20299), .B2(n20748), .ZN(
        n20251) );
  OAI211_X1 U23185 ( .C1(n20263), .C2(n20253), .A(n20252), .B(n20251), .ZN(
        P1_U3037) );
  AOI22_X1 U23186 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20267), .B1(DATAI_21_), 
        .B2(n20266), .ZN(n20757) );
  AOI22_X1 U23187 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20267), .B1(DATAI_29_), 
        .B2(n20266), .ZN(n20702) );
  INV_X1 U23188 ( .A(n20702), .ZN(n20754) );
  AOI22_X1 U23189 ( .A1(n9795), .A2(n20268), .B1(n20761), .B2(n20754), .ZN(
        n20257) );
  NAND2_X1 U23190 ( .A1(n20255), .A2(n20269), .ZN(n20563) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20272), .B1(
        n20752), .B2(n20271), .ZN(n20256) );
  OAI211_X1 U23192 ( .C1(n20757), .C2(n20292), .A(n20257), .B(n20256), .ZN(
        P1_U3038) );
  NOR2_X2 U23193 ( .A1(n20265), .A2(n20258), .ZN(n20759) );
  AOI22_X1 U23194 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20267), .B1(DATAI_30_), 
        .B2(n20266), .ZN(n20765) );
  INV_X1 U23195 ( .A(n20765), .ZN(n20662) );
  AOI22_X1 U23196 ( .A1(n20759), .A2(n20268), .B1(n20761), .B2(n20662), .ZN(
        n20261) );
  NAND2_X1 U23197 ( .A1(n20259), .A2(n20269), .ZN(n20566) );
  AOI22_X1 U23198 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20267), .B1(DATAI_22_), 
        .B2(n20266), .ZN(n20665) );
  INV_X1 U23199 ( .A(n20665), .ZN(n20760) );
  AOI22_X1 U23200 ( .A1(n20758), .A2(n20271), .B1(n20299), .B2(n20760), .ZN(
        n20260) );
  OAI211_X1 U23201 ( .C1(n20263), .C2(n20262), .A(n20261), .B(n20260), .ZN(
        P1_U3039) );
  AOI22_X1 U23202 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20267), .B1(DATAI_23_), 
        .B2(n20266), .ZN(n20776) );
  NOR2_X2 U23203 ( .A1(n20265), .A2(n20264), .ZN(n20769) );
  AOI22_X1 U23204 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20267), .B1(DATAI_31_), 
        .B2(n20266), .ZN(n20712) );
  INV_X1 U23205 ( .A(n20712), .ZN(n20770) );
  AOI22_X1 U23206 ( .A1(n20769), .A2(n20268), .B1(n20761), .B2(n20770), .ZN(
        n20274) );
  NAND2_X1 U23207 ( .A1(n20270), .A2(n20269), .ZN(n20572) );
  AOI22_X1 U23208 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20272), .B1(
        n20767), .B2(n20271), .ZN(n20273) );
  OAI211_X1 U23209 ( .C1(n20776), .C2(n20292), .A(n20274), .B(n20273), .ZN(
        P1_U3040) );
  NOR2_X1 U23210 ( .A1(n20863), .A2(n20278), .ZN(n20298) );
  INV_X1 U23211 ( .A(n20335), .ZN(n20277) );
  INV_X1 U23212 ( .A(n20276), .ZN(n20641) );
  AOI21_X1 U23213 ( .B1(n20277), .B2(n20641), .A(n20298), .ZN(n20279) );
  OAI22_X1 U23214 ( .A1(n20279), .A2(n20859), .B1(n20278), .B2(n20715), .ZN(
        n20297) );
  AOI22_X1 U23215 ( .A1(n20718), .A2(n20298), .B1(n20717), .B2(n20297), .ZN(
        n20283) );
  OAI21_X1 U23216 ( .B1(n20333), .B2(n20847), .A(n20279), .ZN(n20280) );
  OAI221_X1 U23217 ( .B1(n20846), .B2(n20281), .C1(n20859), .C2(n20280), .A(
        n20722), .ZN(n20300) );
  INV_X1 U23218 ( .A(n20649), .ZN(n20724) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20300), .B1(
        n20326), .B2(n20724), .ZN(n20282) );
  OAI211_X1 U23220 ( .C1(n20727), .C2(n20292), .A(n20283), .B(n20282), .ZN(
        P1_U3041) );
  AOI22_X1 U23221 ( .A1(n20729), .A2(n20298), .B1(n20728), .B2(n20297), .ZN(
        n20285) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20300), .B1(
        n20326), .B2(n20685), .ZN(n20284) );
  OAI211_X1 U23223 ( .C1(n20688), .C2(n20292), .A(n20285), .B(n20284), .ZN(
        P1_U3042) );
  AOI22_X1 U23224 ( .A1(n20735), .A2(n20298), .B1(n20734), .B2(n20297), .ZN(
        n20287) );
  INV_X1 U23225 ( .A(n20739), .ZN(n20689) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20300), .B1(
        n20326), .B2(n20689), .ZN(n20286) );
  OAI211_X1 U23227 ( .C1(n20692), .C2(n20292), .A(n20287), .B(n20286), .ZN(
        P1_U3043) );
  AOI22_X1 U23228 ( .A1(n20741), .A2(n20298), .B1(n20740), .B2(n20297), .ZN(
        n20289) );
  INV_X1 U23229 ( .A(n20745), .ZN(n20693) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20300), .B1(
        n20326), .B2(n20693), .ZN(n20288) );
  OAI211_X1 U23231 ( .C1(n20696), .C2(n20292), .A(n20289), .B(n20288), .ZN(
        P1_U3044) );
  AOI22_X1 U23232 ( .A1(n20747), .A2(n20298), .B1(n20746), .B2(n20297), .ZN(
        n20291) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20300), .B1(
        n20326), .B2(n20748), .ZN(n20290) );
  OAI211_X1 U23234 ( .C1(n20751), .C2(n20292), .A(n20291), .B(n20290), .ZN(
        P1_U3045) );
  AOI22_X1 U23235 ( .A1(n9795), .A2(n20298), .B1(n20752), .B2(n20297), .ZN(
        n20294) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20754), .ZN(n20293) );
  OAI211_X1 U23237 ( .C1(n20757), .C2(n20325), .A(n20294), .B(n20293), .ZN(
        P1_U3046) );
  AOI22_X1 U23238 ( .A1(n20759), .A2(n20298), .B1(n20758), .B2(n20297), .ZN(
        n20296) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20662), .ZN(n20295) );
  OAI211_X1 U23240 ( .C1(n20665), .C2(n20325), .A(n20296), .B(n20295), .ZN(
        P1_U3047) );
  AOI22_X1 U23241 ( .A1(n20769), .A2(n20298), .B1(n20767), .B2(n20297), .ZN(
        n20302) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20770), .ZN(n20301) );
  OAI211_X1 U23243 ( .C1(n20776), .C2(n20325), .A(n20302), .B(n20301), .ZN(
        P1_U3048) );
  NAND3_X1 U23244 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20574), .A3(
        n11859), .ZN(n20341) );
  NOR2_X1 U23245 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20341), .ZN(
        n20327) );
  INV_X1 U23246 ( .A(n20333), .ZN(n20303) );
  AOI22_X1 U23247 ( .A1(n20718), .A2(n20327), .B1(n20359), .B2(n20724), .ZN(
        n20312) );
  OAI21_X1 U23248 ( .B1(n20359), .B2(n20326), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20304) );
  NAND2_X1 U23249 ( .A1(n20304), .A2(n20846), .ZN(n20310) );
  NOR2_X1 U23250 ( .A1(n20335), .A2(n20613), .ZN(n20307) );
  INV_X1 U23251 ( .A(n20327), .ZN(n20305) );
  INV_X1 U23252 ( .A(n20536), .ZN(n20478) );
  NOR2_X1 U23253 ( .A1(n20478), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20421) );
  NOR2_X1 U23254 ( .A1(n20421), .A2(n20715), .ZN(n20424) );
  AOI211_X1 U23255 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20305), .A(n20424), 
        .B(n20480), .ZN(n20306) );
  INV_X1 U23256 ( .A(n20307), .ZN(n20309) );
  INV_X1 U23257 ( .A(n20421), .ZN(n20308) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20329), .B1(
        n20717), .B2(n20328), .ZN(n20311) );
  OAI211_X1 U23259 ( .C1(n20727), .C2(n20325), .A(n20312), .B(n20311), .ZN(
        P1_U3049) );
  AOI22_X1 U23260 ( .A1(n20729), .A2(n20327), .B1(n20326), .B2(n20730), .ZN(
        n20314) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20329), .B1(
        n20728), .B2(n20328), .ZN(n20313) );
  OAI211_X1 U23262 ( .C1(n20733), .C2(n20356), .A(n20314), .B(n20313), .ZN(
        P1_U3050) );
  AOI22_X1 U23263 ( .A1(n20735), .A2(n20327), .B1(n20326), .B2(n20736), .ZN(
        n20316) );
  AOI22_X1 U23264 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20329), .B1(
        n20734), .B2(n20328), .ZN(n20315) );
  OAI211_X1 U23265 ( .C1(n20739), .C2(n20356), .A(n20316), .B(n20315), .ZN(
        P1_U3051) );
  AOI22_X1 U23266 ( .A1(n20741), .A2(n20327), .B1(n20326), .B2(n20742), .ZN(
        n20318) );
  AOI22_X1 U23267 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20329), .B1(
        n20740), .B2(n20328), .ZN(n20317) );
  OAI211_X1 U23268 ( .C1(n20745), .C2(n20356), .A(n20318), .B(n20317), .ZN(
        P1_U3052) );
  AOI22_X1 U23269 ( .A1(n20747), .A2(n20327), .B1(n20359), .B2(n20748), .ZN(
        n20320) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20329), .B1(
        n20746), .B2(n20328), .ZN(n20319) );
  OAI211_X1 U23271 ( .C1(n20751), .C2(n20325), .A(n20320), .B(n20319), .ZN(
        P1_U3053) );
  AOI22_X1 U23272 ( .A1(n9795), .A2(n20327), .B1(n20326), .B2(n20754), .ZN(
        n20322) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20329), .B1(
        n20752), .B2(n20328), .ZN(n20321) );
  OAI211_X1 U23274 ( .C1(n20757), .C2(n20356), .A(n20322), .B(n20321), .ZN(
        P1_U3054) );
  AOI22_X1 U23275 ( .A1(n20759), .A2(n20327), .B1(n20359), .B2(n20760), .ZN(
        n20324) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20329), .B1(
        n20758), .B2(n20328), .ZN(n20323) );
  OAI211_X1 U23277 ( .C1(n20765), .C2(n20325), .A(n20324), .B(n20323), .ZN(
        P1_U3055) );
  AOI22_X1 U23278 ( .A1(n20769), .A2(n20327), .B1(n20326), .B2(n20770), .ZN(
        n20331) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20329), .B1(
        n20767), .B2(n20328), .ZN(n20330) );
  OAI211_X1 U23280 ( .C1(n20776), .C2(n20356), .A(n20331), .B(n20330), .ZN(
        P1_U3056) );
  NOR2_X1 U23281 ( .A1(n20575), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20360) );
  AOI22_X1 U23282 ( .A1(n20718), .A2(n20360), .B1(n20390), .B2(n20724), .ZN(
        n20345) );
  INV_X1 U23283 ( .A(n20332), .ZN(n20579) );
  OAI21_X1 U23284 ( .B1(n20333), .B2(n20579), .A(n20846), .ZN(n20342) );
  AND2_X1 U23285 ( .A1(n11939), .A2(n20334), .ZN(n20713) );
  INV_X1 U23286 ( .A(n20713), .ZN(n20451) );
  OR2_X1 U23287 ( .A1(n20335), .A2(n20451), .ZN(n20337) );
  INV_X1 U23288 ( .A(n20360), .ZN(n20336) );
  AND2_X1 U23289 ( .A1(n20337), .A2(n20336), .ZN(n20343) );
  INV_X1 U23290 ( .A(n20343), .ZN(n20340) );
  INV_X1 U23291 ( .A(n20722), .ZN(n20338) );
  AOI21_X1 U23292 ( .B1(n20859), .B2(n20341), .A(n20338), .ZN(n20339) );
  OAI21_X1 U23293 ( .B1(n20342), .B2(n20340), .A(n20339), .ZN(n20362) );
  OAI22_X1 U23294 ( .A1(n20343), .A2(n20342), .B1(n20715), .B2(n20341), .ZN(
        n20361) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20362), .B1(
        n20717), .B2(n20361), .ZN(n20344) );
  OAI211_X1 U23296 ( .C1(n20727), .C2(n20356), .A(n20345), .B(n20344), .ZN(
        P1_U3057) );
  AOI22_X1 U23297 ( .A1(n20729), .A2(n20360), .B1(n20390), .B2(n20685), .ZN(
        n20347) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20362), .B1(
        n20728), .B2(n20361), .ZN(n20346) );
  OAI211_X1 U23299 ( .C1(n20688), .C2(n20356), .A(n20347), .B(n20346), .ZN(
        P1_U3058) );
  AOI22_X1 U23300 ( .A1(n20735), .A2(n20360), .B1(n20359), .B2(n20736), .ZN(
        n20349) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20362), .B1(
        n20734), .B2(n20361), .ZN(n20348) );
  OAI211_X1 U23302 ( .C1(n20739), .C2(n20387), .A(n20349), .B(n20348), .ZN(
        P1_U3059) );
  AOI22_X1 U23303 ( .A1(n20741), .A2(n20360), .B1(n20390), .B2(n20693), .ZN(
        n20351) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20362), .B1(
        n20740), .B2(n20361), .ZN(n20350) );
  OAI211_X1 U23305 ( .C1(n20696), .C2(n20356), .A(n20351), .B(n20350), .ZN(
        P1_U3060) );
  AOI22_X1 U23306 ( .A1(n20747), .A2(n20360), .B1(n20390), .B2(n20748), .ZN(
        n20353) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20362), .B1(
        n20746), .B2(n20361), .ZN(n20352) );
  OAI211_X1 U23308 ( .C1(n20751), .C2(n20356), .A(n20353), .B(n20352), .ZN(
        P1_U3061) );
  INV_X1 U23309 ( .A(n20757), .ZN(n20699) );
  AOI22_X1 U23310 ( .A1(n9795), .A2(n20360), .B1(n20390), .B2(n20699), .ZN(
        n20355) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20362), .B1(
        n20752), .B2(n20361), .ZN(n20354) );
  OAI211_X1 U23312 ( .C1(n20702), .C2(n20356), .A(n20355), .B(n20354), .ZN(
        P1_U3062) );
  AOI22_X1 U23313 ( .A1(n20759), .A2(n20360), .B1(n20359), .B2(n20662), .ZN(
        n20358) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20362), .B1(
        n20758), .B2(n20361), .ZN(n20357) );
  OAI211_X1 U23315 ( .C1(n20665), .C2(n20387), .A(n20358), .B(n20357), .ZN(
        P1_U3063) );
  AOI22_X1 U23316 ( .A1(n20769), .A2(n20360), .B1(n20359), .B2(n20770), .ZN(
        n20364) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20362), .B1(
        n20767), .B2(n20361), .ZN(n20363) );
  OAI211_X1 U23318 ( .C1(n20776), .C2(n20387), .A(n20364), .B(n20363), .ZN(
        P1_U3064) );
  NAND3_X1 U23319 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20574), .A3(
        n20539), .ZN(n20395) );
  NOR2_X1 U23320 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20395), .ZN(
        n20389) );
  NOR2_X1 U23321 ( .A1(n20612), .A2(n20365), .ZN(n20420) );
  NAND2_X1 U23322 ( .A1(n20420), .A2(n20846), .ZN(n20452) );
  OAI22_X1 U23323 ( .A1(n20452), .A2(n20678), .B1(n20673), .B2(n20366), .ZN(
        n20388) );
  AOI22_X1 U23324 ( .A1(n20718), .A2(n20389), .B1(n20717), .B2(n20388), .ZN(
        n20373) );
  AOI21_X1 U23325 ( .B1(n20387), .B2(n20417), .A(n20847), .ZN(n20368) );
  AOI21_X1 U23326 ( .B1(n20420), .B2(n20613), .A(n20368), .ZN(n20369) );
  NOR2_X1 U23327 ( .A1(n20369), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20371) );
  INV_X1 U23328 ( .A(n20417), .ZN(n20384) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20391), .B1(
        n20384), .B2(n20724), .ZN(n20372) );
  OAI211_X1 U23330 ( .C1(n20727), .C2(n20387), .A(n20373), .B(n20372), .ZN(
        P1_U3065) );
  AOI22_X1 U23331 ( .A1(n20729), .A2(n20389), .B1(n20728), .B2(n20388), .ZN(
        n20375) );
  AOI22_X1 U23332 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20730), .ZN(n20374) );
  OAI211_X1 U23333 ( .C1(n20733), .C2(n20417), .A(n20375), .B(n20374), .ZN(
        P1_U3066) );
  AOI22_X1 U23334 ( .A1(n20735), .A2(n20389), .B1(n20734), .B2(n20388), .ZN(
        n20377) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20736), .ZN(n20376) );
  OAI211_X1 U23336 ( .C1(n20739), .C2(n20417), .A(n20377), .B(n20376), .ZN(
        P1_U3067) );
  AOI22_X1 U23337 ( .A1(n20741), .A2(n20389), .B1(n20740), .B2(n20388), .ZN(
        n20379) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20742), .ZN(n20378) );
  OAI211_X1 U23339 ( .C1(n20745), .C2(n20417), .A(n20379), .B(n20378), .ZN(
        P1_U3068) );
  AOI22_X1 U23340 ( .A1(n20747), .A2(n20389), .B1(n20746), .B2(n20388), .ZN(
        n20381) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20391), .B1(
        n20384), .B2(n20748), .ZN(n20380) );
  OAI211_X1 U23342 ( .C1(n20751), .C2(n20387), .A(n20381), .B(n20380), .ZN(
        P1_U3069) );
  AOI22_X1 U23343 ( .A1(n9795), .A2(n20389), .B1(n20752), .B2(n20388), .ZN(
        n20383) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20754), .ZN(n20382) );
  OAI211_X1 U23345 ( .C1(n20757), .C2(n20417), .A(n20383), .B(n20382), .ZN(
        P1_U3070) );
  AOI22_X1 U23346 ( .A1(n20759), .A2(n20389), .B1(n20758), .B2(n20388), .ZN(
        n20386) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20391), .B1(
        n20384), .B2(n20760), .ZN(n20385) );
  OAI211_X1 U23348 ( .C1(n20765), .C2(n20387), .A(n20386), .B(n20385), .ZN(
        P1_U3071) );
  AOI22_X1 U23349 ( .A1(n20769), .A2(n20389), .B1(n20767), .B2(n20388), .ZN(
        n20393) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20391), .B1(
        n20390), .B2(n20770), .ZN(n20392) );
  OAI211_X1 U23351 ( .C1(n20776), .C2(n20417), .A(n20393), .B(n20392), .ZN(
        P1_U3072) );
  NOR2_X1 U23352 ( .A1(n20863), .A2(n20395), .ZN(n20413) );
  INV_X1 U23353 ( .A(n20413), .ZN(n20394) );
  OAI222_X1 U23354 ( .A1(n20394), .A2(n20859), .B1(n20715), .B2(n20395), .C1(
        n20276), .C2(n20452), .ZN(n20412) );
  AOI22_X1 U23355 ( .A1(n20718), .A2(n20413), .B1(n20717), .B2(n20412), .ZN(
        n20399) );
  INV_X1 U23356 ( .A(n20449), .ZN(n20454) );
  OAI21_X1 U23357 ( .B1(n20454), .B2(n20396), .A(n20395), .ZN(n20397) );
  NAND2_X1 U23358 ( .A1(n20397), .A2(n20722), .ZN(n20414) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20414), .B1(
        n20442), .B2(n20724), .ZN(n20398) );
  OAI211_X1 U23360 ( .C1(n20727), .C2(n20417), .A(n20399), .B(n20398), .ZN(
        P1_U3073) );
  AOI22_X1 U23361 ( .A1(n20729), .A2(n20413), .B1(n20728), .B2(n20412), .ZN(
        n20401) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20414), .B1(
        n20442), .B2(n20685), .ZN(n20400) );
  OAI211_X1 U23363 ( .C1(n20688), .C2(n20417), .A(n20401), .B(n20400), .ZN(
        P1_U3074) );
  AOI22_X1 U23364 ( .A1(n20735), .A2(n20413), .B1(n20734), .B2(n20412), .ZN(
        n20403) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20414), .B1(
        n20442), .B2(n20689), .ZN(n20402) );
  OAI211_X1 U23366 ( .C1(n20692), .C2(n20417), .A(n20403), .B(n20402), .ZN(
        P1_U3075) );
  AOI22_X1 U23367 ( .A1(n20741), .A2(n20413), .B1(n20740), .B2(n20412), .ZN(
        n20405) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20414), .B1(
        n20442), .B2(n20693), .ZN(n20404) );
  OAI211_X1 U23369 ( .C1(n20696), .C2(n20417), .A(n20405), .B(n20404), .ZN(
        P1_U3076) );
  AOI22_X1 U23370 ( .A1(n20747), .A2(n20413), .B1(n20746), .B2(n20412), .ZN(
        n20407) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20414), .B1(
        n20442), .B2(n20748), .ZN(n20406) );
  OAI211_X1 U23372 ( .C1(n20751), .C2(n20417), .A(n20407), .B(n20406), .ZN(
        P1_U3077) );
  AOI22_X1 U23373 ( .A1(n9795), .A2(n20413), .B1(n20752), .B2(n20412), .ZN(
        n20409) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20414), .B1(
        n20442), .B2(n20699), .ZN(n20408) );
  OAI211_X1 U23375 ( .C1(n20702), .C2(n20417), .A(n20409), .B(n20408), .ZN(
        P1_U3078) );
  AOI22_X1 U23376 ( .A1(n20759), .A2(n20413), .B1(n20758), .B2(n20412), .ZN(
        n20411) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20414), .B1(
        n20442), .B2(n20760), .ZN(n20410) );
  OAI211_X1 U23378 ( .C1(n20765), .C2(n20417), .A(n20411), .B(n20410), .ZN(
        P1_U3079) );
  AOI22_X1 U23379 ( .A1(n20769), .A2(n20413), .B1(n20767), .B2(n20412), .ZN(
        n20416) );
  INV_X1 U23380 ( .A(n20776), .ZN(n20707) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20414), .B1(
        n20442), .B2(n20707), .ZN(n20415) );
  OAI211_X1 U23382 ( .C1(n20712), .C2(n20417), .A(n20416), .B(n20415), .ZN(
        P1_U3080) );
  INV_X1 U23383 ( .A(n20442), .ZN(n20418) );
  NAND2_X1 U23384 ( .A1(n20418), .A2(n20846), .ZN(n20419) );
  OAI21_X1 U23385 ( .B1(n20419), .B2(n20472), .A(n20609), .ZN(n20426) );
  AND2_X1 U23386 ( .A1(n20420), .A2(n20678), .ZN(n20423) );
  INV_X1 U23387 ( .A(n20673), .ZN(n20422) );
  NOR2_X1 U23388 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20453), .ZN(
        n20443) );
  INV_X1 U23389 ( .A(n20727), .ZN(n20646) );
  AOI22_X1 U23390 ( .A1(n20718), .A2(n20443), .B1(n20442), .B2(n20646), .ZN(
        n20429) );
  INV_X1 U23391 ( .A(n20423), .ZN(n20425) );
  AOI21_X1 U23392 ( .B1(n20426), .B2(n20425), .A(n20424), .ZN(n20427) );
  OAI211_X1 U23393 ( .C1(n20443), .C2(n20615), .A(n20681), .B(n20427), .ZN(
        n20444) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20444), .B1(
        n20472), .B2(n20724), .ZN(n20428) );
  OAI211_X1 U23395 ( .C1(n20447), .C2(n20548), .A(n20429), .B(n20428), .ZN(
        P1_U3081) );
  AOI22_X1 U23396 ( .A1(n20729), .A2(n20443), .B1(n20442), .B2(n20730), .ZN(
        n20431) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20444), .B1(
        n20472), .B2(n20685), .ZN(n20430) );
  OAI211_X1 U23398 ( .C1(n20447), .C2(n20551), .A(n20431), .B(n20430), .ZN(
        P1_U3082) );
  AOI22_X1 U23399 ( .A1(n20735), .A2(n20443), .B1(n20472), .B2(n20689), .ZN(
        n20433) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20444), .B1(
        n20442), .B2(n20736), .ZN(n20432) );
  OAI211_X1 U23401 ( .C1(n20447), .C2(n20554), .A(n20433), .B(n20432), .ZN(
        P1_U3083) );
  AOI22_X1 U23402 ( .A1(n20741), .A2(n20443), .B1(n20472), .B2(n20693), .ZN(
        n20435) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20444), .B1(
        n20442), .B2(n20742), .ZN(n20434) );
  OAI211_X1 U23404 ( .C1(n20447), .C2(n20557), .A(n20435), .B(n20434), .ZN(
        P1_U3084) );
  AOI22_X1 U23405 ( .A1(n20747), .A2(n20443), .B1(n20472), .B2(n20748), .ZN(
        n20437) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20444), .B1(
        n20442), .B2(n20656), .ZN(n20436) );
  OAI211_X1 U23407 ( .C1(n20447), .C2(n20560), .A(n20437), .B(n20436), .ZN(
        P1_U3085) );
  AOI22_X1 U23408 ( .A1(n9795), .A2(n20443), .B1(n20472), .B2(n20699), .ZN(
        n20439) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20444), .B1(
        n20442), .B2(n20754), .ZN(n20438) );
  OAI211_X1 U23410 ( .C1(n20447), .C2(n20563), .A(n20439), .B(n20438), .ZN(
        P1_U3086) );
  AOI22_X1 U23411 ( .A1(n20759), .A2(n20443), .B1(n20472), .B2(n20760), .ZN(
        n20441) );
  AOI22_X1 U23412 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20444), .B1(
        n20442), .B2(n20662), .ZN(n20440) );
  OAI211_X1 U23413 ( .C1(n20447), .C2(n20566), .A(n20441), .B(n20440), .ZN(
        P1_U3087) );
  AOI22_X1 U23414 ( .A1(n20769), .A2(n20443), .B1(n20442), .B2(n20770), .ZN(
        n20446) );
  AOI22_X1 U23415 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20444), .B1(
        n20472), .B2(n20707), .ZN(n20445) );
  OAI211_X1 U23416 ( .C1(n20447), .C2(n20572), .A(n20446), .B(n20445), .ZN(
        P1_U3088) );
  INV_X1 U23417 ( .A(n20448), .ZN(n20583) );
  OAI222_X1 U23418 ( .A1(n20452), .A2(n20451), .B1(n20715), .B2(n20453), .C1(
        n20859), .C2(n20450), .ZN(n20470) );
  AOI22_X1 U23419 ( .A1(n20718), .A2(n20471), .B1(n20717), .B2(n20470), .ZN(
        n20457) );
  INV_X1 U23420 ( .A(n20453), .ZN(n20455) );
  NOR3_X1 U23421 ( .A1(n20454), .A2(n20859), .A3(n20579), .ZN(n20851) );
  OAI21_X1 U23422 ( .B1(n20455), .B2(n20851), .A(n20722), .ZN(n20473) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20646), .ZN(n20456) );
  OAI211_X1 U23424 ( .C1(n20649), .C2(n20507), .A(n20457), .B(n20456), .ZN(
        P1_U3089) );
  AOI22_X1 U23425 ( .A1(n20729), .A2(n20471), .B1(n20728), .B2(n20470), .ZN(
        n20459) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20730), .ZN(n20458) );
  OAI211_X1 U23427 ( .C1(n20733), .C2(n20507), .A(n20459), .B(n20458), .ZN(
        P1_U3090) );
  AOI22_X1 U23428 ( .A1(n20735), .A2(n20471), .B1(n20734), .B2(n20470), .ZN(
        n20461) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20736), .ZN(n20460) );
  OAI211_X1 U23430 ( .C1(n20739), .C2(n20507), .A(n20461), .B(n20460), .ZN(
        P1_U3091) );
  AOI22_X1 U23431 ( .A1(n20741), .A2(n20471), .B1(n20740), .B2(n20470), .ZN(
        n20463) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20742), .ZN(n20462) );
  OAI211_X1 U23433 ( .C1(n20745), .C2(n20507), .A(n20463), .B(n20462), .ZN(
        P1_U3092) );
  AOI22_X1 U23434 ( .A1(n20747), .A2(n20471), .B1(n20746), .B2(n20470), .ZN(
        n20465) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20656), .ZN(n20464) );
  OAI211_X1 U23436 ( .C1(n20659), .C2(n20507), .A(n20465), .B(n20464), .ZN(
        P1_U3093) );
  AOI22_X1 U23437 ( .A1(n9795), .A2(n20471), .B1(n20752), .B2(n20470), .ZN(
        n20467) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20754), .ZN(n20466) );
  OAI211_X1 U23439 ( .C1(n20757), .C2(n20507), .A(n20467), .B(n20466), .ZN(
        P1_U3094) );
  AOI22_X1 U23440 ( .A1(n20759), .A2(n20471), .B1(n20758), .B2(n20470), .ZN(
        n20469) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20662), .ZN(n20468) );
  OAI211_X1 U23442 ( .C1(n20665), .C2(n20507), .A(n20469), .B(n20468), .ZN(
        P1_U3095) );
  AOI22_X1 U23443 ( .A1(n20769), .A2(n20471), .B1(n20767), .B2(n20470), .ZN(
        n20475) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20770), .ZN(n20474) );
  OAI211_X1 U23445 ( .C1(n20776), .C2(n20507), .A(n20475), .B(n20474), .ZN(
        P1_U3096) );
  NOR3_X1 U23446 ( .A1(n20574), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20511) );
  INV_X1 U23447 ( .A(n20511), .ZN(n20508) );
  NOR2_X1 U23448 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20508), .ZN(
        n20502) );
  AND2_X1 U23449 ( .A1(n20476), .A2(n20612), .ZN(n20576) );
  AOI21_X1 U23450 ( .B1(n20576), .B2(n20613), .A(n20502), .ZN(n20484) );
  NAND2_X1 U23451 ( .A1(n20478), .A2(n20477), .ZN(n20617) );
  OAI22_X1 U23452 ( .A1(n20484), .A2(n20859), .B1(n20479), .B2(n20617), .ZN(
        n20501) );
  AOI22_X1 U23453 ( .A1(n20718), .A2(n20502), .B1(n20717), .B2(n20501), .ZN(
        n20488) );
  INV_X1 U23454 ( .A(n20480), .ZN(n20541) );
  INV_X1 U23455 ( .A(n20507), .ZN(n20483) );
  OAI21_X1 U23456 ( .B1(n20503), .B2(n20483), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20485) );
  NAND2_X1 U23457 ( .A1(n20485), .A2(n20484), .ZN(n20486) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20504), .B1(
        n20503), .B2(n20724), .ZN(n20487) );
  OAI211_X1 U23459 ( .C1(n20727), .C2(n20507), .A(n20488), .B(n20487), .ZN(
        P1_U3097) );
  AOI22_X1 U23460 ( .A1(n20729), .A2(n20502), .B1(n20728), .B2(n20501), .ZN(
        n20490) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20504), .B1(
        n20503), .B2(n20685), .ZN(n20489) );
  OAI211_X1 U23462 ( .C1(n20688), .C2(n20507), .A(n20490), .B(n20489), .ZN(
        P1_U3098) );
  AOI22_X1 U23463 ( .A1(n20735), .A2(n20502), .B1(n20734), .B2(n20501), .ZN(
        n20492) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20504), .B1(
        n20503), .B2(n20689), .ZN(n20491) );
  OAI211_X1 U23465 ( .C1(n20692), .C2(n20507), .A(n20492), .B(n20491), .ZN(
        P1_U3099) );
  AOI22_X1 U23466 ( .A1(n20741), .A2(n20502), .B1(n20740), .B2(n20501), .ZN(
        n20494) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20504), .B1(
        n20503), .B2(n20693), .ZN(n20493) );
  OAI211_X1 U23468 ( .C1(n20696), .C2(n20507), .A(n20494), .B(n20493), .ZN(
        P1_U3100) );
  AOI22_X1 U23469 ( .A1(n20747), .A2(n20502), .B1(n20746), .B2(n20501), .ZN(
        n20496) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20504), .B1(
        n20503), .B2(n20748), .ZN(n20495) );
  OAI211_X1 U23471 ( .C1(n20751), .C2(n20507), .A(n20496), .B(n20495), .ZN(
        P1_U3101) );
  AOI22_X1 U23472 ( .A1(n9795), .A2(n20502), .B1(n20752), .B2(n20501), .ZN(
        n20498) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20504), .B1(
        n20503), .B2(n20699), .ZN(n20497) );
  OAI211_X1 U23474 ( .C1(n20702), .C2(n20507), .A(n20498), .B(n20497), .ZN(
        P1_U3102) );
  AOI22_X1 U23475 ( .A1(n20759), .A2(n20502), .B1(n20758), .B2(n20501), .ZN(
        n20500) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20504), .B1(
        n20503), .B2(n20760), .ZN(n20499) );
  OAI211_X1 U23477 ( .C1(n20765), .C2(n20507), .A(n20500), .B(n20499), .ZN(
        P1_U3103) );
  AOI22_X1 U23478 ( .A1(n20769), .A2(n20502), .B1(n20767), .B2(n20501), .ZN(
        n20506) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20504), .B1(
        n20503), .B2(n20707), .ZN(n20505) );
  OAI211_X1 U23480 ( .C1(n20712), .C2(n20507), .A(n20506), .B(n20505), .ZN(
        P1_U3104) );
  NOR2_X1 U23481 ( .A1(n20863), .A2(n20508), .ZN(n20528) );
  AOI21_X1 U23482 ( .B1(n20576), .B2(n20641), .A(n20528), .ZN(n20509) );
  OAI22_X1 U23483 ( .A1(n20509), .A2(n20859), .B1(n20508), .B2(n20715), .ZN(
        n20527) );
  AOI22_X1 U23484 ( .A1(n20718), .A2(n20528), .B1(n20717), .B2(n20527), .ZN(
        n20514) );
  OAI21_X1 U23485 ( .B1(n20580), .B2(n20847), .A(n20509), .ZN(n20510) );
  OAI221_X1 U23486 ( .B1(n20846), .B2(n20511), .C1(n20859), .C2(n20510), .A(
        n20722), .ZN(n20529) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20529), .B1(
        n20568), .B2(n20724), .ZN(n20513) );
  OAI211_X1 U23488 ( .C1(n20727), .C2(n20532), .A(n20514), .B(n20513), .ZN(
        P1_U3105) );
  AOI22_X1 U23489 ( .A1(n20729), .A2(n20528), .B1(n20728), .B2(n20527), .ZN(
        n20516) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20529), .B1(
        n20568), .B2(n20685), .ZN(n20515) );
  OAI211_X1 U23491 ( .C1(n20688), .C2(n20532), .A(n20516), .B(n20515), .ZN(
        P1_U3106) );
  AOI22_X1 U23492 ( .A1(n20735), .A2(n20528), .B1(n20734), .B2(n20527), .ZN(
        n20518) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20529), .B1(
        n20568), .B2(n20689), .ZN(n20517) );
  OAI211_X1 U23494 ( .C1(n20692), .C2(n20532), .A(n20518), .B(n20517), .ZN(
        P1_U3107) );
  AOI22_X1 U23495 ( .A1(n20741), .A2(n20528), .B1(n20740), .B2(n20527), .ZN(
        n20520) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20529), .B1(
        n20568), .B2(n20693), .ZN(n20519) );
  OAI211_X1 U23497 ( .C1(n20696), .C2(n20532), .A(n20520), .B(n20519), .ZN(
        P1_U3108) );
  AOI22_X1 U23498 ( .A1(n20747), .A2(n20528), .B1(n20746), .B2(n20527), .ZN(
        n20522) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20529), .B1(
        n20568), .B2(n20748), .ZN(n20521) );
  OAI211_X1 U23500 ( .C1(n20751), .C2(n20532), .A(n20522), .B(n20521), .ZN(
        P1_U3109) );
  AOI22_X1 U23501 ( .A1(n9795), .A2(n20528), .B1(n20752), .B2(n20527), .ZN(
        n20524) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20529), .B1(
        n20568), .B2(n20699), .ZN(n20523) );
  OAI211_X1 U23503 ( .C1(n20702), .C2(n20532), .A(n20524), .B(n20523), .ZN(
        P1_U3110) );
  AOI22_X1 U23504 ( .A1(n20759), .A2(n20528), .B1(n20758), .B2(n20527), .ZN(
        n20526) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20529), .B1(
        n20568), .B2(n20760), .ZN(n20525) );
  OAI211_X1 U23506 ( .C1(n20765), .C2(n20532), .A(n20526), .B(n20525), .ZN(
        P1_U3111) );
  AOI22_X1 U23507 ( .A1(n20769), .A2(n20528), .B1(n20767), .B2(n20527), .ZN(
        n20531) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20529), .B1(
        n20568), .B2(n20707), .ZN(n20530) );
  OAI211_X1 U23509 ( .C1(n20712), .C2(n20532), .A(n20531), .B(n20530), .ZN(
        P1_U3112) );
  INV_X1 U23510 ( .A(n20533), .ZN(n20675) );
  INV_X1 U23511 ( .A(n20568), .ZN(n20534) );
  NAND3_X1 U23512 ( .A1(n20606), .A2(n20534), .A3(n20846), .ZN(n20535) );
  NAND2_X1 U23513 ( .A1(n20535), .A2(n20609), .ZN(n20544) );
  AND2_X1 U23514 ( .A1(n20576), .A2(n20678), .ZN(n20540) );
  NAND2_X1 U23515 ( .A1(n20536), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20674) );
  INV_X1 U23516 ( .A(n20674), .ZN(n20537) );
  NOR3_X1 U23517 ( .A1(n20574), .A2(n20539), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20582) );
  INV_X1 U23518 ( .A(n20582), .ZN(n20577) );
  NOR2_X1 U23519 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20577), .ZN(
        n20567) );
  AOI22_X1 U23520 ( .A1(n20718), .A2(n20567), .B1(n20568), .B2(n20646), .ZN(
        n20547) );
  INV_X1 U23521 ( .A(n20540), .ZN(n20543) );
  NAND2_X1 U23522 ( .A1(n20674), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20680) );
  OAI211_X1 U23523 ( .C1(n20615), .C2(n20567), .A(n20680), .B(n20541), .ZN(
        n20542) );
  AOI21_X1 U23524 ( .B1(n20544), .B2(n20543), .A(n20542), .ZN(n20545) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20569), .B1(
        n20587), .B2(n20724), .ZN(n20546) );
  OAI211_X1 U23526 ( .C1(n20573), .C2(n20548), .A(n20547), .B(n20546), .ZN(
        P1_U3113) );
  AOI22_X1 U23527 ( .A1(n20729), .A2(n20567), .B1(n20568), .B2(n20730), .ZN(
        n20550) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20569), .B1(
        n20587), .B2(n20685), .ZN(n20549) );
  OAI211_X1 U23529 ( .C1(n20573), .C2(n20551), .A(n20550), .B(n20549), .ZN(
        P1_U3114) );
  AOI22_X1 U23530 ( .A1(n20735), .A2(n20567), .B1(n20568), .B2(n20736), .ZN(
        n20553) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20569), .B1(
        n20587), .B2(n20689), .ZN(n20552) );
  OAI211_X1 U23532 ( .C1(n20573), .C2(n20554), .A(n20553), .B(n20552), .ZN(
        P1_U3115) );
  AOI22_X1 U23533 ( .A1(n20741), .A2(n20567), .B1(n20568), .B2(n20742), .ZN(
        n20556) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20569), .B1(
        n20587), .B2(n20693), .ZN(n20555) );
  OAI211_X1 U23535 ( .C1(n20573), .C2(n20557), .A(n20556), .B(n20555), .ZN(
        P1_U3116) );
  AOI22_X1 U23536 ( .A1(n20747), .A2(n20567), .B1(n20587), .B2(n20748), .ZN(
        n20559) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20569), .B1(
        n20568), .B2(n20656), .ZN(n20558) );
  OAI211_X1 U23538 ( .C1(n20573), .C2(n20560), .A(n20559), .B(n20558), .ZN(
        P1_U3117) );
  AOI22_X1 U23539 ( .A1(n9795), .A2(n20567), .B1(n20568), .B2(n20754), .ZN(
        n20562) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20569), .B1(
        n20587), .B2(n20699), .ZN(n20561) );
  OAI211_X1 U23541 ( .C1(n20573), .C2(n20563), .A(n20562), .B(n20561), .ZN(
        P1_U3118) );
  AOI22_X1 U23542 ( .A1(n20759), .A2(n20567), .B1(n20568), .B2(n20662), .ZN(
        n20565) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20569), .B1(
        n20587), .B2(n20760), .ZN(n20564) );
  OAI211_X1 U23544 ( .C1(n20573), .C2(n20566), .A(n20565), .B(n20564), .ZN(
        P1_U3119) );
  AOI22_X1 U23545 ( .A1(n20769), .A2(n20567), .B1(n20587), .B2(n20707), .ZN(
        n20571) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20569), .B1(
        n20568), .B2(n20770), .ZN(n20570) );
  OAI211_X1 U23547 ( .C1(n20573), .C2(n20572), .A(n20571), .B(n20570), .ZN(
        P1_U3120) );
  NOR2_X1 U23548 ( .A1(n20575), .A2(n20574), .ZN(n20601) );
  AOI21_X1 U23549 ( .B1(n20576), .B2(n20713), .A(n20601), .ZN(n20578) );
  OAI22_X1 U23550 ( .A1(n20578), .A2(n20859), .B1(n20577), .B2(n20715), .ZN(
        n20600) );
  AOI22_X1 U23551 ( .A1(n20718), .A2(n20601), .B1(n20717), .B2(n20600), .ZN(
        n20586) );
  OAI21_X1 U23552 ( .B1(n20580), .B2(n20579), .A(n20578), .ZN(n20581) );
  OAI221_X1 U23553 ( .B1(n20846), .B2(n20582), .C1(n20859), .C2(n20581), .A(
        n20722), .ZN(n20603) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20724), .ZN(n20585) );
  OAI211_X1 U23555 ( .C1(n20727), .C2(n20606), .A(n20586), .B(n20585), .ZN(
        P1_U3121) );
  AOI22_X1 U23556 ( .A1(n20729), .A2(n20601), .B1(n20728), .B2(n20600), .ZN(
        n20589) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20603), .B1(
        n20587), .B2(n20730), .ZN(n20588) );
  OAI211_X1 U23558 ( .C1(n20733), .C2(n20639), .A(n20589), .B(n20588), .ZN(
        P1_U3122) );
  AOI22_X1 U23559 ( .A1(n20735), .A2(n20601), .B1(n20734), .B2(n20600), .ZN(
        n20591) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20689), .ZN(n20590) );
  OAI211_X1 U23561 ( .C1(n20692), .C2(n20606), .A(n20591), .B(n20590), .ZN(
        P1_U3123) );
  AOI22_X1 U23562 ( .A1(n20741), .A2(n20601), .B1(n20740), .B2(n20600), .ZN(
        n20593) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20693), .ZN(n20592) );
  OAI211_X1 U23564 ( .C1(n20696), .C2(n20606), .A(n20593), .B(n20592), .ZN(
        P1_U3124) );
  AOI22_X1 U23565 ( .A1(n20747), .A2(n20601), .B1(n20746), .B2(n20600), .ZN(
        n20595) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20748), .ZN(n20594) );
  OAI211_X1 U23567 ( .C1(n20751), .C2(n20606), .A(n20595), .B(n20594), .ZN(
        P1_U3125) );
  AOI22_X1 U23568 ( .A1(n9795), .A2(n20601), .B1(n20752), .B2(n20600), .ZN(
        n20597) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20699), .ZN(n20596) );
  OAI211_X1 U23570 ( .C1(n20702), .C2(n20606), .A(n20597), .B(n20596), .ZN(
        P1_U3126) );
  AOI22_X1 U23571 ( .A1(n20759), .A2(n20601), .B1(n20758), .B2(n20600), .ZN(
        n20599) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20760), .ZN(n20598) );
  OAI211_X1 U23573 ( .C1(n20765), .C2(n20606), .A(n20599), .B(n20598), .ZN(
        P1_U3127) );
  AOI22_X1 U23574 ( .A1(n20769), .A2(n20601), .B1(n20767), .B2(n20600), .ZN(
        n20605) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20603), .B1(
        n20602), .B2(n20707), .ZN(n20604) );
  OAI211_X1 U23576 ( .C1(n20712), .C2(n20606), .A(n20605), .B(n20604), .ZN(
        P1_U3128) );
  NOR3_X1 U23577 ( .A1(n11859), .A2(n20574), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20645) );
  INV_X1 U23578 ( .A(n20645), .ZN(n20642) );
  NOR2_X1 U23579 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20642), .ZN(
        n20634) );
  OR2_X1 U23580 ( .A1(n20676), .A2(n20607), .ZN(n20608) );
  AOI22_X1 U23581 ( .A1(n20718), .A2(n20634), .B1(n20668), .B2(n20724), .ZN(
        n20621) );
  NAND3_X1 U23582 ( .A1(n20639), .A2(n20846), .A3(n20608), .ZN(n20610) );
  NAND2_X1 U23583 ( .A1(n20610), .A2(n20609), .ZN(n20616) );
  NOR2_X1 U23584 ( .A1(n20612), .A2(n20611), .ZN(n20714) );
  NAND2_X1 U23585 ( .A1(n20714), .A2(n20613), .ZN(n20618) );
  AOI22_X1 U23586 ( .A1(n20616), .A2(n20618), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20617), .ZN(n20614) );
  OAI211_X1 U23587 ( .C1(n20634), .C2(n20615), .A(n20681), .B(n20614), .ZN(
        n20636) );
  INV_X1 U23588 ( .A(n20616), .ZN(n20619) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20636), .B1(
        n20717), .B2(n20635), .ZN(n20620) );
  OAI211_X1 U23590 ( .C1(n20727), .C2(n20639), .A(n20621), .B(n20620), .ZN(
        P1_U3129) );
  AOI22_X1 U23591 ( .A1(n20729), .A2(n20634), .B1(n20668), .B2(n20685), .ZN(
        n20623) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20636), .B1(
        n20728), .B2(n20635), .ZN(n20622) );
  OAI211_X1 U23593 ( .C1(n20688), .C2(n20639), .A(n20623), .B(n20622), .ZN(
        P1_U3130) );
  AOI22_X1 U23594 ( .A1(n20735), .A2(n20634), .B1(n20668), .B2(n20689), .ZN(
        n20625) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20636), .B1(
        n20734), .B2(n20635), .ZN(n20624) );
  OAI211_X1 U23596 ( .C1(n20692), .C2(n20639), .A(n20625), .B(n20624), .ZN(
        P1_U3131) );
  AOI22_X1 U23597 ( .A1(n20741), .A2(n20634), .B1(n20668), .B2(n20693), .ZN(
        n20627) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20636), .B1(
        n20740), .B2(n20635), .ZN(n20626) );
  OAI211_X1 U23599 ( .C1(n20696), .C2(n20639), .A(n20627), .B(n20626), .ZN(
        P1_U3132) );
  AOI22_X1 U23600 ( .A1(n20747), .A2(n20634), .B1(n20668), .B2(n20748), .ZN(
        n20629) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20636), .B1(
        n20746), .B2(n20635), .ZN(n20628) );
  OAI211_X1 U23602 ( .C1(n20751), .C2(n20639), .A(n20629), .B(n20628), .ZN(
        P1_U3133) );
  AOI22_X1 U23603 ( .A1(n9795), .A2(n20634), .B1(n20668), .B2(n20699), .ZN(
        n20631) );
  AOI22_X1 U23604 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20636), .B1(
        n20752), .B2(n20635), .ZN(n20630) );
  OAI211_X1 U23605 ( .C1(n20702), .C2(n20639), .A(n20631), .B(n20630), .ZN(
        P1_U3134) );
  AOI22_X1 U23606 ( .A1(n20759), .A2(n20634), .B1(n20668), .B2(n20760), .ZN(
        n20633) );
  AOI22_X1 U23607 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20636), .B1(
        n20758), .B2(n20635), .ZN(n20632) );
  OAI211_X1 U23608 ( .C1(n20765), .C2(n20639), .A(n20633), .B(n20632), .ZN(
        P1_U3135) );
  AOI22_X1 U23609 ( .A1(n20769), .A2(n20634), .B1(n20668), .B2(n20707), .ZN(
        n20638) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20636), .B1(
        n20767), .B2(n20635), .ZN(n20637) );
  OAI211_X1 U23611 ( .C1(n20712), .C2(n20639), .A(n20638), .B(n20637), .ZN(
        P1_U3136) );
  INV_X1 U23612 ( .A(n20676), .ZN(n20854) );
  NOR2_X1 U23613 ( .A1(n20863), .A2(n20642), .ZN(n20667) );
  AOI21_X1 U23614 ( .B1(n20714), .B2(n20641), .A(n20667), .ZN(n20643) );
  OAI22_X1 U23615 ( .A1(n20643), .A2(n20859), .B1(n20642), .B2(n20715), .ZN(
        n20666) );
  AOI22_X1 U23616 ( .A1(n20718), .A2(n20667), .B1(n20717), .B2(n20666), .ZN(
        n20648) );
  OAI21_X1 U23617 ( .B1(n20676), .B2(n20847), .A(n20643), .ZN(n20644) );
  OAI221_X1 U23618 ( .B1(n20846), .B2(n20645), .C1(n20859), .C2(n20644), .A(
        n20722), .ZN(n20669) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20646), .ZN(n20647) );
  OAI211_X1 U23620 ( .C1(n20649), .C2(n20711), .A(n20648), .B(n20647), .ZN(
        P1_U3137) );
  AOI22_X1 U23621 ( .A1(n20729), .A2(n20667), .B1(n20728), .B2(n20666), .ZN(
        n20651) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20730), .ZN(n20650) );
  OAI211_X1 U23623 ( .C1(n20733), .C2(n20711), .A(n20651), .B(n20650), .ZN(
        P1_U3138) );
  AOI22_X1 U23624 ( .A1(n20735), .A2(n20667), .B1(n20734), .B2(n20666), .ZN(
        n20653) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20736), .ZN(n20652) );
  OAI211_X1 U23626 ( .C1(n20739), .C2(n20711), .A(n20653), .B(n20652), .ZN(
        P1_U3139) );
  AOI22_X1 U23627 ( .A1(n20741), .A2(n20667), .B1(n20740), .B2(n20666), .ZN(
        n20655) );
  AOI22_X1 U23628 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20742), .ZN(n20654) );
  OAI211_X1 U23629 ( .C1(n20745), .C2(n20711), .A(n20655), .B(n20654), .ZN(
        P1_U3140) );
  AOI22_X1 U23630 ( .A1(n20747), .A2(n20667), .B1(n20746), .B2(n20666), .ZN(
        n20658) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20656), .ZN(n20657) );
  OAI211_X1 U23632 ( .C1(n20659), .C2(n20711), .A(n20658), .B(n20657), .ZN(
        P1_U3141) );
  AOI22_X1 U23633 ( .A1(n9795), .A2(n20667), .B1(n20752), .B2(n20666), .ZN(
        n20661) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20754), .ZN(n20660) );
  OAI211_X1 U23635 ( .C1(n20757), .C2(n20711), .A(n20661), .B(n20660), .ZN(
        P1_U3142) );
  AOI22_X1 U23636 ( .A1(n20759), .A2(n20667), .B1(n20758), .B2(n20666), .ZN(
        n20664) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20662), .ZN(n20663) );
  OAI211_X1 U23638 ( .C1(n20665), .C2(n20711), .A(n20664), .B(n20663), .ZN(
        P1_U3143) );
  AOI22_X1 U23639 ( .A1(n20769), .A2(n20667), .B1(n20767), .B2(n20666), .ZN(
        n20671) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20770), .ZN(n20670) );
  OAI211_X1 U23641 ( .C1(n20776), .C2(n20711), .A(n20671), .B(n20670), .ZN(
        P1_U3144) );
  NOR2_X1 U23642 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20716), .ZN(
        n20706) );
  NAND3_X1 U23643 ( .A1(n20714), .A2(n20678), .A3(n20846), .ZN(n20672) );
  OAI21_X1 U23644 ( .B1(n20674), .B2(n20673), .A(n20672), .ZN(n20705) );
  AOI22_X1 U23645 ( .A1(n20718), .A2(n20706), .B1(n20717), .B2(n20705), .ZN(
        n20684) );
  AOI21_X1 U23646 ( .B1(n20711), .B2(n20764), .A(n20847), .ZN(n20677) );
  AOI21_X1 U23647 ( .B1(n20714), .B2(n20678), .A(n20677), .ZN(n20679) );
  NOR2_X1 U23648 ( .A1(n20679), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20682) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20708), .B1(
        n20771), .B2(n20724), .ZN(n20683) );
  OAI211_X1 U23650 ( .C1(n20727), .C2(n20711), .A(n20684), .B(n20683), .ZN(
        P1_U3145) );
  AOI22_X1 U23651 ( .A1(n20729), .A2(n20706), .B1(n20705), .B2(n20728), .ZN(
        n20687) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20708), .B1(
        n20771), .B2(n20685), .ZN(n20686) );
  OAI211_X1 U23653 ( .C1(n20688), .C2(n20711), .A(n20687), .B(n20686), .ZN(
        P1_U3146) );
  AOI22_X1 U23654 ( .A1(n20735), .A2(n20706), .B1(n20705), .B2(n20734), .ZN(
        n20691) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20708), .B1(
        n20771), .B2(n20689), .ZN(n20690) );
  OAI211_X1 U23656 ( .C1(n20692), .C2(n20711), .A(n20691), .B(n20690), .ZN(
        P1_U3147) );
  AOI22_X1 U23657 ( .A1(n20741), .A2(n20706), .B1(n20705), .B2(n20740), .ZN(
        n20695) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20708), .B1(
        n20771), .B2(n20693), .ZN(n20694) );
  OAI211_X1 U23659 ( .C1(n20696), .C2(n20711), .A(n20695), .B(n20694), .ZN(
        P1_U3148) );
  AOI22_X1 U23660 ( .A1(n20747), .A2(n20706), .B1(n20705), .B2(n20746), .ZN(
        n20698) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20708), .B1(
        n20771), .B2(n20748), .ZN(n20697) );
  OAI211_X1 U23662 ( .C1(n20751), .C2(n20711), .A(n20698), .B(n20697), .ZN(
        P1_U3149) );
  AOI22_X1 U23663 ( .A1(n9795), .A2(n20706), .B1(n20705), .B2(n20752), .ZN(
        n20701) );
  AOI22_X1 U23664 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20708), .B1(
        n20771), .B2(n20699), .ZN(n20700) );
  OAI211_X1 U23665 ( .C1(n20702), .C2(n20711), .A(n20701), .B(n20700), .ZN(
        P1_U3150) );
  AOI22_X1 U23666 ( .A1(n20759), .A2(n20706), .B1(n20705), .B2(n20758), .ZN(
        n20704) );
  AOI22_X1 U23667 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20708), .B1(
        n20771), .B2(n20760), .ZN(n20703) );
  OAI211_X1 U23668 ( .C1(n20765), .C2(n20711), .A(n20704), .B(n20703), .ZN(
        P1_U3151) );
  AOI22_X1 U23669 ( .A1(n20769), .A2(n20706), .B1(n20705), .B2(n20767), .ZN(
        n20710) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20708), .B1(
        n20771), .B2(n20707), .ZN(n20709) );
  OAI211_X1 U23671 ( .C1(n20712), .C2(n20711), .A(n20710), .B(n20709), .ZN(
        P1_U3152) );
  AOI21_X1 U23672 ( .B1(n20714), .B2(n20713), .A(n20768), .ZN(n20719) );
  OAI22_X1 U23673 ( .A1(n20719), .A2(n20859), .B1(n20716), .B2(n20715), .ZN(
        n20766) );
  AOI22_X1 U23674 ( .A1(n20718), .A2(n20768), .B1(n20717), .B2(n20766), .ZN(
        n20726) );
  OAI21_X1 U23675 ( .B1(n20851), .B2(n20720), .A(n20719), .ZN(n20721) );
  OAI211_X1 U23676 ( .C1(n20723), .C2(n20846), .A(n20722), .B(n20721), .ZN(
        n20772) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20772), .B1(
        n20761), .B2(n20724), .ZN(n20725) );
  OAI211_X1 U23678 ( .C1(n20727), .C2(n20764), .A(n20726), .B(n20725), .ZN(
        P1_U3153) );
  AOI22_X1 U23679 ( .A1(n20729), .A2(n20768), .B1(n20728), .B2(n20766), .ZN(
        n20732) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20772), .B1(
        n20771), .B2(n20730), .ZN(n20731) );
  OAI211_X1 U23681 ( .C1(n20733), .C2(n20775), .A(n20732), .B(n20731), .ZN(
        P1_U3154) );
  AOI22_X1 U23682 ( .A1(n20735), .A2(n20768), .B1(n20734), .B2(n20766), .ZN(
        n20738) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20772), .B1(
        n20771), .B2(n20736), .ZN(n20737) );
  OAI211_X1 U23684 ( .C1(n20739), .C2(n20775), .A(n20738), .B(n20737), .ZN(
        P1_U3155) );
  AOI22_X1 U23685 ( .A1(n20741), .A2(n20768), .B1(n20740), .B2(n20766), .ZN(
        n20744) );
  AOI22_X1 U23686 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20772), .B1(
        n20771), .B2(n20742), .ZN(n20743) );
  OAI211_X1 U23687 ( .C1(n20745), .C2(n20775), .A(n20744), .B(n20743), .ZN(
        P1_U3156) );
  AOI22_X1 U23688 ( .A1(n20747), .A2(n20768), .B1(n20746), .B2(n20766), .ZN(
        n20750) );
  AOI22_X1 U23689 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20772), .B1(
        n20761), .B2(n20748), .ZN(n20749) );
  OAI211_X1 U23690 ( .C1(n20751), .C2(n20764), .A(n20750), .B(n20749), .ZN(
        P1_U3157) );
  AOI22_X1 U23691 ( .A1(n9795), .A2(n20768), .B1(n20752), .B2(n20766), .ZN(
        n20756) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20772), .B1(
        n20771), .B2(n20754), .ZN(n20755) );
  OAI211_X1 U23693 ( .C1(n20757), .C2(n20775), .A(n20756), .B(n20755), .ZN(
        P1_U3158) );
  AOI22_X1 U23694 ( .A1(n20759), .A2(n20768), .B1(n20758), .B2(n20766), .ZN(
        n20763) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20772), .B1(
        n20761), .B2(n20760), .ZN(n20762) );
  OAI211_X1 U23696 ( .C1(n20765), .C2(n20764), .A(n20763), .B(n20762), .ZN(
        P1_U3159) );
  AOI22_X1 U23697 ( .A1(n20769), .A2(n20768), .B1(n20767), .B2(n20766), .ZN(
        n20774) );
  AOI22_X1 U23698 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20772), .B1(
        n20771), .B2(n20770), .ZN(n20773) );
  OAI211_X1 U23699 ( .C1(n20776), .C2(n20775), .A(n20774), .B(n20773), .ZN(
        P1_U3160) );
  NAND3_X1 U23700 ( .A1(n20779), .A2(n20778), .A3(n20777), .ZN(P1_U3163) );
  AND2_X1 U23701 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20780), .ZN(
        P1_U3164) );
  AND2_X1 U23702 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20780), .ZN(
        P1_U3165) );
  AND2_X1 U23703 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20780), .ZN(
        P1_U3166) );
  AND2_X1 U23704 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20780), .ZN(
        P1_U3167) );
  AND2_X1 U23705 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20780), .ZN(
        P1_U3168) );
  INV_X1 U23706 ( .A(P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n21099) );
  NOR2_X1 U23707 ( .A1(n20844), .A2(n21099), .ZN(P1_U3169) );
  AND2_X1 U23708 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20780), .ZN(
        P1_U3170) );
  AND2_X1 U23709 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20780), .ZN(
        P1_U3171) );
  AND2_X1 U23710 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20780), .ZN(
        P1_U3172) );
  AND2_X1 U23711 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20780), .ZN(
        P1_U3173) );
  AND2_X1 U23712 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20780), .ZN(
        P1_U3174) );
  AND2_X1 U23713 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20780), .ZN(
        P1_U3175) );
  AND2_X1 U23714 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20780), .ZN(
        P1_U3176) );
  AND2_X1 U23715 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20780), .ZN(
        P1_U3177) );
  AND2_X1 U23716 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20780), .ZN(
        P1_U3178) );
  AND2_X1 U23717 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20780), .ZN(
        P1_U3179) );
  AND2_X1 U23718 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20780), .ZN(
        P1_U3180) );
  AND2_X1 U23719 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20780), .ZN(
        P1_U3181) );
  AND2_X1 U23720 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20780), .ZN(
        P1_U3182) );
  AND2_X1 U23721 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20780), .ZN(
        P1_U3183) );
  AND2_X1 U23722 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20780), .ZN(
        P1_U3184) );
  AND2_X1 U23723 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20780), .ZN(
        P1_U3185) );
  AND2_X1 U23724 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20780), .ZN(P1_U3186) );
  AND2_X1 U23725 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20780), .ZN(P1_U3187) );
  AND2_X1 U23726 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20780), .ZN(P1_U3188) );
  AND2_X1 U23727 ( .A1(n20780), .A2(P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(P1_U3189) );
  AND2_X1 U23728 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20780), .ZN(P1_U3190) );
  AND2_X1 U23729 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20780), .ZN(P1_U3191) );
  INV_X1 U23730 ( .A(P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21101) );
  NOR2_X1 U23731 ( .A1(n20844), .A2(n21101), .ZN(P1_U3192) );
  AND2_X1 U23732 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20780), .ZN(P1_U3193) );
  AOI21_X1 U23733 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20781), .A(n21063), 
        .ZN(n20794) );
  NOR2_X1 U23734 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20783) );
  OAI22_X1 U23735 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20786), .B1(n20783), 
        .B2(n20782), .ZN(n20784) );
  NOR2_X1 U23736 ( .A1(n20790), .A2(n20784), .ZN(n20785) );
  OAI22_X1 U23737 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20794), .B1(n20873), 
        .B2(n20785), .ZN(P1_U3194) );
  OAI21_X1 U23738 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20787), .A(n20786), 
        .ZN(n20792) );
  AOI221_X1 U23739 ( .B1(NA), .B2(n20788), .C1(n20880), .C2(n20788), .A(n21063), .ZN(n20789) );
  OAI211_X1 U23740 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20790), .A(HOLD), .B(
        n20789), .ZN(n20791) );
  OAI221_X1 U23741 ( .B1(n20794), .B2(n20793), .C1(n20794), .C2(n20792), .A(
        n20791), .ZN(P1_U3196) );
  INV_X1 U23742 ( .A(n20830), .ZN(n20836) );
  NOR2_X2 U23743 ( .A1(n20795), .A2(n20884), .ZN(n20834) );
  OAI222_X1 U23744 ( .A1(n20836), .A2(n20083), .B1(n20797), .B2(n20873), .C1(
        n20796), .C2(n20832), .ZN(P1_U3197) );
  AOI222_X1 U23745 ( .A1(n20834), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20830), .ZN(n20798) );
  INV_X1 U23746 ( .A(n20798), .ZN(P1_U3198) );
  AOI22_X1 U23747 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(n20884), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(n20830), .ZN(n20799) );
  OAI21_X1 U23748 ( .B1(n13687), .B2(n20832), .A(n20799), .ZN(P1_U3199) );
  AOI222_X1 U23749 ( .A1(n20830), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20834), .ZN(n20800) );
  INV_X1 U23750 ( .A(n20800), .ZN(P1_U3200) );
  AOI222_X1 U23751 ( .A1(n20834), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20830), .ZN(n20801) );
  INV_X1 U23752 ( .A(n20801), .ZN(P1_U3201) );
  AOI222_X1 U23753 ( .A1(n20830), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20834), .ZN(n20802) );
  INV_X1 U23754 ( .A(n20802), .ZN(P1_U3202) );
  AOI22_X1 U23755 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20884), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20830), .ZN(n20803) );
  OAI21_X1 U23756 ( .B1(n20804), .B2(n20832), .A(n20803), .ZN(P1_U3203) );
  AOI22_X1 U23757 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20884), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20834), .ZN(n20805) );
  OAI21_X1 U23758 ( .B1(n20806), .B2(n20836), .A(n20805), .ZN(P1_U3204) );
  AOI222_X1 U23759 ( .A1(n20834), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20830), .ZN(n20807) );
  INV_X1 U23760 ( .A(n20807), .ZN(P1_U3205) );
  AOI222_X1 U23761 ( .A1(n20830), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20834), .ZN(n20808) );
  INV_X1 U23762 ( .A(n20808), .ZN(P1_U3206) );
  AOI222_X1 U23763 ( .A1(n20834), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20830), .ZN(n20809) );
  INV_X1 U23764 ( .A(n20809), .ZN(P1_U3207) );
  AOI222_X1 U23765 ( .A1(n20834), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20830), .ZN(n20810) );
  INV_X1 U23766 ( .A(n20810), .ZN(P1_U3208) );
  AOI222_X1 U23767 ( .A1(n20834), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20830), .ZN(n20811) );
  INV_X1 U23768 ( .A(n20811), .ZN(P1_U3209) );
  AOI222_X1 U23769 ( .A1(n20830), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20834), .ZN(n20812) );
  INV_X1 U23770 ( .A(n20812), .ZN(P1_U3210) );
  INV_X1 U23771 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21165) );
  OAI222_X1 U23772 ( .A1(n20832), .A2(n20813), .B1(n21165), .B2(n20873), .C1(
        n14993), .C2(n20836), .ZN(P1_U3211) );
  AOI22_X1 U23773 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20884), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20830), .ZN(n20814) );
  OAI21_X1 U23774 ( .B1(n14993), .B2(n20832), .A(n20814), .ZN(P1_U3212) );
  AOI222_X1 U23775 ( .A1(n20834), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20830), .ZN(n20815) );
  INV_X1 U23776 ( .A(n20815), .ZN(P1_U3213) );
  AOI222_X1 U23777 ( .A1(n20834), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20830), .ZN(n20816) );
  INV_X1 U23778 ( .A(n20816), .ZN(P1_U3214) );
  AOI222_X1 U23779 ( .A1(n20834), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20830), .ZN(n20817) );
  INV_X1 U23780 ( .A(n20817), .ZN(P1_U3215) );
  AOI22_X1 U23781 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20884), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n20830), .ZN(n20818) );
  OAI21_X1 U23782 ( .B1(n14979), .B2(n20832), .A(n20818), .ZN(P1_U3216) );
  AOI22_X1 U23783 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20884), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20830), .ZN(n20819) );
  OAI21_X1 U23784 ( .B1(n14792), .B2(n20832), .A(n20819), .ZN(P1_U3217) );
  AOI22_X1 U23785 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20884), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20830), .ZN(n20820) );
  OAI21_X1 U23786 ( .B1(n14788), .B2(n20832), .A(n20820), .ZN(P1_U3218) );
  AOI22_X1 U23787 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20884), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20834), .ZN(n20821) );
  OAI21_X1 U23788 ( .B1(n20822), .B2(n20836), .A(n20821), .ZN(P1_U3219) );
  AOI222_X1 U23789 ( .A1(n20834), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20884), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20830), .ZN(n20823) );
  INV_X1 U23790 ( .A(n20823), .ZN(P1_U3220) );
  INV_X1 U23791 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20824) );
  OAI222_X1 U23792 ( .A1(n20832), .A2(n20825), .B1(n20824), .B2(n20873), .C1(
        n14755), .C2(n20836), .ZN(P1_U3221) );
  INV_X1 U23793 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20826) );
  OAI222_X1 U23794 ( .A1(n20832), .A2(n14755), .B1(n20826), .B2(n20873), .C1(
        n20828), .C2(n20836), .ZN(P1_U3222) );
  AOI22_X1 U23795 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20830), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20884), .ZN(n20827) );
  OAI21_X1 U23796 ( .B1(n20828), .B2(n20832), .A(n20827), .ZN(P1_U3223) );
  AOI22_X1 U23797 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20834), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20884), .ZN(n20829) );
  OAI21_X1 U23798 ( .B1(n20833), .B2(n20836), .A(n20829), .ZN(P1_U3224) );
  AOI22_X1 U23799 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20830), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20884), .ZN(n20831) );
  OAI21_X1 U23800 ( .B1(n20833), .B2(n20832), .A(n20831), .ZN(P1_U3225) );
  AOI22_X1 U23801 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20834), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20884), .ZN(n20835) );
  OAI21_X1 U23802 ( .B1(n20837), .B2(n20836), .A(n20835), .ZN(P1_U3226) );
  OAI22_X1 U23803 ( .A1(n20884), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20873), .ZN(n20838) );
  INV_X1 U23804 ( .A(n20838), .ZN(P1_U3458) );
  OAI22_X1 U23805 ( .A1(n20884), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20873), .ZN(n20839) );
  INV_X1 U23806 ( .A(n20839), .ZN(P1_U3459) );
  OAI22_X1 U23807 ( .A1(n20884), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20873), .ZN(n20840) );
  INV_X1 U23808 ( .A(n20840), .ZN(P1_U3460) );
  OAI22_X1 U23809 ( .A1(n20884), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20873), .ZN(n20841) );
  INV_X1 U23810 ( .A(n20841), .ZN(P1_U3461) );
  OAI21_X1 U23811 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20844), .A(n20843), 
        .ZN(n20842) );
  INV_X1 U23812 ( .A(n20842), .ZN(P1_U3464) );
  OAI21_X1 U23813 ( .B1(n20844), .B2(n21065), .A(n20843), .ZN(P1_U3465) );
  INV_X1 U23814 ( .A(n20864), .ZN(n20856) );
  OAI211_X1 U23815 ( .C1(n20848), .C2(n20847), .A(n11914), .B(n20846), .ZN(
        n20849) );
  OAI21_X1 U23816 ( .B1(n20850), .B2(n20858), .A(n20849), .ZN(n20852) );
  AOI211_X1 U23817 ( .C1(n20854), .C2(n20853), .A(n20852), .B(n20851), .ZN(
        n20855) );
  AOI22_X1 U23818 ( .A1(n20856), .A2(n20574), .B1(n20855), .B2(n20864), .ZN(
        P1_U3475) );
  OAI22_X1 U23819 ( .A1(n12694), .A2(n20859), .B1(n20858), .B2(n20857), .ZN(
        n20860) );
  OAI21_X1 U23820 ( .B1(n20861), .B2(n20860), .A(n20864), .ZN(n20862) );
  OAI21_X1 U23821 ( .B1(n20864), .B2(n20863), .A(n20862), .ZN(P1_U3478) );
  AOI211_X1 U23822 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20865) );
  AOI21_X1 U23823 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20865), .ZN(n20867) );
  INV_X1 U23824 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20866) );
  AOI22_X1 U23825 ( .A1(n20871), .A2(n20867), .B1(n20866), .B2(n20868), .ZN(
        P1_U3481) );
  NOR2_X1 U23826 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20870) );
  INV_X1 U23827 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20869) );
  AOI22_X1 U23828 ( .A1(n20871), .A2(n20870), .B1(n20869), .B2(n20868), .ZN(
        P1_U3482) );
  INV_X1 U23829 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20872) );
  AOI22_X1 U23830 ( .A1(n20873), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20872), 
        .B2(n20884), .ZN(P1_U3483) );
  OAI21_X1 U23831 ( .B1(n20874), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20876) );
  OAI21_X1 U23832 ( .B1(n20877), .B2(n20876), .A(n20875), .ZN(n20883) );
  AOI211_X1 U23833 ( .C1(n20121), .C2(n20880), .A(n20879), .B(n20878), .ZN(
        n20882) );
  NAND2_X1 U23834 ( .A1(n20882), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20881) );
  OAI21_X1 U23835 ( .B1(n20883), .B2(n20882), .A(n20881), .ZN(P1_U3485) );
  MUX2_X1 U23836 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20884), .Z(P1_U3486) );
  AOI222_X1 U23837 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n20887), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n20886), .C1(P1_DATAO_REG_1__SCAN_IN), 
        .C2(n20885), .ZN(n21270) );
  AOI22_X1 U23838 ( .A1(P3_UWORD_REG_7__SCAN_IN), .A2(keyinput191), .B1(
        P3_INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput146), .ZN(n20888) );
  OAI221_X1 U23839 ( .B1(P3_UWORD_REG_7__SCAN_IN), .B2(keyinput191), .C1(
        P3_INSTQUEUE_REG_2__3__SCAN_IN), .C2(keyinput146), .A(n20888), .ZN(
        n20895) );
  AOI22_X1 U23840 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(keyinput195), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(keyinput254), .ZN(n20889) );
  OAI221_X1 U23841 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(keyinput195), .C1(
        P1_EBX_REG_20__SCAN_IN), .C2(keyinput254), .A(n20889), .ZN(n20894) );
  AOI22_X1 U23842 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(keyinput242), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(keyinput228), .ZN(n20890) );
  OAI221_X1 U23843 ( .B1(P1_DATAO_REG_6__SCAN_IN), .B2(keyinput242), .C1(
        P1_DATAO_REG_12__SCAN_IN), .C2(keyinput228), .A(n20890), .ZN(n20893)
         );
  AOI22_X1 U23844 ( .A1(P1_EAX_REG_4__SCAN_IN), .A2(keyinput130), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(keyinput240), .ZN(n20891) );
  OAI221_X1 U23845 ( .B1(P1_EAX_REG_4__SCAN_IN), .B2(keyinput130), .C1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .C2(keyinput240), .A(n20891), .ZN(
        n20892) );
  NOR4_X1 U23846 ( .A1(n20895), .A2(n20894), .A3(n20893), .A4(n20892), .ZN(
        n20923) );
  AOI22_X1 U23847 ( .A1(P1_EAX_REG_29__SCAN_IN), .A2(keyinput132), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput154), .ZN(n20896) );
  OAI221_X1 U23848 ( .B1(P1_EAX_REG_29__SCAN_IN), .B2(keyinput132), .C1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(keyinput154), .A(n20896), 
        .ZN(n20903) );
  AOI22_X1 U23849 ( .A1(P3_ADDRESS_REG_2__SCAN_IN), .A2(keyinput139), .B1(
        BUF2_REG_10__SCAN_IN), .B2(keyinput131), .ZN(n20897) );
  OAI221_X1 U23850 ( .B1(P3_ADDRESS_REG_2__SCAN_IN), .B2(keyinput139), .C1(
        BUF2_REG_10__SCAN_IN), .C2(keyinput131), .A(n20897), .ZN(n20902) );
  AOI22_X1 U23851 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(keyinput201), .B1(
        P3_INSTQUEUE_REG_7__2__SCAN_IN), .B2(keyinput251), .ZN(n20898) );
  OAI221_X1 U23852 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(keyinput201), .C1(
        P3_INSTQUEUE_REG_7__2__SCAN_IN), .C2(keyinput251), .A(n20898), .ZN(
        n20901) );
  AOI22_X1 U23853 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput197), 
        .B1(P2_EAX_REG_17__SCAN_IN), .B2(keyinput214), .ZN(n20899) );
  OAI221_X1 U23854 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput197), 
        .C1(P2_EAX_REG_17__SCAN_IN), .C2(keyinput214), .A(n20899), .ZN(n20900)
         );
  NOR4_X1 U23855 ( .A1(n20903), .A2(n20902), .A3(n20901), .A4(n20900), .ZN(
        n20922) );
  AOI22_X1 U23856 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(keyinput150), 
        .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput180), .ZN(n20904) );
  OAI221_X1 U23857 ( .B1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B2(keyinput150), 
        .C1(P1_EBX_REG_27__SCAN_IN), .C2(keyinput180), .A(n20904), .ZN(n20911)
         );
  AOI22_X1 U23858 ( .A1(P2_LWORD_REG_14__SCAN_IN), .A2(keyinput238), .B1(
        BUF1_REG_8__SCAN_IN), .B2(keyinput216), .ZN(n20905) );
  OAI221_X1 U23859 ( .B1(P2_LWORD_REG_14__SCAN_IN), .B2(keyinput238), .C1(
        BUF1_REG_8__SCAN_IN), .C2(keyinput216), .A(n20905), .ZN(n20910) );
  AOI22_X1 U23860 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput215), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(keyinput179), .ZN(n20906) );
  OAI221_X1 U23861 ( .B1(P3_DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput215), .C1(
        P1_EBX_REG_31__SCAN_IN), .C2(keyinput179), .A(n20906), .ZN(n20909) );
  AOI22_X1 U23862 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(keyinput156), 
        .B1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput217), .ZN(n20907) );
  OAI221_X1 U23863 ( .B1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B2(keyinput156), 
        .C1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .C2(keyinput217), .A(n20907), 
        .ZN(n20908) );
  NOR4_X1 U23864 ( .A1(n20911), .A2(n20910), .A3(n20909), .A4(n20908), .ZN(
        n20921) );
  AOI22_X1 U23865 ( .A1(BUF1_REG_18__SCAN_IN), .A2(keyinput223), .B1(
        P3_INSTQUEUE_REG_6__3__SCAN_IN), .B2(keyinput160), .ZN(n20912) );
  OAI221_X1 U23866 ( .B1(BUF1_REG_18__SCAN_IN), .B2(keyinput223), .C1(
        P3_INSTQUEUE_REG_6__3__SCAN_IN), .C2(keyinput160), .A(n20912), .ZN(
        n20919) );
  AOI22_X1 U23867 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(keyinput213), 
        .B1(P2_EAX_REG_9__SCAN_IN), .B2(keyinput248), .ZN(n20913) );
  OAI221_X1 U23868 ( .B1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B2(keyinput213), 
        .C1(P2_EAX_REG_9__SCAN_IN), .C2(keyinput248), .A(n20913), .ZN(n20918)
         );
  AOI22_X1 U23869 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(keyinput135), 
        .B1(P1_ADDRESS_REG_16__SCAN_IN), .B2(keyinput211), .ZN(n20914) );
  OAI221_X1 U23870 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput135), 
        .C1(P1_ADDRESS_REG_16__SCAN_IN), .C2(keyinput211), .A(n20914), .ZN(
        n20917) );
  AOI22_X1 U23871 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(keyinput237), 
        .B1(P2_EBX_REG_13__SCAN_IN), .B2(keyinput246), .ZN(n20915) );
  OAI221_X1 U23872 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput237), 
        .C1(P2_EBX_REG_13__SCAN_IN), .C2(keyinput246), .A(n20915), .ZN(n20916)
         );
  NOR4_X1 U23873 ( .A1(n20919), .A2(n20918), .A3(n20917), .A4(n20916), .ZN(
        n20920) );
  NAND4_X1 U23874 ( .A1(n20923), .A2(n20922), .A3(n20921), .A4(n20920), .ZN(
        n21060) );
  AOI22_X1 U23875 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(keyinput202), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput142), .ZN(n20924) );
  OAI221_X1 U23876 ( .B1(P1_DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput202), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput142), .A(n20924), .ZN(n20931) );
  AOI22_X1 U23877 ( .A1(P2_W_R_N_REG_SCAN_IN), .A2(keyinput143), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(keyinput144), .ZN(n20925) );
  OAI221_X1 U23878 ( .B1(P2_W_R_N_REG_SCAN_IN), .B2(keyinput143), .C1(
        P1_EAX_REG_27__SCAN_IN), .C2(keyinput144), .A(n20925), .ZN(n20930) );
  AOI22_X1 U23879 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(keyinput207), .B1(
        BUF1_REG_7__SCAN_IN), .B2(keyinput159), .ZN(n20926) );
  OAI221_X1 U23880 ( .B1(P1_DATAO_REG_25__SCAN_IN), .B2(keyinput207), .C1(
        BUF1_REG_7__SCAN_IN), .C2(keyinput159), .A(n20926), .ZN(n20929) );
  AOI22_X1 U23881 ( .A1(P1_EBX_REG_23__SCAN_IN), .A2(keyinput134), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(keyinput148), .ZN(n20927) );
  OAI221_X1 U23882 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(keyinput134), .C1(
        P1_STATE_REG_0__SCAN_IN), .C2(keyinput148), .A(n20927), .ZN(n20928) );
  NOR4_X1 U23883 ( .A1(n20931), .A2(n20930), .A3(n20929), .A4(n20928), .ZN(
        n20959) );
  AOI22_X1 U23884 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(keyinput232), .B1(
        P1_INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput226), .ZN(n20932) );
  OAI221_X1 U23885 ( .B1(P1_ADDRESS_REG_3__SCAN_IN), .B2(keyinput232), .C1(
        P1_INSTQUEUE_REG_9__3__SCAN_IN), .C2(keyinput226), .A(n20932), .ZN(
        n20939) );
  AOI22_X1 U23886 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(keyinput178), .B1(
        P2_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput162), .ZN(n20933) );
  OAI221_X1 U23887 ( .B1(P3_DATAWIDTH_REG_29__SCAN_IN), .B2(keyinput178), .C1(
        P2_INSTQUEUE_REG_7__5__SCAN_IN), .C2(keyinput162), .A(n20933), .ZN(
        n20938) );
  AOI22_X1 U23888 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(keyinput147), .B1(
        P2_ADDRESS_REG_15__SCAN_IN), .B2(keyinput129), .ZN(n20934) );
  OAI221_X1 U23889 ( .B1(P2_LWORD_REG_11__SCAN_IN), .B2(keyinput147), .C1(
        P2_ADDRESS_REG_15__SCAN_IN), .C2(keyinput129), .A(n20934), .ZN(n20937)
         );
  AOI22_X1 U23890 ( .A1(P3_BE_N_REG_0__SCAN_IN), .A2(keyinput177), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(keyinput170), .ZN(n20935) );
  OAI221_X1 U23891 ( .B1(P3_BE_N_REG_0__SCAN_IN), .B2(keyinput177), .C1(
        P2_EBX_REG_18__SCAN_IN), .C2(keyinput170), .A(n20935), .ZN(n20936) );
  NOR4_X1 U23892 ( .A1(n20939), .A2(n20938), .A3(n20937), .A4(n20936), .ZN(
        n20958) );
  AOI22_X1 U23893 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(keyinput190), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(keyinput167), .ZN(n20940) );
  OAI221_X1 U23894 ( .B1(P2_DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput190), .C1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .C2(keyinput167), .A(n20940), .ZN(
        n20947) );
  AOI22_X1 U23895 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(keyinput136), 
        .B1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput173), .ZN(n20941) );
  OAI221_X1 U23896 ( .B1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B2(keyinput136), 
        .C1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .C2(keyinput173), .A(n20941), 
        .ZN(n20946) );
  AOI22_X1 U23897 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput239), .B1(
        BUF1_REG_4__SCAN_IN), .B2(keyinput221), .ZN(n20942) );
  OAI221_X1 U23898 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput239), .C1(
        BUF1_REG_4__SCAN_IN), .C2(keyinput221), .A(n20942), .ZN(n20945) );
  AOI22_X1 U23899 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(keyinput250), 
        .B1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B2(keyinput185), .ZN(n20943) );
  OAI221_X1 U23900 ( .B1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(keyinput250), 
        .C1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .C2(keyinput185), .A(n20943), 
        .ZN(n20944) );
  NOR4_X1 U23901 ( .A1(n20947), .A2(n20946), .A3(n20945), .A4(n20944), .ZN(
        n20957) );
  AOI22_X1 U23902 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(keyinput193), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput229), .ZN(n20948) );
  OAI221_X1 U23903 ( .B1(P2_ADDRESS_REG_24__SCAN_IN), .B2(keyinput193), .C1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput229), .A(n20948), .ZN(
        n20955) );
  AOI22_X1 U23904 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput244), 
        .B1(P2_REIP_REG_0__SCAN_IN), .B2(keyinput176), .ZN(n20949) );
  OAI221_X1 U23905 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput244), 
        .C1(P2_REIP_REG_0__SCAN_IN), .C2(keyinput176), .A(n20949), .ZN(n20954)
         );
  AOI22_X1 U23906 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(keyinput233), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(keyinput212), .ZN(n20950) );
  OAI221_X1 U23907 ( .B1(P1_DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput233), .C1(
        P2_M_IO_N_REG_SCAN_IN), .C2(keyinput212), .A(n20950), .ZN(n20953) );
  AOI22_X1 U23908 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(keyinput155), .B1(
        P2_ADDRESS_REG_7__SCAN_IN), .B2(keyinput153), .ZN(n20951) );
  OAI221_X1 U23909 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(keyinput155), .C1(
        P2_ADDRESS_REG_7__SCAN_IN), .C2(keyinput153), .A(n20951), .ZN(n20952)
         );
  NOR4_X1 U23910 ( .A1(n20955), .A2(n20954), .A3(n20953), .A4(n20952), .ZN(
        n20956) );
  NAND4_X1 U23911 ( .A1(n20959), .A2(n20958), .A3(n20957), .A4(n20956), .ZN(
        n21059) );
  INV_X1 U23912 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n20961) );
  AOI22_X1 U23913 ( .A1(n20961), .A2(keyinput140), .B1(keyinput200), .B2(
        n21065), .ZN(n20960) );
  OAI221_X1 U23914 ( .B1(n20961), .B2(keyinput140), .C1(n21065), .C2(
        keyinput200), .A(n20960), .ZN(n20972) );
  AOI22_X1 U23915 ( .A1(n21111), .A2(keyinput219), .B1(keyinput253), .B2(
        n20963), .ZN(n20962) );
  OAI221_X1 U23916 ( .B1(n21111), .B2(keyinput219), .C1(n20963), .C2(
        keyinput253), .A(n20962), .ZN(n20971) );
  INV_X1 U23917 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n20966) );
  AOI22_X1 U23918 ( .A1(n20966), .A2(keyinput206), .B1(n20965), .B2(
        keyinput203), .ZN(n20964) );
  OAI221_X1 U23919 ( .B1(n20966), .B2(keyinput206), .C1(n20965), .C2(
        keyinput203), .A(n20964), .ZN(n20970) );
  XNOR2_X1 U23920 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B(keyinput243), .ZN(
        n20968) );
  XNOR2_X1 U23921 ( .A(keyinput245), .B(P1_EBX_REG_11__SCAN_IN), .ZN(n20967)
         );
  NAND2_X1 U23922 ( .A1(n20968), .A2(n20967), .ZN(n20969) );
  NOR4_X1 U23923 ( .A1(n20972), .A2(n20971), .A3(n20970), .A4(n20969), .ZN(
        n21011) );
  AOI22_X1 U23924 ( .A1(n20974), .A2(keyinput149), .B1(n21115), .B2(
        keyinput174), .ZN(n20973) );
  OAI221_X1 U23925 ( .B1(n20974), .B2(keyinput149), .C1(n21115), .C2(
        keyinput174), .A(n20973), .ZN(n20985) );
  AOI22_X1 U23926 ( .A1(n20977), .A2(keyinput188), .B1(keyinput141), .B2(
        n20976), .ZN(n20975) );
  OAI221_X1 U23927 ( .B1(n20977), .B2(keyinput188), .C1(n20976), .C2(
        keyinput141), .A(n20975), .ZN(n20984) );
  AOI22_X1 U23928 ( .A1(n20979), .A2(keyinput145), .B1(n14638), .B2(
        keyinput198), .ZN(n20978) );
  OAI221_X1 U23929 ( .B1(n20979), .B2(keyinput145), .C1(n14638), .C2(
        keyinput198), .A(n20978), .ZN(n20983) );
  AOI22_X1 U23930 ( .A1(n20981), .A2(keyinput220), .B1(n21132), .B2(
        keyinput218), .ZN(n20980) );
  OAI221_X1 U23931 ( .B1(n20981), .B2(keyinput220), .C1(n21132), .C2(
        keyinput218), .A(n20980), .ZN(n20982) );
  NOR4_X1 U23932 ( .A1(n20985), .A2(n20984), .A3(n20983), .A4(n20982), .ZN(
        n21010) );
  AOI22_X1 U23933 ( .A1(n21086), .A2(keyinput247), .B1(n14269), .B2(
        keyinput175), .ZN(n20986) );
  OAI221_X1 U23934 ( .B1(n21086), .B2(keyinput247), .C1(n14269), .C2(
        keyinput175), .A(n20986), .ZN(n20996) );
  INV_X1 U23935 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n20988) );
  AOI22_X1 U23936 ( .A1(n20988), .A2(keyinput169), .B1(n10847), .B2(
        keyinput186), .ZN(n20987) );
  OAI221_X1 U23937 ( .B1(n20988), .B2(keyinput169), .C1(n10847), .C2(
        keyinput186), .A(n20987), .ZN(n20995) );
  AOI22_X1 U23938 ( .A1(n21095), .A2(keyinput137), .B1(n21130), .B2(
        keyinput204), .ZN(n20989) );
  OAI221_X1 U23939 ( .B1(n21095), .B2(keyinput137), .C1(n21130), .C2(
        keyinput204), .A(n20989), .ZN(n20994) );
  AOI22_X1 U23940 ( .A1(n20992), .A2(keyinput182), .B1(n20991), .B2(
        keyinput164), .ZN(n20990) );
  OAI221_X1 U23941 ( .B1(n20992), .B2(keyinput182), .C1(n20991), .C2(
        keyinput164), .A(n20990), .ZN(n20993) );
  NOR4_X1 U23942 ( .A1(n20996), .A2(n20995), .A3(n20994), .A4(n20993), .ZN(
        n21009) );
  INV_X1 U23943 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n20998) );
  AOI22_X1 U23944 ( .A1(n20998), .A2(keyinput158), .B1(n21165), .B2(
        keyinput165), .ZN(n20997) );
  OAI221_X1 U23945 ( .B1(n20998), .B2(keyinput158), .C1(n21165), .C2(
        keyinput165), .A(n20997), .ZN(n21007) );
  AOI22_X1 U23946 ( .A1(n21000), .A2(keyinput151), .B1(n10485), .B2(
        keyinput225), .ZN(n20999) );
  OAI221_X1 U23947 ( .B1(n21000), .B2(keyinput151), .C1(n10485), .C2(
        keyinput225), .A(n20999), .ZN(n21006) );
  INV_X1 U23948 ( .A(DATAI_26_), .ZN(n21180) );
  AOI22_X1 U23949 ( .A1(n21180), .A2(keyinput249), .B1(keyinput230), .B2(
        n21101), .ZN(n21001) );
  OAI221_X1 U23950 ( .B1(n21180), .B2(keyinput249), .C1(n21101), .C2(
        keyinput230), .A(n21001), .ZN(n21005) );
  AOI22_X1 U23951 ( .A1(n21003), .A2(keyinput133), .B1(n21177), .B2(
        keyinput241), .ZN(n21002) );
  OAI221_X1 U23952 ( .B1(n21003), .B2(keyinput133), .C1(n21177), .C2(
        keyinput241), .A(n21002), .ZN(n21004) );
  NOR4_X1 U23953 ( .A1(n21007), .A2(n21006), .A3(n21005), .A4(n21004), .ZN(
        n21008) );
  NAND4_X1 U23954 ( .A1(n21011), .A2(n21010), .A3(n21009), .A4(n21008), .ZN(
        n21058) );
  INV_X1 U23955 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21068) );
  AOI22_X1 U23956 ( .A1(n10497), .A2(keyinput192), .B1(keyinput231), .B2(
        n21068), .ZN(n21012) );
  OAI221_X1 U23957 ( .B1(n10497), .B2(keyinput192), .C1(n21068), .C2(
        keyinput231), .A(n21012), .ZN(n21020) );
  AOI22_X1 U23958 ( .A1(n15189), .A2(keyinput209), .B1(keyinput152), .B2(
        n21014), .ZN(n21013) );
  OAI221_X1 U23959 ( .B1(n15189), .B2(keyinput209), .C1(n21014), .C2(
        keyinput152), .A(n21013), .ZN(n21019) );
  AOI22_X1 U23960 ( .A1(n21098), .A2(keyinput163), .B1(keyinput183), .B2(
        n21083), .ZN(n21015) );
  OAI221_X1 U23961 ( .B1(n21098), .B2(keyinput163), .C1(n21083), .C2(
        keyinput183), .A(n21015), .ZN(n21018) );
  AOI22_X1 U23962 ( .A1(n21113), .A2(keyinput128), .B1(keyinput189), .B2(
        n14849), .ZN(n21016) );
  OAI221_X1 U23963 ( .B1(n21113), .B2(keyinput128), .C1(n14849), .C2(
        keyinput189), .A(n21016), .ZN(n21017) );
  NOR4_X1 U23964 ( .A1(n21020), .A2(n21019), .A3(n21018), .A4(n21017), .ZN(
        n21056) );
  AOI22_X1 U23965 ( .A1(n21096), .A2(keyinput234), .B1(keyinput210), .B2(
        n21022), .ZN(n21021) );
  OAI221_X1 U23966 ( .B1(n21096), .B2(keyinput234), .C1(n21022), .C2(
        keyinput210), .A(n21021), .ZN(n21032) );
  AOI22_X1 U23967 ( .A1(n21025), .A2(keyinput166), .B1(n21024), .B2(
        keyinput236), .ZN(n21023) );
  OAI221_X1 U23968 ( .B1(n21025), .B2(keyinput166), .C1(n21024), .C2(
        keyinput236), .A(n21023), .ZN(n21031) );
  AOI22_X1 U23969 ( .A1(n21126), .A2(keyinput199), .B1(n9798), .B2(keyinput168), .ZN(n21026) );
  OAI221_X1 U23970 ( .B1(n21126), .B2(keyinput199), .C1(n21179), .C2(
        keyinput168), .A(n21026), .ZN(n21030) );
  AOI22_X1 U23971 ( .A1(n21028), .A2(keyinput194), .B1(keyinput181), .B2(
        n12889), .ZN(n21027) );
  OAI221_X1 U23972 ( .B1(n21028), .B2(keyinput194), .C1(n12889), .C2(
        keyinput181), .A(n21027), .ZN(n21029) );
  NOR4_X1 U23973 ( .A1(n21032), .A2(n21031), .A3(n21030), .A4(n21029), .ZN(
        n21055) );
  INV_X1 U23974 ( .A(DATAI_11_), .ZN(n21145) );
  AOI22_X1 U23975 ( .A1(n21145), .A2(keyinput157), .B1(n21162), .B2(
        keyinput138), .ZN(n21033) );
  OAI221_X1 U23976 ( .B1(n21145), .B2(keyinput157), .C1(n21162), .C2(
        keyinput138), .A(n21033), .ZN(n21042) );
  AOI22_X1 U23977 ( .A1(n21208), .A2(keyinput187), .B1(keyinput205), .B2(
        n21077), .ZN(n21034) );
  OAI221_X1 U23978 ( .B1(n21208), .B2(keyinput187), .C1(n21077), .C2(
        keyinput205), .A(n21034), .ZN(n21041) );
  AOI22_X1 U23979 ( .A1(n21209), .A2(keyinput184), .B1(n10449), .B2(
        keyinput227), .ZN(n21035) );
  OAI221_X1 U23980 ( .B1(n21209), .B2(keyinput184), .C1(n10449), .C2(
        keyinput227), .A(n21035), .ZN(n21040) );
  XNOR2_X1 U23981 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B(keyinput196), .ZN(
        n21037) );
  NAND2_X1 U23982 ( .A1(n21038), .A2(n21037), .ZN(n21039) );
  NOR4_X1 U23983 ( .A1(n21042), .A2(n21041), .A3(n21040), .A4(n21039), .ZN(
        n21054) );
  AOI22_X1 U23984 ( .A1(n21092), .A2(keyinput224), .B1(n21158), .B2(
        keyinput172), .ZN(n21043) );
  OAI221_X1 U23985 ( .B1(n21092), .B2(keyinput224), .C1(n21158), .C2(
        keyinput172), .A(n21043), .ZN(n21052) );
  INV_X1 U23986 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n21172) );
  AOI22_X1 U23987 ( .A1(n21172), .A2(keyinput161), .B1(n21045), .B2(
        keyinput235), .ZN(n21044) );
  OAI221_X1 U23988 ( .B1(n21172), .B2(keyinput161), .C1(n21045), .C2(
        keyinput235), .A(n21044), .ZN(n21051) );
  INV_X1 U23989 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n21110) );
  INV_X1 U23990 ( .A(P3_UWORD_REG_1__SCAN_IN), .ZN(n21135) );
  AOI22_X1 U23991 ( .A1(n21110), .A2(keyinput255), .B1(keyinput208), .B2(
        n21135), .ZN(n21046) );
  OAI221_X1 U23992 ( .B1(n21110), .B2(keyinput255), .C1(n21135), .C2(
        keyinput208), .A(n21046), .ZN(n21050) );
  AOI22_X1 U23993 ( .A1(n21048), .A2(keyinput252), .B1(keyinput222), .B2(
        n21079), .ZN(n21047) );
  OAI221_X1 U23994 ( .B1(n21048), .B2(keyinput252), .C1(n21079), .C2(
        keyinput222), .A(n21047), .ZN(n21049) );
  NOR4_X1 U23995 ( .A1(n21052), .A2(n21051), .A3(n21050), .A4(n21049), .ZN(
        n21053) );
  NAND4_X1 U23996 ( .A1(n21056), .A2(n21055), .A3(n21054), .A4(n21053), .ZN(
        n21057) );
  NOR4_X1 U23997 ( .A1(n21060), .A2(n21059), .A3(n21058), .A4(n21057), .ZN(
        n21268) );
  AOI22_X1 U23998 ( .A1(n21063), .A2(keyinput20), .B1(n21062), .B2(keyinput85), 
        .ZN(n21061) );
  OAI221_X1 U23999 ( .B1(n21063), .B2(keyinput20), .C1(n21062), .C2(keyinput85), .A(n21061), .ZN(n21074) );
  AOI22_X1 U24000 ( .A1(n21066), .A2(keyinput15), .B1(keyinput72), .B2(n21065), 
        .ZN(n21064) );
  OAI221_X1 U24001 ( .B1(n21066), .B2(keyinput15), .C1(n21065), .C2(keyinput72), .A(n21064), .ZN(n21073) );
  AOI22_X1 U24002 ( .A1(n21069), .A2(keyinput6), .B1(n21068), .B2(keyinput103), 
        .ZN(n21067) );
  OAI221_X1 U24003 ( .B1(n21069), .B2(keyinput6), .C1(n21068), .C2(keyinput103), .A(n21067), .ZN(n21072) );
  AOI22_X1 U24004 ( .A1(n12670), .A2(keyinput51), .B1(n14642), .B2(keyinput16), 
        .ZN(n21070) );
  OAI221_X1 U24005 ( .B1(n12670), .B2(keyinput51), .C1(n14642), .C2(keyinput16), .A(n21070), .ZN(n21071) );
  NOR4_X1 U24006 ( .A1(n21074), .A2(n21073), .A3(n21072), .A4(n21071), .ZN(
        n21124) );
  AOI22_X1 U24007 ( .A1(n21077), .A2(keyinput77), .B1(n21076), .B2(keyinput98), 
        .ZN(n21075) );
  OAI221_X1 U24008 ( .B1(n21077), .B2(keyinput77), .C1(n21076), .C2(keyinput98), .A(n21075), .ZN(n21090) );
  AOI22_X1 U24009 ( .A1(n21080), .A2(keyinput122), .B1(n21079), .B2(keyinput94), .ZN(n21078) );
  OAI221_X1 U24010 ( .B1(n21080), .B2(keyinput122), .C1(n21079), .C2(
        keyinput94), .A(n21078), .ZN(n21089) );
  INV_X1 U24011 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21082) );
  AOI22_X1 U24012 ( .A1(n21083), .A2(keyinput55), .B1(n21082), .B2(keyinput57), 
        .ZN(n21081) );
  OAI221_X1 U24013 ( .B1(n21083), .B2(keyinput55), .C1(n21082), .C2(keyinput57), .A(n21081), .ZN(n21088) );
  AOI22_X1 U24014 ( .A1(n21086), .A2(keyinput119), .B1(n21085), .B2(
        keyinput120), .ZN(n21084) );
  OAI221_X1 U24015 ( .B1(n21086), .B2(keyinput119), .C1(n21085), .C2(
        keyinput120), .A(n21084), .ZN(n21087) );
  NOR4_X1 U24016 ( .A1(n21090), .A2(n21089), .A3(n21088), .A4(n21087), .ZN(
        n21123) );
  AOI22_X1 U24017 ( .A1(n21093), .A2(keyinput8), .B1(keyinput96), .B2(n21092), 
        .ZN(n21091) );
  OAI221_X1 U24018 ( .B1(n21093), .B2(keyinput8), .C1(n21092), .C2(keyinput96), 
        .A(n21091), .ZN(n21105) );
  AOI22_X1 U24019 ( .A1(n21096), .A2(keyinput106), .B1(keyinput9), .B2(n21095), 
        .ZN(n21094) );
  OAI221_X1 U24020 ( .B1(n21096), .B2(keyinput106), .C1(n21095), .C2(keyinput9), .A(n21094), .ZN(n21104) );
  AOI22_X1 U24021 ( .A1(n21099), .A2(keyinput74), .B1(n21098), .B2(keyinput35), 
        .ZN(n21097) );
  OAI221_X1 U24022 ( .B1(n21099), .B2(keyinput74), .C1(n21098), .C2(keyinput35), .A(n21097), .ZN(n21103) );
  AOI22_X1 U24023 ( .A1(n21101), .A2(keyinput102), .B1(n10485), .B2(keyinput97), .ZN(n21100) );
  OAI221_X1 U24024 ( .B1(n21101), .B2(keyinput102), .C1(n10485), .C2(
        keyinput97), .A(n21100), .ZN(n21102) );
  NOR4_X1 U24025 ( .A1(n21105), .A2(n21104), .A3(n21103), .A4(n21102), .ZN(
        n21122) );
  AOI22_X1 U24026 ( .A1(n21108), .A2(keyinput109), .B1(n21107), .B2(
        keyinput117), .ZN(n21106) );
  OAI221_X1 U24027 ( .B1(n21108), .B2(keyinput109), .C1(n21107), .C2(
        keyinput117), .A(n21106), .ZN(n21120) );
  AOI22_X1 U24028 ( .A1(n21111), .A2(keyinput91), .B1(keyinput127), .B2(n21110), .ZN(n21109) );
  OAI221_X1 U24029 ( .B1(n21111), .B2(keyinput91), .C1(n21110), .C2(
        keyinput127), .A(n21109), .ZN(n21119) );
  AOI22_X1 U24030 ( .A1(n21113), .A2(keyinput0), .B1(n15021), .B2(keyinput101), 
        .ZN(n21112) );
  OAI221_X1 U24031 ( .B1(n21113), .B2(keyinput0), .C1(n15021), .C2(keyinput101), .A(n21112), .ZN(n21118) );
  AOI22_X1 U24032 ( .A1(n21116), .A2(keyinput100), .B1(n21115), .B2(keyinput46), .ZN(n21114) );
  OAI221_X1 U24033 ( .B1(n21116), .B2(keyinput100), .C1(n21115), .C2(
        keyinput46), .A(n21114), .ZN(n21117) );
  NOR4_X1 U24034 ( .A1(n21120), .A2(n21119), .A3(n21118), .A4(n21117), .ZN(
        n21121) );
  NAND4_X1 U24035 ( .A1(n21124), .A2(n21123), .A3(n21122), .A4(n21121), .ZN(
        n21267) );
  AOI22_X1 U24036 ( .A1(n21127), .A2(keyinput118), .B1(keyinput71), .B2(n21126), .ZN(n21125) );
  OAI221_X1 U24037 ( .B1(n21127), .B2(keyinput118), .C1(n21126), .C2(
        keyinput71), .A(n21125), .ZN(n21140) );
  AOI22_X1 U24038 ( .A1(n21130), .A2(keyinput76), .B1(keyinput111), .B2(n21129), .ZN(n21128) );
  OAI221_X1 U24039 ( .B1(n21130), .B2(keyinput76), .C1(n21129), .C2(
        keyinput111), .A(n21128), .ZN(n21139) );
  AOI22_X1 U24040 ( .A1(n21133), .A2(keyinput86), .B1(keyinput90), .B2(n21132), 
        .ZN(n21131) );
  OAI221_X1 U24041 ( .B1(n21133), .B2(keyinput86), .C1(n21132), .C2(keyinput90), .A(n21131), .ZN(n21138) );
  INV_X1 U24042 ( .A(P3_UWORD_REG_7__SCAN_IN), .ZN(n21136) );
  AOI22_X1 U24043 ( .A1(n21136), .A2(keyinput63), .B1(keyinput80), .B2(n21135), 
        .ZN(n21134) );
  OAI221_X1 U24044 ( .B1(n21136), .B2(keyinput63), .C1(n21135), .C2(keyinput80), .A(n21134), .ZN(n21137) );
  NOR4_X1 U24045 ( .A1(n21140), .A2(n21139), .A3(n21138), .A4(n21137), .ZN(
        n21188) );
  INV_X1 U24046 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n21143) );
  AOI22_X1 U24047 ( .A1(n21143), .A2(keyinput114), .B1(n21142), .B2(keyinput7), 
        .ZN(n21141) );
  OAI221_X1 U24048 ( .B1(n21143), .B2(keyinput114), .C1(n21142), .C2(keyinput7), .A(n21141), .ZN(n21154) );
  AOI22_X1 U24049 ( .A1(n21146), .A2(keyinput62), .B1(n21145), .B2(keyinput29), 
        .ZN(n21144) );
  OAI221_X1 U24050 ( .B1(n21146), .B2(keyinput62), .C1(n21145), .C2(keyinput29), .A(n21144), .ZN(n21153) );
  XOR2_X1 U24051 ( .A(n15189), .B(keyinput81), .Z(n21149) );
  XNOR2_X1 U24052 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B(keyinput68), .ZN(
        n21148) );
  XNOR2_X1 U24053 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B(keyinput115), .ZN(
        n21147) );
  NAND3_X1 U24054 ( .A1(n21149), .A2(n21148), .A3(n21147), .ZN(n21152) );
  XNOR2_X1 U24055 ( .A(n21150), .B(keyinput49), .ZN(n21151) );
  NOR4_X1 U24056 ( .A1(n21154), .A2(n21153), .A3(n21152), .A4(n21151), .ZN(
        n21187) );
  INV_X1 U24057 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n21156) );
  AOI22_X1 U24058 ( .A1(n21156), .A2(keyinput19), .B1(n14849), .B2(keyinput61), 
        .ZN(n21155) );
  OAI221_X1 U24059 ( .B1(n21156), .B2(keyinput19), .C1(n14849), .C2(keyinput61), .A(n21155), .ZN(n21169) );
  INV_X1 U24060 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21159) );
  AOI22_X1 U24061 ( .A1(n21159), .A2(keyinput89), .B1(keyinput44), .B2(n21158), 
        .ZN(n21157) );
  OAI221_X1 U24062 ( .B1(n21159), .B2(keyinput89), .C1(n21158), .C2(keyinput44), .A(n21157), .ZN(n21168) );
  AOI22_X1 U24063 ( .A1(n21162), .A2(keyinput10), .B1(keyinput73), .B2(n21161), 
        .ZN(n21160) );
  OAI221_X1 U24064 ( .B1(n21162), .B2(keyinput10), .C1(n21161), .C2(keyinput73), .A(n21160), .ZN(n21167) );
  INV_X1 U24065 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21164) );
  AOI22_X1 U24066 ( .A1(n21165), .A2(keyinput37), .B1(keyinput83), .B2(n21164), 
        .ZN(n21163) );
  OAI221_X1 U24067 ( .B1(n21165), .B2(keyinput37), .C1(n21164), .C2(keyinput83), .A(n21163), .ZN(n21166) );
  NOR4_X1 U24068 ( .A1(n21169), .A2(n21168), .A3(n21167), .A4(n21166), .ZN(
        n21186) );
  AOI22_X1 U24069 ( .A1(n21172), .A2(keyinput33), .B1(keyinput84), .B2(n21171), 
        .ZN(n21170) );
  OAI221_X1 U24070 ( .B1(n21172), .B2(keyinput33), .C1(n21171), .C2(keyinput84), .A(n21170), .ZN(n21184) );
  INV_X1 U24071 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21174) );
  AOI22_X1 U24072 ( .A1(n21175), .A2(keyinput25), .B1(n21174), .B2(keyinput112), .ZN(n21173) );
  OAI221_X1 U24073 ( .B1(n21175), .B2(keyinput25), .C1(n21174), .C2(
        keyinput112), .A(n21173), .ZN(n21183) );
  AOI22_X1 U24074 ( .A1(n21177), .A2(keyinput113), .B1(keyinput53), .B2(n12889), .ZN(n21176) );
  OAI221_X1 U24075 ( .B1(n21177), .B2(keyinput113), .C1(n12889), .C2(
        keyinput53), .A(n21176), .ZN(n21182) );
  AOI22_X1 U24076 ( .A1(n21180), .A2(keyinput121), .B1(keyinput40), .B2(n21179), .ZN(n21178) );
  OAI221_X1 U24077 ( .B1(n21180), .B2(keyinput121), .C1(n21179), .C2(
        keyinput40), .A(n21178), .ZN(n21181) );
  NOR4_X1 U24078 ( .A1(n21184), .A2(n21183), .A3(n21182), .A4(n21181), .ZN(
        n21185) );
  NAND4_X1 U24079 ( .A1(n21188), .A2(n21187), .A3(n21186), .A4(n21185), .ZN(
        n21266) );
  OAI22_X1 U24080 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(keyinput17), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(keyinput30), .ZN(n21189) );
  AOI221_X1 U24081 ( .B1(P3_REIP_REG_29__SCAN_IN), .B2(keyinput17), .C1(
        keyinput30), .C2(P1_UWORD_REG_1__SCAN_IN), .A(n21189), .ZN(n21196) );
  OAI22_X1 U24082 ( .A1(P1_EBX_REG_30__SCAN_IN), .A2(keyinput14), .B1(
        keyinput92), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n21190) );
  AOI221_X1 U24083 ( .B1(P1_EBX_REG_30__SCAN_IN), .B2(keyinput14), .C1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .C2(keyinput92), .A(n21190), .ZN(
        n21195) );
  OAI22_X1 U24084 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(keyinput60), .B1(
        keyinput24), .B2(P1_EBX_REG_16__SCAN_IN), .ZN(n21191) );
  AOI221_X1 U24085 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(keyinput60), .C1(
        P1_EBX_REG_16__SCAN_IN), .C2(keyinput24), .A(n21191), .ZN(n21194) );
  OAI22_X1 U24086 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(keyinput48), .B1(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput116), .ZN(n21192) );
  AOI221_X1 U24087 ( .B1(P2_REIP_REG_0__SCAN_IN), .B2(keyinput48), .C1(
        keyinput116), .C2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n21192), 
        .ZN(n21193) );
  NAND4_X1 U24088 ( .A1(n21196), .A2(n21195), .A3(n21194), .A4(n21193), .ZN(
        n21226) );
  OAI22_X1 U24089 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(keyinput75), 
        .B1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput43), .ZN(n21197)
         );
  AOI221_X1 U24090 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput75), 
        .C1(keyinput43), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(n21197), 
        .ZN(n21204) );
  OAI22_X1 U24091 ( .A1(P1_EBX_REG_20__SCAN_IN), .A2(keyinput126), .B1(
        P3_DATAWIDTH_REG_29__SCAN_IN), .B2(keyinput50), .ZN(n21198) );
  AOI221_X1 U24092 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(keyinput126), .C1(
        keyinput50), .C2(P3_DATAWIDTH_REG_29__SCAN_IN), .A(n21198), .ZN(n21203) );
  OAI22_X1 U24093 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(keyinput47), 
        .B1(P3_DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput87), .ZN(n21199) );
  AOI221_X1 U24094 ( .B1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput47), 
        .C1(keyinput87), .C2(P3_DATAWIDTH_REG_20__SCAN_IN), .A(n21199), .ZN(
        n21202) );
  OAI22_X1 U24095 ( .A1(BUF1_REG_8__SCAN_IN), .A2(keyinput88), .B1(keyinput31), 
        .B2(BUF1_REG_7__SCAN_IN), .ZN(n21200) );
  AOI221_X1 U24096 ( .B1(BUF1_REG_8__SCAN_IN), .B2(keyinput88), .C1(
        BUF1_REG_7__SCAN_IN), .C2(keyinput31), .A(n21200), .ZN(n21201) );
  NAND4_X1 U24097 ( .A1(n21204), .A2(n21203), .A3(n21202), .A4(n21201), .ZN(
        n21225) );
  OAI22_X1 U24098 ( .A1(P1_EAX_REG_29__SCAN_IN), .A2(keyinput4), .B1(
        keyinput104), .B2(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21205) );
  AOI221_X1 U24099 ( .B1(P1_EAX_REG_29__SCAN_IN), .B2(keyinput4), .C1(
        P1_ADDRESS_REG_3__SCAN_IN), .C2(keyinput104), .A(n21205), .ZN(n21214)
         );
  OAI22_X1 U24100 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(keyinput99), .B1(
        P3_INSTQUEUE_REG_7__2__SCAN_IN), .B2(keyinput123), .ZN(n21206) );
  AOI221_X1 U24101 ( .B1(P2_EBX_REG_11__SCAN_IN), .B2(keyinput99), .C1(
        keyinput123), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(n21206), .ZN(
        n21213) );
  OAI22_X1 U24102 ( .A1(n21209), .A2(keyinput56), .B1(n21208), .B2(keyinput59), 
        .ZN(n21207) );
  AOI221_X1 U24103 ( .B1(n21209), .B2(keyinput56), .C1(keyinput59), .C2(n21208), .A(n21207), .ZN(n21212) );
  OAI22_X1 U24104 ( .A1(P2_ADDRESS_REG_4__SCAN_IN), .A2(keyinput108), .B1(
        P2_LWORD_REG_14__SCAN_IN), .B2(keyinput110), .ZN(n21210) );
  AOI221_X1 U24105 ( .B1(P2_ADDRESS_REG_4__SCAN_IN), .B2(keyinput108), .C1(
        keyinput110), .C2(P2_LWORD_REG_14__SCAN_IN), .A(n21210), .ZN(n21211)
         );
  NAND4_X1 U24106 ( .A1(n21214), .A2(n21213), .A3(n21212), .A4(n21211), .ZN(
        n21224) );
  OAI22_X1 U24107 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(keyinput32), .B1(
        keyinput54), .B2(P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21215) );
  AOI221_X1 U24108 ( .B1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B2(keyinput32), 
        .C1(P2_DATAWIDTH_REG_8__SCAN_IN), .C2(keyinput54), .A(n21215), .ZN(
        n21222) );
  OAI22_X1 U24109 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(keyinput45), .B1(
        keyinput23), .B2(P3_EAX_REG_17__SCAN_IN), .ZN(n21216) );
  AOI221_X1 U24110 ( .B1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput45), 
        .C1(P3_EAX_REG_17__SCAN_IN), .C2(keyinput23), .A(n21216), .ZN(n21221)
         );
  OAI22_X1 U24111 ( .A1(BUF2_REG_10__SCAN_IN), .A2(keyinput3), .B1(keyinput125), .B2(DATAI_17_), .ZN(n21217) );
  AOI221_X1 U24112 ( .B1(BUF2_REG_10__SCAN_IN), .B2(keyinput3), .C1(DATAI_17_), 
        .C2(keyinput125), .A(n21217), .ZN(n21220) );
  OAI22_X1 U24113 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(keyinput36), .B1(
        keyinput67), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n21218) );
  AOI221_X1 U24114 ( .B1(P2_ADDRESS_REG_6__SCAN_IN), .B2(keyinput36), .C1(
        P3_REIP_REG_3__SCAN_IN), .C2(keyinput67), .A(n21218), .ZN(n21219) );
  NAND4_X1 U24115 ( .A1(n21222), .A2(n21221), .A3(n21220), .A4(n21219), .ZN(
        n21223) );
  NOR4_X1 U24116 ( .A1(n21226), .A2(n21225), .A3(n21224), .A4(n21223), .ZN(
        n21264) );
  OAI22_X1 U24117 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(keyinput34), .B1(
        keyinput95), .B2(BUF1_REG_18__SCAN_IN), .ZN(n21227) );
  AOI221_X1 U24118 ( .B1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput34), 
        .C1(BUF1_REG_18__SCAN_IN), .C2(keyinput95), .A(n21227), .ZN(n21234) );
  OAI22_X1 U24119 ( .A1(P1_EAX_REG_28__SCAN_IN), .A2(keyinput70), .B1(
        P2_UWORD_REG_2__SCAN_IN), .B2(keyinput41), .ZN(n21228) );
  AOI221_X1 U24120 ( .B1(P1_EAX_REG_28__SCAN_IN), .B2(keyinput70), .C1(
        keyinput41), .C2(P2_UWORD_REG_2__SCAN_IN), .A(n21228), .ZN(n21233) );
  OAI22_X1 U24121 ( .A1(P2_EBX_REG_7__SCAN_IN), .A2(keyinput58), .B1(
        keyinput22), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n21229) );
  AOI221_X1 U24122 ( .B1(P2_EBX_REG_7__SCAN_IN), .B2(keyinput58), .C1(
        P3_INSTQUEUE_REG_8__0__SCAN_IN), .C2(keyinput22), .A(n21229), .ZN(
        n21232) );
  OAI22_X1 U24123 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(keyinput12), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(keyinput13), .ZN(n21230) );
  AOI221_X1 U24124 ( .B1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput12), 
        .C1(keyinput13), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n21230), 
        .ZN(n21231) );
  NAND4_X1 U24125 ( .A1(n21234), .A2(n21233), .A3(n21232), .A4(n21231), .ZN(
        n21262) );
  OAI22_X1 U24126 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(keyinput64), .B1(
        P1_EBX_REG_27__SCAN_IN), .B2(keyinput52), .ZN(n21235) );
  AOI221_X1 U24127 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(keyinput64), .C1(
        keyinput52), .C2(P1_EBX_REG_27__SCAN_IN), .A(n21235), .ZN(n21242) );
  OAI22_X1 U24128 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(keyinput1), .B1(
        P3_DATAWIDTH_REG_24__SCAN_IN), .B2(keyinput21), .ZN(n21236) );
  AOI221_X1 U24129 ( .B1(P2_ADDRESS_REG_15__SCAN_IN), .B2(keyinput1), .C1(
        keyinput21), .C2(P3_DATAWIDTH_REG_24__SCAN_IN), .A(n21236), .ZN(n21241) );
  OAI22_X1 U24130 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(keyinput28), 
        .B1(keyinput105), .B2(P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n21237) );
  AOI221_X1 U24131 ( .B1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B2(keyinput28), 
        .C1(P1_DATAWIDTH_REG_6__SCAN_IN), .C2(keyinput105), .A(n21237), .ZN(
        n21240) );
  OAI22_X1 U24132 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput5), 
        .B1(P3_ADDRESS_REG_2__SCAN_IN), .B2(keyinput11), .ZN(n21238) );
  AOI221_X1 U24133 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput5), 
        .C1(keyinput11), .C2(P3_ADDRESS_REG_2__SCAN_IN), .A(n21238), .ZN(
        n21239) );
  NAND4_X1 U24134 ( .A1(n21242), .A2(n21241), .A3(n21240), .A4(n21239), .ZN(
        n21261) );
  OAI22_X1 U24135 ( .A1(BUF2_REG_2__SCAN_IN), .A2(keyinput38), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(keyinput27), .ZN(n21243) );
  AOI221_X1 U24136 ( .B1(BUF2_REG_2__SCAN_IN), .B2(keyinput38), .C1(keyinput27), .C2(P1_LWORD_REG_11__SCAN_IN), .A(n21243), .ZN(n21250) );
  OAI22_X1 U24137 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput69), 
        .B1(keyinput18), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n21244) );
  AOI221_X1 U24138 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput69), 
        .C1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .C2(keyinput18), .A(n21244), .ZN(
        n21249) );
  OAI22_X1 U24139 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(keyinput39), 
        .B1(keyinput2), .B2(P1_EAX_REG_4__SCAN_IN), .ZN(n21245) );
  AOI221_X1 U24140 ( .B1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(keyinput39), 
        .C1(P1_EAX_REG_4__SCAN_IN), .C2(keyinput2), .A(n21245), .ZN(n21248) );
  OAI22_X1 U24141 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(keyinput107), 
        .B1(keyinput93), .B2(BUF1_REG_4__SCAN_IN), .ZN(n21246) );
  AOI221_X1 U24142 ( .B1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B2(keyinput107), 
        .C1(BUF1_REG_4__SCAN_IN), .C2(keyinput93), .A(n21246), .ZN(n21247) );
  NAND4_X1 U24143 ( .A1(n21250), .A2(n21249), .A3(n21248), .A4(n21247), .ZN(
        n21260) );
  OAI22_X1 U24144 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(keyinput42), .B1(
        keyinput79), .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n21251) );
  AOI221_X1 U24145 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(keyinput42), .C1(
        P1_DATAO_REG_25__SCAN_IN), .C2(keyinput79), .A(n21251), .ZN(n21258) );
  OAI22_X1 U24146 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(keyinput124), 
        .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput26), .ZN(n21252)
         );
  AOI221_X1 U24147 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput124), 
        .C1(keyinput26), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n21252), 
        .ZN(n21257) );
  OAI22_X1 U24148 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(keyinput66), 
        .B1(keyinput78), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21253) );
  AOI221_X1 U24149 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput66), 
        .C1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .C2(keyinput78), .A(n21253), .ZN(
        n21256) );
  OAI22_X1 U24150 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(keyinput65), .B1(
        P3_STATE2_REG_1__SCAN_IN), .B2(keyinput82), .ZN(n21254) );
  AOI221_X1 U24151 ( .B1(P2_ADDRESS_REG_24__SCAN_IN), .B2(keyinput65), .C1(
        keyinput82), .C2(P3_STATE2_REG_1__SCAN_IN), .A(n21254), .ZN(n21255) );
  NAND4_X1 U24152 ( .A1(n21258), .A2(n21257), .A3(n21256), .A4(n21255), .ZN(
        n21259) );
  NOR4_X1 U24153 ( .A1(n21262), .A2(n21261), .A3(n21260), .A4(n21259), .ZN(
        n21263) );
  NAND2_X1 U24154 ( .A1(n21264), .A2(n21263), .ZN(n21265) );
  NOR4_X1 U24155 ( .A1(n21268), .A2(n21267), .A3(n21266), .A4(n21265), .ZN(
        n21269) );
  XNOR2_X1 U24156 ( .A(n21270), .B(n21269), .ZN(U246) );
  INV_X1 U13361 ( .A(n10540), .ZN(n11555) );
  AND2_X1 U12798 ( .A1(n11337), .A2(n10362), .ZN(n10363) );
  OAI21_X1 U11524 ( .B1(n12694), .B2(n12754), .A(n12693), .ZN(n13086) );
  NAND2_X1 U12795 ( .A1(n15371), .A2(n11608), .ZN(n15511) );
  CLKBUF_X1 U11245 ( .A(n11902), .Z(n11791) );
  AND4_X1 U11263 ( .A1(n11651), .A2(n11650), .A3(n11649), .A4(n11648), .ZN(
        n11652) );
  NOR2_X1 U11276 ( .A1(n13036), .A2(n11555), .ZN(n10353) );
  CLKBUF_X1 U11281 ( .A(n10676), .Z(n14143) );
  NAND2_X1 U11283 ( .A1(n16036), .A2(n16035), .ZN(n16034) );
  INV_X1 U11285 ( .A(n10655), .ZN(n10645) );
  INV_X1 U11318 ( .A(n10931), .ZN(n10959) );
  CLKBUF_X1 U11339 ( .A(n10768), .Z(n13515) );
  CLKBUF_X1 U11361 ( .A(n12530), .Z(n12655) );
  AOI21_X1 U11364 ( .B1(n10071), .B2(n9867), .A(n9829), .ZN(n10069) );
  OR2_X1 U11376 ( .A1(n13010), .A2(n13786), .ZN(n13825) );
  CLKBUF_X1 U11496 ( .A(n13068), .Z(n20613) );
  INV_X1 U11586 ( .A(n13140), .ZN(n10627) );
  CLKBUF_X1 U11763 ( .A(n11938), .Z(n11939) );
  NAND2_X1 U11821 ( .A1(n13691), .A2(n13717), .ZN(n13716) );
  CLKBUF_X1 U11912 ( .A(n14807), .Z(n14813) );
  CLKBUF_X1 U12001 ( .A(n17539), .Z(n17542) );
  OR2_X1 U12032 ( .A1(n20265), .A2(n20254), .ZN(n21271) );
  OR2_X1 U12245 ( .A1(n11013), .A2(n11009), .ZN(n21272) );
  NOR2_X2 U12434 ( .A1(n13317), .A2(n13318), .ZN(n13316) );
  AND2_X2 U12548 ( .A1(n13487), .A2(n13692), .ZN(n13691) );
  NAND2_X2 U12633 ( .A1(n9918), .A2(n12018), .ZN(n12757) );
  NAND2_X4 U12638 ( .A1(n12757), .A2(n12756), .ZN(n12766) );
  OAI21_X2 U12724 ( .B1(n14761), .B2(n12779), .A(n14858), .ZN(n14753) );
  CLKBUF_X1 U12854 ( .A(n11875), .Z(n11793) );
  CLKBUF_X1 U13699 ( .A(n11827), .Z(n12396) );
endmodule

