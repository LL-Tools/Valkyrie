

module b17_C_AntiSAT_k_256_3 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9819, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9839, n9840, n9841,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629;

  INV_X1 U11263 ( .A(n16219), .ZN(n16189) );
  INV_X1 U11264 ( .A(n14592), .ZN(n11183) );
  INV_X2 U11265 ( .A(n17157), .ZN(n17065) );
  INV_X2 U11266 ( .A(n16194), .ZN(n14999) );
  NOR2_X1 U11267 ( .A1(n10750), .A2(n10749), .ZN(n10776) );
  INV_X1 U11268 ( .A(n17612), .ZN(n18545) );
  NAND2_X1 U11269 ( .A1(n11848), .A2(n11847), .ZN(n12016) );
  NOR2_X1 U11270 ( .A1(n11840), .A2(n19533), .ZN(n19977) );
  BUF_X2 U11271 ( .A(n13288), .Z(n11832) );
  BUF_X2 U11272 ( .A(n13270), .Z(n14338) );
  INV_X1 U11273 ( .A(n13375), .ZN(n13430) );
  INV_X1 U11274 ( .A(n13371), .ZN(n13427) );
  CLKBUF_X1 U11275 ( .A(n10551), .Z(n20517) );
  CLKBUF_X2 U11276 ( .A(n10471), .Z(n9836) );
  CLKBUF_X2 U11277 ( .A(n10500), .Z(n9862) );
  INV_X2 U11278 ( .A(n10551), .ZN(n13974) );
  INV_X1 U11279 ( .A(n12916), .ZN(n17473) );
  AND2_X1 U11280 ( .A1(n10032), .A2(n10061), .ZN(n9924) );
  INV_X1 U11281 ( .A(n9911), .ZN(n17451) );
  CLKBUF_X3 U11283 ( .A(n10479), .Z(n11213) );
  NAND2_X1 U11284 ( .A1(n11695), .A2(n11694), .ZN(n11886) );
  AND2_X1 U11285 ( .A1(n14044), .A2(n13839), .ZN(n11058) );
  CLKBUF_X1 U11286 ( .A(n9839), .Z(n9830) );
  AND2_X1 U11287 ( .A1(n10401), .A2(n10405), .ZN(n10471) );
  AND2_X2 U11288 ( .A1(n14064), .A2(n14045), .ZN(n10479) );
  AND2_X1 U11289 ( .A1(n10394), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10401) );
  BUF_X1 U11290 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11784) );
  CLKBUF_X1 U11291 ( .A(n10707), .Z(n9819) );
  NOR2_X1 U11292 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10707) );
  AND2_X1 U11294 ( .A1(n10405), .A2(n14045), .ZN(n9839) );
  BUF_X1 U11295 ( .A(n9839), .Z(n9825) );
  CLKBUF_X2 U11296 ( .A(n11058), .Z(n9856) );
  AND4_X1 U11297 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10430) );
  INV_X1 U11298 ( .A(n13447), .ZN(n12661) );
  AND3_X1 U11299 ( .A1(n20534), .A2(n20501), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11289) );
  NAND2_X1 U11300 ( .A1(n11702), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12690) );
  NOR2_X1 U11301 ( .A1(n11832), .A2(n11831), .ZN(n19579) );
  OR2_X1 U11302 ( .A1(n12885), .A2(n12887), .ZN(n12956) );
  NAND2_X1 U11303 ( .A1(n19108), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12887) );
  INV_X1 U11304 ( .A(n11725), .ZN(n12226) );
  NAND2_X1 U11305 ( .A1(n11816), .A2(n11782), .ZN(n11813) );
  INV_X1 U11307 ( .A(n10029), .ZN(n17481) );
  NAND2_X1 U11308 ( .A1(n11886), .A2(n14199), .ZN(n12362) );
  AND4_X1 U11309 ( .A1(n12121), .A2(n12120), .A3(n12119), .A4(n12118), .ZN(
        n12320) );
  NOR2_X2 U11310 ( .A1(n13205), .A2(n15439), .ZN(n13183) );
  XNOR2_X1 U11311 ( .A(n11813), .B(n11812), .ZN(n13270) );
  INV_X1 U11312 ( .A(n12320), .ZN(n12787) );
  BUF_X1 U11313 ( .A(n11814), .Z(n11820) );
  INV_X1 U11314 ( .A(n13982), .ZN(n10288) );
  NOR2_X1 U11315 ( .A1(n15208), .A2(n13590), .ZN(n13617) );
  INV_X1 U11317 ( .A(n12916), .ZN(n17458) );
  NAND2_X1 U11318 ( .A1(n18375), .A2(n18956), .ZN(n18393) );
  INV_X1 U11319 ( .A(n20307), .ZN(n20294) );
  INV_X1 U11320 ( .A(n20350), .ZN(n20333) );
  NAND2_X2 U11321 ( .A1(n20561), .A2(n10608), .ZN(n14077) );
  INV_X1 U11322 ( .A(n20435), .ZN(n20258) );
  NOR2_X1 U11323 ( .A1(n18511), .A2(n18393), .ZN(n18945) );
  INV_X1 U11324 ( .A(n10887), .ZN(n9829) );
  AOI22_X2 U11325 ( .A1(n13006), .A2(n10064), .B1(n10376), .B2(n9916), .ZN(
        n13249) );
  NOR2_X1 U11326 ( .A1(n15992), .A2(n16684), .ZN(n15991) );
  AND3_X1 U11327 ( .A1(n11733), .A2(n11725), .A3(n12202), .ZN(n11726) );
  NOR2_X2 U11328 ( .A1(n18030), .A2(n17806), .ZN(n16702) );
  AND2_X2 U11329 ( .A1(n10273), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10406) );
  OAI21_X2 U11330 ( .B1(n12229), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10013), .ZN(n14392) );
  INV_X8 U11331 ( .A(n10391), .ZN(n17449) );
  AND2_X1 U11332 ( .A1(n11438), .A2(n10546), .ZN(n13771) );
  NAND2_X2 U11333 ( .A1(n9918), .A2(n9885), .ZN(n10546) );
  INV_X2 U11334 ( .A(n10602), .ZN(n10543) );
  XNOR2_X2 U11335 ( .A(n12969), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18155) );
  XNOR2_X2 U11336 ( .A(n12100), .B(n12101), .ZN(n12250) );
  NAND2_X2 U11337 ( .A1(n12051), .A2(n12050), .ZN(n12100) );
  NAND2_X2 U11339 ( .A1(n11338), .A2(n11337), .ZN(n11343) );
  NOR2_X2 U11340 ( .A1(n15241), .A2(n13479), .ZN(n13501) );
  CLKBUF_X1 U11342 ( .A(n10471), .Z(n9837) );
  XNOR2_X2 U11343 ( .A(n13526), .B(n9981), .ZN(n15228) );
  NAND2_X2 U11344 ( .A1(n15234), .A2(n13504), .ZN(n13526) );
  OAI221_X2 U11345 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18030), 
        .C1(n21488), .C2(n17840), .A(n17839), .ZN(n17818) );
  NOR3_X1 U11347 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19108), .A3(
        n17153), .ZN(n12957) );
  NOR4_X2 U11348 ( .A1(n17649), .A2(n16702), .A3(n17794), .A4(n18942), .ZN(
        n16709) );
  INV_X4 U11349 ( .A(n9915), .ZN(n9822) );
  INV_X1 U11350 ( .A(n9915), .ZN(n9823) );
  AND2_X4 U11351 ( .A1(n11855), .A2(n11784), .ZN(n11866) );
  XNOR2_X1 U11352 ( .A(n12843), .B(n12842), .ZN(n12861) );
  AND2_X1 U11353 ( .A1(n10091), .A2(n10090), .ZN(n14857) );
  OR2_X1 U11354 ( .A1(n13000), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17807) );
  AND2_X1 U11355 ( .A1(n12867), .A2(n12825), .ZN(n13640) );
  AND2_X1 U11356 ( .A1(n15303), .A2(n15302), .ZN(n16389) );
  CLKBUF_X1 U11357 ( .A(n17857), .Z(n17928) );
  OR3_X1 U11358 ( .A1(n12354), .A2(n12320), .A3(n15596), .ZN(n15426) );
  AND2_X1 U11360 ( .A1(n11844), .A2(n15836), .ZN(n19736) );
  NAND2_X1 U11362 ( .A1(n12288), .A2(n12287), .ZN(n12309) );
  OR2_X1 U11363 ( .A1(n12292), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12294) );
  INV_X1 U11364 ( .A(n18965), .ZN(n18956) );
  CLKBUF_X2 U11366 ( .A(n12389), .Z(n12795) );
  AND2_X1 U11367 ( .A1(n12809), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13204) );
  CLKBUF_X2 U11368 ( .A(n11789), .Z(n12844) );
  OR2_X1 U11369 ( .A1(n13197), .A2(n10161), .ZN(n10160) );
  CLKBUF_X2 U11370 ( .A(n11732), .Z(n19557) );
  NAND2_X1 U11371 ( .A1(n9859), .A2(n16637), .ZN(n12148) );
  CLKBUF_X3 U11372 ( .A(n12226), .Z(n12227) );
  CLKBUF_X3 U11373 ( .A(n11886), .Z(n14211) );
  INV_X2 U11374 ( .A(n14199), .ZN(n16637) );
  INV_X2 U11375 ( .A(n12944), .ZN(n17343) );
  CLKBUF_X2 U11376 ( .A(n10717), .Z(n11001) );
  CLKBUF_X2 U11377 ( .A(n10489), .Z(n10989) );
  INV_X2 U11378 ( .A(n12690), .ZN(n13431) );
  CLKBUF_X2 U11379 ( .A(n11043), .Z(n11144) );
  INV_X2 U11380 ( .A(n9917), .ZN(n17432) );
  CLKBUF_X1 U11383 ( .A(n9839), .Z(n9841) );
  CLKBUF_X1 U11384 ( .A(n9913), .Z(n10533) );
  CLKBUF_X2 U11385 ( .A(n10479), .Z(n9855) );
  OR2_X1 U11386 ( .A1(n12888), .A2(n12880), .ZN(n15920) );
  CLKBUF_X1 U11387 ( .A(n10630), .Z(n9826) );
  CLKBUF_X2 U11388 ( .A(n11861), .Z(n13606) );
  NOR2_X2 U11389 ( .A1(n13017), .A2(n19121), .ZN(n18957) );
  INV_X4 U11390 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16617) );
  OAI21_X1 U11391 ( .B1(n12861), .B2(n16543), .A(n10381), .ZN(n12857) );
  OR2_X1 U11392 ( .A1(n12829), .A2(n16543), .ZN(n12816) );
  AOI21_X1 U11393 ( .B1(n12835), .B2(n12834), .A(n12833), .ZN(n12841) );
  AOI21_X1 U11394 ( .B1(n10232), .B2(n10231), .A(n12781), .ZN(n15396) );
  NAND2_X1 U11395 ( .A1(n12777), .A2(n12356), .ZN(n15406) );
  NAND2_X1 U11396 ( .A1(n14857), .A2(n11414), .ZN(n14849) );
  OAI21_X1 U11397 ( .B1(n14898), .B2(n20496), .A(n10046), .ZN(n10045) );
  OR2_X1 U11398 ( .A1(n15054), .A2(n20258), .ZN(n10048) );
  NAND2_X1 U11399 ( .A1(n10018), .A2(n15527), .ZN(n15522) );
  NAND2_X1 U11400 ( .A1(n14620), .A2(n10047), .ZN(n14898) );
  AND2_X1 U11401 ( .A1(n10250), .A2(n10248), .ZN(n15427) );
  OR2_X1 U11402 ( .A1(n14621), .A2(n14619), .ZN(n10047) );
  OR2_X1 U11403 ( .A1(n15528), .A2(n15461), .ZN(n10018) );
  NOR2_X1 U11404 ( .A1(n16516), .A2(n15724), .ZN(n15753) );
  CLKBUF_X1 U11405 ( .A(n14592), .Z(n14593) );
  NOR2_X1 U11406 ( .A1(n14618), .A2(n11137), .ZN(n14607) );
  OAI21_X1 U11407 ( .B1(n10259), .B2(n9960), .A(n10007), .ZN(n15454) );
  INV_X1 U11408 ( .A(n10080), .ZN(n16510) );
  CLKBUF_X1 U11409 ( .A(n14659), .Z(n14660) );
  NAND2_X1 U11410 ( .A1(n10096), .A2(n16172), .ZN(n11409) );
  NAND2_X1 U11411 ( .A1(n14988), .A2(n10282), .ZN(n16173) );
  NAND2_X1 U11412 ( .A1(n10012), .A2(n12267), .ZN(n13655) );
  OAI22_X1 U11413 ( .A1(n19492), .A2(n19491), .B1(n14285), .B2(n19502), .ZN(
        n14393) );
  OAI21_X1 U11414 ( .B1(n10282), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16194), .ZN(n10281) );
  AND2_X1 U11415 ( .A1(n10283), .A2(n9950), .ZN(n10282) );
  INV_X1 U11416 ( .A(n14395), .ZN(n12048) );
  AND2_X1 U11417 ( .A1(n12047), .A2(n14403), .ZN(n14395) );
  AOI21_X1 U11418 ( .B1(n12229), .B2(n9897), .A(n9959), .ZN(n10013) );
  NAND2_X1 U11419 ( .A1(n10025), .A2(n10023), .ZN(n16204) );
  AND2_X1 U11420 ( .A1(n10024), .A2(n16210), .ZN(n10023) );
  OR2_X1 U11421 ( .A1(n14991), .A2(n11399), .ZN(n14978) );
  AOI22_X1 U11422 ( .A1(n9932), .A2(n10255), .B1(n10253), .B2(n10252), .ZN(
        n10251) );
  AND2_X1 U11423 ( .A1(n12046), .A2(n12045), .ZN(n12050) );
  AND2_X1 U11424 ( .A1(n12093), .A2(n12092), .ZN(n12101) );
  AND2_X1 U11425 ( .A1(n11964), .A2(n11963), .ZN(n11965) );
  OR2_X1 U11426 ( .A1(n11407), .A2(n21526), .ZN(n14977) );
  AND4_X1 U11427 ( .A1(n12014), .A2(n12013), .A3(n12012), .A4(n12011), .ZN(
        n12023) );
  NAND2_X1 U11428 ( .A1(n11389), .A2(n11388), .ZN(n11407) );
  AND3_X1 U11429 ( .A1(n11835), .A2(n11834), .A3(n11833), .ZN(n11836) );
  INV_X1 U11430 ( .A(n16566), .ZN(n15381) );
  OAI21_X1 U11431 ( .B1(n18067), .B2(n10068), .A(n10067), .ZN(n17996) );
  AND2_X1 U11432 ( .A1(n10226), .A2(n10225), .ZN(n11834) );
  OAI21_X1 U11433 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n15966), .A(n16814), 
        .ZN(n18164) );
  NOR2_X2 U11434 ( .A1(n10315), .A2(n15836), .ZN(n12015) );
  AND2_X1 U11435 ( .A1(n11848), .A2(n9935), .ZN(n20022) );
  NOR2_X1 U11436 ( .A1(n14746), .A2(n11524), .ZN(n14735) );
  NAND2_X1 U11437 ( .A1(n9887), .A2(n14338), .ZN(n14262) );
  NAND2_X1 U11438 ( .A1(n13286), .A2(n13285), .ZN(n13890) );
  NAND2_X1 U11439 ( .A1(n11848), .A2(n11845), .ZN(n19824) );
  NOR2_X1 U11440 ( .A1(n11840), .A2(n14338), .ZN(n14228) );
  NOR2_X2 U11441 ( .A1(n14036), .A2(n20497), .ZN(n11311) );
  NAND2_X1 U11442 ( .A1(n9887), .A2(n19533), .ZN(n19911) );
  NOR2_X1 U11443 ( .A1(n11839), .A2(n19533), .ZN(n11844) );
  NOR2_X2 U11444 ( .A1(n11832), .A2(n11825), .ZN(n14202) );
  OR2_X1 U11445 ( .A1(n15793), .A2(n10289), .ZN(n15761) );
  AND2_X1 U11446 ( .A1(n13285), .A2(n13276), .ZN(n13828) );
  XNOR2_X1 U11447 ( .A(n10606), .B(n10605), .ZN(n10019) );
  NAND2_X1 U11448 ( .A1(n18079), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18078) );
  CLKBUF_X1 U11449 ( .A(n14076), .Z(n9870) );
  AOI21_X1 U11450 ( .B1(n10661), .B2(n10662), .A(n10655), .ZN(n10656) );
  NAND2_X1 U11451 ( .A1(n15795), .A2(n15794), .ZN(n15793) );
  NAND2_X1 U11452 ( .A1(n12294), .A2(n12357), .ZN(n12288) );
  AOI21_X1 U11453 ( .B1(n13749), .B2(n13750), .A(n13284), .ZN(n13829) );
  NAND2_X1 U11454 ( .A1(n10328), .A2(n11799), .ZN(n12375) );
  NOR2_X1 U11455 ( .A1(n9878), .A2(n10149), .ZN(n19261) );
  NAND2_X1 U11456 ( .A1(n11813), .A2(n11812), .ZN(n10328) );
  INV_X1 U11457 ( .A(n9871), .ZN(n9878) );
  NOR2_X1 U11458 ( .A1(n13991), .A2(n14194), .ZN(n19387) );
  NAND2_X1 U11459 ( .A1(n13281), .A2(n13280), .ZN(n15819) );
  NAND2_X1 U11460 ( .A1(n10021), .A2(n10589), .ZN(n10020) );
  AND2_X1 U11461 ( .A1(n11798), .A2(n11799), .ZN(n11812) );
  AOI22_X1 U11462 ( .A1(n13179), .A2(n16656), .B1(n12842), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10150) );
  NOR2_X2 U11463 ( .A1(n19548), .A2(n19981), .ZN(n19549) );
  NOR2_X2 U11464 ( .A1(n19451), .A2(n19981), .ZN(n14206) );
  NOR2_X2 U11465 ( .A1(n19441), .A2(n19981), .ZN(n14210) );
  AND2_X1 U11466 ( .A1(n12376), .A2(n11808), .ZN(n12378) );
  AOI22_X1 U11467 ( .A1(n13179), .A2(n16656), .B1(n12842), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n9871) );
  NOR2_X2 U11468 ( .A1(n14354), .A2(n19981), .ZN(n14355) );
  AND2_X1 U11469 ( .A1(n11817), .A2(n11811), .ZN(n19365) );
  NAND2_X1 U11470 ( .A1(n18938), .A2(n9929), .ZN(n15971) );
  AND2_X1 U11471 ( .A1(n10670), .A2(n10668), .ZN(n10607) );
  NOR2_X1 U11472 ( .A1(n12496), .A2(n10285), .ZN(n10287) );
  NOR2_X1 U11473 ( .A1(n19152), .A2(n17781), .ZN(n17773) );
  NAND2_X1 U11474 ( .A1(n11765), .A2(n11782), .ZN(n11814) );
  NOR2_X2 U11475 ( .A1(n13118), .A2(n15974), .ZN(n18938) );
  NAND2_X1 U11476 ( .A1(n10351), .A2(n10350), .ZN(n11817) );
  NAND2_X1 U11477 ( .A1(n18119), .A2(n12974), .ZN(n12976) );
  NAND2_X1 U11478 ( .A1(n11809), .A2(n11810), .ZN(n11811) );
  NOR2_X1 U11479 ( .A1(n16813), .A2(n13124), .ZN(n15974) );
  NAND2_X1 U11480 ( .A1(n11771), .A2(n11800), .ZN(n11809) );
  AOI21_X1 U11481 ( .B1(n11783), .B2(n16615), .A(n11785), .ZN(n11794) );
  INV_X1 U11482 ( .A(n10274), .ZN(n12495) );
  OAI21_X1 U11483 ( .B1(n11775), .B2(n12743), .A(n11774), .ZN(n11780) );
  NOR4_X1 U11484 ( .A1(n19152), .A2(n18508), .A3(n16069), .A4(n19149), .ZN(
        n17519) );
  OAI21_X1 U11485 ( .B1(n13985), .B2(n13984), .A(n9930), .ZN(n10274) );
  XNOR2_X1 U11486 ( .A(n12486), .B(n12485), .ZN(n13985) );
  NAND2_X1 U11487 ( .A1(n17533), .A2(n13125), .ZN(n17721) );
  NAND2_X1 U11488 ( .A1(n11776), .A2(n11756), .ZN(n11787) );
  AND3_X1 U11489 ( .A1(n13117), .A2(n13116), .A3(n17683), .ZN(n13125) );
  AND2_X1 U11490 ( .A1(n13807), .A2(n13806), .ZN(n12486) );
  OAI21_X1 U11491 ( .B1(n12698), .B2(n13763), .A(n12471), .ZN(n13807) );
  CLKBUF_X1 U11492 ( .A(n12458), .Z(n15813) );
  OR2_X1 U11493 ( .A1(n11548), .A2(n11449), .ZN(n11544) );
  AND2_X1 U11494 ( .A1(n12488), .A2(n12470), .ZN(n12471) );
  AND2_X1 U11495 ( .A1(n10570), .A2(n10555), .ZN(n11561) );
  AND2_X1 U11497 ( .A1(n11759), .A2(n11758), .ZN(n11789) );
  INV_X1 U11498 ( .A(n11449), .ZN(n10210) );
  AND3_X1 U11499 ( .A1(n10304), .A2(n11881), .A3(n9931), .ZN(n12497) );
  NAND2_X1 U11500 ( .A1(n12743), .A2(n12742), .ZN(n12744) );
  NAND2_X1 U11501 ( .A1(n12743), .A2(n11757), .ZN(n11801) );
  NOR2_X1 U11502 ( .A1(n11921), .A2(n11920), .ZN(n13763) );
  NOR2_X1 U11503 ( .A1(n13626), .A2(n11732), .ZN(n11721) );
  NAND2_X1 U11504 ( .A1(n12148), .A2(n12362), .ZN(n12729) );
  BUF_X1 U11505 ( .A(n10544), .Z(n20550) );
  AND2_X1 U11506 ( .A1(n13621), .A2(n12149), .ZN(n12743) );
  NAND4_X2 U11507 ( .A1(n10541), .A2(n10540), .A3(n10539), .A4(n10538), .ZN(
        n10551) );
  INV_X1 U11508 ( .A(n19152), .ZN(n18511) );
  AND2_X2 U11509 ( .A1(n11730), .A2(n11726), .ZN(n15985) );
  NAND3_X1 U11510 ( .A1(n13071), .A2(n13070), .A3(n13069), .ZN(n17683) );
  CLKBUF_X1 U11511 ( .A(n12149), .Z(n13214) );
  AOI22_X1 U11512 ( .A1(DATAI_23_), .A2(n20498), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20552), .ZN(n21056) );
  OAI21_X1 U11513 ( .B1(n12472), .B2(n19557), .A(n11681), .ZN(n11751) );
  INV_X2 U11514 ( .A(n12227), .ZN(n19552) );
  AND3_X2 U11515 ( .A1(n9891), .A2(n9879), .A3(n10519), .ZN(n14309) );
  AND4_X1 U11516 ( .A1(n10528), .A2(n10527), .A3(n10526), .A4(n10525), .ZN(
        n10540) );
  INV_X2 U11517 ( .A(n16767), .ZN(n16764) );
  AND2_X1 U11518 ( .A1(n12730), .A2(n11741), .ZN(n13621) );
  AND2_X2 U11519 ( .A1(n14211), .A2(n16669), .ZN(n12491) );
  AND2_X1 U11520 ( .A1(n19570), .A2(n16669), .ZN(n12481) );
  NOR2_X1 U11521 ( .A1(n13641), .A2(n12226), .ZN(n11717) );
  NAND2_X1 U11522 ( .A1(n13198), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13197) );
  AND3_X1 U11523 ( .A1(n12730), .A2(n11716), .A3(n19547), .ZN(n11720) );
  OR2_X1 U11524 ( .A1(n10495), .A2(n10494), .ZN(n10547) );
  NAND4_X1 U11525 ( .A1(n12226), .A2(n19547), .A3(n11732), .A4(n11655), .ZN(
        n12734) );
  INV_X1 U11526 ( .A(n11741), .ZN(n12727) );
  NOR2_X2 U11527 ( .A1(n20497), .A2(n20496), .ZN(n20498) );
  INV_X2 U11528 ( .A(U212), .ZN(n16759) );
  NAND2_X1 U11529 ( .A1(n11668), .A2(n11667), .ZN(n11741) );
  NAND2_X1 U11530 ( .A1(n11654), .A2(n11653), .ZN(n12202) );
  AND4_X1 U11531 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10514) );
  AND4_X1 U11532 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n10428) );
  AND4_X1 U11533 ( .A1(n10532), .A2(n10531), .A3(n10530), .A4(n10529), .ZN(
        n10539) );
  AND4_X1 U11534 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10541) );
  AND4_X1 U11535 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10469) );
  AND4_X1 U11536 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10470) );
  AND4_X1 U11537 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n10435), .ZN(
        n10449) );
  AND4_X1 U11538 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10450) );
  AND4_X1 U11539 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10468) );
  AND4_X1 U11540 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10467) );
  BUF_X2 U11541 ( .A(n9924), .Z(n17368) );
  AND4_X1 U11542 ( .A1(n10442), .A2(n10441), .A3(n10440), .A4(n10439), .ZN(
        n10448) );
  AND4_X1 U11543 ( .A1(n10426), .A2(n10425), .A3(n10424), .A4(n10423), .ZN(
        n10427) );
  AND4_X1 U11544 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10513) );
  AND4_X1 U11545 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10519) );
  AND4_X1 U11546 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10538) );
  AND4_X1 U11547 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10447) );
  AND2_X2 U11548 ( .A1(n13591), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13444) );
  INV_X2 U11549 ( .A(n21166), .ZN(n9827) );
  AND4_X1 U11550 ( .A1(n10418), .A2(n10417), .A3(n10416), .A4(n10415), .ZN(
        n10429) );
  INV_X2 U11551 ( .A(n16800), .ZN(U215) );
  INV_X2 U11552 ( .A(n12515), .ZN(n13437) );
  AND2_X2 U11553 ( .A1(n13591), .A2(n16617), .ZN(n13443) );
  NAND2_X2 U11554 ( .A1(n20246), .A2(n20130), .ZN(n20185) );
  BUF_X4 U11555 ( .A(n10476), .Z(n11145) );
  NAND2_X2 U11556 ( .A1(n19140), .A2(n19034), .ZN(n19083) );
  AND2_X1 U11557 ( .A1(n11634), .A2(n11633), .ZN(n11637) );
  CLKBUF_X1 U11558 ( .A(n13708), .Z(n14196) );
  NAND2_X2 U11559 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20246), .ZN(n20186) );
  NAND2_X1 U11560 ( .A1(n10162), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10161) );
  INV_X2 U11561 ( .A(n15920), .ZN(n17456) );
  AND2_X1 U11562 ( .A1(n9886), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9889) );
  NAND2_X1 U11563 ( .A1(n10031), .A2(n10061), .ZN(n12944) );
  INV_X2 U11564 ( .A(n19027), .ZN(n19090) );
  AND4_X1 U11565 ( .A1(n11631), .A2(n11630), .A3(n11629), .A4(n11628), .ZN(
        n11632) );
  CLKBUF_X2 U11566 ( .A(n9863), .Z(n9865) );
  NOR2_X4 U11567 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12190), .ZN(
        n12595) );
  AND2_X2 U11568 ( .A1(n13606), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13438) );
  AND2_X2 U11569 ( .A1(n10405), .A2(n14044), .ZN(n11208) );
  OR2_X1 U11570 ( .A1(n12886), .A2(n17182), .ZN(n9915) );
  OR2_X1 U11571 ( .A1(n12888), .A2(n12887), .ZN(n9917) );
  INV_X1 U11572 ( .A(n10163), .ZN(n10162) );
  NAND3_X1 U11573 ( .A1(n10155), .A2(n10153), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13191) );
  AND2_X1 U11574 ( .A1(n10156), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9886) );
  AND2_X1 U11575 ( .A1(n10395), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10407) );
  NAND2_X1 U11576 ( .A1(n19121), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12888) );
  NAND2_X1 U11577 ( .A1(n13017), .A2(n19108), .ZN(n12880) );
  AND2_X2 U11578 ( .A1(n10577), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10405) );
  OR2_X1 U11579 ( .A1(n18976), .A2(n12886), .ZN(n12916) );
  AND2_X2 U11580 ( .A1(n11855), .A2(n12135), .ZN(n9858) );
  NAND2_X1 U11581 ( .A1(n19121), .A2(n19128), .ZN(n17182) );
  NOR2_X1 U11582 ( .A1(n16548), .A2(n10154), .ZN(n10153) );
  NOR2_X1 U11583 ( .A1(n16508), .A2(n10157), .ZN(n10156) );
  INV_X1 U11584 ( .A(n13188), .ZN(n10155) );
  OR2_X1 U11585 ( .A1(n10164), .A2(n19235), .ZN(n10163) );
  AND2_X2 U11586 ( .A1(n13839), .A2(n14045), .ZN(n10990) );
  NAND2_X2 U11587 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18976) );
  INV_X2 U11588 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19108) );
  INV_X2 U11589 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19128) );
  AND2_X2 U11590 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13839) );
  AND2_X2 U11591 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14045) );
  INV_X1 U11592 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10577) );
  NAND2_X1 U11593 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13188) );
  INV_X1 U11594 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15550) );
  NOR2_X2 U11595 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14044) );
  AND2_X1 U11596 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11602) );
  INV_X1 U11597 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15839) );
  INV_X1 U11598 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11603) );
  INV_X1 U11599 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12135) );
  NAND2_X1 U11600 ( .A1(n18108), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18107) );
  XNOR2_X2 U11601 ( .A(n12867), .B(n12866), .ZN(n16379) );
  NOR2_X2 U11602 ( .A1(n15729), .A2(n15731), .ZN(n15730) );
  NOR2_X2 U11603 ( .A1(n9909), .A2(n12722), .ZN(n12819) );
  NAND2_X1 U11604 ( .A1(n14478), .A2(n11395), .ZN(n9831) );
  NOR2_X1 U11605 ( .A1(n10277), .A2(n10275), .ZN(n9832) );
  CLKBUF_X1 U11606 ( .A(n14132), .Z(n9833) );
  NAND2_X1 U11607 ( .A1(n14478), .A2(n11395), .ZN(n14998) );
  NOR2_X1 U11608 ( .A1(n10277), .A2(n10275), .ZN(n14893) );
  XNOR2_X1 U11609 ( .A(n11325), .B(n11324), .ZN(n14132) );
  NAND2_X2 U11610 ( .A1(n12128), .A2(n12127), .ZN(n13651) );
  OAI21_X2 U11611 ( .B1(n10075), .B2(n15545), .A(n10071), .ZN(n12128) );
  AND2_X1 U11612 ( .A1(n13839), .A2(n14045), .ZN(n9834) );
  AND2_X2 U11613 ( .A1(n13839), .A2(n14045), .ZN(n9835) );
  NAND2_X1 U11614 ( .A1(n19489), .A2(n19502), .ZN(n10076) );
  NOR2_X4 U11615 ( .A1(n18976), .A2(n12880), .ZN(n17478) );
  AND2_X1 U11616 ( .A1(n10405), .A2(n14045), .ZN(n9840) );
  AND2_X1 U11621 ( .A1(n10405), .A2(n14045), .ZN(n11143) );
  NOR2_X4 U11622 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15845) );
  NOR2_X2 U11623 ( .A1(n14361), .A2(n14414), .ZN(n14415) );
  NAND2_X1 U11624 ( .A1(n11615), .A2(n11614), .ZN(n9848) );
  OAI211_X1 U11625 ( .C1(n20628), .C2(n10022), .A(n10020), .B(n10587), .ZN(
        n10681) );
  OR2_X2 U11626 ( .A1(n20628), .A2(n10607), .ZN(n20561) );
  AOI21_X2 U11627 ( .B1(n12123), .B2(n10074), .A(n10073), .ZN(n10071) );
  NAND2_X1 U11628 ( .A1(n12468), .A2(n9848), .ZN(n12698) );
  INV_X1 U11629 ( .A(n17435), .ZN(n9849) );
  BUF_X8 U11630 ( .A(n11208), .Z(n9850) );
  OR2_X1 U11631 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  NAND2_X1 U11632 ( .A1(n11966), .A2(n11965), .ZN(n11996) );
  NAND2_X1 U11633 ( .A1(n11966), .A2(n9884), .ZN(n12049) );
  BUF_X4 U11634 ( .A(n11142), .Z(n9851) );
  BUF_X4 U11635 ( .A(n11142), .Z(n9852) );
  AND2_X2 U11636 ( .A1(n10406), .A2(n14045), .ZN(n11142) );
  NAND2_X1 U11637 ( .A1(n11884), .A2(n11883), .ZN(n11966) );
  NAND2_X2 U11638 ( .A1(n11354), .A2(n11353), .ZN(n16218) );
  INV_X2 U11639 ( .A(n14975), .ZN(n14988) );
  NAND2_X2 U11640 ( .A1(n14998), .A2(n11396), .ZN(n14975) );
  AND2_X2 U11641 ( .A1(n15452), .A2(n10324), .ZN(n15394) );
  NOR2_X2 U11642 ( .A1(n15623), .A2(n15617), .ZN(n15452) );
  MUX2_X2 U11643 ( .A(n10496), .B(n10499), .S(n10547), .Z(n10497) );
  INV_X1 U11644 ( .A(n11449), .ZN(n9854) );
  OR2_X2 U11645 ( .A1(n10482), .A2(n10566), .ZN(n10556) );
  OR2_X1 U11646 ( .A1(n13288), .A2(n19365), .ZN(n11839) );
  OR2_X1 U11647 ( .A1(n13288), .A2(n11828), .ZN(n12007) );
  AND2_X1 U11648 ( .A1(n11855), .A2(n12135), .ZN(n9857) );
  AND2_X1 U11649 ( .A1(n11855), .A2(n12135), .ZN(n11702) );
  OAI21_X2 U11650 ( .B1(n14443), .B2(n11393), .A(n11394), .ZN(n14478) );
  NAND2_X2 U11651 ( .A1(n11385), .A2(n11384), .ZN(n14443) );
  INV_X1 U11652 ( .A(n11886), .ZN(n9859) );
  XNOR2_X2 U11653 ( .A(n11336), .B(n20470), .ZN(n14121) );
  NOR2_X2 U11654 ( .A1(n14932), .A2(n14999), .ZN(n10277) );
  AND2_X1 U11655 ( .A1(n14211), .A2(n16669), .ZN(n9860) );
  AND2_X1 U11656 ( .A1(n14211), .A2(n16669), .ZN(n9861) );
  AND2_X1 U11657 ( .A1(n10401), .A2(n14064), .ZN(n9863) );
  CLKBUF_X1 U11658 ( .A(n9863), .Z(n9864) );
  AND2_X1 U11659 ( .A1(n10401), .A2(n14064), .ZN(n10630) );
  NAND2_X2 U11660 ( .A1(n10207), .A2(n10560), .ZN(n14066) );
  NOR2_X4 U11661 ( .A1(n10498), .A2(n10497), .ZN(n10560) );
  AND2_X1 U11662 ( .A1(n14044), .A2(n14064), .ZN(n9867) );
  AND2_X1 U11663 ( .A1(n14044), .A2(n14064), .ZN(n9868) );
  INV_X2 U11664 ( .A(n9829), .ZN(n9869) );
  AND2_X1 U11665 ( .A1(n10406), .A2(n14044), .ZN(n10887) );
  NOR2_X4 U11666 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14064) );
  INV_X1 U11670 ( .A(n9824), .ZN(n9875) );
  INV_X1 U11671 ( .A(n9824), .ZN(n9876) );
  INV_X1 U11672 ( .A(n9824), .ZN(n9877) );
  NAND2_X1 U11673 ( .A1(n10203), .A2(n10202), .ZN(n10201) );
  NOR2_X1 U11674 ( .A1(n14309), .A2(n11427), .ZN(n10202) );
  NAND2_X1 U11675 ( .A1(n10544), .A2(n10602), .ZN(n10482) );
  NOR2_X1 U11676 ( .A1(n13913), .A2(n14360), .ZN(n13271) );
  AOI22_X1 U11677 ( .A1(n11556), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n10604), 
        .B2(n10568), .ZN(n10561) );
  INV_X1 U11678 ( .A(n12362), .ZN(n12149) );
  AND2_X1 U11679 ( .A1(n16656), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13287) );
  NAND2_X1 U11680 ( .A1(n21487), .A2(n16615), .ZN(n12138) );
  AND2_X1 U11681 ( .A1(n12204), .A2(n12202), .ZN(n11729) );
  OR2_X1 U11682 ( .A1(n10687), .A2(n11378), .ZN(n10651) );
  NAND2_X1 U11683 ( .A1(n10193), .A2(n9953), .ZN(n14592) );
  NOR2_X1 U11684 ( .A1(n10196), .A2(n11137), .ZN(n10195) );
  INV_X1 U11685 ( .A(n14608), .ZN(n10196) );
  AND2_X1 U11686 ( .A1(n20980), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11229) );
  NAND2_X1 U11687 ( .A1(n10114), .A2(n14761), .ZN(n10113) );
  INV_X1 U11688 ( .A(n14508), .ZN(n10114) );
  INV_X1 U11689 ( .A(n11544), .ZN(n11531) );
  OR2_X1 U11690 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20494), .ZN(
        n11239) );
  AND2_X1 U11691 ( .A1(n9945), .A2(n10340), .ZN(n10339) );
  INV_X1 U11692 ( .A(n15290), .ZN(n10340) );
  NAND2_X1 U11693 ( .A1(n15427), .A2(n15428), .ZN(n12777) );
  AND2_X1 U11694 ( .A1(n10256), .A2(n10258), .ZN(n10255) );
  NAND2_X1 U11695 ( .A1(n10257), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10256) );
  NOR2_X1 U11696 ( .A1(n10257), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10253) );
  OR2_X1 U11697 ( .A1(n15163), .A2(n12320), .ZN(n12328) );
  NAND2_X1 U11698 ( .A1(n10011), .A2(n10010), .ZN(n10080) );
  INV_X1 U11699 ( .A(n13653), .ZN(n10010) );
  INV_X1 U11700 ( .A(n13655), .ZN(n10011) );
  NAND2_X1 U11701 ( .A1(n12102), .A2(n12101), .ZN(n12124) );
  NAND2_X1 U11702 ( .A1(n14398), .A2(n12094), .ZN(n12098) );
  NAND2_X1 U11703 ( .A1(n15180), .A2(n10286), .ZN(n10285) );
  INV_X1 U11704 ( .A(n14281), .ZN(n10286) );
  NAND2_X1 U11705 ( .A1(n11967), .A2(n11968), .ZN(n10323) );
  INV_X1 U11706 ( .A(n11965), .ZN(n11968) );
  NAND2_X1 U11707 ( .A1(n11780), .A2(n11779), .ZN(n11810) );
  NAND2_X1 U11708 ( .A1(n13269), .A2(n13271), .ZN(n13285) );
  NAND2_X1 U11709 ( .A1(n11848), .A2(n14338), .ZN(n10315) );
  INV_X1 U11710 ( .A(n17182), .ZN(n10031) );
  AND2_X1 U11711 ( .A1(n17948), .A2(n10143), .ZN(n10142) );
  NOR2_X1 U11712 ( .A1(n10144), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10143) );
  INV_X1 U11713 ( .A(n9947), .ZN(n10144) );
  NAND2_X1 U11714 ( .A1(n17996), .A2(n13250), .ZN(n12993) );
  NAND2_X1 U11715 ( .A1(n12979), .A2(n18089), .ZN(n12982) );
  NAND2_X1 U11716 ( .A1(n18095), .A2(n18096), .ZN(n18094) );
  NAND2_X1 U11717 ( .A1(n17668), .A2(n12969), .ZN(n12955) );
  OR2_X1 U11718 ( .A1(n14066), .A2(n11429), .ZN(n13850) );
  NOR2_X1 U11719 ( .A1(n16010), .A2(n20251), .ZN(n14120) );
  AND2_X1 U11720 ( .A1(n10520), .A2(n13974), .ZN(n10207) );
  INV_X1 U11721 ( .A(n12783), .ZN(n10301) );
  NAND2_X1 U11722 ( .A1(n10290), .A2(n15168), .ZN(n10289) );
  INV_X1 U11723 ( .A(n10291), .ZN(n10290) );
  NOR3_X1 U11724 ( .A1(n9893), .A2(n10337), .A3(n10336), .ZN(n15205) );
  NOR2_X1 U11725 ( .A1(n9893), .A2(n10336), .ZN(n15137) );
  INV_X1 U11726 ( .A(n10008), .ZN(n10007) );
  OAI21_X1 U11727 ( .B1(n10260), .B2(n9960), .A(n12337), .ZN(n10008) );
  AND2_X1 U11728 ( .A1(n12217), .A2(n16665), .ZN(n12755) );
  AOI21_X1 U11729 ( .B1(n15836), .B2(n13287), .A(n13279), .ZN(n13749) );
  NAND2_X1 U11730 ( .A1(n12163), .A2(n12162), .ZN(n16642) );
  INV_X1 U11731 ( .A(n16811), .ZN(n18941) );
  NAND2_X1 U11732 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n13162), .ZN(
        n16670) );
  INV_X1 U11733 ( .A(n16670), .ZN(n16688) );
  NAND2_X1 U11734 ( .A1(n10065), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10064) );
  INV_X1 U11735 ( .A(n16054), .ZN(n10065) );
  INV_X1 U11736 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20233) );
  NOR2_X1 U11737 ( .A1(n12894), .A2(n12893), .ZN(n17649) );
  NAND2_X1 U11738 ( .A1(n14202), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10225) );
  NAND2_X1 U11739 ( .A1(n19708), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10226) );
  NAND2_X1 U11740 ( .A1(n12734), .A2(n11681), .ZN(n11682) );
  NAND2_X1 U11741 ( .A1(n20022), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12013) );
  NOR2_X1 U11742 ( .A1(n12459), .A2(n16656), .ZN(n11752) );
  NAND2_X1 U11743 ( .A1(n12152), .A2(n12134), .ZN(n12147) );
  XNOR2_X1 U11744 ( .A(n9848), .B(n11723), .ZN(n12200) );
  AOI22_X1 U11745 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9858), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11648) );
  NAND2_X1 U11746 ( .A1(n14975), .A2(n16262), .ZN(n10278) );
  OR2_X1 U11747 ( .A1(n10687), .A2(n11390), .ZN(n11387) );
  INV_X1 U11748 ( .A(n10687), .ZN(n10191) );
  INV_X1 U11749 ( .A(n10402), .ZN(n10403) );
  NAND2_X1 U11750 ( .A1(n14309), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10686) );
  NAND2_X1 U11751 ( .A1(n15985), .A2(n16637), .ZN(n12196) );
  INV_X1 U11752 ( .A(n11741), .ZN(n11716) );
  NOR2_X1 U11753 ( .A1(n12955), .A2(n13136), .ZN(n12954) );
  NOR2_X1 U11754 ( .A1(n17655), .A2(n12975), .ZN(n12979) );
  AOI21_X1 U11755 ( .B1(n18969), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13019), .ZN(n13029) );
  AND2_X1 U11756 ( .A1(n13126), .A2(n13018), .ZN(n13019) );
  INV_X1 U11757 ( .A(n14043), .ZN(n10557) );
  NAND2_X1 U11758 ( .A1(n15125), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11199) );
  NOR2_X1 U11759 ( .A1(n10211), .A2(n14685), .ZN(n10051) );
  NAND2_X1 U11760 ( .A1(n10212), .A2(n10378), .ZN(n10211) );
  INV_X1 U11761 ( .A(n10214), .ZN(n10212) );
  NOR2_X1 U11762 ( .A1(n10119), .A2(n10118), .ZN(n10117) );
  INV_X1 U11763 ( .A(n14600), .ZN(n10118) );
  INV_X1 U11764 ( .A(n10120), .ZN(n10119) );
  NOR2_X1 U11765 ( .A1(n14978), .A2(n11400), .ZN(n10283) );
  INV_X1 U11766 ( .A(n14461), .ZN(n10102) );
  NOR2_X1 U11767 ( .A1(n14418), .A2(n10104), .ZN(n10103) );
  INV_X1 U11768 ( .A(n14364), .ZN(n10104) );
  OR2_X1 U11769 ( .A1(n10640), .A2(n10639), .ZN(n11378) );
  INV_X1 U11770 ( .A(n11362), .ZN(n10027) );
  NOR2_X1 U11771 ( .A1(n14085), .A2(n14023), .ZN(n10111) );
  NAND2_X1 U11772 ( .A1(n10543), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10687) );
  NAND4_X2 U11773 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        n10602) );
  NAND2_X1 U11774 ( .A1(n10687), .A2(n10686), .ZN(n11275) );
  AND2_X1 U11775 ( .A1(n20517), .A2(n11248), .ZN(n11422) );
  AOI21_X1 U11776 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20209), .A(
        n12141), .ZN(n12143) );
  NOR2_X1 U11777 ( .A1(n12140), .A2(n12144), .ZN(n12141) );
  INV_X1 U11778 ( .A(n11880), .ZN(n10304) );
  NOR2_X1 U11779 ( .A1(n12350), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12359) );
  INV_X1 U11780 ( .A(n12308), .ZN(n10312) );
  NOR2_X1 U11781 ( .A1(n10307), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10306) );
  INV_X1 U11782 ( .A(n12259), .ZN(n10307) );
  AND2_X1 U11783 ( .A1(n12258), .A2(n12257), .ZN(n12262) );
  AND2_X1 U11784 ( .A1(n9859), .A2(n14199), .ZN(n13220) );
  NOR2_X1 U11785 ( .A1(n12734), .A2(n16656), .ZN(n11757) );
  AND2_X1 U11786 ( .A1(n13526), .A2(n9981), .ZN(n13527) );
  INV_X1 U11787 ( .A(n15343), .ZN(n10298) );
  INV_X1 U11788 ( .A(n13913), .ZN(n13546) );
  INV_X1 U11789 ( .A(n12612), .ZN(n13432) );
  NAND2_X1 U11790 ( .A1(n10295), .A2(n13658), .ZN(n10294) );
  INV_X1 U11791 ( .A(n14293), .ZN(n10295) );
  AND2_X1 U11792 ( .A1(n11727), .A2(n11852), .ZN(n12737) );
  NAND2_X1 U11793 ( .A1(n11723), .A2(n12202), .ZN(n13641) );
  OR3_X1 U11794 ( .A1(n15225), .A2(n15236), .A3(n10338), .ZN(n10336) );
  INV_X1 U11795 ( .A(n14155), .ZN(n10347) );
  NOR2_X1 U11796 ( .A1(n15397), .A2(n12776), .ZN(n10229) );
  NOR2_X1 U11797 ( .A1(n15141), .A2(n12320), .ZN(n15408) );
  NOR2_X1 U11798 ( .A1(n16401), .A2(n12320), .ZN(n15405) );
  OR2_X1 U11799 ( .A1(n16000), .A2(n12320), .ZN(n12336) );
  NAND2_X1 U11800 ( .A1(n9880), .A2(n15526), .ZN(n10081) );
  INV_X1 U11801 ( .A(n15527), .ZN(n10083) );
  INV_X1 U11802 ( .A(n15463), .ZN(n10088) );
  INV_X1 U11803 ( .A(n14456), .ZN(n10341) );
  NOR2_X1 U11804 ( .A1(n15985), .A2(n14199), .ZN(n11737) );
  AOI21_X1 U11805 ( .B1(n11725), .B2(n19557), .A(n11733), .ZN(n11734) );
  AND3_X1 U11806 ( .A1(n19547), .A2(n11741), .A3(n11723), .ZN(n11730) );
  INV_X1 U11807 ( .A(n11903), .ZN(n19671) );
  AOI22_X1 U11809 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9857), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U11810 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11633) );
  NOR2_X1 U11811 ( .A1(n10042), .A2(n10039), .ZN(n10038) );
  INV_X1 U11812 ( .A(n13077), .ZN(n10042) );
  INV_X1 U11813 ( .A(n10135), .ZN(n10134) );
  OAI21_X1 U11814 ( .B1(n12916), .B2(n17518), .A(n10136), .ZN(n10135) );
  NAND2_X1 U11815 ( .A1(n12922), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10136) );
  NAND2_X1 U11816 ( .A1(n12915), .A2(n12920), .ZN(n10130) );
  INV_X1 U11817 ( .A(n12918), .ZN(n10131) );
  NAND2_X1 U11818 ( .A1(n12923), .A2(n12919), .ZN(n10137) );
  INV_X1 U11819 ( .A(n10390), .ZN(n17470) );
  INV_X1 U11820 ( .A(n13164), .ZN(n13162) );
  XNOR2_X1 U11821 ( .A(n17659), .B(n10066), .ZN(n12973) );
  INV_X1 U11822 ( .A(n12954), .ZN(n10066) );
  NOR2_X1 U11823 ( .A1(n17817), .A2(n12998), .ZN(n13000) );
  NAND2_X1 U11824 ( .A1(n18078), .A2(n10138), .ZN(n12987) );
  NOR2_X1 U11825 ( .A1(n10139), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10138) );
  INV_X1 U11826 ( .A(n12985), .ZN(n10139) );
  NOR2_X1 U11827 ( .A1(n12983), .A2(n10059), .ZN(n10058) );
  INV_X1 U11828 ( .A(n12981), .ZN(n10059) );
  NOR2_X1 U11829 ( .A1(n12984), .A2(n10056), .ZN(n10055) );
  INV_X1 U11830 ( .A(n18096), .ZN(n10056) );
  NAND2_X1 U11831 ( .A1(n18107), .A2(n12978), .ZN(n18095) );
  XNOR2_X1 U11832 ( .A(n12969), .B(n17668), .ZN(n12970) );
  AOI21_X1 U11833 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18502), .A(
        n13025), .ZN(n13128) );
  NAND2_X1 U11834 ( .A1(n14676), .A2(n16076), .ZN(n20324) );
  NOR3_X1 U11835 ( .A1(n14521), .A2(n10115), .A3(n14508), .ZN(n14762) );
  NAND2_X1 U11836 ( .A1(n14836), .A2(n10204), .ZN(n14036) );
  NOR2_X1 U11837 ( .A1(n10224), .A2(n10222), .ZN(n10221) );
  INV_X1 U11838 ( .A(n10223), .ZN(n10222) );
  OR2_X1 U11839 ( .A1(n11201), .A2(n14873), .ZN(n11202) );
  NAND2_X1 U11840 ( .A1(n11160), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11201) );
  NAND2_X1 U11841 ( .A1(n11076), .A2(n11075), .ZN(n14647) );
  INV_X1 U11842 ( .A(n14661), .ZN(n11075) );
  NAND2_X1 U11843 ( .A1(n11070), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11111) );
  OR2_X1 U11844 ( .A1(n16172), .A2(n10094), .ZN(n10093) );
  AND2_X1 U11845 ( .A1(n10726), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10752) );
  AOI21_X1 U11846 ( .B1(n10660), .B2(n10912), .A(n10200), .ZN(n10199) );
  INV_X1 U11847 ( .A(n10680), .ZN(n10200) );
  NOR2_X1 U11848 ( .A1(n14999), .A2(n15029), .ZN(n10090) );
  INV_X1 U11849 ( .A(n14880), .ZN(n10091) );
  NAND2_X1 U11850 ( .A1(n14923), .A2(n15076), .ZN(n14902) );
  OR3_X1 U11851 ( .A1(n10115), .A2(n10113), .A3(n14756), .ZN(n10112) );
  NAND2_X1 U11852 ( .A1(n14497), .A2(n14496), .ZN(n14519) );
  AND2_X1 U11853 ( .A1(n11467), .A2(n11466), .ZN(n14164) );
  NAND2_X1 U11854 ( .A1(n21189), .A2(n20500), .ZN(n14124) );
  NAND2_X1 U11855 ( .A1(n10203), .A2(n9854), .ZN(n10206) );
  AND2_X1 U11856 ( .A1(n11440), .A2(n11439), .ZN(n11573) );
  INV_X1 U11857 ( .A(n13834), .ZN(n10205) );
  XNOR2_X1 U11858 ( .A(n10654), .B(n10652), .ZN(n10662) );
  XNOR2_X1 U11859 ( .A(n10019), .B(n10656), .ZN(n15119) );
  NAND2_X1 U11860 ( .A1(n10097), .A2(n10700), .ZN(n10737) );
  NAND2_X1 U11861 ( .A1(n20502), .A2(n10701), .ZN(n10054) );
  NOR2_X1 U11862 ( .A1(n20523), .A2(n10546), .ZN(n14043) );
  INV_X1 U11863 ( .A(n10589), .ZN(n10022) );
  NAND2_X1 U11864 ( .A1(n13858), .A2(n13857), .ZN(n16014) );
  AND2_X1 U11865 ( .A1(n21012), .A2(n20505), .ZN(n20856) );
  INV_X1 U11866 ( .A(n21195), .ZN(n20890) );
  AND2_X1 U11867 ( .A1(n9870), .A2(n21207), .ZN(n20889) );
  NAND2_X1 U11868 ( .A1(n20500), .A2(n20499), .ZN(n20670) );
  AND2_X1 U11869 ( .A1(n11238), .A2(n11239), .ZN(n11251) );
  OR2_X1 U11870 ( .A1(n11240), .A2(n11237), .ZN(n11238) );
  NAND2_X1 U11871 ( .A1(n11289), .A2(n11422), .ZN(n11255) );
  AND2_X1 U11872 ( .A1(n16040), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16049) );
  XNOR2_X1 U11873 ( .A(n12837), .B(n12785), .ZN(n13231) );
  NAND2_X1 U11874 ( .A1(n16418), .A2(n9877), .ZN(n16407) );
  OR2_X1 U11875 ( .A1(n12309), .A2(n10310), .ZN(n12315) );
  OR2_X1 U11876 ( .A1(n16638), .A2(n13210), .ZN(n13219) );
  NAND2_X1 U11877 ( .A1(n12247), .A2(n12246), .ZN(n12252) );
  NAND2_X1 U11878 ( .A1(n10359), .A2(n13304), .ZN(n10358) );
  INV_X1 U11879 ( .A(n10360), .ZN(n10359) );
  NAND2_X1 U11880 ( .A1(n10293), .A2(n10292), .ZN(n10291) );
  INV_X1 U11881 ( .A(n16578), .ZN(n10292) );
  INV_X1 U11882 ( .A(n10294), .ZN(n10293) );
  INV_X1 U11883 ( .A(n13708), .ZN(n14194) );
  AND2_X1 U11884 ( .A1(n13187), .A2(n9889), .ZN(n13198) );
  INV_X1 U11885 ( .A(n12123), .ZN(n10075) );
  NOR2_X1 U11886 ( .A1(n13191), .A2(n15550), .ZN(n13193) );
  NAND2_X1 U11887 ( .A1(n13193), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13192) );
  XNOR2_X1 U11888 ( .A(n12125), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16536) );
  NOR2_X1 U11889 ( .A1(n13918), .A2(n10329), .ZN(n13965) );
  NAND2_X1 U11890 ( .A1(n9943), .A2(n10330), .ZN(n10329) );
  INV_X1 U11891 ( .A(n9982), .ZN(n10330) );
  NAND2_X1 U11892 ( .A1(n10241), .A2(n10238), .ZN(n19492) );
  INV_X1 U11893 ( .A(n10239), .ZN(n10238) );
  OAI21_X1 U11894 ( .B1(n10246), .B2(n10240), .A(n10245), .ZN(n10239) );
  INV_X1 U11895 ( .A(n10382), .ZN(n10236) );
  INV_X1 U11896 ( .A(n15455), .ZN(n10252) );
  NAND2_X1 U11897 ( .A1(n10009), .A2(n9927), .ZN(n10250) );
  OR3_X1 U11898 ( .A1(n10344), .A2(n10343), .A3(n15246), .ZN(n10342) );
  INV_X1 U11899 ( .A(n10261), .ZN(n10260) );
  OAI21_X1 U11900 ( .B1(n12331), .B2(n10262), .A(n12330), .ZN(n10261) );
  NAND2_X1 U11901 ( .A1(n10265), .A2(n10267), .ZN(n10262) );
  NOR2_X1 U11902 ( .A1(n12331), .A2(n10264), .ZN(n10263) );
  INV_X1 U11903 ( .A(n10265), .ZN(n10264) );
  OR2_X1 U11904 ( .A1(n19223), .A2(n12326), .ZN(n15674) );
  NAND2_X1 U11905 ( .A1(n10087), .A2(n15504), .ZN(n10086) );
  NAND2_X1 U11906 ( .A1(n10088), .A2(n15521), .ZN(n10087) );
  NAND2_X1 U11907 ( .A1(n15522), .A2(n10088), .ZN(n10017) );
  AND2_X1 U11908 ( .A1(n12703), .A2(n12702), .ZN(n15373) );
  NOR2_X1 U11909 ( .A1(n15775), .A2(n10272), .ZN(n10271) );
  INV_X1 U11910 ( .A(n16512), .ZN(n10272) );
  NAND2_X1 U11911 ( .A1(n12256), .A2(n9925), .ZN(n10012) );
  AND3_X1 U11912 ( .A1(n12505), .A2(n12504), .A3(n12503), .ZN(n14281) );
  CLKBUF_X1 U11913 ( .A(n12462), .Z(n12463) );
  OAI21_X1 U11914 ( .B1(n12233), .B2(n12787), .A(n15183), .ZN(n10247) );
  NAND2_X1 U11915 ( .A1(n13270), .A2(n13287), .ZN(n13275) );
  AND2_X1 U11916 ( .A1(n20202), .A2(n20228), .ZN(n19675) );
  NAND2_X1 U11917 ( .A1(n20202), .A2(n19447), .ZN(n19780) );
  NAND2_X1 U11918 ( .A1(n19677), .A2(n20221), .ZN(n19779) );
  NOR2_X1 U11919 ( .A1(n19677), .A2(n19676), .ZN(n20199) );
  AND2_X1 U11920 ( .A1(n19677), .A2(n19676), .ZN(n19986) );
  NOR2_X1 U11921 ( .A1(n20202), .A2(n20228), .ZN(n19987) );
  OAI21_X2 U11922 ( .B1(n16660), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12805), 
        .ZN(n20020) );
  INV_X1 U11923 ( .A(n20020), .ZN(n19981) );
  INV_X1 U11924 ( .A(n17721), .ZN(n13118) );
  NOR2_X1 U11925 ( .A1(n16869), .A2(n16870), .ZN(n16868) );
  INV_X2 U11926 ( .A(n13062), .ZN(n17433) );
  NAND2_X1 U11927 ( .A1(n12930), .A2(n12929), .ZN(n10123) );
  NAND2_X1 U11928 ( .A1(n12931), .A2(n12928), .ZN(n10127) );
  AOI22_X1 U11929 ( .A1(n15978), .A2(n15979), .B1(n15873), .B2(n15872), .ZN(
        n16069) );
  AOI21_X1 U11930 ( .B1(n18939), .B2(n9919), .A(n15976), .ZN(n16071) );
  INV_X1 U11931 ( .A(n17674), .ZN(n16072) );
  AOI211_X1 U11932 ( .C1(n17458), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n13068), .B(n13067), .ZN(n13069) );
  NOR2_X1 U11933 ( .A1(n18017), .A2(n16968), .ZN(n17989) );
  AOI21_X1 U11934 ( .B1(n18446), .B2(n18128), .A(n12972), .ZN(n18118) );
  NAND2_X1 U11935 ( .A1(n10141), .A2(n10140), .ZN(n17852) );
  NAND2_X1 U11936 ( .A1(n12994), .A2(n18068), .ZN(n10140) );
  AND2_X1 U11937 ( .A1(n10142), .A2(n10146), .ZN(n17932) );
  OAI21_X1 U11938 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n12990), .A(
        n18030), .ZN(n17948) );
  NAND2_X1 U11939 ( .A1(n18078), .A2(n12985), .ZN(n12986) );
  OR2_X1 U11940 ( .A1(n18067), .A2(n18068), .ZN(n10069) );
  XNOR2_X1 U11941 ( .A(n12976), .B(n10147), .ZN(n18108) );
  INV_X1 U11942 ( .A(n12977), .ZN(n10147) );
  OR2_X1 U11943 ( .A1(n13815), .A2(n20251), .ZN(n14549) );
  NOR2_X1 U11944 ( .A1(n10551), .A2(n20501), .ZN(n14306) );
  INV_X1 U11945 ( .A(n20345), .ZN(n20301) );
  AOI21_X1 U11946 ( .B1(n16189), .B2(n14900), .A(n14899), .ZN(n10046) );
  INV_X1 U11947 ( .A(n20432), .ZN(n16209) );
  CLKBUF_X1 U11948 ( .A(n15119), .Z(n15120) );
  NOR2_X1 U11949 ( .A1(n20931), .A2(n16010), .ZN(n21188) );
  INV_X1 U11950 ( .A(n20800), .ZN(n20821) );
  INV_X1 U11951 ( .A(n19343), .ZN(n19364) );
  AND2_X1 U11952 ( .A1(n12602), .A2(n12601), .ZN(n14152) );
  CLKBUF_X1 U11953 ( .A(n13968), .Z(n13969) );
  INV_X1 U11954 ( .A(n15289), .ZN(n15294) );
  NAND2_X1 U11955 ( .A1(n13920), .A2(n19570), .ZN(n15289) );
  INV_X1 U11956 ( .A(n20228), .ZN(n19447) );
  INV_X1 U11957 ( .A(n11811), .ZN(n11815) );
  NAND2_X1 U11958 ( .A1(n12755), .A2(n12461), .ZN(n19534) );
  INV_X1 U11959 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20209) );
  NAND2_X1 U11960 ( .A1(n19365), .A2(n13287), .ZN(n13281) );
  NAND2_X1 U11961 ( .A1(n19008), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19149) );
  OR2_X1 U11962 ( .A1(n16868), .A2(n17065), .ZN(n10188) );
  NAND2_X1 U11963 ( .A1(n10186), .A2(n10185), .ZN(n10184) );
  NAND2_X1 U11964 ( .A1(n16854), .A2(n16853), .ZN(n10185) );
  INV_X1 U11965 ( .A(n16852), .ZN(n10186) );
  NAND2_X1 U11966 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16688), .ZN(
        n13161) );
  NAND2_X1 U11967 ( .A1(n17197), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17184) );
  INV_X1 U11968 ( .A(n17183), .ZN(n17197) );
  NAND4_X1 U11969 ( .A1(n16833), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n18511), 
        .A4(n16832), .ZN(n17194) );
  NOR2_X2 U11970 ( .A1(n17522), .A2(n17612), .ZN(n17523) );
  INV_X1 U11971 ( .A(n17544), .ZN(n17539) );
  INV_X1 U11972 ( .A(n18422), .ZN(n18489) );
  NAND2_X1 U11973 ( .A1(n11885), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U11974 ( .A1(n19775), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11891) );
  NOR2_X1 U11975 ( .A1(n19911), .A2(n11819), .ZN(n11822) );
  AND4_X1 U11976 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12069) );
  OAI21_X1 U11977 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13017), .A(
        n13020), .ZN(n13021) );
  OR2_X1 U11978 ( .A1(n13028), .A2(n13029), .ZN(n13020) );
  NOR2_X1 U11979 ( .A1(n9974), .A2(n14648), .ZN(n10194) );
  NAND3_X1 U11980 ( .A1(n10097), .A2(n10700), .A3(n10738), .ZN(n10750) );
  OR2_X1 U11981 ( .A1(n10768), .A2(n10767), .ZN(n11376) );
  OR2_X1 U11982 ( .A1(n10723), .A2(n10722), .ZN(n11365) );
  INV_X1 U11983 ( .A(n13771), .ZN(n11562) );
  OR2_X1 U11984 ( .A1(n10618), .A2(n10617), .ZN(n11328) );
  NOR2_X1 U11985 ( .A1(n10542), .A2(n10548), .ZN(n10496) );
  OR2_X1 U11986 ( .A1(n10697), .A2(n10696), .ZN(n11347) );
  NAND2_X1 U11987 ( .A1(n12139), .A2(n12138), .ZN(n12145) );
  XNOR2_X1 U11988 ( .A(n16617), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12144) );
  NOR2_X1 U11989 ( .A1(n12298), .A2(n10309), .ZN(n10308) );
  INV_X1 U11990 ( .A(n12279), .ZN(n10309) );
  OR2_X1 U11991 ( .A1(n12151), .A2(n12150), .ZN(n12152) );
  NOR2_X1 U11992 ( .A1(n16615), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13409) );
  NAND2_X1 U11993 ( .A1(n11882), .A2(n11852), .ZN(n11883) );
  OAI21_X1 U11994 ( .B1(n11854), .B2(n11853), .A(n14211), .ZN(n11884) );
  NAND2_X1 U11995 ( .A1(n11745), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11746) );
  NAND3_X1 U11996 ( .A1(n11751), .A2(n11750), .A3(n12729), .ZN(n12458) );
  CLKBUF_X1 U11997 ( .A(n12200), .Z(n12201) );
  AND2_X1 U11998 ( .A1(n12174), .A2(n12175), .ZN(n12182) );
  NAND2_X1 U11999 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10040) );
  INV_X1 U12000 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10041) );
  INV_X1 U12001 ( .A(n12885), .ZN(n10062) );
  NAND2_X1 U12002 ( .A1(n19128), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12885) );
  NAND2_X1 U12003 ( .A1(n10061), .A2(n10062), .ZN(n10390) );
  NOR2_X1 U12004 ( .A1(n14581), .A2(n14595), .ZN(n10223) );
  NAND2_X1 U12005 ( .A1(n14753), .A2(n10215), .ZN(n10214) );
  INV_X1 U12006 ( .A(n14759), .ZN(n10215) );
  AND2_X1 U12007 ( .A1(n10216), .A2(n14459), .ZN(n10052) );
  AND2_X1 U12008 ( .A1(n10881), .A2(n10217), .ZN(n10216) );
  OR2_X1 U12009 ( .A1(n14483), .A2(n14491), .ZN(n10217) );
  NOR2_X1 U12010 ( .A1(n10832), .A2(n20277), .ZN(n10836) );
  XNOR2_X1 U12011 ( .A(n11389), .B(n10779), .ZN(n11373) );
  NAND2_X1 U12012 ( .A1(n10542), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10912) );
  AND2_X1 U12013 ( .A1(n10204), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10729) );
  NOR2_X1 U12014 ( .A1(n14609), .A2(n10121), .ZN(n10120) );
  INV_X1 U12015 ( .A(n14622), .ZN(n10121) );
  INV_X1 U12016 ( .A(n10281), .ZN(n10280) );
  NAND2_X1 U12017 ( .A1(n14121), .A2(n14122), .ZN(n11338) );
  NAND2_X1 U12018 ( .A1(n10210), .A2(n11525), .ZN(n11539) );
  NAND2_X1 U12019 ( .A1(n10646), .A2(n10645), .ZN(n10676) );
  INV_X1 U12020 ( .A(n11328), .ZN(n10648) );
  NAND2_X1 U12021 ( .A1(n10603), .A2(n10191), .ZN(n10190) );
  INV_X1 U12022 ( .A(n10701), .ZN(n10097) );
  NAND2_X1 U12023 ( .A1(n10656), .A2(n10019), .ZN(n10701) );
  NOR2_X1 U12024 ( .A1(n10546), .A2(n20501), .ZN(n10208) );
  AOI21_X1 U12025 ( .B1(n10581), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10582), .ZN(n10590) );
  NOR2_X1 U12026 ( .A1(n10404), .A2(n10403), .ZN(n10410) );
  INV_X1 U12027 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20922) );
  NAND2_X1 U12028 ( .A1(n11962), .A2(n11961), .ZN(n12170) );
  NOR2_X1 U12029 ( .A1(n12774), .A2(n12773), .ZN(n10302) );
  NAND2_X1 U12030 ( .A1(n12836), .A2(n12360), .ZN(n12774) );
  NOR2_X1 U12031 ( .A1(n12338), .A2(n10314), .ZN(n10313) );
  NAND2_X1 U12032 ( .A1(n12333), .A2(n9985), .ZN(n10314) );
  OR2_X1 U12033 ( .A1(n12309), .A2(n12308), .ZN(n12311) );
  NAND2_X1 U12034 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U12035 ( .A1(n12280), .A2(n10308), .ZN(n12301) );
  NAND2_X1 U12036 ( .A1(n12227), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n12224) );
  OR2_X1 U12037 ( .A1(n11860), .A2(n16617), .ZN(n13371) );
  OR2_X1 U12038 ( .A1(n13407), .A2(n16617), .ZN(n12515) );
  OR2_X1 U12039 ( .A1(n13408), .A2(n16617), .ZN(n13375) );
  INV_X1 U12040 ( .A(n11860), .ZN(n13607) );
  INV_X1 U12041 ( .A(n13408), .ZN(n13609) );
  NAND2_X1 U12042 ( .A1(n13503), .A2(n13498), .ZN(n13504) );
  INV_X1 U12043 ( .A(n15335), .ZN(n10297) );
  AND2_X1 U12044 ( .A1(n10373), .A2(n13349), .ZN(n10372) );
  NOR2_X1 U12045 ( .A1(n14451), .A2(n10374), .ZN(n10373) );
  INV_X1 U12046 ( .A(n14387), .ZN(n10374) );
  NOR2_X1 U12047 ( .A1(n16400), .A2(n10159), .ZN(n10158) );
  NOR2_X1 U12048 ( .A1(n19196), .A2(n10152), .ZN(n10151) );
  INV_X1 U12049 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10152) );
  INV_X1 U12050 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10157) );
  INV_X1 U12051 ( .A(n15546), .ZN(n10074) );
  INV_X1 U12052 ( .A(n16536), .ZN(n10073) );
  INV_X1 U12053 ( .A(n12124), .ZN(n12126) );
  INV_X1 U12054 ( .A(n13936), .ZN(n10331) );
  AND2_X1 U12055 ( .A1(n10334), .A2(n13904), .ZN(n10333) );
  INV_X1 U12056 ( .A(n13885), .ZN(n10334) );
  INV_X1 U12057 ( .A(n13918), .ZN(n10332) );
  NOR2_X1 U12058 ( .A1(n12245), .A2(n16611), .ZN(n10246) );
  NAND2_X1 U12059 ( .A1(n12245), .A2(n16611), .ZN(n10245) );
  NAND2_X1 U12060 ( .A1(n15183), .A2(n12787), .ZN(n10240) );
  NOR2_X1 U12061 ( .A1(n10246), .A2(n10243), .ZN(n10242) );
  INV_X1 U12062 ( .A(n15183), .ZN(n10243) );
  INV_X1 U12063 ( .A(n12170), .ZN(n12489) );
  OR2_X1 U12064 ( .A1(n16413), .A2(n12320), .ZN(n12355) );
  NOR2_X1 U12065 ( .A1(n15596), .A2(n21537), .ZN(n10327) );
  INV_X1 U12066 ( .A(n15255), .ZN(n10343) );
  NAND2_X1 U12067 ( .A1(n10346), .A2(n10345), .ZN(n10344) );
  INV_X1 U12068 ( .A(n15270), .ZN(n10345) );
  NOR2_X1 U12069 ( .A1(n10322), .A2(n15655), .ZN(n10320) );
  NAND2_X1 U12070 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10322) );
  INV_X1 U12071 ( .A(n12278), .ZN(n10269) );
  AOI21_X1 U12072 ( .B1(n10268), .B2(n10266), .A(n9977), .ZN(n10265) );
  INV_X1 U12073 ( .A(n10271), .ZN(n10266) );
  AND4_X1 U12074 ( .A1(n12074), .A2(n12073), .A3(n12072), .A4(n12071), .ZN(
        n12090) );
  NOR2_X1 U12075 ( .A1(n12097), .A2(n14397), .ZN(n10319) );
  INV_X1 U12076 ( .A(n19350), .ZN(n10014) );
  AND2_X1 U12077 ( .A1(n12044), .A2(n12043), .ZN(n12506) );
  INV_X1 U12078 ( .A(n13621), .ZN(n12459) );
  AND2_X1 U12079 ( .A1(n11941), .A2(n11940), .ZN(n12482) );
  INV_X1 U12080 ( .A(n11810), .ZN(n10351) );
  INV_X1 U12081 ( .A(n11809), .ZN(n10350) );
  NOR2_X2 U12082 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11858) );
  CLKBUF_X1 U12083 ( .A(n12196), .Z(n12197) );
  NAND2_X1 U12084 ( .A1(n11832), .A2(n11829), .ZN(n11840) );
  NAND2_X1 U12085 ( .A1(n11647), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11654) );
  NAND2_X1 U12086 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12886) );
  INV_X1 U12087 ( .A(n12888), .ZN(n10032) );
  NOR2_X1 U12088 ( .A1(n12944), .A2(n21467), .ZN(n10125) );
  AND3_X1 U12089 ( .A1(n10061), .A2(n10062), .A3(
        P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10063) );
  INV_X1 U12090 ( .A(n12917), .ZN(n13062) );
  NAND2_X1 U12091 ( .A1(n10061), .A2(n10030), .ZN(n10029) );
  INV_X1 U12092 ( .A(n18976), .ZN(n10030) );
  NOR2_X1 U12093 ( .A1(n17807), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13001) );
  NOR2_X1 U12094 ( .A1(n18976), .A2(n12887), .ZN(n12922) );
  INV_X1 U12095 ( .A(n18957), .ZN(n17153) );
  NOR2_X1 U12096 ( .A1(n18949), .A2(n13122), .ZN(n15972) );
  NOR2_X1 U12097 ( .A1(n13050), .A2(n13049), .ZN(n13117) );
  AOI221_X1 U12098 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19109), .C1(n19005), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n19122), .ZN(n18506) );
  AND2_X1 U12099 ( .A1(n11534), .A2(n11533), .ZN(n14649) );
  AND2_X1 U12100 ( .A1(n11024), .A2(n11023), .ZN(n14732) );
  OR2_X1 U12101 ( .A1(n16098), .A2(n10728), .ZN(n11023) );
  AND2_X1 U12102 ( .A1(n11159), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11160) );
  AND2_X1 U12103 ( .A1(n14900), .A2(n9819), .ZN(n11134) );
  AND2_X1 U12104 ( .A1(n11112), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11113) );
  INV_X1 U12105 ( .A(n11111), .ZN(n11112) );
  OR2_X1 U12106 ( .A1(n14924), .A2(n10728), .ZN(n11073) );
  AND2_X1 U12107 ( .A1(n9819), .A2(n16099), .ZN(n10998) );
  NOR2_X1 U12108 ( .A1(n10050), .A2(n14748), .ZN(n10049) );
  INV_X1 U12109 ( .A(n10051), .ZN(n10050) );
  NOR2_X1 U12110 ( .A1(n10979), .A2(n14956), .ZN(n10980) );
  NAND2_X1 U12111 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n10980), .ZN(
        n11017) );
  NAND2_X1 U12112 ( .A1(n10948), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10979) );
  AND2_X1 U12113 ( .A1(n10935), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10948) );
  NOR2_X1 U12114 ( .A1(n10918), .A2(n14690), .ZN(n10935) );
  NAND2_X1 U12115 ( .A1(n10899), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10918) );
  INV_X1 U12116 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14690) );
  NOR2_X1 U12117 ( .A1(n10882), .A2(n14526), .ZN(n10899) );
  INV_X1 U12118 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16147) );
  AND2_X1 U12119 ( .A1(n10836), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10837) );
  NAND2_X1 U12120 ( .A1(n10837), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10876) );
  OR2_X1 U12121 ( .A1(n10806), .A2(n20289), .ZN(n10832) );
  INV_X1 U12122 ( .A(n10780), .ZN(n10781) );
  NAND2_X1 U12123 ( .A1(n10770), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10780) );
  AND2_X1 U12124 ( .A1(n10752), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10770) );
  AND2_X1 U12125 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10702), .ZN(
        n10726) );
  NAND2_X1 U12126 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10703) );
  INV_X1 U12127 ( .A(n14021), .ZN(n10679) );
  INV_X1 U12128 ( .A(n14589), .ZN(n10116) );
  NAND2_X1 U12129 ( .A1(n14640), .A2(n10117), .ZN(n14602) );
  AND2_X1 U12130 ( .A1(n14640), .A2(n10120), .ZN(n14611) );
  NAND2_X1 U12131 ( .A1(n14640), .A2(n14622), .ZN(n14624) );
  NOR2_X1 U12132 ( .A1(n14662), .A2(n14649), .ZN(n14651) );
  AND2_X1 U12133 ( .A1(n14651), .A2(n14642), .ZN(n14640) );
  OR2_X1 U12134 ( .A1(n14728), .A2(n14664), .ZN(n14662) );
  INV_X1 U12135 ( .A(n11411), .ZN(n10276) );
  NAND2_X1 U12136 ( .A1(n14735), .A2(n14726), .ZN(n14728) );
  OR2_X1 U12137 ( .A1(n9908), .A2(n11517), .ZN(n14746) );
  NOR2_X1 U12138 ( .A1(n11409), .A2(n14954), .ZN(n16244) );
  NAND2_X1 U12139 ( .A1(n10279), .A2(n10283), .ZN(n14965) );
  AND2_X1 U12140 ( .A1(n11502), .A2(n11501), .ZN(n14508) );
  NOR2_X1 U12141 ( .A1(n14521), .A2(n14508), .ZN(n14687) );
  OR2_X1 U12142 ( .A1(n14519), .A2(n14518), .ZN(n14521) );
  AND2_X1 U12143 ( .A1(n14365), .A2(n9964), .ZN(n14497) );
  INV_X1 U12144 ( .A(n9984), .ZN(n10101) );
  NAND2_X1 U12145 ( .A1(n14365), .A2(n10103), .ZN(n14462) );
  NAND2_X1 U12146 ( .A1(n14365), .A2(n14364), .ZN(n14419) );
  OR2_X1 U12147 ( .A1(n14221), .A2(n14219), .ZN(n14342) );
  NOR2_X1 U12148 ( .A1(n14342), .A2(n14341), .ZN(n14365) );
  NAND2_X1 U12149 ( .A1(n16218), .A2(n10026), .ZN(n10025) );
  NAND2_X1 U12150 ( .A1(n10027), .A2(n16211), .ZN(n10024) );
  OR2_X1 U12151 ( .A1(n20470), .A2(n20471), .ZN(n16336) );
  OR2_X1 U12152 ( .A1(n11573), .A2(n11557), .ZN(n16333) );
  NAND2_X1 U12153 ( .A1(n10106), .A2(n10111), .ZN(n14221) );
  NOR2_X1 U12154 ( .A1(n14024), .A2(n10107), .ZN(n10106) );
  NAND2_X1 U12155 ( .A1(n14183), .A2(n10108), .ZN(n10107) );
  INV_X1 U12156 ( .A(n14164), .ZN(n10108) );
  NOR2_X1 U12157 ( .A1(n9973), .A2(n10109), .ZN(n14184) );
  INV_X1 U12158 ( .A(n10111), .ZN(n10109) );
  NAND2_X1 U12159 ( .A1(n10110), .A2(n10111), .ZN(n14163) );
  INV_X1 U12160 ( .A(n14024), .ZN(n10110) );
  OR2_X1 U12161 ( .A1(n11573), .A2(n11572), .ZN(n15083) );
  OR2_X1 U12162 ( .A1(n14024), .A2(n14023), .ZN(n14086) );
  NAND2_X1 U12163 ( .A1(n11513), .A2(n11525), .ZN(n14138) );
  XNOR2_X1 U12164 ( .A(n10677), .B(n10676), .ZN(n20588) );
  NAND2_X1 U12165 ( .A1(n10565), .A2(n10643), .ZN(n10670) );
  INV_X1 U12166 ( .A(n10556), .ZN(n15125) );
  NAND2_X1 U12167 ( .A1(n21200), .A2(n15120), .ZN(n20631) );
  OR2_X1 U12168 ( .A1(n15120), .A2(n10700), .ZN(n20764) );
  BUF_X1 U12169 ( .A(n10602), .Z(n20534) );
  AND3_X1 U12170 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20500), .A3(n20499), 
        .ZN(n20551) );
  NOR2_X1 U12171 ( .A1(n20671), .A2(n20670), .ZN(n21021) );
  OR2_X1 U12172 ( .A1(n15120), .A2(n20502), .ZN(n21069) );
  AOI21_X1 U12173 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21214), .A(n20670), 
        .ZN(n21070) );
  INV_X1 U12174 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16040) );
  AOI221_X1 U12175 ( .B1(n12143), .B2(n15989), .C1(n12143), .C2(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n12142), .ZN(n12186) );
  OAI21_X1 U12176 ( .B1(n12497), .B2(n12362), .A(n10303), .ZN(n12225) );
  NAND2_X1 U12177 ( .A1(n12362), .A2(n12175), .ZN(n10303) );
  NAND2_X1 U12178 ( .A1(n12358), .A2(n12357), .ZN(n12836) );
  INV_X1 U12179 ( .A(n10302), .ZN(n12784) );
  NOR3_X1 U12180 ( .A1(n12339), .A2(n12338), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n12349) );
  NAND2_X1 U12181 ( .A1(n15627), .A2(n15628), .ZN(n15630) );
  OR2_X1 U12182 ( .A1(n12339), .A2(n12338), .ZN(n12345) );
  NAND2_X1 U12183 ( .A1(n9912), .A2(n12357), .ZN(n12332) );
  NOR2_X1 U12184 ( .A1(n13197), .A2(n15530), .ZN(n13199) );
  NAND2_X1 U12185 ( .A1(n12280), .A2(n12279), .ZN(n12299) );
  NAND2_X1 U12186 ( .A1(n12270), .A2(n9955), .ZN(n12281) );
  NAND2_X1 U12187 ( .A1(n12270), .A2(n10306), .ZN(n12272) );
  NAND2_X1 U12188 ( .A1(n12270), .A2(n12259), .ZN(n12269) );
  AND2_X2 U12189 ( .A1(n12262), .A2(n12261), .ZN(n12270) );
  NOR2_X1 U12190 ( .A1(n12252), .A2(n12251), .ZN(n12258) );
  NOR2_X1 U12191 ( .A1(n12240), .A2(n12230), .ZN(n12247) );
  MUX2_X1 U12192 ( .A(n12220), .B(n11792), .S(n12227), .Z(n12242) );
  NAND2_X1 U12193 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  INV_X1 U12194 ( .A(n10363), .ZN(n10362) );
  NAND2_X1 U12195 ( .A1(n14170), .A2(n10364), .ZN(n10363) );
  INV_X1 U12196 ( .A(n14152), .ZN(n10364) );
  INV_X1 U12197 ( .A(n15221), .ZN(n10370) );
  NAND2_X1 U12198 ( .A1(n13552), .A2(n9905), .ZN(n10365) );
  NAND2_X1 U12199 ( .A1(n15627), .A2(n9968), .ZN(n15345) );
  AND2_X1 U12200 ( .A1(n15627), .A2(n9970), .ZN(n15337) );
  AND2_X1 U12201 ( .A1(n10357), .A2(n10354), .ZN(n10353) );
  INV_X1 U12202 ( .A(n15253), .ZN(n10354) );
  OR2_X1 U12203 ( .A1(n15261), .A2(n13475), .ZN(n10352) );
  AND3_X1 U12205 ( .A1(n12629), .A2(n12628), .A3(n12627), .ZN(n15760) );
  AND3_X1 U12206 ( .A1(n12581), .A2(n12580), .A3(n12579), .ZN(n16578) );
  OR2_X1 U12207 ( .A1(n15793), .A2(n10294), .ZN(n16579) );
  NAND2_X1 U12208 ( .A1(n13268), .A2(n13757), .ZN(n13913) );
  XNOR2_X1 U12209 ( .A(n12852), .B(n12851), .ZN(n13179) );
  AND2_X1 U12210 ( .A1(n13183), .A2(n9898), .ZN(n13208) );
  NAND2_X1 U12211 ( .A1(n13183), .A2(n10158), .ZN(n13206) );
  NAND2_X1 U12212 ( .A1(n13204), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13205) );
  NOR2_X1 U12213 ( .A1(n15271), .A2(n10344), .ZN(n15259) );
  NAND2_X1 U12214 ( .A1(n13186), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13202) );
  AND2_X1 U12215 ( .A1(n14389), .A2(n9902), .ZN(n15286) );
  NOR2_X1 U12216 ( .A1(n13197), .A2(n10163), .ZN(n13201) );
  INV_X1 U12217 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19235) );
  NAND2_X1 U12218 ( .A1(n13187), .A2(n9886), .ZN(n13195) );
  NAND2_X1 U12219 ( .A1(n14093), .A2(n9899), .ZN(n14256) );
  AND2_X1 U12220 ( .A1(n13187), .A2(n10156), .ZN(n13196) );
  NAND2_X1 U12221 ( .A1(n13187), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13194) );
  NAND2_X1 U12222 ( .A1(n10332), .A2(n10333), .ZN(n13935) );
  NAND2_X1 U12223 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10154) );
  NOR2_X1 U12224 ( .A1(n13918), .A2(n13885), .ZN(n13903) );
  NOR2_X1 U12225 ( .A1(n13188), .A2(n16562), .ZN(n13190) );
  OR2_X1 U12226 ( .A1(n12832), .A2(n15398), .ZN(n12833) );
  OAI21_X1 U12227 ( .B1(n12786), .B2(n12320), .A(n12870), .ZN(n12834) );
  NAND2_X1 U12228 ( .A1(n10228), .A2(n9923), .ZN(n12835) );
  NAND2_X1 U12229 ( .A1(n10232), .A2(n10229), .ZN(n10228) );
  AND3_X1 U12230 ( .A1(n13231), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12787), .ZN(n12832) );
  NOR2_X1 U12231 ( .A1(n10325), .A2(n12750), .ZN(n10324) );
  NAND2_X1 U12232 ( .A1(n10327), .A2(n10326), .ZN(n10325) );
  AND2_X1 U12233 ( .A1(n10251), .A2(n10249), .ZN(n10248) );
  INV_X1 U12234 ( .A(n15435), .ZN(n10249) );
  NOR2_X1 U12235 ( .A1(n10100), .A2(n9987), .ZN(n10098) );
  INV_X1 U12236 ( .A(n10327), .ZN(n10100) );
  OR3_X1 U12237 ( .A1(n15632), .A2(n15617), .A3(n15636), .ZN(n15601) );
  NAND2_X1 U12238 ( .A1(n15473), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15623) );
  CLKBUF_X1 U12239 ( .A(n15470), .Z(n15471) );
  NAND2_X1 U12240 ( .A1(n10084), .A2(n10082), .ZN(n15493) );
  NOR2_X1 U12241 ( .A1(n10085), .A2(n9958), .ZN(n10082) );
  AND2_X1 U12242 ( .A1(n10086), .A2(n15674), .ZN(n10085) );
  INV_X1 U12243 ( .A(n15511), .ZN(n10321) );
  INV_X1 U12244 ( .A(n15373), .ZN(n10296) );
  NAND2_X1 U12245 ( .A1(n14389), .A2(n9945), .ZN(n15291) );
  NAND2_X1 U12246 ( .A1(n14389), .A2(n14388), .ZN(n14455) );
  OR2_X1 U12247 ( .A1(n19251), .A2(n12295), .ZN(n15505) );
  NAND2_X1 U12248 ( .A1(n15381), .A2(n15382), .ZN(n15384) );
  NOR2_X1 U12249 ( .A1(n14380), .A2(n14374), .ZN(n14389) );
  AND2_X1 U12250 ( .A1(n15538), .A2(n15536), .ZN(n15716) );
  NAND2_X1 U12251 ( .A1(n14093), .A2(n9956), .ZN(n14378) );
  INV_X1 U12252 ( .A(n14255), .ZN(n10348) );
  OR2_X1 U12253 ( .A1(n14378), .A2(n14377), .ZN(n14380) );
  NAND2_X1 U12254 ( .A1(n10079), .A2(n10265), .ZN(n15538) );
  NAND2_X1 U12255 ( .A1(n10080), .A2(n10268), .ZN(n10079) );
  NAND2_X1 U12256 ( .A1(n16510), .A2(n16512), .ZN(n15774) );
  AND2_X1 U12257 ( .A1(n13965), .A2(n13656), .ZN(n14093) );
  NAND2_X1 U12258 ( .A1(n14093), .A2(n14092), .ZN(n14154) );
  AND2_X1 U12259 ( .A1(n14401), .A2(n12756), .ZN(n15781) );
  AND3_X1 U12260 ( .A1(n12536), .A2(n12535), .A3(n12534), .ZN(n14293) );
  NOR2_X1 U12261 ( .A1(n15793), .A2(n14293), .ZN(n14292) );
  NAND2_X1 U12262 ( .A1(n12256), .A2(n12255), .ZN(n15547) );
  NAND2_X1 U12263 ( .A1(n12229), .A2(n19350), .ZN(n12248) );
  AOI21_X1 U12264 ( .B1(n12375), .B2(n12378), .A(n12377), .ZN(n13917) );
  NAND2_X1 U12265 ( .A1(n13265), .A2(n19873), .ZN(n13292) );
  CLKBUF_X1 U12266 ( .A(n11855), .Z(n11856) );
  CLKBUF_X1 U12267 ( .A(n12456), .Z(n12457) );
  OR2_X1 U12268 ( .A1(n11832), .A2(n11826), .ZN(n12006) );
  INV_X1 U12269 ( .A(n12006), .ZN(n19708) );
  OR2_X1 U12270 ( .A1(n20202), .A2(n19447), .ZN(n19948) );
  NAND2_X2 U12271 ( .A1(n11680), .A2(n11679), .ZN(n14199) );
  NAND2_X1 U12272 ( .A1(n11678), .A2(n16617), .ZN(n11679) );
  OAI21_X1 U12273 ( .B1(n11713), .B2(n11712), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11714) );
  CLKBUF_X1 U12274 ( .A(n11741), .Z(n11681) );
  NAND2_X2 U12275 ( .A1(n11640), .A2(n11639), .ZN(n19547) );
  NAND4_X1 U12276 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11639) );
  INV_X1 U12277 ( .A(n19568), .ZN(n19561) );
  INV_X1 U12278 ( .A(n19567), .ZN(n19559) );
  NOR2_X2 U12279 ( .A1(n14196), .A2(n14195), .ZN(n19568) );
  NOR2_X2 U12280 ( .A1(n14194), .A2(n14195), .ZN(n19567) );
  INV_X1 U12281 ( .A(n19948), .ZN(n14270) );
  INV_X1 U12282 ( .A(n19779), .ZN(n14269) );
  INV_X1 U12283 ( .A(n19546), .ZN(n19569) );
  CLKBUF_X1 U12284 ( .A(n12179), .Z(n12180) );
  INV_X1 U12285 ( .A(n19163), .ZN(n19155) );
  NOR2_X1 U12286 ( .A1(n19075), .A2(n16937), .ZN(n16837) );
  NOR2_X1 U12287 ( .A1(n17873), .A2(n17889), .ZN(n10174) );
  INV_X1 U12288 ( .A(n17873), .ZN(n10173) );
  NOR2_X1 U12289 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17036), .ZN(n17019) );
  NOR2_X1 U12290 ( .A1(n17745), .A2(n10034), .ZN(n10033) );
  NOR2_X1 U12291 ( .A1(n13079), .A2(n10037), .ZN(n17533) );
  INV_X1 U12292 ( .A(n17608), .ZN(n17574) );
  NOR2_X1 U12293 ( .A1(n13089), .A2(n13088), .ZN(n17526) );
  NOR2_X1 U12294 ( .A1(n10137), .A2(n10133), .ZN(n10132) );
  NOR2_X1 U12295 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  NOR2_X1 U12296 ( .A1(n17720), .A2(n17682), .ZN(n17701) );
  NOR2_X1 U12297 ( .A1(n17721), .A2(n17720), .ZN(n17722) );
  AND2_X1 U12298 ( .A1(n10166), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10165) );
  NOR2_X1 U12299 ( .A1(n17801), .A2(n10169), .ZN(n10166) );
  NAND2_X1 U12300 ( .A1(n17832), .A2(n10168), .ZN(n17786) );
  NOR2_X1 U12301 ( .A1(n17819), .A2(n16842), .ZN(n17832) );
  AND2_X1 U12302 ( .A1(n17941), .A2(n10176), .ZN(n17874) );
  NOR2_X1 U12303 ( .A1(n10177), .A2(n17900), .ZN(n10176) );
  INV_X1 U12304 ( .A(n10178), .ZN(n10177) );
  NOR3_X1 U12305 ( .A1(n10180), .A2(n10181), .A3(n10182), .ZN(n10178) );
  NOR2_X1 U12306 ( .A1(n17973), .A2(n17974), .ZN(n17941) );
  NOR4_X1 U12307 ( .A1(n21455), .A2(n18064), .A3(n18048), .A4(n17070), .ZN(
        n18019) );
  INV_X1 U12308 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18048) );
  NAND2_X1 U12309 ( .A1(n18106), .A2(n9926), .ZN(n18017) );
  NOR2_X1 U12310 ( .A1(n18098), .A2(n10171), .ZN(n10170) );
  NOR2_X1 U12311 ( .A1(n13148), .A2(n18103), .ZN(n18087) );
  INV_X1 U12312 ( .A(n18139), .ZN(n17144) );
  INV_X1 U12313 ( .A(n18164), .ZN(n18117) );
  AOI21_X1 U12314 ( .B1(n13002), .B2(n18030), .A(n13258), .ZN(n10148) );
  NAND2_X1 U12315 ( .A1(n15991), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16054) );
  OAI21_X1 U12316 ( .B1(n16702), .B2(n13001), .A(n16698), .ZN(n15992) );
  NOR2_X1 U12317 ( .A1(n16058), .A2(n13157), .ZN(n16683) );
  INV_X1 U12318 ( .A(n17807), .ZN(n16696) );
  NOR2_X1 U12319 ( .A1(n17818), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17817) );
  NAND2_X1 U12320 ( .A1(n17852), .A2(n17856), .ZN(n17851) );
  NOR2_X1 U12321 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17887), .ZN(
        n17880) );
  INV_X1 U12322 ( .A(n17932), .ZN(n10070) );
  INV_X1 U12323 ( .A(n17879), .ZN(n17896) );
  OR3_X1 U12324 ( .A1(n18030), .A2(n17926), .A3(n17886), .ZN(n17907) );
  NAND2_X1 U12325 ( .A1(n17995), .A2(n13250), .ZN(n18306) );
  NOR2_X1 U12326 ( .A1(n17962), .A2(n18362), .ZN(n17995) );
  OR2_X1 U12327 ( .A1(n18068), .A2(n17962), .ZN(n10068) );
  NAND2_X1 U12328 ( .A1(n18024), .A2(n18321), .ZN(n10067) );
  NOR2_X1 U12329 ( .A1(n18360), .A2(n17962), .ZN(n18341) );
  NOR2_X1 U12330 ( .A1(n18967), .A2(n18958), .ZN(n18375) );
  INV_X1 U12331 ( .A(n18023), .ZN(n18362) );
  INV_X1 U12332 ( .A(n12987), .ZN(n12988) );
  NAND2_X1 U12333 ( .A1(n10060), .A2(n10057), .ZN(n18079) );
  AOI21_X1 U12334 ( .B1(n10055), .B2(n18095), .A(n9933), .ZN(n10060) );
  NAND2_X1 U12335 ( .A1(n18094), .A2(n10058), .ZN(n10057) );
  NOR2_X1 U12336 ( .A1(n18105), .A2(n18104), .ZN(n18103) );
  INV_X1 U12337 ( .A(n18981), .ZN(n18958) );
  OAI21_X1 U12338 ( .B1(n13131), .B2(n13129), .A(n13128), .ZN(n16811) );
  NAND2_X1 U12339 ( .A1(n19155), .A2(n15979), .ZN(n18981) );
  INV_X1 U12340 ( .A(n15971), .ZN(n18950) );
  INV_X1 U12341 ( .A(n12922), .ZN(n17435) );
  NOR2_X1 U12342 ( .A1(n13100), .A2(n13099), .ZN(n18516) );
  INV_X1 U12343 ( .A(n17683), .ZN(n18508) );
  NOR2_X1 U12344 ( .A1(n13040), .A2(n13039), .ZN(n18521) );
  INV_X1 U12345 ( .A(n17533), .ZN(n18531) );
  INV_X1 U12346 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18968) );
  OAI21_X1 U12347 ( .B1(n13636), .B2(n13635), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13708) );
  NAND2_X1 U12348 ( .A1(n21225), .A2(n14310), .ZN(n14676) );
  INV_X1 U12349 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14526) );
  OR2_X1 U12350 ( .A1(n14676), .A2(n14553), .ZN(n20279) );
  NAND2_X1 U12351 ( .A1(n21225), .A2(n14312), .ZN(n20330) );
  INV_X1 U12352 ( .A(n20351), .ZN(n20342) );
  AND2_X1 U12353 ( .A1(n21225), .A2(n14314), .ZN(n20345) );
  INV_X1 U12354 ( .A(n20330), .ZN(n20344) );
  INV_X1 U12355 ( .A(n14772), .ZN(n14511) );
  INV_X1 U12356 ( .A(n14770), .ZN(n14720) );
  AND2_X1 U12357 ( .A1(n14770), .A2(n13878), .ZN(n14721) );
  AND2_X1 U12358 ( .A1(n13877), .A2(n13876), .ZN(n14770) );
  INV_X1 U12359 ( .A(n14511), .ZN(n14767) );
  INV_X1 U12360 ( .A(n14721), .ZN(n14768) );
  INV_X1 U12361 ( .A(n14805), .ZN(n14833) );
  AOI21_X1 U12362 ( .B1(n13850), .B2(n11249), .A(n20251), .ZN(n11299) );
  AND2_X1 U12363 ( .A1(n13853), .A2(n14120), .ZN(n11298) );
  AND2_X1 U12364 ( .A1(n14831), .A2(n14036), .ZN(n14838) );
  NOR2_X1 U12365 ( .A1(n14303), .A2(n14853), .ZN(n14304) );
  OAI211_X1 U12366 ( .C1(n11183), .C2(n11230), .A(n10220), .B(n10218), .ZN(
        n14845) );
  OR2_X1 U12367 ( .A1(n10221), .A2(n11230), .ZN(n10220) );
  AND2_X1 U12368 ( .A1(n10221), .A2(n11230), .ZN(n10219) );
  AND2_X1 U12369 ( .A1(n14303), .A2(n11203), .ZN(n14859) );
  AOI21_X1 U12370 ( .B1(n14595), .B2(n14593), .A(n14594), .ZN(n14871) );
  INV_X1 U12371 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20289) );
  AND2_X1 U12372 ( .A1(n21206), .A2(n14123), .ZN(n16214) );
  NAND2_X1 U12373 ( .A1(n20258), .A2(n14125), .ZN(n20432) );
  INV_X1 U12374 ( .A(n16214), .ZN(n20496) );
  XNOR2_X1 U12375 ( .A(n10089), .B(n11414), .ZN(n15026) );
  OAI21_X1 U12376 ( .B1(n14857), .B2(n11408), .A(n9890), .ZN(n10089) );
  NAND2_X1 U12377 ( .A1(n10028), .A2(n11362), .ZN(n16213) );
  NAND2_X1 U12378 ( .A1(n16218), .A2(n16217), .ZN(n10028) );
  OR2_X1 U12379 ( .A1(n11573), .A2(n11445), .ZN(n20449) );
  NAND2_X1 U12380 ( .A1(n14066), .A2(n10206), .ZN(n11443) );
  NOR2_X1 U12381 ( .A1(n15097), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20475) );
  OR2_X1 U12382 ( .A1(n11573), .A2(n11554), .ZN(n20479) );
  INV_X1 U12383 ( .A(n20479), .ZN(n20486) );
  INV_X1 U12384 ( .A(n20588), .ZN(n21207) );
  NOR2_X2 U12385 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21206) );
  INV_X1 U12386 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20850) );
  INV_X1 U12387 ( .A(n10662), .ZN(n10663) );
  NAND2_X1 U12388 ( .A1(n10681), .A2(n10591), .ZN(n13832) );
  INV_X1 U12389 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21205) );
  OR2_X1 U12390 ( .A1(n21200), .A2(n20796), .ZN(n21195) );
  INV_X1 U12391 ( .A(n21206), .ZN(n21194) );
  INV_X1 U12392 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20494) );
  OR2_X1 U12393 ( .A1(n14075), .A2(n20505), .ZN(n21212) );
  NAND2_X1 U12394 ( .A1(n10053), .A2(n20665), .ZN(n14065) );
  INV_X1 U12395 ( .A(n10681), .ZN(n10053) );
  NOR2_X1 U12396 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21189) );
  INV_X1 U12397 ( .A(n20673), .ZN(n20716) );
  OR2_X1 U12398 ( .A1(n20764), .A2(n20987), .ZN(n20762) );
  OAI211_X1 U12399 ( .C1(n20820), .C2(n20931), .A(n20856), .B(n20804), .ZN(
        n20822) );
  INV_X1 U12400 ( .A(n20901), .ZN(n20918) );
  INV_X1 U12401 ( .A(n20925), .ZN(n21065) );
  INV_X1 U12402 ( .A(n20940), .ZN(n21079) );
  INV_X1 U12403 ( .A(n20945), .ZN(n21084) );
  INV_X1 U12404 ( .A(n20950), .ZN(n21089) );
  INV_X1 U12405 ( .A(n20955), .ZN(n21094) );
  INV_X1 U12406 ( .A(n20960), .ZN(n21099) );
  INV_X1 U12407 ( .A(n20965), .ZN(n21104) );
  INV_X1 U12408 ( .A(n21073), .ZN(n21113) );
  INV_X1 U12409 ( .A(n20971), .ZN(n21111) );
  AND2_X1 U12410 ( .A1(n11297), .A2(n11296), .ZN(n16010) );
  OR2_X1 U12411 ( .A1(n11255), .A2(n11250), .ZN(n11297) );
  XOR2_X1 U12412 ( .A(n12783), .B(n12784), .Z(n16388) );
  NOR3_X1 U12413 ( .A1(n12309), .A2(n12308), .A3(n12306), .ZN(n12313) );
  AND2_X1 U12414 ( .A1(n19270), .A2(n19271), .ZN(n10149) );
  INV_X1 U12415 ( .A(n19368), .ZN(n19353) );
  AND2_X1 U12416 ( .A1(n13219), .A2(n13218), .ZN(n19369) );
  NAND2_X1 U12417 ( .A1(n19170), .A2(n16653), .ZN(n19371) );
  OR4_X1 U12418 ( .A1(n15818), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .A4(P2_STATEBS16_REG_SCAN_IN), .ZN(n19334)
         );
  NAND2_X1 U12419 ( .A1(n19170), .A2(n13211), .ZN(n19343) );
  XNOR2_X1 U12420 ( .A(n9939), .B(n12848), .ZN(n16380) );
  CLKBUF_X1 U12421 ( .A(n14370), .Z(n14371) );
  AND2_X1 U12422 ( .A1(n12672), .A2(n12671), .ZN(n14382) );
  CLKBUF_X1 U12423 ( .A(n14368), .Z(n14369) );
  CLKBUF_X1 U12424 ( .A(n14089), .Z(n14090) );
  CLKBUF_X1 U12425 ( .A(n14029), .Z(n14030) );
  CLKBUF_X1 U12426 ( .A(n13883), .Z(n13884) );
  NAND2_X1 U12427 ( .A1(n15213), .A2(n10366), .ZN(n10369) );
  NAND2_X1 U12428 ( .A1(n13552), .A2(n10370), .ZN(n10366) );
  NOR2_X1 U12429 ( .A1(n15793), .A2(n10291), .ZN(n15167) );
  AND2_X1 U12430 ( .A1(n13624), .A2(n16665), .ZN(n19415) );
  NOR2_X1 U12431 ( .A1(n19444), .A2(n19443), .ZN(n19423) );
  AND2_X1 U12432 ( .A1(n19415), .A2(n11655), .ZN(n19443) );
  INV_X1 U12433 ( .A(n19415), .ZN(n19442) );
  CLKBUF_X1 U12435 ( .A(n19484), .Z(n19475) );
  NOR2_X1 U12436 ( .A1(n19452), .A2(n19466), .ZN(n19484) );
  CLKBUF_X1 U12437 ( .A(n13710), .Z(n13745) );
  OR2_X1 U12438 ( .A1(n15205), .A2(n15138), .ZN(n15573) );
  INV_X1 U12439 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16527) );
  NAND2_X1 U12440 ( .A1(n15545), .A2(n15546), .ZN(n10072) );
  NAND2_X1 U12441 ( .A1(n10076), .A2(n12001), .ZN(n14394) );
  CLKBUF_X1 U12442 ( .A(n19489), .Z(n19490) );
  INV_X1 U12443 ( .A(n16550), .ZN(n19499) );
  NAND2_X1 U12444 ( .A1(n19173), .A2(n12806), .ZN(n16561) );
  AND2_X1 U12445 ( .A1(n16561), .A2(n13765), .ZN(n16550) );
  INV_X1 U12446 ( .A(n16561), .ZN(n19488) );
  OR2_X1 U12447 ( .A1(n19173), .A2(n14211), .ZN(n16543) );
  NAND2_X1 U12448 ( .A1(n13640), .A2(n19517), .ZN(n10299) );
  INV_X1 U12449 ( .A(n10300), .ZN(n10077) );
  OAI211_X1 U12450 ( .C1(n14545), .C2(n19534), .A(n9957), .B(n9900), .ZN(
        n10300) );
  OAI211_X1 U12451 ( .C1(n12363), .C2(n10237), .A(n10235), .B(n10233), .ZN(
        n15580) );
  NAND2_X1 U12452 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10237) );
  OAI21_X1 U12453 ( .B1(n15407), .B2(n10382), .A(n10234), .ZN(n10233) );
  NAND2_X1 U12454 ( .A1(n10250), .A2(n10251), .ZN(n15436) );
  AND2_X1 U12455 ( .A1(n10254), .A2(n9882), .ZN(n15447) );
  NAND2_X1 U12456 ( .A1(n15454), .A2(n15455), .ZN(n10254) );
  NAND2_X1 U12457 ( .A1(n10259), .A2(n10260), .ZN(n15626) );
  NAND2_X1 U12458 ( .A1(n10017), .A2(n10016), .ZN(n15676) );
  INV_X1 U12459 ( .A(n10086), .ZN(n10016) );
  NAND2_X1 U12460 ( .A1(n10270), .A2(n12278), .ZN(n15766) );
  NAND2_X1 U12461 ( .A1(n16510), .A2(n10271), .ZN(n10270) );
  AND2_X1 U12462 ( .A1(n14399), .A2(n12757), .ZN(n15780) );
  CLKBUF_X1 U12463 ( .A(n14421), .Z(n14422) );
  INV_X1 U12464 ( .A(n19526), .ZN(n16587) );
  NAND2_X1 U12465 ( .A1(n10288), .A2(n9975), .ZN(n14280) );
  INV_X1 U12466 ( .A(n12496), .ZN(n10284) );
  INV_X1 U12467 ( .A(n12233), .ZN(n16557) );
  NAND2_X1 U12468 ( .A1(n12755), .A2(n12467), .ZN(n16603) );
  NOR2_X1 U12469 ( .A1(n13982), .A2(n12496), .ZN(n15181) );
  NAND2_X1 U12470 ( .A1(n10244), .A2(n16611), .ZN(n16552) );
  INV_X1 U12471 ( .A(n19534), .ZN(n19500) );
  AND2_X1 U12472 ( .A1(n19523), .A2(n19512), .ZN(n15726) );
  INV_X1 U12473 ( .A(n19365), .ZN(n13805) );
  OR2_X1 U12474 ( .A1(n15819), .A2(n13758), .ZN(n20228) );
  INV_X1 U12475 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21540) );
  INV_X1 U12476 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21487) );
  XNOR2_X1 U12477 ( .A(n13749), .B(n13751), .ZN(n19676) );
  XNOR2_X1 U12478 ( .A(n13828), .B(n13830), .ZN(n19677) );
  INV_X1 U12479 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15989) );
  CLKBUF_X1 U12480 ( .A(n12148), .Z(n16632) );
  INV_X1 U12481 ( .A(n19659), .ZN(n19670) );
  OAI21_X1 U12482 ( .B1(n19682), .B2(n19681), .A(n19680), .ZN(n19701) );
  INV_X1 U12483 ( .A(n19765), .ZN(n19755) );
  OR2_X1 U12484 ( .A1(n19738), .A2(n19737), .ZN(n19762) );
  INV_X1 U12485 ( .A(n19870), .ZN(n19857) );
  AND2_X1 U12486 ( .A1(n19987), .A2(n19583), .ZN(n19903) );
  INV_X1 U12487 ( .A(n19889), .ZN(n19904) );
  OAI21_X1 U12488 ( .B1(n19971), .B2(n19873), .A(n19953), .ZN(n19973) );
  NOR2_X1 U12489 ( .A1(n19948), .A2(n19947), .ZN(n19999) );
  OAI22_X1 U12490 ( .A1(n16726), .A2(n19561), .B1(n21500), .B2(n19559), .ZN(
        n20033) );
  INV_X1 U12491 ( .A(n20050), .ZN(n20032) );
  OAI21_X1 U12492 ( .B1(n20025), .B2(n20024), .A(n20023), .ZN(n20046) );
  INV_X1 U12493 ( .A(n20096), .ZN(n20054) );
  AND2_X1 U12494 ( .A1(n11724), .A2(n19569), .ZN(n20059) );
  OAI22_X1 U12495 ( .A1(n15358), .A2(n19561), .B1(n15357), .B2(n19559), .ZN(
        n20077) );
  AND2_X1 U12496 ( .A1(n19552), .A2(n19569), .ZN(n20075) );
  NAND2_X1 U12497 ( .A1(n14270), .A2(n14269), .ZN(n20096) );
  AND2_X1 U12498 ( .A1(n19987), .A2(n14269), .ZN(n20092) );
  AOI21_X1 U12499 ( .B1(n18938), .B2(n18939), .A(n17720), .ZN(n19168) );
  NAND2_X1 U12500 ( .A1(n19002), .A2(n18941), .ZN(n17720) );
  INV_X1 U12501 ( .A(n10188), .ZN(n16859) );
  AND2_X1 U12502 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16837), .ZN(n16914) );
  NOR2_X1 U12503 ( .A1(n16938), .A2(n17018), .ZN(n16952) );
  NOR2_X1 U12504 ( .A1(n16950), .A2(n17889), .ZN(n16949) );
  NOR2_X1 U12505 ( .A1(n16961), .A2(n17065), .ZN(n16950) );
  NOR2_X1 U12506 ( .A1(n17187), .A2(n16835), .ZN(n17023) );
  NOR2_X1 U12507 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17059), .ZN(n17044) );
  NOR2_X1 U12508 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17136), .ZN(n17116) );
  INV_X1 U12509 ( .A(n19011), .ZN(n17147) );
  INV_X1 U12510 ( .A(n17194), .ZN(n17176) );
  INV_X1 U12511 ( .A(n17187), .ZN(n17173) );
  NAND2_X1 U12512 ( .A1(n16833), .A2(n18995), .ZN(n17187) );
  NOR4_X2 U12513 ( .A1(n18479), .A2(n19168), .A3(n17147), .A4(n19000), .ZN(
        n17183) );
  NOR2_X1 U12514 ( .A1(n17183), .A2(n17173), .ZN(n17201) );
  INV_X1 U12515 ( .A(n17154), .ZN(n17193) );
  NOR2_X1 U12516 ( .A1(n17429), .A2(n17428), .ZN(n17411) );
  NAND2_X1 U12517 ( .A1(n17556), .A2(n9906), .ZN(n17544) );
  NAND2_X1 U12518 ( .A1(n17556), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17552) );
  NOR2_X1 U12519 ( .A1(n17742), .A2(n17563), .ZN(n17556) );
  OR2_X1 U12520 ( .A1(n17740), .A2(n17562), .ZN(n17563) );
  NOR2_X1 U12521 ( .A1(n17738), .A2(n17569), .ZN(n17568) );
  NOR2_X1 U12522 ( .A1(n17726), .A2(n17599), .ZN(n17600) );
  INV_X1 U12523 ( .A(n17663), .ZN(n17614) );
  NAND2_X1 U12524 ( .A1(n9921), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17608) );
  INV_X1 U12525 ( .A(n17589), .ZN(n17607) );
  NOR2_X1 U12526 ( .A1(n17643), .A2(n10035), .ZN(n17613) );
  NAND2_X1 U12527 ( .A1(n17618), .A2(n10036), .ZN(n10035) );
  NOR2_X1 U12528 ( .A1(n17528), .A2(n17772), .ZN(n10036) );
  NOR2_X2 U12529 ( .A1(n13060), .A2(n13059), .ZN(n17612) );
  NOR2_X1 U12530 ( .A1(n12904), .A2(n12903), .ZN(n17655) );
  NAND2_X1 U12531 ( .A1(n18545), .A2(n16072), .ZN(n17663) );
  NOR2_X1 U12532 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  NOR2_X1 U12533 ( .A1(n10124), .A2(n10123), .ZN(n10122) );
  INV_X1 U12534 ( .A(n12927), .ZN(n10128) );
  NOR2_X1 U12535 ( .A1(n18964), .A2(n17663), .ZN(n17675) );
  OAI21_X1 U12536 ( .B1(n16071), .B2(n16070), .A(n19002), .ZN(n17674) );
  NAND2_X1 U12537 ( .A1(n18964), .A2(n16072), .ZN(n17680) );
  CLKBUF_X1 U12538 ( .A(n17698), .Z(n17717) );
  OAI21_X1 U12539 ( .B1(n19152), .B2(n19153), .A(n17722), .ZN(n17776) );
  CLKBUF_X1 U12540 ( .A(n17776), .Z(n17781) );
  NOR2_X2 U12542 ( .A1(n18541), .A2(n18847), .ZN(n18883) );
  NAND2_X1 U12543 ( .A1(n17941), .A2(n10178), .ZN(n17901) );
  NAND2_X1 U12544 ( .A1(n17941), .A2(n9896), .ZN(n17935) );
  NAND3_X1 U12545 ( .A1(n18164), .A2(n19151), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n17944) );
  INV_X1 U12546 ( .A(n17944), .ZN(n18006) );
  AND2_X1 U12547 ( .A1(n18106), .A2(n10170), .ZN(n18074) );
  NAND2_X1 U12548 ( .A1(n18106), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18097) );
  INV_X1 U12549 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18098) );
  NOR2_X1 U12550 ( .A1(n18139), .A2(n18122), .ZN(n18106) );
  INV_X1 U12551 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18122) );
  CLKBUF_X1 U12552 ( .A(n18118), .Z(n18120) );
  NAND2_X1 U12553 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18139) );
  INV_X1 U12554 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18135) );
  INV_X1 U12555 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18153) );
  INV_X2 U12556 ( .A(n18883), .ZN(n18540) );
  NOR2_X1 U12557 ( .A1(n18195), .A2(n18275), .ZN(n18246) );
  NAND2_X1 U12558 ( .A1(n10146), .A2(n10145), .ZN(n17933) );
  AND2_X1 U12559 ( .A1(n17948), .A2(n9947), .ZN(n10145) );
  INV_X1 U12560 ( .A(n10069), .ZN(n18066) );
  INV_X1 U12561 ( .A(n18490), .ZN(n18473) );
  NOR2_X1 U12562 ( .A1(n15981), .A2(n15980), .ZN(n19129) );
  INV_X1 U12563 ( .A(n19129), .ZN(n19126) );
  NOR2_X1 U12564 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19102), .ZN(
        n19122) );
  NOR2_X1 U12565 ( .A1(n19099), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19008) );
  INV_X1 U12566 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19102) );
  AND2_X1 U12567 ( .A1(n11309), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20497)
         );
  NAND2_X1 U12569 ( .A1(n10048), .A2(n10044), .ZN(P1_U2973) );
  INV_X1 U12570 ( .A(n10045), .ZN(n10044) );
  CLKBUF_X1 U12571 ( .A(n13966), .Z(n13967) );
  INV_X1 U12572 ( .A(n12876), .ZN(n12877) );
  AOI21_X1 U12573 ( .B1(n10188), .B2(n10187), .A(n10184), .ZN(n16855) );
  NOR2_X1 U12574 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  AOI21_X1 U12575 ( .B1(n13262), .B2(n18489), .A(n13261), .ZN(n13263) );
  OAI21_X1 U12576 ( .B1(n13260), .B2(n18335), .A(n13259), .ZN(n13261) );
  INV_X1 U12577 ( .A(n11702), .ZN(n13602) );
  INV_X1 U12578 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16562) );
  AND2_X4 U12579 ( .A1(n12473), .A2(n12481), .ZN(n12719) );
  INV_X1 U12580 ( .A(n14338), .ZN(n19533) );
  AND4_X1 U12581 ( .A1(n10518), .A2(n10517), .A3(n10516), .A4(n10515), .ZN(
        n9879) );
  AND2_X1 U12582 ( .A1(n15674), .A2(n10088), .ZN(n9880) );
  AND4_X1 U12583 ( .A1(n10155), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9881) );
  AND2_X2 U12584 ( .A1(n13409), .A2(n11857), .ZN(n11914) );
  INV_X1 U12585 ( .A(n11705), .ZN(n13600) );
  NAND2_X1 U12586 ( .A1(n10544), .A2(n10553), .ZN(n10549) );
  OR3_X1 U12587 ( .A1(n12342), .A2(n12320), .A3(n15617), .ZN(n9882) );
  NOR2_X1 U12588 ( .A1(n15438), .A2(n15596), .ZN(n15425) );
  NAND2_X1 U12589 ( .A1(n14731), .A2(n14732), .ZN(n14723) );
  NOR2_X1 U12590 ( .A1(n14683), .A2(n10214), .ZN(n9883) );
  AND2_X1 U12591 ( .A1(n11964), .A2(n9954), .ZN(n9884) );
  AND3_X1 U12592 ( .A1(n10392), .A2(n10481), .A3(n10480), .ZN(n9885) );
  NAND2_X1 U12593 ( .A1(n10321), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15496) );
  AND2_X1 U12594 ( .A1(n11832), .A2(n11827), .ZN(n9887) );
  INV_X1 U12595 ( .A(n11248), .ZN(n10548) );
  OR2_X1 U12596 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9888) );
  NOR2_X1 U12597 ( .A1(n15219), .A2(n15221), .ZN(n15220) );
  NAND2_X1 U12598 ( .A1(n10551), .A2(n20501), .ZN(n11449) );
  OR2_X1 U12599 ( .A1(n14858), .A2(n14999), .ZN(n9890) );
  AND2_X1 U12600 ( .A1(n10514), .A2(n10513), .ZN(n9891) );
  INV_X1 U12601 ( .A(n10213), .ZN(n14754) );
  INV_X1 U12602 ( .A(n15623), .ZN(n10099) );
  NAND2_X1 U12603 ( .A1(n12270), .A2(n9948), .ZN(n9892) );
  INV_X1 U12604 ( .A(n19547), .ZN(n12204) );
  OR2_X1 U12605 ( .A1(n15271), .A2(n10342), .ZN(n9893) );
  INV_X1 U12606 ( .A(n11788), .ZN(n12389) );
  AND2_X1 U12607 ( .A1(n14370), .A2(n10372), .ZN(n9894) );
  AND2_X1 U12608 ( .A1(n14092), .A2(n10347), .ZN(n9895) );
  AND2_X1 U12609 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9896) );
  AND2_X1 U12610 ( .A1(n19350), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9897) );
  AND2_X1 U12611 ( .A1(n10158), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9898) );
  AND2_X1 U12612 ( .A1(n9895), .A2(n14167), .ZN(n9899) );
  OR2_X1 U12613 ( .A1(n12864), .A2(n12870), .ZN(n9900) );
  OR3_X1 U12614 ( .A1(n12321), .A2(n12320), .A3(n16570), .ZN(n15526) );
  AND2_X1 U12615 ( .A1(n10308), .A2(n9969), .ZN(n9901) );
  AND2_X1 U12616 ( .A1(n10339), .A2(n15284), .ZN(n9902) );
  AND2_X1 U12617 ( .A1(n9898), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9903) );
  NOR2_X1 U12618 ( .A1(n14089), .A2(n14152), .ZN(n9904) );
  AND2_X1 U12619 ( .A1(n10367), .A2(n10370), .ZN(n9905) );
  AND2_X1 U12620 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15846) );
  AND2_X1 U12621 ( .A1(n10033), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9906) );
  AND2_X2 U12622 ( .A1(n13409), .A2(n11856), .ZN(n11913) );
  OR2_X1 U12623 ( .A1(n19570), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9907) );
  OR2_X1 U12624 ( .A1(n14521), .A2(n10112), .ZN(n9908) );
  OR2_X1 U12625 ( .A1(n15319), .A2(n15320), .ZN(n9909) );
  OR2_X1 U12626 ( .A1(n15522), .A2(n15521), .ZN(n9910) );
  OR2_X1 U12627 ( .A1(n12888), .A2(n12886), .ZN(n9911) );
  OR3_X1 U12628 ( .A1(n12309), .A2(n10310), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n9912) );
  AND2_X2 U12629 ( .A1(n14044), .A2(n14064), .ZN(n9913) );
  NOR2_X1 U12630 ( .A1(n14647), .A2(n14648), .ZN(n14633) );
  NOR2_X1 U12631 ( .A1(n15511), .A2(n10322), .ZN(n15486) );
  OR2_X1 U12632 ( .A1(n14647), .A2(n10192), .ZN(n14618) );
  AND2_X1 U12633 ( .A1(n17556), .A2(n10033), .ZN(n9914) );
  NAND2_X1 U12634 ( .A1(n11409), .A2(n14954), .ZN(n14939) );
  NAND2_X1 U12635 ( .A1(n16054), .A2(n10148), .ZN(n9916) );
  AND4_X1 U12636 ( .A1(n10475), .A2(n10474), .A3(n10473), .A4(n10472), .ZN(
        n9918) );
  NAND2_X1 U12637 ( .A1(n10917), .A2(n10916), .ZN(n14683) );
  NAND2_X1 U12638 ( .A1(n10917), .A2(n10051), .ZN(n14672) );
  AND2_X1 U12639 ( .A1(n10917), .A2(n10049), .ZN(n14738) );
  OR2_X1 U12640 ( .A1(n17721), .A2(n19152), .ZN(n9919) );
  INV_X1 U12641 ( .A(n10542), .ZN(n10553) );
  NAND2_X1 U12642 ( .A1(n10072), .A2(n12123), .ZN(n16535) );
  AND2_X1 U12643 ( .A1(n12280), .A2(n9901), .ZN(n9920) );
  AND2_X1 U12644 ( .A1(n17613), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n9921) );
  AND2_X1 U12645 ( .A1(n14415), .A2(n14459), .ZN(n9922) );
  NAND3_X1 U12646 ( .A1(n10380), .A2(n13771), .A3(n10545), .ZN(n13852) );
  INV_X1 U12647 ( .A(n13852), .ZN(n10203) );
  OR2_X1 U12648 ( .A1(n10230), .A2(n15397), .ZN(n9923) );
  NAND2_X1 U12649 ( .A1(n13651), .A2(n15680), .ZN(n15511) );
  NAND2_X1 U12650 ( .A1(n15233), .A2(n15235), .ZN(n15234) );
  NAND2_X1 U12651 ( .A1(n10369), .A2(n15215), .ZN(n15209) );
  NAND2_X1 U12652 ( .A1(n12281), .A2(n12357), .ZN(n12280) );
  OR2_X1 U12653 ( .A1(n14683), .A2(n14759), .ZN(n10213) );
  AND2_X1 U12654 ( .A1(n12255), .A2(n10227), .ZN(n9925) );
  AND2_X1 U12655 ( .A1(n10170), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9926) );
  OR2_X1 U12656 ( .A1(n10255), .A2(n10253), .ZN(n9927) );
  INV_X1 U12657 ( .A(n10180), .ZN(n10179) );
  NAND2_X1 U12658 ( .A1(n9896), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10180) );
  AND2_X1 U12659 ( .A1(n10299), .A2(n10077), .ZN(n9928) );
  NAND3_X1 U12660 ( .A1(n13114), .A2(n15873), .A3(n19152), .ZN(n9929) );
  INV_X1 U12661 ( .A(n14397), .ZN(n12094) );
  AND2_X1 U12662 ( .A1(n12219), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14397) );
  OR2_X1 U12663 ( .A1(n12486), .A2(n12485), .ZN(n9930) );
  AND4_X1 U12664 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n9931) );
  NAND2_X1 U12665 ( .A1(n15455), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9932) );
  NAND4_X1 U12666 ( .A1(n10393), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10544) );
  AND2_X1 U12667 ( .A1(n14738), .A2(n14740), .ZN(n14731) );
  NAND2_X1 U12668 ( .A1(n10099), .A2(n10098), .ZN(n12815) );
  NAND2_X1 U12669 ( .A1(n9922), .A2(n14483), .ZN(n14482) );
  NOR2_X1 U12670 ( .A1(n12984), .A2(n12981), .ZN(n9933) );
  INV_X1 U12671 ( .A(n12781), .ZN(n10230) );
  NAND2_X1 U12672 ( .A1(n12356), .A2(n12780), .ZN(n12781) );
  AND2_X1 U12673 ( .A1(n11470), .A2(n11469), .ZN(n14183) );
  AND2_X1 U12674 ( .A1(n15366), .A2(n15156), .ZN(n15155) );
  INV_X1 U12676 ( .A(n10547), .ZN(n11438) );
  NOR2_X1 U12677 ( .A1(n10125), .A2(n10063), .ZN(n9934) );
  AND2_X1 U12678 ( .A1(n15836), .A2(n14338), .ZN(n9935) );
  AND2_X1 U12679 ( .A1(n10093), .A2(n14999), .ZN(n9936) );
  AND2_X1 U12680 ( .A1(n14397), .A2(n12095), .ZN(n9937) );
  AND2_X1 U12681 ( .A1(n10078), .A2(n9928), .ZN(n9938) );
  INV_X1 U12682 ( .A(n10095), .ZN(n10094) );
  AND2_X1 U12683 ( .A1(n14954), .A2(n9988), .ZN(n10095) );
  AND2_X2 U12684 ( .A1(n11858), .A2(n13409), .ZN(n12109) );
  INV_X1 U12685 ( .A(n12719), .ZN(n12490) );
  AND2_X1 U12686 ( .A1(n10560), .A2(n10520), .ZN(n11420) );
  OR2_X1 U12687 ( .A1(n15207), .A2(n12803), .ZN(n9939) );
  INV_X1 U12688 ( .A(n10549), .ZN(n10204) );
  NAND2_X1 U12689 ( .A1(n14370), .A2(n14387), .ZN(n14386) );
  AND2_X1 U12690 ( .A1(n14389), .A2(n10339), .ZN(n9940) );
  NAND2_X1 U12691 ( .A1(n14415), .A2(n10052), .ZN(n14501) );
  NOR2_X1 U12692 ( .A1(n13192), .A2(n16527), .ZN(n13187) );
  OR2_X1 U12693 ( .A1(n14089), .A2(n10360), .ZN(n9941) );
  XNOR2_X1 U12694 ( .A(n11320), .B(n10663), .ZN(n14076) );
  INV_X1 U12695 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16656) );
  AND2_X1 U12696 ( .A1(n10103), .A2(n10102), .ZN(n9942) );
  AND2_X1 U12697 ( .A1(n10333), .A2(n10331), .ZN(n9943) );
  OR2_X1 U12698 ( .A1(n17949), .A2(n18303), .ZN(n10146) );
  OR2_X1 U12699 ( .A1(n9893), .A2(n15236), .ZN(n9944) );
  AND2_X1 U12700 ( .A1(n14388), .A2(n10341), .ZN(n9945) );
  OR2_X1 U12701 ( .A1(n15271), .A2(n15270), .ZN(n9946) );
  OR2_X1 U12702 ( .A1(n18030), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9947) );
  NAND2_X1 U12703 ( .A1(n10015), .A2(n12249), .ZN(n14423) );
  NOR2_X1 U12704 ( .A1(n14160), .A2(n14181), .ZN(n14180) );
  AND2_X1 U12705 ( .A1(n10306), .A2(n10305), .ZN(n9948) );
  NAND2_X1 U12706 ( .A1(n14370), .A2(n10373), .ZN(n9949) );
  AND2_X1 U12707 ( .A1(n14967), .A2(n15106), .ZN(n9950) );
  OR3_X1 U12708 ( .A1(n15271), .A2(n10344), .A3(n10343), .ZN(n9951) );
  OR3_X1 U12709 ( .A1(n14521), .A2(n10115), .A3(n10113), .ZN(n9952) );
  NAND2_X1 U12710 ( .A1(n13294), .A2(n13293), .ZN(n13892) );
  NAND2_X1 U12711 ( .A1(n10699), .A2(n10698), .ZN(n10700) );
  OR2_X1 U12712 ( .A1(n13892), .A2(n13893), .ZN(n13891) );
  INV_X1 U12713 ( .A(n10268), .ZN(n10267) );
  NOR2_X1 U12714 ( .A1(n15764), .A2(n10269), .ZN(n10268) );
  AND2_X1 U12715 ( .A1(n10195), .A2(n10194), .ZN(n9953) );
  AND2_X1 U12716 ( .A1(n11963), .A2(n12173), .ZN(n9954) );
  AND2_X1 U12717 ( .A1(n9948), .A2(n14159), .ZN(n9955) );
  AND2_X1 U12718 ( .A1(n9899), .A2(n10348), .ZN(n9956) );
  NOR2_X1 U12719 ( .A1(n12827), .A2(n12828), .ZN(n9957) );
  INV_X1 U12720 ( .A(n14595), .ZN(n11182) );
  INV_X1 U12721 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15541) );
  AND2_X1 U12722 ( .A1(n9880), .A2(n10083), .ZN(n9958) );
  INV_X1 U12723 ( .A(n10169), .ZN(n10168) );
  NAND3_X1 U12724 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10169) );
  AND2_X1 U12725 ( .A1(n10014), .A2(n14403), .ZN(n9959) );
  OR2_X1 U12726 ( .A1(n10601), .A2(n10600), .ZN(n10603) );
  INV_X1 U12727 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15530) );
  AND2_X1 U12728 ( .A1(n12336), .A2(n15636), .ZN(n9960) );
  AND2_X1 U12729 ( .A1(n10151), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9961) );
  AND2_X1 U12730 ( .A1(n10296), .A2(n15382), .ZN(n9962) );
  AND2_X1 U12731 ( .A1(n10372), .A2(n15283), .ZN(n9963) );
  AND2_X1 U12732 ( .A1(n9942), .A2(n10101), .ZN(n9964) );
  INV_X1 U12733 ( .A(n9882), .ZN(n10257) );
  AND2_X1 U12734 ( .A1(n9901), .A2(n12304), .ZN(n9965) );
  AND2_X1 U12735 ( .A1(n11042), .A2(n14732), .ZN(n9966) );
  INV_X1 U12736 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16548) );
  INV_X1 U12737 ( .A(n14015), .ZN(n20397) );
  INV_X1 U12738 ( .A(n11703), .ZN(n13407) );
  BUF_X1 U12739 ( .A(n10855), .Z(n11002) );
  NAND2_X1 U12740 ( .A1(n10203), .A2(n20501), .ZN(n11551) );
  NAND2_X1 U12741 ( .A1(n13753), .A2(n16665), .ZN(n13754) );
  OR2_X1 U12742 ( .A1(n14089), .A2(n10363), .ZN(n14169) );
  NAND2_X1 U12743 ( .A1(n13183), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13182) );
  NOR2_X1 U12744 ( .A1(n10160), .A2(n15497), .ZN(n13186) );
  AND2_X1 U12745 ( .A1(n13186), .A2(n10151), .ZN(n9967) );
  AND2_X1 U12746 ( .A1(n10298), .A2(n15628), .ZN(n9968) );
  INV_X1 U12747 ( .A(n12306), .ZN(n10311) );
  OR2_X1 U12748 ( .A1(n19552), .A2(n12408), .ZN(n9969) );
  AND2_X1 U12749 ( .A1(n9968), .A2(n10297), .ZN(n9970) );
  NAND2_X1 U12750 ( .A1(n12986), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18360) );
  NAND2_X1 U12751 ( .A1(n14019), .A2(n10680), .ZN(n14081) );
  OR2_X1 U12752 ( .A1(n13197), .A2(n10164), .ZN(n9971) );
  AND2_X1 U12753 ( .A1(n10288), .A2(n10287), .ZN(n9972) );
  OR2_X1 U12754 ( .A1(n14024), .A2(n14164), .ZN(n9973) );
  NAND2_X1 U12755 ( .A1(n11117), .A2(n11116), .ZN(n9974) );
  NAND2_X1 U12756 ( .A1(n10332), .A2(n9943), .ZN(n10335) );
  NAND2_X1 U12757 ( .A1(n14365), .A2(n9942), .ZN(n10105) );
  AND2_X1 U12758 ( .A1(n10284), .A2(n15180), .ZN(n9975) );
  AND2_X1 U12759 ( .A1(n10069), .A2(n18360), .ZN(n9976) );
  AND2_X1 U12760 ( .A1(n12283), .A2(n15756), .ZN(n9977) );
  AND2_X1 U12761 ( .A1(n10117), .A2(n10116), .ZN(n9978) );
  AND2_X1 U12762 ( .A1(n9970), .A2(n15328), .ZN(n9979) );
  NAND2_X1 U12763 ( .A1(n14093), .A2(n9895), .ZN(n10349) );
  AND2_X1 U12764 ( .A1(n10052), .A2(n10898), .ZN(n9980) );
  INV_X1 U12765 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20500) );
  INV_X1 U12766 ( .A(n10368), .ZN(n10367) );
  OR2_X1 U12767 ( .A1(n15210), .A2(n10371), .ZN(n10368) );
  INV_X1 U12768 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10305) );
  INV_X1 U12769 ( .A(n17889), .ZN(n10175) );
  INV_X1 U12770 ( .A(n18068), .ZN(n18030) );
  NOR2_X2 U12771 ( .A1(n17649), .A2(n12982), .ZN(n18068) );
  INV_X1 U12772 ( .A(n11866), .ZN(n13482) );
  INV_X2 U12773 ( .A(n12379), .ZN(n12453) );
  INV_X1 U12774 ( .A(n11801), .ZN(n12379) );
  AND2_X1 U12775 ( .A1(n13524), .A2(n13545), .ZN(n9981) );
  AND2_X1 U12776 ( .A1(n12374), .A2(n12373), .ZN(n9982) );
  AND2_X1 U12777 ( .A1(n17832), .A2(n10166), .ZN(n9983) );
  NAND2_X1 U12778 ( .A1(n11492), .A2(n11491), .ZN(n9984) );
  NAND2_X1 U12779 ( .A1(n17941), .A2(n10179), .ZN(n10183) );
  NOR2_X1 U12780 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(P2_EBX_REG_24__SCAN_IN), 
        .ZN(n9985) );
  AND2_X1 U12781 ( .A1(n15680), .A2(n10320), .ZN(n9986) );
  NAND2_X1 U12782 ( .A1(n10205), .A2(n10204), .ZN(n10209) );
  INV_X1 U12783 ( .A(n15215), .ZN(n10371) );
  INV_X1 U12784 ( .A(n19247), .ZN(n19348) );
  INV_X1 U12785 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10273) );
  INV_X1 U12786 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10167) );
  AND2_X1 U12787 ( .A1(n12556), .A2(n12555), .ZN(n14028) );
  INV_X1 U12788 ( .A(n14028), .ZN(n13300) );
  AND2_X1 U12789 ( .A1(n12649), .A2(n12648), .ZN(n14253) );
  INV_X1 U12790 ( .A(n14253), .ZN(n10361) );
  OR2_X1 U12791 ( .A1(n15617), .A2(n12750), .ZN(n9987) );
  AND2_X1 U12792 ( .A1(n15087), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9988) );
  NOR2_X1 U12793 ( .A1(n11412), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9989) );
  INV_X1 U12794 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10181) );
  INV_X1 U12795 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10034) );
  INV_X1 U12796 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10182) );
  INV_X1 U12797 ( .A(n15557), .ZN(n10326) );
  INV_X1 U12798 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10159) );
  INV_X1 U12799 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10171) );
  NOR2_X2 U12800 ( .A1(n20496), .A2(n20495), .ZN(n20552) );
  INV_X1 U12801 ( .A(n9990), .ZN(n21041) );
  NAND2_X1 U12802 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20552), .ZN(n9991) );
  NAND2_X1 U12803 ( .A1(DATAI_20_), .A2(n20498), .ZN(n9992) );
  NAND2_X1 U12804 ( .A1(n9991), .A2(n9992), .ZN(n9990) );
  INV_X1 U12805 ( .A(n21097), .ZN(n9993) );
  INV_X1 U12806 ( .A(n9993), .ZN(n9994) );
  INV_X1 U12807 ( .A(n21118), .ZN(n9995) );
  INV_X1 U12808 ( .A(n9995), .ZN(n9996) );
  INV_X1 U12809 ( .A(n21049), .ZN(n9997) );
  INV_X1 U12810 ( .A(n9997), .ZN(n9998) );
  INV_X1 U12811 ( .A(n21030), .ZN(n9999) );
  INV_X1 U12812 ( .A(n9999), .ZN(n10000) );
  INV_X1 U12813 ( .A(n21034), .ZN(n10001) );
  INV_X1 U12814 ( .A(n10001), .ZN(n10002) );
  INV_X1 U12815 ( .A(n21038), .ZN(n10003) );
  INV_X1 U12816 ( .A(n10003), .ZN(n10004) );
  INV_X1 U12817 ( .A(n21045), .ZN(n10005) );
  INV_X1 U12818 ( .A(n10005), .ZN(n10006) );
  INV_X1 U12819 ( .A(n15258), .ZN(n10346) );
  INV_X1 U12820 ( .A(n10194), .ZN(n10192) );
  AOI22_X2 U12821 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20552), .B1(DATAI_16_), 
        .B2(n20498), .ZN(n21026) );
  AND2_X2 U12822 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11855) );
  OR2_X2 U12823 ( .A1(n12363), .A2(n12779), .ZN(n15417) );
  XNOR2_X2 U12824 ( .A(n15406), .B(n15405), .ZN(n12363) );
  INV_X1 U12825 ( .A(n15454), .ZN(n10009) );
  NAND2_X1 U12826 ( .A1(n14393), .A2(n14392), .ZN(n10015) );
  OAI21_X1 U12827 ( .B1(n15119), .B2(n11386), .A(n11335), .ZN(n14122) );
  NAND2_X1 U12828 ( .A1(n20628), .A2(n10607), .ZN(n10608) );
  XNOR2_X2 U12829 ( .A(n10043), .B(n10576), .ZN(n20628) );
  INV_X1 U12830 ( .A(n10607), .ZN(n10021) );
  AND2_X1 U12831 ( .A1(n16217), .A2(n16211), .ZN(n10026) );
  NOR2_X2 U12832 ( .A1(n11409), .A2(n11410), .ZN(n14932) );
  NOR2_X2 U12833 ( .A1(n10277), .A2(n10276), .ZN(n14923) );
  AND2_X2 U12834 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13017), .ZN(
        n10061) );
  INV_X2 U12835 ( .A(n10029), .ZN(n15918) );
  NAND3_X1 U12836 ( .A1(n13076), .A2(n13078), .A3(n10038), .ZN(n10037) );
  OAI21_X1 U12837 ( .B1(n10029), .B2(n10041), .A(n10040), .ZN(n10039) );
  NAND2_X1 U12838 ( .A1(n18950), .A2(n15972), .ZN(n18939) );
  NAND2_X1 U12839 ( .A1(n10564), .A2(n10563), .ZN(n10043) );
  NAND2_X1 U12840 ( .A1(n14415), .A2(n9980), .ZN(n14500) );
  XNOR2_X1 U12841 ( .A(n10681), .B(n20665), .ZN(n14039) );
  NAND3_X1 U12842 ( .A1(n10054), .A2(n10737), .A3(n10863), .ZN(n10712) );
  NAND2_X1 U12843 ( .A1(n10737), .A2(n10054), .ZN(n21200) );
  NAND2_X1 U12844 ( .A1(n18094), .A2(n12981), .ZN(n17961) );
  INV_X2 U12845 ( .A(n10390), .ZN(n15908) );
  NAND2_X2 U12846 ( .A1(n10122), .A2(n10126), .ZN(n17668) );
  NAND2_X2 U12847 ( .A1(n10070), .A2(n18030), .ZN(n17879) );
  XNOR2_X2 U12848 ( .A(n12122), .B(n16596), .ZN(n15545) );
  NAND3_X2 U12849 ( .A1(n10076), .A2(n12048), .A3(n12001), .ZN(n14398) );
  OR2_X1 U12850 ( .A1(n12829), .A2(n16604), .ZN(n10078) );
  OR2_X1 U12851 ( .A1(n15528), .A2(n10081), .ZN(n10084) );
  NAND2_X1 U12852 ( .A1(n11403), .A2(n11404), .ZN(n10096) );
  NAND2_X1 U12853 ( .A1(n10092), .A2(n9936), .ZN(n14931) );
  NAND3_X1 U12854 ( .A1(n11403), .A2(n11404), .A3(n10095), .ZN(n10092) );
  INV_X4 U12855 ( .A(n14309), .ZN(n20501) );
  NAND2_X1 U12856 ( .A1(n10551), .A2(n14309), .ZN(n14319) );
  OR2_X1 U12857 ( .A1(n15623), .A2(n9987), .ZN(n15438) );
  NAND2_X1 U12858 ( .A1(n13651), .A2(n9986), .ZN(n15470) );
  INV_X1 U12859 ( .A(n15470), .ZN(n12130) );
  INV_X1 U12860 ( .A(n10105), .ZN(n14484) );
  INV_X1 U12861 ( .A(n14686), .ZN(n10115) );
  NAND2_X1 U12862 ( .A1(n14640), .A2(n9978), .ZN(n14587) );
  NAND3_X1 U12863 ( .A1(n12932), .A2(n12925), .A3(n9934), .ZN(n10124) );
  NAND2_X2 U12864 ( .A1(n10132), .A2(n10129), .ZN(n12969) );
  NAND3_X1 U12865 ( .A1(n12924), .A2(n12921), .A3(n10134), .ZN(n10133) );
  NAND3_X1 U12866 ( .A1(n10142), .A2(n10146), .A3(n12994), .ZN(n10141) );
  INV_X2 U12867 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19121) );
  NAND2_X1 U12868 ( .A1(n13186), .A2(n9961), .ZN(n13203) );
  INV_X1 U12869 ( .A(n13203), .ZN(n12809) );
  NAND3_X1 U12870 ( .A1(n10155), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13189) );
  NAND2_X1 U12871 ( .A1(n13183), .A2(n9903), .ZN(n12849) );
  NAND2_X1 U12872 ( .A1(n17832), .A2(n10165), .ZN(n13164) );
  AOI22_X1 U12873 ( .A1(n16961), .A2(n10174), .B1(n17065), .B2(n10173), .ZN(
        n10172) );
  INV_X1 U12874 ( .A(n10172), .ZN(n16939) );
  AOI21_X1 U12875 ( .B1(n16961), .B2(n10175), .A(n17065), .ZN(n16940) );
  INV_X1 U12876 ( .A(n10183), .ZN(n17918) );
  NOR3_X1 U12877 ( .A1(n17065), .A2(n16860), .A3(n17186), .ZN(n10187) );
  NAND2_X1 U12878 ( .A1(n10189), .A2(n10190), .ZN(n10606) );
  NAND3_X1 U12879 ( .A1(n10681), .A2(n20500), .A3(n10591), .ZN(n10189) );
  INV_X1 U12880 ( .A(n14647), .ZN(n10193) );
  NAND2_X1 U12881 ( .A1(n15119), .A2(n10660), .ZN(n10197) );
  NAND2_X1 U12882 ( .A1(n10197), .A2(n10199), .ZN(n14022) );
  INV_X1 U12883 ( .A(n14022), .ZN(n10198) );
  NAND2_X1 U12884 ( .A1(n10198), .A2(n10679), .ZN(n14019) );
  NAND4_X1 U12885 ( .A1(n14066), .A2(n10206), .A3(n10209), .A4(n10201), .ZN(
        n10550) );
  NAND4_X1 U12886 ( .A1(n11438), .A2(n10548), .A3(n10208), .A4(n13974), .ZN(
        n13834) );
  INV_X1 U12887 ( .A(n10209), .ZN(n11552) );
  NAND2_X1 U12888 ( .A1(n14731), .A2(n9966), .ZN(n14659) );
  INV_X1 U12889 ( .A(n14659), .ZN(n11076) );
  AND2_X1 U12890 ( .A1(n11183), .A2(n10223), .ZN(n14580) );
  NAND2_X1 U12891 ( .A1(n11183), .A2(n10219), .ZN(n10218) );
  NAND2_X1 U12892 ( .A1(n11183), .A2(n11182), .ZN(n14579) );
  INV_X1 U12893 ( .A(n14566), .ZN(n10224) );
  INV_X1 U12894 ( .A(n14228), .ZN(n12017) );
  NAND2_X1 U12895 ( .A1(n14228), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11895) );
  NOR2_X1 U12896 ( .A1(n16532), .A2(n16528), .ZN(n10227) );
  INV_X1 U12897 ( .A(n12776), .ZN(n10231) );
  INV_X1 U12898 ( .A(n12777), .ZN(n10232) );
  NAND2_X1 U12899 ( .A1(n15407), .A2(n9888), .ZN(n10234) );
  NAND3_X1 U12900 ( .A1(n12363), .A2(n15407), .A3(n10236), .ZN(n10235) );
  NAND2_X1 U12901 ( .A1(n12233), .A2(n10242), .ZN(n10241) );
  NAND2_X1 U12902 ( .A1(n10247), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16551) );
  INV_X1 U12903 ( .A(n10247), .ZN(n10244) );
  INV_X1 U12904 ( .A(n15445), .ZN(n10258) );
  NAND2_X1 U12905 ( .A1(n16510), .A2(n10263), .ZN(n10259) );
  NAND2_X1 U12906 ( .A1(n11411), .A2(n9989), .ZN(n10275) );
  NAND2_X1 U12907 ( .A1(n11411), .A2(n14999), .ZN(n14891) );
  NAND2_X1 U12908 ( .A1(n10278), .A2(n10280), .ZN(n11402) );
  CLKBUF_X1 U12909 ( .A(n14988), .Z(n10279) );
  NAND3_X1 U12910 ( .A1(n10288), .A2(n10287), .A3(n14408), .ZN(n14407) );
  NAND2_X1 U12911 ( .A1(n15381), .A2(n9962), .ZN(n15682) );
  NAND2_X1 U12912 ( .A1(n15627), .A2(n9979), .ZN(n15319) );
  NAND2_X1 U12913 ( .A1(n10302), .A2(n10301), .ZN(n12837) );
  NAND2_X1 U12914 ( .A1(n12280), .A2(n9965), .ZN(n12292) );
  NAND3_X1 U12915 ( .A1(n10312), .A2(n10311), .A3(n12428), .ZN(n10310) );
  NAND2_X1 U12916 ( .A1(n12332), .A2(n10313), .ZN(n12350) );
  NAND2_X1 U12917 ( .A1(n12332), .A2(n12333), .ZN(n12339) );
  NAND2_X1 U12918 ( .A1(n12096), .A2(n12097), .ZN(n10317) );
  NAND2_X2 U12919 ( .A1(n10316), .A2(n12099), .ZN(n12122) );
  NAND2_X1 U12920 ( .A1(n14421), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10316) );
  NAND2_X1 U12921 ( .A1(n10317), .A2(n10318), .ZN(n14421) );
  AOI21_X1 U12922 ( .B1(n14398), .B2(n10319), .A(n9937), .ZN(n10318) );
  NAND2_X1 U12923 ( .A1(n10323), .A2(n11996), .ZN(n12233) );
  NAND3_X1 U12924 ( .A1(n10323), .A2(n11996), .A3(n16556), .ZN(n16555) );
  AND3_X4 U12925 ( .A1(n11603), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11704) );
  INV_X1 U12926 ( .A(n10335), .ZN(n13964) );
  NOR3_X1 U12927 ( .A1(n9893), .A2(n15236), .A3(n15225), .ZN(n15226) );
  INV_X1 U12928 ( .A(n15136), .ZN(n10337) );
  INV_X1 U12929 ( .A(n12454), .ZN(n10338) );
  INV_X1 U12930 ( .A(n10349), .ZN(n14166) );
  NAND3_X1 U12931 ( .A1(n10352), .A2(n10353), .A3(n10355), .ZN(n15251) );
  NAND2_X1 U12932 ( .A1(n15261), .A2(n10356), .ZN(n10355) );
  NAND3_X1 U12933 ( .A1(n10355), .A2(n10357), .A3(n10352), .ZN(n15250) );
  AND2_X2 U12934 ( .A1(n13454), .A2(n15251), .ZN(n15240) );
  AND2_X1 U12935 ( .A1(n15261), .A2(n13406), .ZN(n13453) );
  AND2_X1 U12936 ( .A1(n13475), .A2(n13406), .ZN(n10356) );
  OR2_X1 U12937 ( .A1(n13475), .A2(n13406), .ZN(n10357) );
  NOR2_X2 U12938 ( .A1(n14089), .A2(n10358), .ZN(n14368) );
  OAI21_X1 U12939 ( .B1(n15213), .B2(n10368), .A(n10365), .ZN(n15208) );
  NAND2_X1 U12940 ( .A1(n15213), .A2(n13552), .ZN(n15219) );
  AND2_X2 U12941 ( .A1(n14370), .A2(n9963), .ZN(n15277) );
  INV_X1 U12942 ( .A(n12100), .ZN(n12102) );
  INV_X1 U12943 ( .A(n12049), .ZN(n12051) );
  INV_X1 U12944 ( .A(n14500), .ZN(n10917) );
  NAND2_X1 U12945 ( .A1(n14081), .A2(n14083), .ZN(n14082) );
  AOI21_X1 U12946 ( .B1(n11866), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n11664), .ZN(n11666) );
  NAND2_X1 U12947 ( .A1(n10769), .A2(n10774), .ZN(n11363) );
  AOI21_X1 U12948 ( .B1(n11705), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n16617), .ZN(n11634) );
  AOI22_X1 U12949 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11662) );
  INV_X1 U12950 ( .A(n12491), .ZN(n12513) );
  NAND2_X1 U12951 ( .A1(n15301), .A2(n15300), .ZN(n15303) );
  NAND2_X1 U12952 ( .A1(n10542), .A2(n11248), .ZN(n10566) );
  XNOR2_X1 U12953 ( .A(n11419), .B(n11418), .ZN(n14847) );
  XNOR2_X1 U12954 ( .A(n13501), .B(n13498), .ZN(n15233) );
  NAND2_X1 U12955 ( .A1(n13890), .A2(n13896), .ZN(n13909) );
  INV_X1 U12956 ( .A(n14326), .ZN(n10805) );
  NAND2_X1 U12957 ( .A1(n15205), .A2(n15204), .ZN(n15207) );
  AND2_X1 U12958 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13297) );
  NAND2_X1 U12959 ( .A1(n12456), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U12960 ( .A1(n11747), .A2(n11746), .ZN(n11748) );
  NAND2_X1 U12961 ( .A1(n10805), .A2(n10379), .ZN(n14361) );
  NAND2_X1 U12962 ( .A1(n10776), .A2(n10775), .ZN(n11389) );
  NAND2_X1 U12963 ( .A1(n15286), .A2(n15153), .ZN(n15271) );
  INV_X1 U12964 ( .A(n14082), .ZN(n10736) );
  INV_X1 U12965 ( .A(n11966), .ZN(n11967) );
  CLKBUF_X1 U12966 ( .A(n13288), .Z(n16601) );
  XNOR2_X1 U12967 ( .A(n15819), .B(n13282), .ZN(n13750) );
  INV_X1 U12968 ( .A(n11783), .ZN(n11800) );
  AND2_X1 U12969 ( .A1(n14211), .A2(n19569), .ZN(n20051) );
  AND2_X1 U12970 ( .A1(n14211), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13268) );
  INV_X1 U12971 ( .A(n11787), .ZN(n11788) );
  AOI21_X1 U12972 ( .B1(n14845), .B2(n16214), .A(n14844), .ZN(n14846) );
  NAND2_X1 U12973 ( .A1(n14845), .A2(n10377), .ZN(n11316) );
  NAND2_X1 U12974 ( .A1(n13551), .A2(n13549), .ZN(n13552) );
  NAND2_X1 U12975 ( .A1(n12830), .A2(n19526), .ZN(n12831) );
  AOI22_X1 U12976 ( .A1(n11866), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U12977 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U12978 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U12979 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U12980 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11604) );
  INV_X1 U12981 ( .A(n10400), .ZN(n10404) );
  NOR2_X1 U12982 ( .A1(n11299), .A2(n11298), .ZN(n14801) );
  INV_X2 U12983 ( .A(n14801), .ZN(n14836) );
  AND3_X1 U12984 ( .A1(n21205), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10375) );
  INV_X1 U12985 ( .A(n12202), .ZN(n11655) );
  NOR2_X1 U12986 ( .A1(n13005), .A2(n13004), .ZN(n10376) );
  AND2_X1 U12987 ( .A1(n14836), .A2(n13878), .ZN(n10377) );
  AND2_X1 U12988 ( .A1(n10964), .A2(n10963), .ZN(n10378) );
  NAND3_X1 U12989 ( .A1(n10804), .A2(n10803), .A3(n10802), .ZN(n10379) );
  AND2_X1 U12990 ( .A1(n10542), .A2(n10543), .ZN(n10380) );
  AND2_X1 U12991 ( .A1(n12856), .A2(n12855), .ZN(n10381) );
  INV_X1 U12992 ( .A(n12926), .ZN(n17370) );
  INV_X1 U12993 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13003) );
  INV_X1 U12994 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11418) );
  INV_X1 U12995 ( .A(n13502), .ZN(n13498) );
  XOR2_X1 U12996 ( .A(n15408), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Z(
        n10382) );
  INV_X2 U12997 ( .A(n17523), .ZN(n17517) );
  AND2_X1 U12998 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10383) );
  INV_X1 U12999 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11414) );
  AND4_X1 U13000 ( .A1(n12526), .A2(n12525), .A3(n12524), .A4(n12523), .ZN(
        n10384) );
  NAND2_X1 U13001 ( .A1(n16656), .A2(n15818), .ZN(n16651) );
  INV_X1 U13002 ( .A(n16651), .ZN(n11745) );
  OR2_X1 U13003 ( .A1(n20122), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n20247) );
  AND3_X1 U13004 ( .A1(n11663), .A2(n11662), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10385) );
  INV_X1 U13005 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20980) );
  XNOR2_X1 U13006 ( .A(n12840), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10386) );
  INV_X1 U13007 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12842) );
  CLKBUF_X1 U13008 ( .A(n16804), .Z(n16805) );
  INV_X1 U13009 ( .A(n18157), .ZN(n13159) );
  INV_X1 U13010 ( .A(n10912), .ZN(n10863) );
  INV_X1 U13011 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20277) );
  OR4_X1 U13012 ( .A1(n15566), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12870), .A4(n15557), .ZN(n10387) );
  OR2_X1 U13013 ( .A1(n15424), .A2(n16604), .ZN(n10388) );
  AND2_X1 U13014 ( .A1(n12772), .A2(n12771), .ZN(n10389) );
  OR2_X2 U13015 ( .A1(n17182), .A2(n12887), .ZN(n10391) );
  INV_X1 U13016 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15818) );
  INV_X1 U13017 ( .A(n17478), .ZN(n17220) );
  INV_X1 U13018 ( .A(n16541), .ZN(n19493) );
  AND2_X1 U13019 ( .A1(n10478), .A2(n10477), .ZN(n10392) );
  AND4_X1 U13021 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10393) );
  NAND2_X1 U13022 ( .A1(n14202), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11890) );
  AND2_X1 U13023 ( .A1(n11891), .A2(n11890), .ZN(n11896) );
  AND2_X1 U13024 ( .A1(n11286), .A2(n11264), .ZN(n11268) );
  NOR2_X1 U13025 ( .A1(n13641), .A2(n9848), .ZN(n11742) );
  INV_X1 U13026 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10394) );
  OR2_X1 U13027 ( .A1(n10748), .A2(n10747), .ZN(n11364) );
  OR2_X1 U13028 ( .A1(n10687), .A2(n10648), .ZN(n10619) );
  OR2_X1 U13029 ( .A1(n11263), .A2(n13974), .ZN(n11286) );
  AND2_X1 U13030 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  AND2_X1 U13031 ( .A1(n11742), .A2(n13621), .ZN(n11743) );
  AND2_X1 U13032 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11664) );
  INV_X1 U13033 ( .A(n11253), .ZN(n11241) );
  AND2_X1 U13034 ( .A1(n14513), .A2(n14514), .ZN(n10881) );
  INV_X1 U13035 ( .A(n10686), .ZN(n10604) );
  INV_X1 U13036 ( .A(n10560), .ZN(n10568) );
  AND3_X1 U13037 ( .A1(n10651), .A2(n10650), .A3(n10649), .ZN(n10652) );
  NAND2_X1 U13038 ( .A1(n11236), .A2(n11235), .ZN(n11240) );
  NOR2_X1 U13039 ( .A1(n12362), .A2(n16656), .ZN(n11758) );
  INV_X1 U13041 ( .A(n11711), .ZN(n11712) );
  AOI22_X1 U13042 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11660) );
  NOR2_X1 U13043 ( .A1(n11240), .A2(n11239), .ZN(n11287) );
  INV_X1 U13044 ( .A(n14162), .ZN(n10735) );
  INV_X1 U13045 ( .A(n14724), .ZN(n11042) );
  INV_X1 U13046 ( .A(n14685), .ZN(n10916) );
  INV_X1 U13047 ( .A(n14502), .ZN(n10898) );
  INV_X1 U13048 ( .A(n14327), .ZN(n10786) );
  NAND2_X1 U13049 ( .A1(n10543), .A2(n11248), .ZN(n10499) );
  OR2_X1 U13050 ( .A1(n10629), .A2(n10628), .ZN(n11329) );
  NAND2_X1 U13051 ( .A1(n15408), .A2(n15567), .ZN(n12780) );
  NAND2_X1 U13052 ( .A1(n11846), .A2(n11845), .ZN(n11899) );
  INV_X1 U13053 ( .A(n14621), .ZN(n11137) );
  NAND2_X1 U13054 ( .A1(n10736), .A2(n10735), .ZN(n14160) );
  OR2_X1 U13055 ( .A1(n11202), .A2(n14861), .ZN(n14303) );
  NOR2_X1 U13056 ( .A1(n11069), .A2(n14935), .ZN(n11070) );
  INV_X1 U13057 ( .A(n10603), .ZN(n11331) );
  NAND2_X1 U13058 ( .A1(n13878), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10784) );
  AND2_X1 U13059 ( .A1(n11490), .A2(n11489), .ZN(n14461) );
  INV_X1 U13060 ( .A(n11329), .ZN(n10644) );
  NAND2_X1 U13061 ( .A1(n10685), .A2(n10684), .ZN(n20665) );
  INV_X1 U13062 ( .A(n14382), .ZN(n13304) );
  INV_X1 U13063 ( .A(n14088), .ZN(n13302) );
  INV_X1 U13064 ( .A(n13429), .ZN(n13374) );
  AND4_X1 U13065 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12119) );
  OR2_X1 U13066 ( .A1(n19297), .A2(n12320), .ZN(n12283) );
  OAI21_X1 U13067 ( .B1(n12225), .B2(n12227), .A(n12224), .ZN(n12230) );
  NOR2_X1 U13068 ( .A1(n18531), .A2(n17526), .ZN(n13115) );
  INV_X1 U13069 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n21366) );
  AOI22_X1 U13070 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9823), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12919) );
  AND2_X1 U13071 ( .A1(n12997), .A2(n18068), .ZN(n12998) );
  INV_X1 U13072 ( .A(n11017), .ZN(n11018) );
  OR2_X1 U13073 ( .A1(n13873), .A2(n13768), .ZN(n11249) );
  AND2_X1 U13074 ( .A1(n14851), .A2(n9819), .ZN(n11226) );
  AOI21_X1 U13075 ( .B1(n11373), .B2(n10863), .A(n10785), .ZN(n14327) );
  AND2_X1 U13076 ( .A1(n11475), .A2(n11474), .ZN(n14219) );
  INV_X1 U13077 ( .A(n16283), .ZN(n15097) );
  AND2_X1 U13078 ( .A1(n20632), .A2(n21206), .ZN(n20634) );
  OAI21_X1 U13079 ( .B1(n21235), .B2(n16043), .A(n15129), .ZN(n20499) );
  AND4_X1 U13080 ( .A1(n12078), .A2(n12077), .A3(n12076), .A4(n12075), .ZN(
        n12089) );
  OAI211_X1 U13081 ( .C1(n12872), .C2(n12842), .A(n12871), .B(n10387), .ZN(
        n12873) );
  INV_X1 U13082 ( .A(n15779), .ZN(n12766) );
  AND2_X1 U13083 ( .A1(n12296), .A2(n15505), .ZN(n15462) );
  INV_X1 U13084 ( .A(n16641), .ZN(n13620) );
  AND2_X1 U13085 ( .A1(n20202), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19704) );
  INV_X1 U13086 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19873) );
  NAND2_X1 U13087 ( .A1(n17879), .A2(n17886), .ZN(n17857) );
  INV_X1 U13088 ( .A(n18321), .ZN(n17962) );
  AND2_X1 U13089 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n11018), .ZN(
        n11019) );
  OR2_X1 U13090 ( .A1(n10876), .A2(n16147), .ZN(n10882) );
  OR2_X1 U13091 ( .A1(n21225), .A2(n14302), .ZN(n16076) );
  INV_X1 U13092 ( .A(n20324), .ZN(n14558) );
  AND2_X1 U13093 ( .A1(n11504), .A2(n11503), .ZN(n14686) );
  NAND2_X1 U13094 ( .A1(n11113), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11158) );
  INV_X1 U13095 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14956) );
  AND2_X1 U13096 ( .A1(n11441), .A2(n11565), .ZN(n16032) );
  OR3_X1 U13097 ( .A1(n15075), .A2(n14894), .A3(n15048), .ZN(n15039) );
  AND2_X1 U13098 ( .A1(n15077), .A2(n11586), .ZN(n15063) );
  OR4_X1 U13099 ( .A1(n11579), .A2(n20490), .A3(n11591), .A4(n16235), .ZN(
        n11580) );
  INV_X1 U13100 ( .A(n16358), .ZN(n16290) );
  INV_X1 U13101 ( .A(n20458), .ZN(n16292) );
  OR2_X1 U13102 ( .A1(n11573), .A2(n16012), .ZN(n16283) );
  INV_X1 U13103 ( .A(n21188), .ZN(n15129) );
  OR2_X1 U13104 ( .A1(n20764), .A2(n20923), .ZN(n20673) );
  OR2_X1 U13105 ( .A1(n21069), .A2(n20763), .ZN(n21073) );
  OR2_X1 U13106 ( .A1(n12748), .A2(n12747), .ZN(n16641) );
  INV_X1 U13107 ( .A(n19369), .ZN(n19349) );
  INV_X1 U13108 ( .A(n19356), .ZN(n19378) );
  AND2_X1 U13109 ( .A1(n12578), .A2(n12577), .ZN(n14088) );
  NAND2_X1 U13110 ( .A1(n19415), .A2(n13627), .ZN(n15386) );
  AND2_X1 U13111 ( .A1(n15726), .A2(n19513), .ZN(n15779) );
  OR3_X1 U13112 ( .A1(n19584), .A2(n19768), .A3(n19581), .ZN(n19612) );
  INV_X1 U13113 ( .A(n19675), .ZN(n19732) );
  NAND3_X1 U13114 ( .A1(n20206), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20020), 
        .ZN(n14195) );
  NOR2_X1 U13115 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16953), .ZN(n16941) );
  NOR2_X1 U13116 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16988), .ZN(n16982) );
  NOR2_X1 U13117 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17011), .ZN(n16998) );
  INV_X1 U13118 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17070) );
  NOR2_X1 U13119 ( .A1(n17337), .A2(n15875), .ZN(n17323) );
  NOR2_X1 U13120 ( .A1(n13113), .A2(n18952), .ZN(n15873) );
  NOR2_X1 U13121 ( .A1(n12914), .A2(n12913), .ZN(n13136) );
  INV_X1 U13122 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n21440) );
  INV_X1 U13123 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17973) );
  NAND2_X1 U13124 ( .A1(n17986), .A2(n18164), .ZN(n17898) );
  NOR2_X1 U13125 ( .A1(n18179), .A2(n16058), .ZN(n16681) );
  INV_X1 U13126 ( .A(n18945), .ZN(n18227) );
  NAND2_X1 U13127 ( .A1(n12988), .A2(n18030), .ZN(n18043) );
  INV_X1 U13128 ( .A(n12984), .ZN(n12983) );
  INV_X1 U13129 ( .A(n18396), .ZN(n18459) );
  INV_X1 U13130 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18969) );
  NOR2_X1 U13131 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18506), .ZN(n18850) );
  INV_X1 U13132 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19109) );
  NAND2_X1 U13133 ( .A1(n16049), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20251) );
  NAND2_X1 U13134 ( .A1(n11019), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11069) );
  AND2_X1 U13135 ( .A1(n16076), .A2(n14305), .ZN(n20307) );
  AND2_X1 U13136 ( .A1(n16076), .A2(n14315), .ZN(n20350) );
  AND2_X1 U13137 ( .A1(n16076), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20351) );
  INV_X1 U13138 ( .A(n20550), .ZN(n13878) );
  AND2_X1 U13139 ( .A1(n11164), .A2(n11163), .ZN(n14608) );
  NAND2_X1 U13140 ( .A1(n10712), .A2(n10711), .ZN(n14083) );
  INV_X2 U13141 ( .A(n20379), .ZN(n20386) );
  INV_X1 U13142 ( .A(n14097), .ZN(n20426) );
  NOR2_X1 U13143 ( .A1(n14517), .A2(n14516), .ZN(n14996) );
  NAND2_X1 U13144 ( .A1(n10781), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10806) );
  AND2_X1 U13145 ( .A1(n16032), .A2(n14120), .ZN(n20435) );
  OR2_X1 U13146 ( .A1(n16239), .A2(n11583), .ZN(n16229) );
  NAND2_X1 U13147 ( .A1(n11574), .A2(n16283), .ZN(n20474) );
  NOR2_X1 U13148 ( .A1(n16290), .A2(n16317), .ZN(n16352) );
  NOR2_X1 U13149 ( .A1(n20475), .A2(n16292), .ZN(n16299) );
  INV_X1 U13150 ( .A(n20449), .ZN(n20489) );
  INV_X1 U13151 ( .A(n20587), .ZN(n20578) );
  OAI21_X1 U13152 ( .B1(n20689), .B2(n20672), .A(n21021), .ZN(n20690) );
  INV_X1 U13153 ( .A(n20775), .ZN(n20792) );
  INV_X1 U13154 ( .A(n20889), .ZN(n20763) );
  INV_X1 U13155 ( .A(n20883), .ZN(n20845) );
  OR2_X1 U13156 ( .A1(n9870), .A2(n20588), .ZN(n20987) );
  NAND2_X1 U13157 ( .A1(n9870), .A2(n20588), .ZN(n21008) );
  OAI22_X1 U13158 ( .A1(n20936), .A2(n20935), .B1(n21012), .B2(n20934), .ZN(
        n20973) );
  OR2_X1 U13159 ( .A1(n9870), .A2(n21207), .ZN(n20923) );
  OAI211_X1 U13160 ( .C1(n21051), .C2(n21022), .A(n21021), .B(n21020), .ZN(
        n21053) );
  INV_X1 U13161 ( .A(n21224), .ZN(n21132) );
  OAI21_X1 U13162 ( .B1(n20240), .B2(n12218), .A(n12193), .ZN(n12791) );
  OR2_X1 U13163 ( .A1(n14545), .A2(n19343), .ZN(n13233) );
  NAND2_X1 U13164 ( .A1(n16443), .A2(n9875), .ZN(n16431) );
  INV_X1 U13165 ( .A(n15627), .ZN(n15354) );
  INV_X1 U13166 ( .A(n19371), .ZN(n19275) );
  INV_X1 U13167 ( .A(n19676), .ZN(n20221) );
  INV_X1 U13168 ( .A(n13750), .ZN(n13751) );
  INV_X1 U13169 ( .A(n19419), .ZN(n19444) );
  INV_X1 U13170 ( .A(n13680), .ZN(n13681) );
  AND2_X1 U13171 ( .A1(n13887), .A2(n13886), .ZN(n19360) );
  INV_X1 U13172 ( .A(n16543), .ZN(n19495) );
  INV_X1 U13173 ( .A(n16604), .ZN(n12862) );
  INV_X1 U13174 ( .A(n16603), .ZN(n19517) );
  AND2_X1 U13175 ( .A1(n12755), .A2(n20237), .ZN(n19526) );
  NOR2_X2 U13176 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20206) );
  NAND2_X1 U13177 ( .A1(n16642), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16660) );
  OAI21_X1 U13178 ( .B1(n14247), .B2(n14246), .A(n14245), .ZN(n19573) );
  INV_X1 U13179 ( .A(n19617), .ZN(n19605) );
  NOR2_X1 U13180 ( .A1(n19589), .A2(n19780), .ZN(n19646) );
  AND2_X1 U13181 ( .A1(n19675), .A2(n20199), .ZN(n19659) );
  AND2_X1 U13182 ( .A1(n14198), .A2(n20199), .ZN(n19700) );
  NOR2_X1 U13183 ( .A1(n19732), .A2(n19947), .ZN(n19718) );
  INV_X1 U13184 ( .A(n19986), .ZN(n19947) );
  NOR2_X1 U13185 ( .A1(n19779), .A2(n19732), .ZN(n19791) );
  INV_X1 U13186 ( .A(n19846), .ZN(n19848) );
  NOR2_X1 U13187 ( .A1(n19677), .A2(n20221), .ZN(n19583) );
  NOR2_X1 U13188 ( .A1(n19948), .A2(n19871), .ZN(n19939) );
  INV_X1 U13189 ( .A(n19976), .ZN(n19965) );
  INV_X1 U13190 ( .A(n20069), .ZN(n19994) );
  INV_X1 U13191 ( .A(n19943), .ZN(n20091) );
  AND2_X1 U13192 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13216), .ZN(n16665) );
  NAND2_X1 U13193 ( .A1(n18508), .A2(n18511), .ZN(n13124) );
  NOR2_X1 U13194 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16931), .ZN(n16921) );
  NOR2_X1 U13195 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16970), .ZN(n16957) );
  INV_X1 U13196 ( .A(n17201), .ZN(n16973) );
  NOR2_X1 U13197 ( .A1(n17201), .A2(n17021), .ZN(n17024) );
  NOR2_X1 U13198 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17084), .ZN(n17069) );
  NOR2_X1 U13199 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17110), .ZN(n17093) );
  INV_X1 U13200 ( .A(n17184), .ZN(n17115) );
  INV_X1 U13201 ( .A(n19166), .ZN(n16833) );
  INV_X1 U13202 ( .A(n17250), .ZN(n17243) );
  NOR2_X1 U13203 ( .A1(n18545), .A2(n17295), .ZN(n17297) );
  NOR3_X1 U13204 ( .A1(n17085), .A2(n17502), .A3(n15874), .ZN(n17431) );
  INV_X1 U13205 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17499) );
  NOR2_X1 U13206 ( .A1(n17730), .A2(n17595), .ZN(n17590) );
  INV_X1 U13207 ( .A(n17680), .ZN(n17665) );
  NOR2_X1 U13208 ( .A1(n17931), .A2(n18245), .ZN(n17916) );
  INV_X1 U13209 ( .A(n18360), .ZN(n18024) );
  NOR2_X2 U13210 ( .A1(n17649), .A2(n18168), .ZN(n18069) );
  INV_X1 U13211 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18064) );
  NOR2_X2 U13212 ( .A1(n13016), .A2(n13015), .ZN(n19152) );
  NAND2_X1 U13213 ( .A1(n13170), .A2(n13251), .ZN(n18305) );
  INV_X1 U13214 ( .A(n18474), .ZN(n18456) );
  INV_X1 U13215 ( .A(n18850), .ZN(n18541) );
  INV_X2 U13216 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13017) );
  INV_X1 U13217 ( .A(n18632), .ZN(n18625) );
  INV_X1 U13218 ( .A(n18655), .ZN(n18648) );
  INV_X1 U13219 ( .A(n18678), .ZN(n18671) );
  INV_X1 U13220 ( .A(n18701), .ZN(n18694) );
  INV_X1 U13221 ( .A(n18854), .ZN(n18871) );
  INV_X1 U13222 ( .A(n17526), .ZN(n18535) );
  INV_X1 U13223 ( .A(n19149), .ZN(n19002) );
  INV_X1 U13224 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19034) );
  NOR2_X1 U13225 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13650), .ZN(n16785)
         );
  NAND2_X1 U13226 ( .A1(n14120), .A2(n13816), .ZN(n14550) );
  NAND2_X1 U13227 ( .A1(n14549), .A2(n14550), .ZN(n21225) );
  NAND2_X1 U13228 ( .A1(n21136), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21222) );
  OR2_X1 U13229 ( .A1(n14720), .A2(n13878), .ZN(n14772) );
  OR2_X1 U13230 ( .A1(n20389), .A2(n14309), .ZN(n20365) );
  NAND2_X1 U13231 ( .A1(n20389), .A2(n20380), .ZN(n20379) );
  NAND2_X1 U13232 ( .A1(n13941), .A2(n14120), .ZN(n20389) );
  NOR2_X1 U13233 ( .A1(n14550), .A2(n13973), .ZN(n14015) );
  NAND2_X1 U13234 ( .A1(n20432), .A2(n14127), .ZN(n16219) );
  INV_X1 U13235 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21214) );
  INV_X1 U13236 ( .A(n21192), .ZN(n13869) );
  OR2_X1 U13237 ( .A1(n20631), .A2(n20923), .ZN(n20587) );
  OR2_X1 U13238 ( .A1(n20631), .A2(n20987), .ZN(n20625) );
  OR2_X1 U13239 ( .A1(n20631), .A2(n21008), .ZN(n20664) );
  OR2_X1 U13240 ( .A1(n20631), .A2(n20763), .ZN(n20693) );
  OR2_X1 U13241 ( .A1(n20764), .A2(n21008), .ZN(n20775) );
  OR2_X1 U13242 ( .A1(n20764), .A2(n20763), .ZN(n20800) );
  NAND2_X1 U13243 ( .A1(n20890), .A2(n20797), .ZN(n20849) );
  OR2_X1 U13244 ( .A1(n21195), .A2(n20987), .ZN(n20883) );
  OR2_X1 U13245 ( .A1(n21195), .A2(n21008), .ZN(n20901) );
  NAND2_X1 U13246 ( .A1(n20890), .A2(n20889), .ZN(n20977) );
  OR2_X1 U13247 ( .A1(n21069), .A2(n20923), .ZN(n21007) );
  NAND2_X1 U13248 ( .A1(n21018), .A2(n21009), .ZN(n21117) );
  INV_X1 U13249 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20931) );
  INV_X1 U13250 ( .A(n21186), .ZN(n21122) );
  INV_X1 U13251 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21136) );
  OR2_X1 U13252 ( .A1(n16638), .A2(n13222), .ZN(n13680) );
  INV_X1 U13253 ( .A(n13219), .ZN(n19170) );
  NAND2_X1 U13254 ( .A1(n12791), .A2(n13221), .ZN(n19173) );
  AND2_X1 U13255 ( .A1(n13233), .A2(n13232), .ZN(n13234) );
  INV_X1 U13256 ( .A(n19367), .ZN(n19351) );
  INV_X1 U13257 ( .A(n13920), .ZN(n15273) );
  NAND2_X1 U13258 ( .A1(n13897), .A2(n13909), .ZN(n20202) );
  NAND2_X1 U13259 ( .A1(n19415), .A2(n13625), .ZN(n19419) );
  INV_X1 U13260 ( .A(n19409), .ZN(n19450) );
  INV_X1 U13261 ( .A(n19452), .ZN(n19487) );
  NAND2_X1 U13262 ( .A1(n13681), .A2(n9859), .ZN(n13781) );
  OR2_X1 U13263 ( .A1(n19173), .A2(n11852), .ZN(n16541) );
  INV_X1 U13264 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16508) );
  INV_X1 U13265 ( .A(n15836), .ZN(n15197) );
  NAND2_X1 U13266 ( .A1(n12755), .A2(n20239), .ZN(n16604) );
  INV_X1 U13267 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21356) );
  INV_X1 U13268 ( .A(n19574), .ZN(n19566) );
  INV_X1 U13269 ( .A(n19646), .ZN(n19643) );
  INV_X1 U13270 ( .A(n19667), .ZN(n19664) );
  INV_X1 U13271 ( .A(n19700), .ZN(n19697) );
  INV_X1 U13272 ( .A(n19718), .ZN(n19731) );
  OR2_X1 U13273 ( .A1(n19947), .A2(n19780), .ZN(n19765) );
  INV_X1 U13274 ( .A(n19791), .ZN(n19821) );
  OR2_X1 U13275 ( .A1(n19780), .A2(n19779), .ZN(n19846) );
  NAND2_X1 U13276 ( .A1(n14270), .A2(n19583), .ZN(n19870) );
  INV_X1 U13277 ( .A(n19903), .ZN(n19900) );
  INV_X1 U13278 ( .A(n19939), .ZN(n19935) );
  INV_X1 U13279 ( .A(n20077), .ZN(n19968) );
  INV_X1 U13280 ( .A(n19999), .ZN(n20011) );
  NAND2_X1 U13281 ( .A1(n19987), .A2(n19986), .ZN(n20050) );
  INV_X1 U13282 ( .A(n19660), .ZN(n20086) );
  INV_X1 U13283 ( .A(n20196), .ZN(n20107) );
  NAND2_X1 U13284 ( .A1(n19002), .A2(n18947), .ZN(n16814) );
  NAND2_X1 U13285 ( .A1(n21390), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19161) );
  INV_X1 U13286 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17900) );
  NAND2_X1 U13287 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17023), .ZN(n17018) );
  INV_X1 U13288 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n21455) );
  INV_X1 U13289 ( .A(n17248), .ZN(n17263) );
  AND2_X1 U13290 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17627), .ZN(n17630) );
  INV_X1 U13291 ( .A(n17675), .ZN(n17673) );
  NOR2_X1 U13292 ( .A1(n18997), .A2(n17701), .ZN(n17698) );
  INV_X1 U13293 ( .A(n17701), .ZN(n17719) );
  INV_X1 U13294 ( .A(n18070), .ZN(n18025) );
  INV_X1 U13295 ( .A(n17951), .ZN(n17931) );
  INV_X1 U13296 ( .A(n18069), .ZN(n18057) );
  INV_X1 U13297 ( .A(n18158), .ZN(n18150) );
  OR2_X1 U13298 ( .A1(n19152), .A2(n16814), .ZN(n18168) );
  OAI21_X2 U13299 ( .B1(n13248), .B2(n13247), .A(n19002), .ZN(n18490) );
  INV_X1 U13300 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21466) );
  INV_X1 U13301 ( .A(n18404), .ZN(n18390) );
  INV_X1 U13302 ( .A(n18487), .ZN(n18482) );
  INV_X1 U13303 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18497) );
  INV_X1 U13304 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18502) );
  INV_X1 U13305 ( .A(n18721), .ZN(n18715) );
  INV_X1 U13306 ( .A(n18896), .ZN(n18806) );
  INV_X1 U13307 ( .A(n18862), .ZN(n18912) );
  INV_X1 U13308 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19099) );
  INV_X1 U13309 ( .A(n19097), .ZN(n21240) );
  NAND2_X1 U13310 ( .A1(n11316), .A2(n11315), .ZN(P1_U2873) );
  OR4_X1 U13311 ( .A1(n13667), .A2(n13666), .A3(n13665), .A4(n13664), .ZN(
        P2_U3037) );
  AND2_X2 U13312 ( .A1(n10406), .A2(n10401), .ZN(n11043) );
  AOI22_X1 U13313 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10887), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10399) );
  INV_X1 U13314 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10395) );
  AND2_X2 U13315 ( .A1(n10405), .A2(n10407), .ZN(n10717) );
  AND2_X2 U13316 ( .A1(n10407), .A2(n13839), .ZN(n10500) );
  AOI22_X1 U13317 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10500), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10398) );
  AND2_X2 U13318 ( .A1(n10401), .A2(n13839), .ZN(n10489) );
  AOI22_X1 U13319 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9868), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13320 ( .A1(n11058), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13321 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10479), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U13322 ( .A1(n10471), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9863), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10402) );
  AND2_X2 U13323 ( .A1(n10406), .A2(n10407), .ZN(n10855) );
  AOI22_X1 U13324 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10409) );
  AND2_X2 U13325 ( .A1(n10407), .A2(n14064), .ZN(n10476) );
  AOI22_X1 U13326 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U13327 ( .A1(n9863), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10414) );
  NAND2_X1 U13328 ( .A1(n10471), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10413) );
  NAND2_X1 U13329 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10412) );
  NAND2_X1 U13330 ( .A1(n11208), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10411) );
  NAND2_X1 U13331 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10418) );
  NAND2_X1 U13332 ( .A1(n10887), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10417) );
  NAND2_X1 U13333 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10416) );
  NAND2_X1 U13334 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10415) );
  NAND2_X1 U13335 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10422) );
  NAND2_X1 U13336 ( .A1(n9841), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10421) );
  NAND2_X1 U13337 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10420) );
  NAND2_X1 U13338 ( .A1(n10479), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10419) );
  NAND2_X1 U13339 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10426) );
  NAND2_X1 U13340 ( .A1(n10500), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10425) );
  NAND2_X1 U13341 ( .A1(n11058), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10424) );
  NAND2_X1 U13342 ( .A1(n9834), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10423) );
  NAND2_X1 U13343 ( .A1(n11208), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10434) );
  NAND2_X1 U13344 ( .A1(n10471), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10433) );
  NAND2_X1 U13345 ( .A1(n9830), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10432) );
  NAND2_X1 U13346 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10431) );
  NAND2_X1 U13347 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10438) );
  NAND2_X1 U13348 ( .A1(n10630), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10437) );
  NAND2_X1 U13349 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10436) );
  NAND2_X1 U13350 ( .A1(n10479), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10435) );
  NAND2_X1 U13351 ( .A1(n10887), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10442) );
  NAND2_X1 U13352 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10441) );
  NAND2_X1 U13353 ( .A1(n10500), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10440) );
  NAND2_X1 U13354 ( .A1(n9867), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10439) );
  NAND2_X1 U13355 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10446) );
  NAND2_X1 U13356 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10445) );
  NAND2_X1 U13357 ( .A1(n11058), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10444) );
  NAND2_X1 U13358 ( .A1(n10990), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10443) );
  AND4_X4 U13359 ( .A1(n10450), .A2(n10449), .A3(n10448), .A4(n10447), .ZN(
        n10542) );
  NAND2_X1 U13360 ( .A1(n11208), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10454) );
  NAND2_X1 U13361 ( .A1(n10471), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10453) );
  NAND2_X1 U13362 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10452) );
  NAND2_X1 U13363 ( .A1(n11142), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10451) );
  NAND2_X1 U13364 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10458) );
  NAND2_X1 U13365 ( .A1(n10630), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10457) );
  NAND2_X1 U13366 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10456) );
  NAND2_X1 U13367 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10455) );
  NAND2_X1 U13368 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13369 ( .A1(n10887), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10461) );
  NAND2_X1 U13370 ( .A1(n10479), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10460) );
  NAND2_X1 U13371 ( .A1(n9835), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10459) );
  NAND2_X1 U13372 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10466) );
  NAND2_X1 U13373 ( .A1(n10500), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10465) );
  NAND2_X1 U13374 ( .A1(n11058), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13375 ( .A1(n9868), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10463) );
  NAND4_X4 U13376 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n11248) );
  AOI22_X1 U13377 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9826), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13378 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9851), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13379 ( .A1(n9840), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10887), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13380 ( .A1(n10500), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9913), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13381 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U13382 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U13383 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9855), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13384 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10480) );
  NAND2_X1 U13385 ( .A1(n10556), .A2(n10546), .ZN(n10484) );
  NAND2_X1 U13386 ( .A1(n10549), .A2(n10482), .ZN(n10483) );
  NAND2_X1 U13387 ( .A1(n10484), .A2(n10483), .ZN(n10498) );
  AOI22_X1 U13388 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9826), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13389 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13390 ( .A1(n10887), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10479), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13391 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11058), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10485) );
  NAND4_X1 U13392 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10495) );
  AOI22_X1 U13393 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13394 ( .A1(n9830), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10489), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13395 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10500), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13396 ( .A1(n9913), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9835), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10490) );
  NAND4_X1 U13397 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        n10494) );
  NAND2_X1 U13398 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10504) );
  NAND2_X1 U13399 ( .A1(n10500), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10503) );
  NAND2_X1 U13400 ( .A1(n11058), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10502) );
  NAND2_X1 U13401 ( .A1(n10990), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10501) );
  NAND2_X1 U13402 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10508) );
  NAND2_X1 U13403 ( .A1(n9840), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10507) );
  NAND2_X1 U13404 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10506) );
  NAND2_X1 U13405 ( .A1(n10479), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10505) );
  NAND2_X1 U13406 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10512) );
  NAND2_X1 U13407 ( .A1(n10887), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10511) );
  NAND2_X1 U13408 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10510) );
  NAND2_X1 U13409 ( .A1(n9913), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10509) );
  NAND2_X1 U13410 ( .A1(n10630), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10518) );
  NAND2_X1 U13411 ( .A1(n10471), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10517) );
  NAND2_X1 U13412 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10516) );
  NAND2_X1 U13413 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10515) );
  NOR2_X1 U13414 ( .A1(n10499), .A2(n20501), .ZN(n10520) );
  NAND2_X1 U13415 ( .A1(n9863), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10524) );
  NAND2_X1 U13416 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10523) );
  NAND2_X1 U13417 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10522) );
  NAND2_X1 U13418 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10521) );
  NAND2_X1 U13419 ( .A1(n10887), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10528) );
  NAND2_X1 U13420 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10527) );
  NAND2_X1 U13421 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10526) );
  NAND2_X1 U13422 ( .A1(n10500), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10525) );
  NAND2_X1 U13423 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10532) );
  NAND2_X1 U13424 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10531) );
  NAND2_X1 U13425 ( .A1(n9840), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10530) );
  NAND2_X1 U13426 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10529) );
  NAND2_X1 U13427 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10537) );
  NAND2_X1 U13428 ( .A1(n9913), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10536) );
  NAND2_X1 U13429 ( .A1(n11058), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10535) );
  NAND2_X1 U13430 ( .A1(n9835), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10534) );
  NAND2_X1 U13431 ( .A1(n10548), .A2(n10544), .ZN(n14035) );
  INV_X1 U13432 ( .A(n14035), .ZN(n10545) );
  XNOR2_X1 U13433 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n11427) );
  NAND2_X2 U13434 ( .A1(n10550), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10576) );
  NAND2_X1 U13435 ( .A1(n10546), .A2(n10551), .ZN(n11447) );
  OR2_X1 U13436 ( .A1(n11447), .A2(n10499), .ZN(n13833) );
  NAND2_X1 U13437 ( .A1(n20523), .A2(n20501), .ZN(n11563) );
  AND2_X1 U13438 ( .A1(n14319), .A2(n11563), .ZN(n10552) );
  OAI211_X1 U13439 ( .C1(n21231), .C2(n10543), .A(n13833), .B(n10552), .ZN(
        n10571) );
  INV_X1 U13440 ( .A(n10571), .ZN(n10559) );
  NAND2_X1 U13441 ( .A1(n10548), .A2(n10553), .ZN(n10554) );
  AND2_X1 U13442 ( .A1(n10554), .A2(n20550), .ZN(n10570) );
  OR2_X1 U13443 ( .A1(n10499), .A2(n10553), .ZN(n10555) );
  NAND2_X1 U13444 ( .A1(n11561), .A2(n10543), .ZN(n11424) );
  NAND2_X1 U13445 ( .A1(n11424), .A2(n10556), .ZN(n10558) );
  NAND3_X1 U13446 ( .A1(n10559), .A2(n10558), .A3(n10557), .ZN(n11556) );
  NAND2_X1 U13447 ( .A1(n10576), .A2(n10561), .ZN(n10581) );
  NAND2_X1 U13448 ( .A1(n10581), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10564) );
  NAND2_X1 U13449 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10584) );
  OAI21_X1 U13450 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10584), .ZN(n20853) );
  OR2_X1 U13451 ( .A1(n16049), .A2(n20850), .ZN(n10578) );
  OAI21_X1 U13452 ( .B1(n14124), .B2(n20853), .A(n10578), .ZN(n10562) );
  INV_X1 U13453 ( .A(n10562), .ZN(n10563) );
  NAND2_X1 U13454 ( .A1(n10581), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10565) );
  MUX2_X1 U13455 ( .A(n16049), .B(n14124), .S(n21214), .Z(n10643) );
  INV_X1 U13456 ( .A(n14306), .ZN(n13768) );
  NAND3_X1 U13457 ( .A1(n13768), .A2(n10566), .A3(n10546), .ZN(n10567) );
  NAND2_X1 U13458 ( .A1(n10568), .A2(n10567), .ZN(n10575) );
  INV_X1 U13459 ( .A(n21189), .ZN(n15134) );
  NOR2_X1 U13460 ( .A1(n15134), .A2(n20500), .ZN(n10569) );
  NAND2_X1 U13461 ( .A1(n14043), .A2(n10542), .ZN(n11570) );
  OAI211_X1 U13462 ( .C1(n10570), .C2(n21231), .A(n10569), .B(n11570), .ZN(
        n10572) );
  NOR2_X1 U13463 ( .A1(n10572), .A2(n10571), .ZN(n10574) );
  NAND3_X1 U13464 ( .A1(n11424), .A2(n20517), .A3(n10556), .ZN(n10573) );
  NAND3_X1 U13465 ( .A1(n10575), .A2(n10574), .A3(n10573), .ZN(n10668) );
  INV_X1 U13466 ( .A(n10576), .ZN(n10580) );
  NAND2_X1 U13467 ( .A1(n10578), .A2(n10577), .ZN(n10579) );
  NAND2_X1 U13468 ( .A1(n10580), .A2(n10579), .ZN(n10589) );
  NOR2_X1 U13469 ( .A1(n16049), .A2(n20922), .ZN(n10582) );
  INV_X1 U13470 ( .A(n10584), .ZN(n10583) );
  NAND2_X1 U13471 ( .A1(n10583), .A2(n20922), .ZN(n20891) );
  NAND2_X1 U13472 ( .A1(n10584), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10585) );
  NAND2_X1 U13473 ( .A1(n20891), .A2(n10585), .ZN(n20512) );
  INV_X1 U13474 ( .A(n14124), .ZN(n10586) );
  NAND2_X1 U13475 ( .A1(n20512), .A2(n10586), .ZN(n10588) );
  NAND2_X1 U13476 ( .A1(n10590), .A2(n10588), .ZN(n10587) );
  NAND4_X1 U13477 ( .A1(n10608), .A2(n10590), .A3(n10589), .A4(n10588), .ZN(
        n10591) );
  AOI22_X1 U13478 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13479 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13480 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13481 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10592) );
  NAND4_X1 U13482 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10601) );
  AOI22_X1 U13483 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10599) );
  INV_X1 U13484 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n21509) );
  AOI22_X1 U13485 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13486 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9913), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13487 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10596) );
  NAND4_X1 U13488 ( .A1(n10599), .A2(n10598), .A3(n10597), .A4(n10596), .ZN(
        n10600) );
  AOI22_X1 U13489 ( .A1(n10604), .A2(n10603), .B1(n11289), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13490 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13491 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13492 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13493 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10609) );
  NAND4_X1 U13494 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n10618) );
  AOI22_X1 U13495 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13496 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13497 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13498 ( .A1(n9913), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9835), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10613) );
  NAND4_X1 U13499 ( .A1(n10616), .A2(n10615), .A3(n10614), .A4(n10613), .ZN(
        n10617) );
  OAI21_X2 U13500 ( .B1(n14077), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10619), 
        .ZN(n11320) );
  INV_X1 U13501 ( .A(n11320), .ZN(n10661) );
  AOI22_X1 U13502 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13503 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13504 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9913), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13505 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9856), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10620) );
  NAND4_X1 U13506 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(
        n10629) );
  AOI22_X1 U13507 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13508 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13509 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13510 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10624) );
  NAND4_X1 U13511 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .ZN(
        n10628) );
  NAND2_X1 U13512 ( .A1(n11289), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10642) );
  AOI22_X1 U13513 ( .A1(n9864), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9850), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13514 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13515 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13516 ( .A1(n9913), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9835), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10631) );
  NAND4_X1 U13517 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10640) );
  AOI22_X1 U13518 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13519 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13520 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13521 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10635) );
  NAND4_X1 U13522 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n10639) );
  AOI21_X1 U13523 ( .B1(n10543), .B2(n11378), .A(n20500), .ZN(n10641) );
  OAI211_X1 U13524 ( .C1(n10644), .C2(n20501), .A(n10642), .B(n10641), .ZN(
        n10677) );
  NAND2_X1 U13525 ( .A1(n10643), .A2(n20500), .ZN(n10646) );
  INV_X1 U13526 ( .A(n11378), .ZN(n11390) );
  MUX2_X1 U13527 ( .A(n10651), .B(n11387), .S(n10644), .Z(n10645) );
  NAND2_X1 U13528 ( .A1(n10677), .A2(n10676), .ZN(n10647) );
  NAND2_X1 U13529 ( .A1(n10647), .A2(n11387), .ZN(n10654) );
  NAND2_X1 U13530 ( .A1(n11289), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10650) );
  OR2_X1 U13531 ( .A1(n10686), .A2(n10648), .ZN(n10649) );
  INV_X1 U13532 ( .A(n10652), .ZN(n10653) );
  NOR2_X1 U13533 ( .A1(n10654), .A2(n10653), .ZN(n10655) );
  INV_X1 U13534 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n10658) );
  XNOR2_X1 U13535 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14701) );
  AOI21_X1 U13536 ( .B1(n9819), .B2(n14701), .A(n11229), .ZN(n10657) );
  OAI21_X1 U13537 ( .B1(n10784), .B2(n10658), .A(n10657), .ZN(n10659) );
  AOI21_X1 U13538 ( .B1(n10729), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10659), .ZN(n10660) );
  NAND2_X1 U13539 ( .A1(n11229), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10680) );
  NAND2_X1 U13540 ( .A1(n14076), .A2(n10863), .ZN(n10667) );
  INV_X1 U13541 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n10664) );
  INV_X1 U13542 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14135) );
  OAI22_X1 U13543 ( .A1(n10784), .A2(n10664), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14135), .ZN(n10665) );
  AOI21_X1 U13544 ( .B1(n10729), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10665), .ZN(n10666) );
  NAND2_X1 U13545 ( .A1(n10667), .A2(n10666), .ZN(n13872) );
  INV_X1 U13546 ( .A(n10668), .ZN(n10669) );
  XNOR2_X1 U13547 ( .A(n10670), .B(n10669), .ZN(n21209) );
  NAND2_X1 U13548 ( .A1(n21209), .A2(n10863), .ZN(n10675) );
  INV_X1 U13549 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n10672) );
  INV_X1 U13550 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10671) );
  OAI22_X1 U13551 ( .A1(n10784), .A2(n10672), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n10671), .ZN(n10673) );
  AOI21_X1 U13552 ( .B1(n10729), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10673), .ZN(n10674) );
  NAND2_X1 U13553 ( .A1(n10675), .A2(n10674), .ZN(n14143) );
  AOI21_X1 U13554 ( .B1(n20588), .B2(n10542), .A(n20980), .ZN(n14142) );
  NAND2_X1 U13555 ( .A1(n14143), .A2(n14142), .ZN(n14141) );
  INV_X1 U13556 ( .A(n9819), .ZN(n10728) );
  OR2_X1 U13557 ( .A1(n14143), .A2(n10728), .ZN(n10678) );
  NAND2_X1 U13558 ( .A1(n14141), .A2(n10678), .ZN(n13871) );
  NAND2_X1 U13559 ( .A1(n13872), .A2(n13871), .ZN(n14021) );
  NAND2_X1 U13560 ( .A1(n10581), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10685) );
  NAND2_X1 U13561 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10375), .ZN(
        n20766) );
  NAND2_X1 U13562 ( .A1(n21205), .A2(n20766), .ZN(n10682) );
  NOR3_X1 U13563 ( .A1(n21205), .A2(n20922), .A3(n20850), .ZN(n21072) );
  NAND2_X1 U13564 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21072), .ZN(
        n21060) );
  NAND2_X1 U13565 ( .A1(n10682), .A2(n21060), .ZN(n20798) );
  OAI22_X1 U13566 ( .A1(n14124), .A2(n20798), .B1(n16049), .B2(n21205), .ZN(
        n10683) );
  INV_X1 U13567 ( .A(n10683), .ZN(n10684) );
  NAND2_X1 U13568 ( .A1(n14039), .A2(n20500), .ZN(n10699) );
  AOI22_X1 U13569 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13570 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13571 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13572 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10688) );
  NAND4_X1 U13573 ( .A1(n10691), .A2(n10690), .A3(n10689), .A4(n10688), .ZN(
        n10697) );
  AOI22_X1 U13574 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13575 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13576 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9913), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13577 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9834), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10692) );
  NAND4_X1 U13578 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(
        n10696) );
  AOI22_X1 U13579 ( .A1(n11275), .A2(n11347), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n11289), .ZN(n10698) );
  INV_X1 U13580 ( .A(n10700), .ZN(n20502) );
  INV_X1 U13581 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n10709) );
  INV_X1 U13582 ( .A(n10703), .ZN(n10702) );
  INV_X1 U13583 ( .A(n10726), .ZN(n10706) );
  INV_X1 U13584 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10704) );
  NAND2_X1 U13585 ( .A1(n10704), .A2(n10703), .ZN(n10705) );
  NAND2_X1 U13586 ( .A1(n10706), .A2(n10705), .ZN(n20348) );
  AOI22_X1 U13587 ( .A1(n20348), .A2(n9819), .B1(n11229), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10708) );
  OAI21_X1 U13588 ( .B1(n10784), .B2(n10709), .A(n10708), .ZN(n10710) );
  AOI21_X1 U13589 ( .B1(n10729), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10710), .ZN(n10711) );
  AOI22_X1 U13590 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13591 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13592 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13593 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11143), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10713) );
  NAND4_X1 U13594 ( .A1(n10716), .A2(n10715), .A3(n10714), .A4(n10713), .ZN(
        n10723) );
  AOI22_X1 U13595 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13596 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11001), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13597 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10989), .B1(
        n9913), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13598 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9835), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10718) );
  NAND4_X1 U13599 ( .A1(n10721), .A2(n10720), .A3(n10719), .A4(n10718), .ZN(
        n10722) );
  NAND2_X1 U13600 ( .A1(n11275), .A2(n11365), .ZN(n10725) );
  NAND2_X1 U13601 ( .A1(n11289), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10724) );
  NAND2_X1 U13602 ( .A1(n10725), .A2(n10724), .ZN(n10738) );
  XNOR2_X1 U13603 ( .A(n10737), .B(n10738), .ZN(n11346) );
  NOR2_X1 U13604 ( .A1(n10726), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10727) );
  NOR2_X1 U13605 ( .A1(n10752), .A2(n10727), .ZN(n14175) );
  INV_X1 U13606 ( .A(n10729), .ZN(n10731) );
  INV_X1 U13607 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14067) );
  INV_X2 U13608 ( .A(n10784), .ZN(n10788) );
  AOI22_X1 U13609 ( .A1(n10788), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20980), .ZN(n10730) );
  OAI21_X1 U13610 ( .B1(n10731), .B2(n14067), .A(n10730), .ZN(n10732) );
  NAND2_X1 U13611 ( .A1(n10732), .A2(n10728), .ZN(n10733) );
  OAI21_X1 U13612 ( .B1(n14175), .B2(n10728), .A(n10733), .ZN(n10734) );
  AOI21_X1 U13613 ( .B1(n11346), .B2(n10863), .A(n10734), .ZN(n14162) );
  AOI22_X1 U13614 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13615 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13616 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13617 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10739) );
  NAND4_X1 U13618 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n10748) );
  AOI22_X1 U13619 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13620 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10500), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13621 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9913), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10744) );
  INV_X1 U13622 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n21429) );
  AOI22_X1 U13623 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10743) );
  NAND4_X1 U13624 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n10747) );
  AOI22_X1 U13625 ( .A1(n11275), .A2(n11364), .B1(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n11289), .ZN(n10749) );
  INV_X1 U13626 ( .A(n10776), .ZN(n10769) );
  NAND2_X1 U13627 ( .A1(n10750), .A2(n10749), .ZN(n10751) );
  NAND2_X1 U13628 ( .A1(n10769), .A2(n10751), .ZN(n11359) );
  INV_X1 U13629 ( .A(n11359), .ZN(n10758) );
  INV_X1 U13630 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n14187) );
  INV_X1 U13631 ( .A(n10770), .ZN(n10755) );
  INV_X1 U13632 ( .A(n10752), .ZN(n10753) );
  INV_X1 U13633 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20316) );
  NAND2_X1 U13634 ( .A1(n10753), .A2(n20316), .ZN(n10754) );
  NAND2_X1 U13635 ( .A1(n10755), .A2(n10754), .ZN(n20328) );
  AOI22_X1 U13636 ( .A1(n20328), .A2(n9819), .B1(n11229), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10756) );
  OAI21_X1 U13637 ( .B1(n10784), .B2(n14187), .A(n10756), .ZN(n10757) );
  AOI21_X1 U13638 ( .B1(n10758), .B2(n10863), .A(n10757), .ZN(n14181) );
  INV_X1 U13639 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13640 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13641 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13642 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13643 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10759) );
  NAND4_X1 U13644 ( .A1(n10762), .A2(n10761), .A3(n10760), .A4(n10759), .ZN(
        n10768) );
  AOI22_X1 U13645 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13646 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13647 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9913), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13648 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9834), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10763) );
  NAND4_X1 U13649 ( .A1(n10766), .A2(n10765), .A3(n10764), .A4(n10763), .ZN(
        n10767) );
  AOI22_X1 U13650 ( .A1(n11275), .A2(n11376), .B1(n11289), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U13651 ( .A1(n11363), .A2(n10863), .ZN(n10772) );
  OAI21_X1 U13652 ( .B1(n10770), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n10780), .ZN(n20304) );
  AOI22_X1 U13653 ( .A1(n20304), .A2(n9819), .B1(n11229), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10771) );
  OAI211_X1 U13654 ( .C1(n10784), .C2(n10773), .A(n10772), .B(n10771), .ZN(
        n14217) );
  NAND2_X1 U13655 ( .A1(n14180), .A2(n14217), .ZN(n14216) );
  INV_X1 U13656 ( .A(n14216), .ZN(n10787) );
  INV_X1 U13657 ( .A(n10774), .ZN(n10775) );
  NAND2_X1 U13658 ( .A1(n11275), .A2(n11378), .ZN(n10778) );
  NAND2_X1 U13659 ( .A1(n11289), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10777) );
  NAND2_X1 U13660 ( .A1(n10778), .A2(n10777), .ZN(n10779) );
  INV_X1 U13661 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10783) );
  OAI21_X1 U13662 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10781), .A(
        n10806), .ZN(n16208) );
  AOI22_X1 U13663 ( .A1(n9819), .A2(n16208), .B1(n11229), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10782) );
  OAI21_X1 U13664 ( .B1(n10784), .B2(n10783), .A(n10782), .ZN(n10785) );
  NAND2_X1 U13665 ( .A1(n10787), .A2(n10786), .ZN(n14326) );
  NAND2_X1 U13666 ( .A1(n10788), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10804) );
  XNOR2_X1 U13667 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10806), .ZN(
        n20297) );
  INV_X1 U13668 ( .A(n11229), .ZN(n10789) );
  OAI22_X1 U13669 ( .A1(n20297), .A2(n10728), .B1(n10789), .B2(n20289), .ZN(
        n10790) );
  INV_X1 U13670 ( .A(n10790), .ZN(n10803) );
  AOI22_X1 U13671 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13672 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13673 ( .A1(n9841), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13674 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9856), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10791) );
  NAND4_X1 U13675 ( .A1(n10794), .A2(n10793), .A3(n10792), .A4(n10791), .ZN(
        n10800) );
  AOI22_X1 U13676 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U13677 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U13678 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9913), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13679 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9834), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10795) );
  NAND4_X1 U13680 ( .A1(n10798), .A2(n10797), .A3(n10796), .A4(n10795), .ZN(
        n10799) );
  NOR2_X1 U13681 ( .A1(n10800), .A2(n10799), .ZN(n10801) );
  OR2_X1 U13682 ( .A1(n10912), .A2(n10801), .ZN(n10802) );
  XOR2_X1 U13683 ( .A(n20277), .B(n10832), .Z(n20284) );
  INV_X1 U13684 ( .A(n20284), .ZN(n10821) );
  AOI22_X1 U13685 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13686 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13687 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10500), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13688 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9835), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10807) );
  NAND4_X1 U13689 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n10816) );
  AOI22_X1 U13690 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13691 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13692 ( .A1(n9840), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9855), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13693 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10811) );
  NAND4_X1 U13694 ( .A1(n10814), .A2(n10813), .A3(n10812), .A4(n10811), .ZN(
        n10815) );
  NOR2_X1 U13695 ( .A1(n10816), .A2(n10815), .ZN(n10819) );
  NAND2_X1 U13696 ( .A1(n10788), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10818) );
  NAND2_X1 U13697 ( .A1(n11229), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10817) );
  OAI211_X1 U13698 ( .C1(n10819), .C2(n10912), .A(n10818), .B(n10817), .ZN(
        n10820) );
  AOI21_X1 U13699 ( .B1(n10821), .B2(n9819), .A(n10820), .ZN(n14414) );
  AOI22_X1 U13700 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13701 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13702 ( .A1(n9840), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13703 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9834), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10822) );
  NAND4_X1 U13704 ( .A1(n10825), .A2(n10824), .A3(n10823), .A4(n10822), .ZN(
        n10831) );
  AOI22_X1 U13705 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13706 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13707 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13708 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9856), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10826) );
  NAND4_X1 U13709 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10830) );
  NOR2_X1 U13710 ( .A1(n10831), .A2(n10830), .ZN(n10835) );
  XNOR2_X1 U13711 ( .A(n10836), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14470) );
  NAND2_X1 U13712 ( .A1(n14470), .A2(n9819), .ZN(n10834) );
  AOI22_X1 U13713 ( .A1(n10788), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n11229), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10833) );
  OAI211_X1 U13714 ( .C1(n10835), .C2(n10912), .A(n10834), .B(n10833), .ZN(
        n14459) );
  NAND2_X1 U13715 ( .A1(n10788), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n10839) );
  OAI21_X1 U13716 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10837), .A(
        n10876), .ZN(n16201) );
  AOI22_X1 U13717 ( .A1(n9819), .A2(n16201), .B1(n11229), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10838) );
  NAND2_X1 U13718 ( .A1(n10839), .A2(n10838), .ZN(n14483) );
  AOI22_X1 U13719 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13720 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13721 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10500), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13722 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10840) );
  NAND4_X1 U13723 ( .A1(n10843), .A2(n10842), .A3(n10841), .A4(n10840), .ZN(
        n10849) );
  AOI22_X1 U13724 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13725 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13726 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9867), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13727 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10844) );
  NAND4_X1 U13728 ( .A1(n10847), .A2(n10846), .A3(n10845), .A4(n10844), .ZN(
        n10848) );
  NOR2_X1 U13729 ( .A1(n10849), .A2(n10848), .ZN(n10850) );
  NOR2_X1 U13730 ( .A1(n10912), .A2(n10850), .ZN(n14491) );
  XOR2_X1 U13731 ( .A(n14526), .B(n10882), .Z(n14523) );
  AOI22_X1 U13732 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13733 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13734 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13735 ( .A1(n10500), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9835), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10851) );
  NAND4_X1 U13736 ( .A1(n10854), .A2(n10853), .A3(n10852), .A4(n10851), .ZN(
        n10861) );
  AOI22_X1 U13737 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13738 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13739 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9867), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13740 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10856) );
  NAND4_X1 U13741 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(
        n10860) );
  OR2_X1 U13742 ( .A1(n10861), .A2(n10860), .ZN(n10862) );
  AOI22_X1 U13743 ( .A1(n10863), .A2(n10862), .B1(n11229), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10865) );
  NAND2_X1 U13744 ( .A1(n10788), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10864) );
  OAI211_X1 U13745 ( .C1(n14523), .C2(n10728), .A(n10865), .B(n10864), .ZN(
        n14513) );
  AOI22_X1 U13746 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13747 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11144), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13748 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11001), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13749 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10989), .B1(
        n9913), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10866) );
  NAND4_X1 U13750 ( .A1(n10869), .A2(n10868), .A3(n10867), .A4(n10866), .ZN(
        n10875) );
  AOI22_X1 U13751 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13752 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U13753 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9869), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13754 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10870) );
  NAND4_X1 U13755 ( .A1(n10873), .A2(n10872), .A3(n10871), .A4(n10870), .ZN(
        n10874) );
  NOR2_X1 U13756 ( .A1(n10875), .A2(n10874), .ZN(n10880) );
  NAND2_X1 U13757 ( .A1(n10788), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10879) );
  XOR2_X1 U13758 ( .A(n16147), .B(n10876), .Z(n16190) );
  INV_X1 U13759 ( .A(n16190), .ZN(n10877) );
  AOI22_X1 U13760 ( .A1(n11229), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n9819), .B2(n10877), .ZN(n10878) );
  OAI211_X1 U13761 ( .C1(n10912), .C2(n10880), .A(n10879), .B(n10878), .ZN(
        n14514) );
  XNOR2_X1 U13762 ( .A(n10899), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16140) );
  AOI22_X1 U13763 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U13764 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9825), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U13765 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U13766 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9856), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10883) );
  NAND4_X1 U13767 ( .A1(n10886), .A2(n10885), .A3(n10884), .A4(n10883), .ZN(
        n10893) );
  AOI22_X1 U13768 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13769 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13770 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U13771 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9835), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10888) );
  NAND4_X1 U13772 ( .A1(n10891), .A2(n10890), .A3(n10889), .A4(n10888), .ZN(
        n10892) );
  NOR2_X1 U13773 ( .A1(n10893), .A2(n10892), .ZN(n10896) );
  NAND2_X1 U13774 ( .A1(n10788), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10895) );
  NAND2_X1 U13775 ( .A1(n11229), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10894) );
  OAI211_X1 U13776 ( .C1(n10896), .C2(n10912), .A(n10895), .B(n10894), .ZN(
        n10897) );
  AOI21_X1 U13777 ( .B1(n16140), .B2(n9819), .A(n10897), .ZN(n14502) );
  XOR2_X1 U13778 ( .A(n14690), .B(n10918), .Z(n16181) );
  INV_X1 U13779 ( .A(n16181), .ZN(n10915) );
  AOI22_X1 U13780 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13781 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9830), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13782 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9834), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U13783 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10900) );
  NAND4_X1 U13784 ( .A1(n10903), .A2(n10902), .A3(n10901), .A4(n10900), .ZN(
        n10909) );
  AOI22_X1 U13785 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U13786 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13787 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9855), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U13788 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10904) );
  NAND4_X1 U13789 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n10908) );
  NOR2_X1 U13790 ( .A1(n10909), .A2(n10908), .ZN(n10913) );
  NAND2_X1 U13791 ( .A1(n10788), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10911) );
  NAND2_X1 U13792 ( .A1(n11229), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10910) );
  OAI211_X1 U13793 ( .C1(n10913), .C2(n10912), .A(n10911), .B(n10910), .ZN(
        n10914) );
  AOI21_X1 U13794 ( .B1(n10915), .B2(n9819), .A(n10914), .ZN(n14685) );
  INV_X1 U13795 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14971) );
  XNOR2_X1 U13796 ( .A(n10935), .B(n14971), .ZN(n16126) );
  NAND2_X1 U13797 ( .A1(n16126), .A2(n9819), .ZN(n10934) );
  AOI22_X1 U13798 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9830), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13799 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U13800 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13801 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9855), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10919) );
  NAND4_X1 U13802 ( .A1(n10922), .A2(n10921), .A3(n10920), .A4(n10919), .ZN(
        n10930) );
  NAND2_X1 U13803 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10924) );
  NAND2_X1 U13804 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10923) );
  AND3_X1 U13805 ( .A1(n10924), .A2(n10923), .A3(n10728), .ZN(n10928) );
  AOI22_X1 U13806 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13807 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U13808 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9835), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10925) );
  NAND4_X1 U13809 ( .A1(n10928), .A2(n10927), .A3(n10926), .A4(n10925), .ZN(
        n10929) );
  NAND2_X1 U13810 ( .A1(n11199), .A2(n10728), .ZN(n11035) );
  OAI21_X1 U13811 ( .B1(n10930), .B2(n10929), .A(n11035), .ZN(n10932) );
  AOI22_X1 U13812 ( .A1(n10788), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20980), .ZN(n10931) );
  NAND2_X1 U13813 ( .A1(n10932), .A2(n10931), .ZN(n10933) );
  NAND2_X1 U13814 ( .A1(n10934), .A2(n10933), .ZN(n14759) );
  XOR2_X1 U13815 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10948), .Z(
        n16177) );
  AOI22_X1 U13816 ( .A1(n10788), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n11229), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13817 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U13818 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13819 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13820 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9835), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10936) );
  NAND4_X1 U13821 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(
        n10945) );
  AOI22_X1 U13822 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13823 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9825), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13824 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13825 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10940) );
  NAND4_X1 U13826 ( .A1(n10943), .A2(n10942), .A3(n10941), .A4(n10940), .ZN(
        n10944) );
  INV_X1 U13827 ( .A(n11199), .ZN(n11222) );
  OAI21_X1 U13828 ( .B1(n10945), .B2(n10944), .A(n11222), .ZN(n10946) );
  OAI211_X1 U13829 ( .C1(n16177), .C2(n10728), .A(n10947), .B(n10946), .ZN(
        n14753) );
  XNOR2_X1 U13830 ( .A(n10979), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14958) );
  NAND2_X1 U13831 ( .A1(n14958), .A2(n9819), .ZN(n10964) );
  AOI22_X1 U13832 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U13833 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U13834 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U13835 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9835), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10949) );
  NAND4_X1 U13836 ( .A1(n10952), .A2(n10951), .A3(n10950), .A4(n10949), .ZN(
        n10960) );
  AOI22_X1 U13837 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9840), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10958) );
  NAND2_X1 U13838 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10954) );
  NAND2_X1 U13839 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10953) );
  AND3_X1 U13840 ( .A1(n10954), .A2(n10953), .A3(n10728), .ZN(n10957) );
  AOI22_X1 U13841 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13842 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9856), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10955) );
  NAND4_X1 U13843 ( .A1(n10958), .A2(n10957), .A3(n10956), .A4(n10955), .ZN(
        n10959) );
  OAI21_X1 U13844 ( .B1(n10960), .B2(n10959), .A(n11035), .ZN(n10962) );
  AOI22_X1 U13845 ( .A1(n10788), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20980), .ZN(n10961) );
  NAND2_X1 U13846 ( .A1(n10962), .A2(n10961), .ZN(n10963) );
  AOI22_X1 U13847 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U13848 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U13849 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9855), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10966) );
  AOI22_X1 U13850 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10965) );
  NAND4_X1 U13851 ( .A1(n10968), .A2(n10967), .A3(n10966), .A4(n10965), .ZN(
        n10974) );
  AOI22_X1 U13852 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U13853 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U13854 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U13855 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9834), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10969) );
  NAND4_X1 U13856 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10973) );
  NOR2_X1 U13857 ( .A1(n10974), .A2(n10973), .ZN(n10978) );
  INV_X1 U13858 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10975) );
  OAI21_X1 U13859 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n10975), .A(n10728), 
        .ZN(n10976) );
  AOI21_X1 U13860 ( .B1(n10788), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10976), .ZN(
        n10977) );
  OAI21_X1 U13861 ( .B1(n11199), .B2(n10978), .A(n10977), .ZN(n10982) );
  OAI21_X1 U13862 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n10980), .A(
        n11017), .ZN(n16171) );
  OR2_X1 U13863 ( .A1(n10728), .A2(n16171), .ZN(n10981) );
  NAND2_X1 U13864 ( .A1(n10982), .A2(n10981), .ZN(n14748) );
  AOI22_X1 U13865 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11001), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U13866 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10984) );
  NAND2_X1 U13867 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10983) );
  AND3_X1 U13868 ( .A1(n10984), .A2(n10983), .A3(n10728), .ZN(n10987) );
  AOI22_X1 U13869 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U13870 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n9852), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10985) );
  NAND4_X1 U13871 ( .A1(n10988), .A2(n10987), .A3(n10986), .A4(n10985), .ZN(
        n10996) );
  AOI22_X1 U13872 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13873 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10989), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U13874 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U13875 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10991) );
  NAND4_X1 U13876 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n10995) );
  OR2_X1 U13877 ( .A1(n10996), .A2(n10995), .ZN(n10997) );
  NAND2_X1 U13878 ( .A1(n11035), .A2(n10997), .ZN(n11000) );
  AOI22_X1 U13879 ( .A1(n10788), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20980), .ZN(n10999) );
  XNOR2_X1 U13880 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11017), .ZN(
        n16099) );
  AOI21_X1 U13881 ( .B1(n11000), .B2(n10999), .A(n10998), .ZN(n14740) );
  AOI22_X1 U13882 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U13883 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U13884 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11001), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U13885 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11003) );
  NAND4_X1 U13886 ( .A1(n11006), .A2(n11005), .A3(n11004), .A4(n11003), .ZN(
        n11012) );
  AOI22_X1 U13887 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U13888 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9855), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U13889 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U13890 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9835), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11007) );
  NAND4_X1 U13891 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n11011) );
  NOR2_X1 U13892 ( .A1(n11012), .A2(n11011), .ZN(n11016) );
  INV_X1 U13893 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20927) );
  OAI21_X1 U13894 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20927), .A(
        n20980), .ZN(n11013) );
  INV_X1 U13895 ( .A(n11013), .ZN(n11014) );
  AOI21_X1 U13896 ( .B1(n10788), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11014), .ZN(
        n11015) );
  OAI21_X1 U13897 ( .B1(n11199), .B2(n11016), .A(n11015), .ZN(n11024) );
  INV_X1 U13898 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11021) );
  INV_X1 U13899 ( .A(n11019), .ZN(n11020) );
  NAND2_X1 U13900 ( .A1(n11021), .A2(n11020), .ZN(n11022) );
  NAND2_X1 U13901 ( .A1(n11069), .A2(n11022), .ZN(n16098) );
  AOI22_X1 U13902 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U13903 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U13904 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9856), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U13905 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9834), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11025) );
  NAND4_X1 U13906 ( .A1(n11028), .A2(n11027), .A3(n11026), .A4(n11025), .ZN(
        n11037) );
  AOI22_X1 U13907 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11001), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11034) );
  NAND2_X1 U13908 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11030) );
  NAND2_X1 U13909 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11029) );
  AND3_X1 U13910 ( .A1(n11030), .A2(n11029), .A3(n10728), .ZN(n11033) );
  AOI22_X1 U13911 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9855), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U13912 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11031) );
  NAND4_X1 U13913 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n11036) );
  OAI21_X1 U13914 ( .B1(n11037), .B2(n11036), .A(n11035), .ZN(n11039) );
  AOI22_X1 U13915 ( .A1(n10788), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20980), .ZN(n11038) );
  NAND2_X1 U13916 ( .A1(n11039), .A2(n11038), .ZN(n11041) );
  XNOR2_X1 U13917 ( .A(n11069), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16083) );
  NAND2_X1 U13918 ( .A1(n16083), .A2(n9819), .ZN(n11040) );
  NAND2_X1 U13919 ( .A1(n11041), .A2(n11040), .ZN(n14724) );
  AOI22_X1 U13920 ( .A1(n9865), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U13921 ( .A1(n11043), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U13922 ( .A1(n11001), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U13923 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11044) );
  NAND4_X1 U13924 ( .A1(n11047), .A2(n11046), .A3(n11045), .A4(n11044), .ZN(
        n11053) );
  AOI22_X1 U13925 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11051) );
  AOI22_X1 U13926 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U13927 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9855), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U13928 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9867), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11048) );
  NAND4_X1 U13929 ( .A1(n11051), .A2(n11050), .A3(n11049), .A4(n11048), .ZN(
        n11052) );
  NOR2_X1 U13930 ( .A1(n11053), .A2(n11052), .ZN(n11077) );
  AOI22_X1 U13931 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U13932 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U13933 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U13934 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9867), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11054) );
  NAND4_X1 U13935 ( .A1(n11057), .A2(n11056), .A3(n11055), .A4(n11054), .ZN(
        n11064) );
  AOI22_X1 U13936 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U13937 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U13938 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U13939 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11059) );
  NAND4_X1 U13940 ( .A1(n11062), .A2(n11061), .A3(n11060), .A4(n11059), .ZN(
        n11063) );
  NOR2_X1 U13941 ( .A1(n11064), .A2(n11063), .ZN(n11078) );
  XNOR2_X1 U13942 ( .A(n11077), .B(n11078), .ZN(n11068) );
  NAND2_X1 U13943 ( .A1(n20980), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11065) );
  NAND2_X1 U13944 ( .A1(n10728), .A2(n11065), .ZN(n11066) );
  AOI21_X1 U13945 ( .B1(n10788), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11066), .ZN(
        n11067) );
  OAI21_X1 U13946 ( .B1(n11199), .B2(n11068), .A(n11067), .ZN(n11074) );
  INV_X1 U13947 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14935) );
  INV_X1 U13948 ( .A(n11070), .ZN(n11071) );
  INV_X1 U13949 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14926) );
  NAND2_X1 U13950 ( .A1(n11071), .A2(n14926), .ZN(n11072) );
  NAND2_X1 U13951 ( .A1(n11111), .A2(n11072), .ZN(n14924) );
  NAND2_X1 U13952 ( .A1(n11074), .A2(n11073), .ZN(n14661) );
  NOR2_X1 U13953 ( .A1(n11078), .A2(n11077), .ZN(n11106) );
  AOI22_X1 U13954 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U13955 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U13956 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U13957 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9855), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11079) );
  NAND4_X1 U13958 ( .A1(n11082), .A2(n11081), .A3(n11080), .A4(n11079), .ZN(
        n11088) );
  AOI22_X1 U13959 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U13960 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U13961 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U13962 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11083) );
  NAND4_X1 U13963 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n11087) );
  OR2_X1 U13964 ( .A1(n11088), .A2(n11087), .ZN(n11105) );
  XNOR2_X1 U13965 ( .A(n11106), .B(n11105), .ZN(n11092) );
  NAND2_X1 U13966 ( .A1(n20980), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U13967 ( .A1(n10728), .A2(n11089), .ZN(n11090) );
  AOI21_X1 U13968 ( .B1(n10788), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11090), .ZN(
        n11091) );
  OAI21_X1 U13969 ( .B1(n11092), .B2(n11199), .A(n11091), .ZN(n11094) );
  XNOR2_X1 U13970 ( .A(n11111), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14916) );
  NAND2_X1 U13971 ( .A1(n14916), .A2(n9819), .ZN(n11093) );
  NAND2_X1 U13972 ( .A1(n11094), .A2(n11093), .ZN(n14648) );
  AOI22_X1 U13973 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U13974 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U13975 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9852), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U13976 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11095) );
  NAND4_X1 U13977 ( .A1(n11098), .A2(n11097), .A3(n11096), .A4(n11095), .ZN(
        n11104) );
  AOI22_X1 U13978 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U13979 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9855), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U13980 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U13981 ( .A1(n10489), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11099) );
  NAND4_X1 U13982 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n11099), .ZN(
        n11103) );
  NOR2_X1 U13983 ( .A1(n11104), .A2(n11103), .ZN(n11119) );
  NAND2_X1 U13984 ( .A1(n11106), .A2(n11105), .ZN(n11118) );
  XNOR2_X1 U13985 ( .A(n11119), .B(n11118), .ZN(n11110) );
  NAND2_X1 U13986 ( .A1(n20980), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11107) );
  NAND2_X1 U13987 ( .A1(n10728), .A2(n11107), .ZN(n11108) );
  AOI21_X1 U13988 ( .B1(n10788), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11108), .ZN(
        n11109) );
  OAI21_X1 U13989 ( .B1(n11110), .B2(n11199), .A(n11109), .ZN(n11117) );
  INV_X1 U13990 ( .A(n11113), .ZN(n11114) );
  INV_X1 U13991 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U13992 ( .A1(n11114), .A2(n14907), .ZN(n11115) );
  NAND2_X1 U13993 ( .A1(n11158), .A2(n11115), .ZN(n14905) );
  OR2_X1 U13994 ( .A1(n14905), .A2(n10728), .ZN(n11116) );
  NOR2_X1 U13995 ( .A1(n11119), .A2(n11118), .ZN(n11153) );
  AOI22_X1 U13996 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11123) );
  AOI22_X1 U13997 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11122) );
  AOI22_X1 U13998 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11121) );
  AOI22_X1 U13999 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11120) );
  NAND4_X1 U14000 ( .A1(n11123), .A2(n11122), .A3(n11121), .A4(n11120), .ZN(
        n11129) );
  AOI22_X1 U14001 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11127) );
  AOI22_X1 U14002 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11126) );
  AOI22_X1 U14003 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U14004 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9835), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11124) );
  NAND4_X1 U14005 ( .A1(n11127), .A2(n11126), .A3(n11125), .A4(n11124), .ZN(
        n11128) );
  OR2_X1 U14006 ( .A1(n11129), .A2(n11128), .ZN(n11152) );
  INV_X1 U14007 ( .A(n11152), .ZN(n11130) );
  XNOR2_X1 U14008 ( .A(n11153), .B(n11130), .ZN(n11131) );
  NAND2_X1 U14009 ( .A1(n11131), .A2(n11222), .ZN(n11136) );
  NAND2_X1 U14010 ( .A1(n20980), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14011 ( .A1(n10728), .A2(n11132), .ZN(n11133) );
  AOI21_X1 U14012 ( .B1(n10788), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11133), .ZN(
        n11135) );
  XNOR2_X1 U14013 ( .A(n11158), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14900) );
  AOI21_X1 U14014 ( .B1(n11136), .B2(n11135), .A(n11134), .ZN(n14621) );
  AOI22_X1 U14015 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11141) );
  AOI22_X1 U14016 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11001), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11140) );
  AOI22_X1 U14017 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9855), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14018 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9834), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11138) );
  NAND4_X1 U14019 ( .A1(n11141), .A2(n11140), .A3(n11139), .A4(n11138), .ZN(
        n11151) );
  AOI22_X1 U14020 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11143), .B1(
        n9851), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14021 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11144), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14022 ( .A1(n9864), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14023 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10533), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11146) );
  NAND4_X1 U14024 ( .A1(n11149), .A2(n11148), .A3(n11147), .A4(n11146), .ZN(
        n11150) );
  NOR2_X1 U14025 ( .A1(n11151), .A2(n11150), .ZN(n11166) );
  NAND2_X1 U14026 ( .A1(n11153), .A2(n11152), .ZN(n11165) );
  XNOR2_X1 U14027 ( .A(n11166), .B(n11165), .ZN(n11157) );
  NAND2_X1 U14028 ( .A1(n20980), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11154) );
  NAND2_X1 U14029 ( .A1(n10728), .A2(n11154), .ZN(n11155) );
  AOI21_X1 U14030 ( .B1(n10788), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11155), .ZN(
        n11156) );
  OAI21_X1 U14031 ( .B1(n11157), .B2(n11199), .A(n11156), .ZN(n11164) );
  INV_X1 U14032 ( .A(n11158), .ZN(n11159) );
  INV_X1 U14033 ( .A(n11160), .ZN(n11161) );
  INV_X1 U14034 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14886) );
  NAND2_X1 U14035 ( .A1(n11161), .A2(n14886), .ZN(n11162) );
  NAND2_X1 U14036 ( .A1(n11201), .A2(n11162), .ZN(n14884) );
  OR2_X1 U14037 ( .A1(n14884), .A2(n10728), .ZN(n11163) );
  NOR2_X1 U14038 ( .A1(n11166), .A2(n11165), .ZN(n11195) );
  AOI22_X1 U14039 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9864), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11170) );
  AOI22_X1 U14040 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U14041 ( .A1(n9853), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U14042 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11167) );
  NAND4_X1 U14043 ( .A1(n11170), .A2(n11169), .A3(n11168), .A4(n11167), .ZN(
        n11176) );
  AOI22_X1 U14044 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11174) );
  AOI22_X1 U14045 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11173) );
  AOI22_X1 U14046 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14047 ( .A1(n9856), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10990), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11171) );
  NAND4_X1 U14048 ( .A1(n11174), .A2(n11173), .A3(n11172), .A4(n11171), .ZN(
        n11175) );
  OR2_X1 U14049 ( .A1(n11176), .A2(n11175), .ZN(n11194) );
  XNOR2_X1 U14050 ( .A(n11195), .B(n11194), .ZN(n11179) );
  INV_X1 U14051 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14873) );
  AOI21_X1 U14052 ( .B1(n14873), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11177) );
  AOI21_X1 U14053 ( .B1(n10788), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11177), .ZN(
        n11178) );
  OAI21_X1 U14054 ( .B1(n11179), .B2(n11199), .A(n11178), .ZN(n11181) );
  XNOR2_X1 U14055 ( .A(n11201), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14875) );
  NAND2_X1 U14056 ( .A1(n14875), .A2(n9819), .ZN(n11180) );
  NAND2_X1 U14057 ( .A1(n11181), .A2(n11180), .ZN(n14595) );
  AOI22_X1 U14058 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14059 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U14060 ( .A1(n9869), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10479), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14061 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11184) );
  NAND4_X1 U14062 ( .A1(n11187), .A2(n11186), .A3(n11185), .A4(n11184), .ZN(
        n11193) );
  AOI22_X1 U14063 ( .A1(n9864), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9850), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14064 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14065 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9834), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14066 ( .A1(n9862), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11188) );
  NAND4_X1 U14067 ( .A1(n11191), .A2(n11190), .A3(n11189), .A4(n11188), .ZN(
        n11192) );
  NOR2_X1 U14068 ( .A1(n11193), .A2(n11192), .ZN(n11207) );
  NAND2_X1 U14069 ( .A1(n11195), .A2(n11194), .ZN(n11206) );
  XNOR2_X1 U14070 ( .A(n11207), .B(n11206), .ZN(n11200) );
  NAND2_X1 U14071 ( .A1(n20980), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11196) );
  NAND2_X1 U14072 ( .A1(n10728), .A2(n11196), .ZN(n11197) );
  AOI21_X1 U14073 ( .B1(n10788), .B2(P1_EAX_REG_29__SCAN_IN), .A(n11197), .ZN(
        n11198) );
  OAI21_X1 U14074 ( .B1(n11200), .B2(n11199), .A(n11198), .ZN(n11205) );
  INV_X1 U14075 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14861) );
  NAND2_X1 U14076 ( .A1(n11202), .A2(n14861), .ZN(n11203) );
  NAND2_X1 U14077 ( .A1(n14859), .A2(n9819), .ZN(n11204) );
  NAND2_X1 U14078 ( .A1(n11205), .A2(n11204), .ZN(n14581) );
  NOR2_X1 U14079 ( .A1(n11207), .A2(n11206), .ZN(n11221) );
  AOI22_X1 U14080 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9865), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14081 ( .A1(n9850), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14082 ( .A1(n10717), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9862), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14083 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9856), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11209) );
  NAND4_X1 U14084 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11219) );
  AOI22_X1 U14085 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9869), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14086 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14087 ( .A1(n9851), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9855), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14088 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9834), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11214) );
  NAND4_X1 U14089 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(
        n11218) );
  NOR2_X1 U14090 ( .A1(n11219), .A2(n11218), .ZN(n11220) );
  XNOR2_X1 U14091 ( .A(n11221), .B(n11220), .ZN(n11223) );
  NAND2_X1 U14092 ( .A1(n11223), .A2(n11222), .ZN(n11228) );
  NAND2_X1 U14093 ( .A1(n20980), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11224) );
  NAND2_X1 U14094 ( .A1(n10728), .A2(n11224), .ZN(n11225) );
  AOI21_X1 U14095 ( .B1(n10788), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11225), .ZN(
        n11227) );
  XNOR2_X1 U14096 ( .A(n14303), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14851) );
  AOI21_X1 U14097 ( .B1(n11228), .B2(n11227), .A(n11226), .ZN(n14566) );
  AOI22_X1 U14098 ( .A1(n10788), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11229), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11230) );
  XNOR2_X1 U14099 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11242) );
  NAND2_X1 U14100 ( .A1(n21214), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11253) );
  NAND2_X1 U14101 ( .A1(n11242), .A2(n11241), .ZN(n11232) );
  NAND2_X1 U14102 ( .A1(n20850), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11231) );
  NAND2_X1 U14103 ( .A1(n11232), .A2(n11231), .ZN(n11244) );
  XNOR2_X1 U14104 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11243) );
  NAND2_X1 U14105 ( .A1(n11244), .A2(n11243), .ZN(n11234) );
  NAND2_X1 U14106 ( .A1(n20922), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11233) );
  NAND2_X1 U14107 ( .A1(n11234), .A2(n11233), .ZN(n11246) );
  XNOR2_X1 U14108 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11245) );
  NAND2_X1 U14109 ( .A1(n11246), .A2(n11245), .ZN(n11236) );
  NAND2_X1 U14110 ( .A1(n21205), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11235) );
  NOR2_X1 U14111 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14067), .ZN(
        n11237) );
  XNOR2_X1 U14112 ( .A(n11242), .B(n11241), .ZN(n11264) );
  XNOR2_X1 U14113 ( .A(n11244), .B(n11243), .ZN(n11278) );
  XNOR2_X1 U14114 ( .A(n11246), .B(n11245), .ZN(n11283) );
  NOR4_X1 U14115 ( .A1(n11287), .A2(n11264), .A3(n11278), .A4(n11283), .ZN(
        n11247) );
  NOR2_X1 U14116 ( .A1(n11251), .A2(n11247), .ZN(n13777) );
  NAND2_X1 U14117 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21224) );
  NAND2_X1 U14118 ( .A1(n13777), .A2(n21224), .ZN(n11429) );
  NOR2_X1 U14119 ( .A1(n20534), .A2(n11248), .ZN(n13770) );
  NAND4_X1 U14120 ( .A1(n14043), .A2(n13878), .A3(n13770), .A4(n10553), .ZN(
        n13873) );
  OR2_X1 U14121 ( .A1(n13852), .A2(n21132), .ZN(n11436) );
  AOI21_X1 U14122 ( .B1(n10556), .B2(n14309), .A(n11562), .ZN(n11421) );
  NAND2_X1 U14123 ( .A1(n11421), .A2(n14306), .ZN(n13837) );
  OAI21_X1 U14124 ( .B1(n11436), .B2(n11545), .A(n13837), .ZN(n13853) );
  INV_X1 U14125 ( .A(n11251), .ZN(n11250) );
  NAND2_X1 U14126 ( .A1(n11251), .A2(n11275), .ZN(n11295) );
  INV_X1 U14127 ( .A(n11255), .ZN(n11284) );
  INV_X1 U14128 ( .A(n11289), .ZN(n11252) );
  NAND2_X1 U14129 ( .A1(n11252), .A2(n11283), .ZN(n11282) );
  OAI21_X1 U14130 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21214), .A(
        n11253), .ZN(n11254) );
  INV_X1 U14131 ( .A(n11254), .ZN(n11258) );
  NAND2_X1 U14132 ( .A1(n11275), .A2(n11258), .ZN(n11256) );
  NAND2_X1 U14133 ( .A1(n11256), .A2(n11255), .ZN(n11260) );
  NAND2_X1 U14134 ( .A1(n10548), .A2(n20501), .ZN(n11257) );
  NAND2_X1 U14135 ( .A1(n11257), .A2(n13974), .ZN(n11272) );
  OAI211_X1 U14136 ( .C1(n10499), .C2(n14309), .A(n11272), .B(n11258), .ZN(
        n11259) );
  NAND2_X1 U14137 ( .A1(n11260), .A2(n11259), .ZN(n11267) );
  INV_X1 U14138 ( .A(n11267), .ZN(n11271) );
  NAND2_X1 U14139 ( .A1(n11275), .A2(n20517), .ZN(n11262) );
  NAND2_X1 U14140 ( .A1(n10548), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11261) );
  NAND2_X1 U14141 ( .A1(n11262), .A2(n11261), .ZN(n11263) );
  INV_X1 U14142 ( .A(n11268), .ZN(n11270) );
  INV_X1 U14143 ( .A(n11263), .ZN(n11266) );
  NAND2_X1 U14144 ( .A1(n11289), .A2(n11264), .ZN(n11265) );
  AOI22_X1 U14145 ( .A1(n11268), .A2(n11267), .B1(n11266), .B2(n11265), .ZN(
        n11269) );
  AOI21_X1 U14146 ( .B1(n11271), .B2(n11270), .A(n11269), .ZN(n11280) );
  INV_X1 U14147 ( .A(n11272), .ZN(n11276) );
  INV_X1 U14148 ( .A(n11275), .ZN(n11273) );
  NOR2_X1 U14149 ( .A1(n11273), .A2(n11278), .ZN(n11274) );
  AOI211_X1 U14150 ( .C1(n11289), .C2(n11278), .A(n11276), .B(n11274), .ZN(
        n11279) );
  NAND2_X1 U14151 ( .A1(n11276), .A2(n11275), .ZN(n11277) );
  OAI22_X1 U14152 ( .A1(n11280), .A2(n11279), .B1(n11278), .B2(n11277), .ZN(
        n11281) );
  AOI22_X1 U14153 ( .A1(n11284), .A2(n11283), .B1(n11282), .B2(n11281), .ZN(
        n11292) );
  INV_X1 U14154 ( .A(n11287), .ZN(n11285) );
  NOR2_X1 U14155 ( .A1(n11289), .A2(n11285), .ZN(n11291) );
  INV_X1 U14156 ( .A(n11286), .ZN(n11288) );
  NAND3_X1 U14157 ( .A1(n11289), .A2(n11288), .A3(n11287), .ZN(n11290) );
  OAI21_X1 U14158 ( .B1(n11292), .B2(n11291), .A(n11290), .ZN(n11293) );
  AOI21_X1 U14159 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20500), .A(
        n11293), .ZN(n11294) );
  NAND2_X1 U14160 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  INV_X1 U14161 ( .A(n14036), .ZN(n11310) );
  NOR4_X1 U14162 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11303) );
  NOR4_X1 U14163 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n11302) );
  NOR4_X1 U14164 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11301) );
  NOR4_X1 U14165 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11300) );
  AND4_X1 U14166 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n11308) );
  NOR4_X1 U14167 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n11306) );
  NOR4_X1 U14168 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n11305) );
  NOR4_X1 U14169 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n11304) );
  INV_X1 U14170 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21141) );
  AND4_X1 U14171 ( .A1(n11306), .A2(n11305), .A3(n11304), .A4(n21141), .ZN(
        n11307) );
  NAND2_X1 U14172 ( .A1(n11308), .A2(n11307), .ZN(n11309) );
  NAND2_X1 U14173 ( .A1(n11310), .A2(n20497), .ZN(n14805) );
  INV_X1 U14174 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16718) );
  NOR2_X1 U14175 ( .A1(n14805), .A2(n16718), .ZN(n11314) );
  AOI22_X1 U14176 ( .A1(n11311), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14801), .ZN(n11312) );
  INV_X1 U14177 ( .A(n11312), .ZN(n11313) );
  NOR2_X1 U14178 ( .A1(n11314), .A2(n11313), .ZN(n11315) );
  XNOR2_X1 U14179 ( .A(n11329), .B(n11328), .ZN(n11317) );
  OAI211_X1 U14180 ( .C1(n11317), .C2(n21231), .A(n13771), .B(n11248), .ZN(
        n11318) );
  INV_X1 U14181 ( .A(n11318), .ZN(n11319) );
  OAI21_X2 U14182 ( .B1(n11320), .B2(n13974), .A(n11319), .ZN(n11325) );
  NAND2_X1 U14183 ( .A1(n21207), .A2(n11422), .ZN(n11323) );
  NAND2_X1 U14184 ( .A1(n14309), .A2(n10546), .ZN(n11332) );
  OAI21_X1 U14185 ( .B1(n21231), .B2(n11329), .A(n11332), .ZN(n11321) );
  INV_X1 U14186 ( .A(n11321), .ZN(n11322) );
  NAND2_X1 U14187 ( .A1(n11323), .A2(n11322), .ZN(n20429) );
  NAND2_X1 U14188 ( .A1(n20429), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11324) );
  NAND2_X1 U14189 ( .A1(n14132), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11327) );
  INV_X1 U14190 ( .A(n11324), .ZN(n20430) );
  NAND2_X1 U14191 ( .A1(n11325), .A2(n20430), .ZN(n11326) );
  NAND2_X2 U14192 ( .A1(n11327), .A2(n11326), .ZN(n11336) );
  INV_X1 U14193 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20470) );
  INV_X1 U14194 ( .A(n11422), .ZN(n11386) );
  NAND2_X1 U14195 ( .A1(n11329), .A2(n11328), .ZN(n11330) );
  NAND2_X1 U14196 ( .A1(n11330), .A2(n11331), .ZN(n11348) );
  OAI21_X1 U14197 ( .B1(n11331), .B2(n11330), .A(n11348), .ZN(n11334) );
  INV_X1 U14198 ( .A(n21231), .ZN(n11379) );
  INV_X1 U14199 ( .A(n11332), .ZN(n11333) );
  AOI21_X1 U14200 ( .B1(n11334), .B2(n11379), .A(n11333), .ZN(n11335) );
  NAND2_X1 U14201 ( .A1(n11336), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11337) );
  INV_X1 U14202 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20455) );
  OR2_X1 U14203 ( .A1(n21200), .A2(n11386), .ZN(n11342) );
  INV_X1 U14204 ( .A(n11347), .ZN(n11339) );
  XNOR2_X1 U14205 ( .A(n11348), .B(n11339), .ZN(n11340) );
  NAND2_X1 U14206 ( .A1(n11340), .A2(n11379), .ZN(n11341) );
  NAND2_X1 U14207 ( .A1(n11342), .A2(n11341), .ZN(n14146) );
  NAND2_X1 U14208 ( .A1(n14147), .A2(n14146), .ZN(n11345) );
  NAND2_X1 U14209 ( .A1(n11343), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11344) );
  NAND2_X1 U14210 ( .A1(n11345), .A2(n11344), .ZN(n14174) );
  NAND2_X1 U14211 ( .A1(n11346), .A2(n11422), .ZN(n11351) );
  NAND2_X1 U14212 ( .A1(n11348), .A2(n11347), .ZN(n11367) );
  XNOR2_X1 U14213 ( .A(n11367), .B(n11365), .ZN(n11349) );
  NAND2_X1 U14214 ( .A1(n11349), .A2(n11379), .ZN(n11350) );
  NAND2_X1 U14215 ( .A1(n11351), .A2(n11350), .ZN(n11352) );
  INV_X1 U14216 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20441) );
  XNOR2_X1 U14217 ( .A(n11352), .B(n20441), .ZN(n14173) );
  NAND2_X1 U14218 ( .A1(n14174), .A2(n14173), .ZN(n11354) );
  NAND2_X1 U14219 ( .A1(n11352), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11353) );
  INV_X1 U14220 ( .A(n11365), .ZN(n11355) );
  OR2_X1 U14221 ( .A1(n11367), .A2(n11355), .ZN(n11357) );
  INV_X1 U14222 ( .A(n11364), .ZN(n11356) );
  XNOR2_X1 U14223 ( .A(n11357), .B(n11356), .ZN(n11358) );
  OAI22_X1 U14224 ( .A1(n11359), .A2(n11386), .B1(n11358), .B2(n21231), .ZN(
        n11361) );
  INV_X1 U14225 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11360) );
  XNOR2_X1 U14226 ( .A(n11361), .B(n11360), .ZN(n16217) );
  NAND2_X1 U14227 ( .A1(n11361), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11362) );
  NAND3_X1 U14228 ( .A1(n11389), .A2(n11422), .A3(n11363), .ZN(n11370) );
  NAND2_X1 U14229 ( .A1(n11365), .A2(n11364), .ZN(n11366) );
  OR2_X1 U14230 ( .A1(n11367), .A2(n11366), .ZN(n11375) );
  XNOR2_X1 U14231 ( .A(n11375), .B(n11376), .ZN(n11368) );
  NAND2_X1 U14232 ( .A1(n11368), .A2(n11379), .ZN(n11369) );
  AND2_X1 U14233 ( .A1(n11370), .A2(n11369), .ZN(n11371) );
  INV_X1 U14234 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16337) );
  NAND2_X1 U14235 ( .A1(n11371), .A2(n16337), .ZN(n16211) );
  INV_X1 U14236 ( .A(n11371), .ZN(n11372) );
  NAND2_X1 U14237 ( .A1(n11372), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16210) );
  INV_X1 U14238 ( .A(n11373), .ZN(n11374) );
  OR2_X1 U14239 ( .A1(n11374), .A2(n11386), .ZN(n11382) );
  INV_X1 U14240 ( .A(n11375), .ZN(n11377) );
  NAND2_X1 U14241 ( .A1(n11377), .A2(n11376), .ZN(n11391) );
  XNOR2_X1 U14242 ( .A(n11391), .B(n11378), .ZN(n11380) );
  NAND2_X1 U14243 ( .A1(n11380), .A2(n11379), .ZN(n11381) );
  NAND2_X1 U14244 ( .A1(n11382), .A2(n11381), .ZN(n16202) );
  OR2_X1 U14245 ( .A1(n16202), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11383) );
  NAND2_X1 U14246 ( .A1(n16204), .A2(n11383), .ZN(n11385) );
  NAND2_X1 U14247 ( .A1(n16202), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11384) );
  NOR2_X1 U14248 ( .A1(n11387), .A2(n11386), .ZN(n11388) );
  OR3_X1 U14249 ( .A1(n11391), .A2(n11390), .A3(n21231), .ZN(n11392) );
  NAND2_X1 U14250 ( .A1(n11407), .A2(n11392), .ZN(n14441) );
  AND2_X1 U14251 ( .A1(n14441), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11393) );
  OR2_X1 U14252 ( .A1(n14441), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11394) );
  INV_X1 U14253 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16332) );
  OR2_X1 U14254 ( .A1(n15002), .A2(n16332), .ZN(n11395) );
  NAND2_X1 U14255 ( .A1(n14999), .A2(n16332), .ZN(n11396) );
  INV_X1 U14256 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15112) );
  AND2_X1 U14257 ( .A1(n15002), .A2(n15112), .ZN(n11400) );
  INV_X1 U14258 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21526) );
  NAND2_X1 U14259 ( .A1(n15002), .A2(n21526), .ZN(n11397) );
  NAND2_X1 U14260 ( .A1(n14977), .A2(n11397), .ZN(n14991) );
  INV_X1 U14261 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16305) );
  NAND2_X1 U14262 ( .A1(n14999), .A2(n16305), .ZN(n14990) );
  NAND2_X1 U14263 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11398) );
  NAND2_X1 U14264 ( .A1(n14999), .A2(n11398), .ZN(n14987) );
  NAND2_X1 U14265 ( .A1(n14990), .A2(n14987), .ZN(n11399) );
  XNOR2_X1 U14266 ( .A(n15002), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14967) );
  INV_X1 U14267 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15114) );
  NAND2_X1 U14268 ( .A1(n14999), .A2(n15114), .ZN(n15106) );
  INV_X1 U14269 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16262) );
  INV_X1 U14270 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11401) );
  NAND2_X1 U14271 ( .A1(n11402), .A2(n11401), .ZN(n11404) );
  NAND2_X1 U14272 ( .A1(n16173), .A2(n14999), .ZN(n11403) );
  OR2_X1 U14273 ( .A1(n15002), .A2(n16305), .ZN(n14989) );
  NOR2_X1 U14274 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11405) );
  OR2_X1 U14275 ( .A1(n15002), .A2(n11405), .ZN(n14985) );
  NAND2_X1 U14276 ( .A1(n14989), .A2(n14985), .ZN(n14976) );
  OR2_X1 U14277 ( .A1(n15002), .A2(n15114), .ZN(n15107) );
  OAI211_X1 U14278 ( .C1(n15002), .C2(n15112), .A(n15107), .B(n14977), .ZN(
        n11406) );
  NOR2_X1 U14279 ( .A1(n14976), .A2(n11406), .ZN(n16172) );
  XNOR2_X1 U14280 ( .A(n15002), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14954) );
  AND2_X1 U14281 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15087) );
  NAND2_X1 U14282 ( .A1(n14931), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11411) );
  NAND2_X1 U14283 ( .A1(n14891), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11413) );
  NAND3_X1 U14284 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15048) );
  NOR2_X2 U14285 ( .A1(n11413), .A2(n15048), .ZN(n14878) );
  AND2_X1 U14286 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11595) );
  NAND2_X1 U14287 ( .A1(n14878), .A2(n11595), .ZN(n14858) );
  INV_X1 U14288 ( .A(n14858), .ZN(n11408) );
  NAND3_X1 U14289 ( .A1(n11408), .A2(n11407), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14848) );
  NAND2_X1 U14290 ( .A1(n14848), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11417) );
  INV_X1 U14291 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14940) );
  INV_X1 U14292 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14949) );
  INV_X1 U14293 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16246) );
  INV_X1 U14294 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16225) );
  NAND4_X1 U14295 ( .A1(n14940), .A2(n14949), .A3(n16246), .A4(n16225), .ZN(
        n11410) );
  INV_X1 U14296 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15076) );
  INV_X1 U14297 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15055) );
  INV_X1 U14298 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15065) );
  NAND2_X1 U14299 ( .A1(n15055), .A2(n15065), .ZN(n11412) );
  NAND2_X1 U14300 ( .A1(n14893), .A2(n11413), .ZN(n14880) );
  INV_X1 U14301 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14881) );
  INV_X1 U14302 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14869) );
  NAND2_X1 U14303 ( .A1(n14881), .A2(n14869), .ZN(n15029) );
  INV_X1 U14304 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11415) );
  NAND2_X1 U14305 ( .A1(n14849), .A2(n11415), .ZN(n11416) );
  NAND2_X1 U14306 ( .A1(n11417), .A2(n11416), .ZN(n11419) );
  AND2_X1 U14307 ( .A1(n11421), .A2(n11561), .ZN(n11441) );
  OR2_X1 U14308 ( .A1(n11420), .A2(n11441), .ZN(n11425) );
  NAND2_X1 U14309 ( .A1(n11422), .A2(n10542), .ZN(n11555) );
  AND2_X1 U14310 ( .A1(n11555), .A2(n20501), .ZN(n11423) );
  NAND2_X1 U14311 ( .A1(n11424), .A2(n11423), .ZN(n11568) );
  NAND2_X1 U14312 ( .A1(n11425), .A2(n11568), .ZN(n13847) );
  INV_X1 U14313 ( .A(n11555), .ZN(n11426) );
  NAND2_X1 U14314 ( .A1(n16010), .A2(n11426), .ZN(n11433) );
  INV_X1 U14315 ( .A(n11427), .ZN(n11428) );
  NAND2_X1 U14316 ( .A1(n11428), .A2(n21136), .ZN(n16066) );
  NAND2_X1 U14317 ( .A1(n20517), .A2(n16066), .ZN(n11431) );
  INV_X1 U14318 ( .A(n11429), .ZN(n11430) );
  NAND3_X1 U14319 ( .A1(n11431), .A2(n20523), .A3(n11430), .ZN(n11432) );
  NAND2_X1 U14320 ( .A1(n11433), .A2(n11432), .ZN(n11434) );
  INV_X1 U14321 ( .A(n20251), .ZN(n13876) );
  OAI21_X1 U14322 ( .B1(n13847), .B2(n11434), .A(n13876), .ZN(n11440) );
  INV_X1 U14323 ( .A(n16066), .ZN(n21230) );
  OR2_X1 U14324 ( .A1(n20517), .A2(n21230), .ZN(n14308) );
  INV_X1 U14325 ( .A(n14308), .ZN(n11435) );
  OAI211_X1 U14326 ( .C1(n11436), .C2(n11435), .A(n20501), .B(n10549), .ZN(
        n11437) );
  NAND3_X1 U14327 ( .A1(n14120), .A2(n11438), .A3(n11437), .ZN(n11439) );
  INV_X1 U14328 ( .A(n10499), .ZN(n11565) );
  INV_X1 U14329 ( .A(n16032), .ZN(n11442) );
  OAI211_X1 U14330 ( .C1(n10543), .C2(n10209), .A(n11442), .B(n13837), .ZN(
        n11444) );
  NOR2_X1 U14331 ( .A1(n11444), .A2(n11443), .ZN(n11445) );
  INV_X1 U14332 ( .A(n10546), .ZN(n11446) );
  NAND2_X1 U14333 ( .A1(n11446), .A2(n20501), .ZN(n11513) );
  INV_X1 U14334 ( .A(n11447), .ZN(n11476) );
  INV_X1 U14335 ( .A(n10210), .ZN(n11545) );
  AND2_X1 U14336 ( .A1(n11545), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11448) );
  AOI21_X1 U14337 ( .B1(n14138), .B2(P1_EBX_REG_30__SCAN_IN), .A(n11448), .ZN(
        n14570) );
  INV_X1 U14338 ( .A(n11476), .ZN(n11548) );
  INV_X1 U14339 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14133) );
  NAND2_X1 U14340 ( .A1(n11513), .A2(n14133), .ZN(n11452) );
  INV_X1 U14341 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U14342 ( .A1(n10210), .A2(n11450), .ZN(n11451) );
  NAND3_X1 U14343 ( .A1(n11452), .A2(n11451), .A3(n11525), .ZN(n11453) );
  OAI21_X1 U14344 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(n11544), .A(n11453), .ZN(
        n11456) );
  NAND2_X1 U14345 ( .A1(n11513), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11455) );
  INV_X1 U14346 ( .A(n11476), .ZN(n11525) );
  INV_X1 U14347 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14144) );
  NAND2_X1 U14348 ( .A1(n11525), .A2(n14144), .ZN(n11454) );
  NAND2_X1 U14349 ( .A1(n11455), .A2(n11454), .ZN(n14139) );
  XNOR2_X1 U14350 ( .A(n11456), .B(n14139), .ZN(n14538) );
  NAND2_X1 U14351 ( .A1(n14538), .A2(n10210), .ZN(n13880) );
  NAND2_X1 U14352 ( .A1(n13880), .A2(n11456), .ZN(n14024) );
  INV_X1 U14353 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U14354 ( .A1(n11531), .A2(n11457), .ZN(n11461) );
  NAND2_X1 U14355 ( .A1(n11513), .A2(n20470), .ZN(n11459) );
  NAND2_X1 U14356 ( .A1(n10210), .A2(n11457), .ZN(n11458) );
  NAND3_X1 U14357 ( .A1(n11459), .A2(n11458), .A3(n11525), .ZN(n11460) );
  AND2_X1 U14358 ( .A1(n11461), .A2(n11460), .ZN(n14023) );
  MUX2_X1 U14359 ( .A(n11539), .B(n11525), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11462) );
  OAI21_X1 U14360 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14138), .A(
        n11462), .ZN(n14085) );
  INV_X1 U14361 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n11463) );
  NAND2_X1 U14362 ( .A1(n11531), .A2(n11463), .ZN(n11467) );
  NAND2_X1 U14363 ( .A1(n11525), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11464) );
  NAND2_X1 U14364 ( .A1(n11513), .A2(n11464), .ZN(n11465) );
  OAI21_X1 U14365 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n11545), .A(n11465), .ZN(
        n11466) );
  OR2_X1 U14366 ( .A1(n11539), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14367 ( .A1(n11525), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11468) );
  OAI211_X1 U14368 ( .C1(n11545), .C2(P1_EBX_REG_5__SCAN_IN), .A(n11513), .B(
        n11468), .ZN(n11469) );
  INV_X1 U14369 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U14370 ( .A1(n11531), .A2(n11471), .ZN(n11475) );
  NAND2_X1 U14371 ( .A1(n11525), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11472) );
  NAND2_X1 U14372 ( .A1(n11513), .A2(n11472), .ZN(n11473) );
  OAI21_X1 U14373 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n11545), .A(n11473), .ZN(
        n11474) );
  OR2_X1 U14374 ( .A1(n11539), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11479) );
  NAND2_X1 U14375 ( .A1(n11525), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11477) );
  OAI211_X1 U14376 ( .C1(n11545), .C2(P1_EBX_REG_7__SCAN_IN), .A(n11513), .B(
        n11477), .ZN(n11478) );
  NAND2_X1 U14377 ( .A1(n11479), .A2(n11478), .ZN(n14341) );
  NAND2_X1 U14378 ( .A1(n11525), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11480) );
  NAND2_X1 U14379 ( .A1(n11513), .A2(n11480), .ZN(n11482) );
  OR2_X1 U14380 ( .A1(n11545), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14381 ( .A1(n11482), .A2(n11481), .ZN(n11483) );
  OAI21_X1 U14382 ( .B1(n11544), .B2(P1_EBX_REG_8__SCAN_IN), .A(n11483), .ZN(
        n14364) );
  OR2_X1 U14383 ( .A1(n11539), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n11486) );
  NAND2_X1 U14384 ( .A1(n11525), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11484) );
  OAI211_X1 U14385 ( .C1(n11545), .C2(P1_EBX_REG_9__SCAN_IN), .A(n11513), .B(
        n11484), .ZN(n11485) );
  NAND2_X1 U14386 ( .A1(n11486), .A2(n11485), .ZN(n14418) );
  INV_X1 U14387 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14464) );
  NAND2_X1 U14388 ( .A1(n11531), .A2(n14464), .ZN(n11490) );
  INV_X1 U14389 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16325) );
  NAND2_X1 U14390 ( .A1(n11513), .A2(n16325), .ZN(n11488) );
  NAND2_X1 U14391 ( .A1(n10210), .A2(n14464), .ZN(n11487) );
  NAND3_X1 U14392 ( .A1(n11488), .A2(n11487), .A3(n11525), .ZN(n11489) );
  OR2_X1 U14393 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11492) );
  MUX2_X1 U14394 ( .A(n11539), .B(n11525), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11491) );
  NAND2_X1 U14395 ( .A1(n11525), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11493) );
  NAND2_X1 U14396 ( .A1(n11513), .A2(n11493), .ZN(n11495) );
  OR2_X1 U14397 ( .A1(n11545), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U14398 ( .A1(n11495), .A2(n11494), .ZN(n11496) );
  OAI21_X1 U14399 ( .B1(n11544), .B2(P1_EBX_REG_12__SCAN_IN), .A(n11496), .ZN(
        n14496) );
  MUX2_X1 U14400 ( .A(n11539), .B(n11548), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11498) );
  OR2_X1 U14401 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11497) );
  NAND2_X1 U14402 ( .A1(n11498), .A2(n11497), .ZN(n14518) );
  INV_X1 U14403 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n21404) );
  NAND2_X1 U14404 ( .A1(n11531), .A2(n21404), .ZN(n11502) );
  NAND2_X1 U14405 ( .A1(n11513), .A2(n15112), .ZN(n11500) );
  NAND2_X1 U14406 ( .A1(n10210), .A2(n21404), .ZN(n11499) );
  NAND3_X1 U14407 ( .A1(n11500), .A2(n11499), .A3(n11548), .ZN(n11501) );
  MUX2_X1 U14408 ( .A(n11539), .B(n11548), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11504) );
  OR2_X1 U14409 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11503) );
  NAND2_X1 U14410 ( .A1(n11513), .A2(n16262), .ZN(n11506) );
  INV_X1 U14411 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14764) );
  NAND2_X1 U14412 ( .A1(n10210), .A2(n14764), .ZN(n11505) );
  NAND3_X1 U14413 ( .A1(n11506), .A2(n11505), .A3(n11548), .ZN(n11507) );
  OAI21_X1 U14414 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(n11544), .A(n11507), .ZN(
        n14761) );
  MUX2_X1 U14415 ( .A(n11539), .B(n11525), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11509) );
  OR2_X1 U14416 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14417 ( .A1(n11509), .A2(n11508), .ZN(n14756) );
  OR2_X1 U14418 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11512) );
  INV_X1 U14419 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n11510) );
  MUX2_X1 U14420 ( .A(n11525), .B(n11539), .S(n11510), .Z(n11511) );
  AND2_X1 U14421 ( .A1(n11512), .A2(n11511), .ZN(n14743) );
  NAND2_X1 U14422 ( .A1(n11513), .A2(n16246), .ZN(n11515) );
  INV_X1 U14423 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14750) );
  NAND2_X1 U14424 ( .A1(n10210), .A2(n14750), .ZN(n11514) );
  NAND3_X1 U14425 ( .A1(n11515), .A2(n11514), .A3(n11525), .ZN(n11516) );
  OAI21_X1 U14426 ( .B1(P1_EBX_REG_18__SCAN_IN), .B2(n11544), .A(n11516), .ZN(
        n14674) );
  NAND2_X1 U14427 ( .A1(n14743), .A2(n14674), .ZN(n11517) );
  MUX2_X1 U14428 ( .A(n11539), .B(n11525), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11519) );
  OR2_X1 U14429 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11518) );
  AND2_X1 U14430 ( .A1(n11519), .A2(n11518), .ZN(n14733) );
  NAND2_X1 U14431 ( .A1(n11548), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11520) );
  NAND2_X1 U14432 ( .A1(n11513), .A2(n11520), .ZN(n11522) );
  OR2_X1 U14433 ( .A1(n11545), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n11521) );
  NAND2_X1 U14434 ( .A1(n11522), .A2(n11521), .ZN(n11523) );
  OAI21_X1 U14435 ( .B1(n11544), .B2(P1_EBX_REG_20__SCAN_IN), .A(n11523), .ZN(
        n14741) );
  NAND2_X1 U14436 ( .A1(n14733), .A2(n14741), .ZN(n11524) );
  INV_X1 U14437 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16224) );
  NAND2_X1 U14438 ( .A1(n11513), .A2(n16224), .ZN(n11527) );
  INV_X1 U14439 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U14440 ( .A1(n10210), .A2(n16079), .ZN(n11526) );
  NAND3_X1 U14441 ( .A1(n11527), .A2(n11526), .A3(n11525), .ZN(n11528) );
  OAI21_X1 U14442 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(n11544), .A(n11528), .ZN(
        n14726) );
  MUX2_X1 U14443 ( .A(n11539), .B(n11525), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11530) );
  OR2_X1 U14444 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11529) );
  NAND2_X1 U14445 ( .A1(n11530), .A2(n11529), .ZN(n14664) );
  INV_X1 U14446 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14719) );
  NAND2_X1 U14447 ( .A1(n11531), .A2(n14719), .ZN(n11534) );
  NAND2_X1 U14448 ( .A1(n11513), .A2(n15065), .ZN(n11532) );
  OAI211_X1 U14449 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n11545), .A(n11532), .B(
        n11548), .ZN(n11533) );
  MUX2_X1 U14450 ( .A(n11539), .B(n11525), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11536) );
  OR2_X1 U14451 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11535) );
  AND2_X1 U14452 ( .A1(n11536), .A2(n11535), .ZN(n14642) );
  INV_X1 U14453 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14894) );
  NAND2_X1 U14454 ( .A1(n11513), .A2(n14894), .ZN(n11537) );
  OAI211_X1 U14455 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n11545), .A(n11537), .B(
        n11548), .ZN(n11538) );
  OAI21_X1 U14456 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(n11544), .A(n11538), .ZN(
        n14622) );
  MUX2_X1 U14457 ( .A(n11539), .B(n11525), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11541) );
  OR2_X1 U14458 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11540) );
  NAND2_X1 U14459 ( .A1(n11541), .A2(n11540), .ZN(n14609) );
  NAND2_X1 U14460 ( .A1(n11513), .A2(n14869), .ZN(n11542) );
  OAI211_X1 U14461 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n11545), .A(n11542), .B(
        n11548), .ZN(n11543) );
  OAI21_X1 U14462 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(n11544), .A(n11543), .ZN(
        n14600) );
  OR2_X1 U14463 ( .A1(n11545), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n11547) );
  OR2_X1 U14464 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11546) );
  NAND2_X1 U14465 ( .A1(n11546), .A2(n11547), .ZN(n14567) );
  MUX2_X1 U14466 ( .A(n11547), .B(n14567), .S(n11525), .Z(n14589) );
  MUX2_X1 U14467 ( .A(n14570), .B(n11548), .S(n14587), .Z(n11550) );
  AOI22_X1 U14468 ( .A1(n14138), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11545), .ZN(n11549) );
  XNOR2_X1 U14469 ( .A(n11550), .B(n11549), .ZN(n14710) );
  INV_X1 U14470 ( .A(n14710), .ZN(n11600) );
  OR2_X1 U14471 ( .A1(n11551), .A2(n20517), .ZN(n13939) );
  NAND2_X1 U14472 ( .A1(n11552), .A2(n10543), .ZN(n11553) );
  AND2_X1 U14473 ( .A1(n13939), .A2(n11553), .ZN(n11554) );
  NOR2_X1 U14474 ( .A1(n11556), .A2(n11555), .ZN(n13848) );
  INV_X1 U14475 ( .A(n13848), .ZN(n11557) );
  INV_X1 U14476 ( .A(n16333), .ZN(n20463) );
  NAND2_X1 U14477 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20439) );
  NOR2_X1 U14478 ( .A1(n11360), .A2(n20439), .ZN(n16334) );
  INV_X1 U14479 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20473) );
  OAI21_X1 U14480 ( .B1(n20473), .B2(n14133), .A(n20470), .ZN(n20460) );
  NAND2_X1 U14481 ( .A1(n16334), .A2(n20460), .ZN(n16317) );
  INV_X1 U14482 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21502) );
  INV_X1 U14483 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16343) );
  INV_X1 U14484 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16350) );
  NOR3_X1 U14485 ( .A1(n16343), .A2(n16350), .A3(n16337), .ZN(n16318) );
  NAND3_X1 U14486 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16318), .ZN(n16308) );
  NOR2_X1 U14487 ( .A1(n21502), .A2(n16308), .ZN(n16291) );
  NAND2_X1 U14488 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16291), .ZN(
        n11575) );
  NOR2_X1 U14489 ( .A1(n16317), .A2(n11575), .ZN(n11578) );
  NAND2_X1 U14490 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11578), .ZN(
        n16272) );
  NAND2_X1 U14491 ( .A1(n10542), .A2(n20523), .ZN(n11558) );
  NAND2_X1 U14492 ( .A1(n11558), .A2(n20550), .ZN(n11559) );
  OAI21_X1 U14493 ( .B1(n14043), .B2(n11559), .A(n20517), .ZN(n11560) );
  OAI21_X1 U14494 ( .B1(n11561), .B2(n11525), .A(n11560), .ZN(n11567) );
  NAND2_X1 U14495 ( .A1(n14138), .A2(n11562), .ZN(n11564) );
  OAI211_X1 U14496 ( .C1(n11565), .C2(n14319), .A(n11564), .B(n11563), .ZN(
        n11566) );
  NOR2_X1 U14497 ( .A1(n11567), .A2(n11566), .ZN(n11569) );
  OAI211_X1 U14498 ( .C1(n10560), .C2(n13768), .A(n11569), .B(n11568), .ZN(
        n13836) );
  OAI21_X1 U14499 ( .B1(n13833), .B2(n20501), .A(n11570), .ZN(n11571) );
  NOR2_X1 U14500 ( .A1(n13836), .A2(n11571), .ZN(n11572) );
  OR2_X2 U14501 ( .A1(n14124), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20447) );
  NAND2_X1 U14502 ( .A1(n11573), .A2(n20447), .ZN(n20484) );
  OAI21_X1 U14503 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15083), .A(
        n20484), .ZN(n20457) );
  AOI21_X1 U14504 ( .B1(n20463), .B2(n16272), .A(n20457), .ZN(n15110) );
  NAND2_X1 U14505 ( .A1(n16333), .A2(n15083), .ZN(n20472) );
  INV_X1 U14506 ( .A(n20472), .ZN(n11574) );
  NAND2_X1 U14507 ( .A1(n11420), .A2(n20517), .ZN(n16012) );
  NOR3_X1 U14508 ( .A1(n15114), .A2(n15112), .A3(n16262), .ZN(n16253) );
  NAND2_X1 U14509 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n16253), .ZN(
        n16252) );
  NOR2_X1 U14510 ( .A1(n16246), .A2(n16252), .ZN(n11593) );
  NAND2_X1 U14511 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11593), .ZN(
        n16235) );
  INV_X1 U14512 ( .A(n11575), .ZN(n11576) );
  AND3_X1 U14513 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n16334), .ZN(n16294) );
  NAND2_X1 U14514 ( .A1(n11576), .A2(n16294), .ZN(n16282) );
  OR2_X1 U14515 ( .A1(n16235), .A2(n16282), .ZN(n15085) );
  NAND2_X1 U14516 ( .A1(n20474), .A2(n15085), .ZN(n11577) );
  NAND2_X1 U14517 ( .A1(n15110), .A2(n11577), .ZN(n11581) );
  INV_X1 U14518 ( .A(n15083), .ZN(n11579) );
  NAND2_X1 U14519 ( .A1(n16283), .A2(n20484), .ZN(n20490) );
  INV_X1 U14520 ( .A(n11578), .ZN(n11591) );
  AND2_X1 U14521 ( .A1(n11581), .A2(n11580), .ZN(n16239) );
  INV_X1 U14522 ( .A(n15087), .ZN(n11582) );
  AND2_X1 U14523 ( .A1(n20474), .A2(n11582), .ZN(n11583) );
  AND2_X1 U14524 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16223) );
  INV_X1 U14525 ( .A(n16223), .ZN(n11584) );
  AND2_X1 U14526 ( .A1(n20474), .A2(n11584), .ZN(n11585) );
  NOR2_X1 U14527 ( .A1(n16229), .A2(n11585), .ZN(n15077) );
  NAND2_X1 U14528 ( .A1(n20463), .A2(n15076), .ZN(n11586) );
  NAND2_X1 U14529 ( .A1(n20474), .A2(n15048), .ZN(n11587) );
  AND2_X1 U14530 ( .A1(n15063), .A2(n11587), .ZN(n15047) );
  NAND2_X1 U14531 ( .A1(n15047), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15043) );
  INV_X1 U14532 ( .A(n11595), .ZN(n15028) );
  OR2_X1 U14533 ( .A1(n15043), .A2(n15028), .ZN(n11589) );
  INV_X1 U14534 ( .A(n15063), .ZN(n11588) );
  OR2_X1 U14535 ( .A1(n11588), .A2(n20474), .ZN(n15042) );
  NAND2_X1 U14536 ( .A1(n11589), .A2(n15042), .ZN(n15023) );
  AOI21_X1 U14537 ( .B1(n20474), .B2(n11414), .A(n11415), .ZN(n11590) );
  NAND2_X1 U14538 ( .A1(n15023), .A2(n11590), .ZN(n15014) );
  NAND3_X1 U14539 ( .A1(n15014), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15042), .ZN(n11598) );
  INV_X2 U14540 ( .A(n20447), .ZN(n20487) );
  NAND2_X1 U14541 ( .A1(n20487), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14842) );
  NOR2_X1 U14542 ( .A1(n16333), .A2(n11591), .ZN(n16234) );
  NAND2_X1 U14543 ( .A1(n16234), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11592) );
  NOR2_X1 U14544 ( .A1(n21526), .A2(n16282), .ZN(n15111) );
  NAND2_X1 U14545 ( .A1(n16283), .A2(n15083), .ZN(n20458) );
  NAND2_X1 U14546 ( .A1(n15111), .A2(n16299), .ZN(n15064) );
  NAND2_X1 U14547 ( .A1(n11592), .A2(n15064), .ZN(n16268) );
  AND3_X1 U14548 ( .A1(n11593), .A2(n15087), .A3(n16223), .ZN(n11594) );
  NAND2_X1 U14549 ( .A1(n16268), .A2(n11594), .ZN(n15075) );
  NAND2_X1 U14550 ( .A1(n11595), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11596) );
  NOR2_X1 U14551 ( .A1(n15039), .A2(n11596), .ZN(n15015) );
  NAND3_X1 U14552 ( .A1(n15015), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n11418), .ZN(n11597) );
  NAND3_X1 U14553 ( .A1(n11598), .A2(n14842), .A3(n11597), .ZN(n11599) );
  AOI21_X1 U14554 ( .B1(n11600), .B2(n20486), .A(n11599), .ZN(n11601) );
  OAI21_X1 U14555 ( .B1(n14847), .B2(n20449), .A(n11601), .ZN(P1_U3000) );
  AND2_X4 U14556 ( .A1(n11858), .A2(n11784), .ZN(n11703) );
  AOI22_X1 U14557 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11607) );
  AND2_X4 U14558 ( .A1(n11602), .A2(n15839), .ZN(n11705) );
  AND3_X4 U14559 ( .A1(n12135), .A2(n11603), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14560 ( .A1(n11705), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11861), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11606) );
  INV_X1 U14561 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15815) );
  AND2_X4 U14562 ( .A1(n15845), .A2(n15815), .ZN(n11710) );
  AND2_X4 U14563 ( .A1(n15845), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11709) );
  AOI22_X1 U14564 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11605) );
  NAND4_X1 U14565 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n11608) );
  NAND2_X1 U14566 ( .A1(n11608), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11615) );
  AOI22_X1 U14567 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14568 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14569 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11609) );
  NAND4_X1 U14570 ( .A1(n11612), .A2(n11611), .A3(n11610), .A4(n11609), .ZN(
        n11613) );
  NAND2_X1 U14571 ( .A1(n11613), .A2(n16617), .ZN(n11614) );
  NAND2_X2 U14572 ( .A1(n11615), .A2(n11614), .ZN(n11725) );
  AOI22_X1 U14573 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14574 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14575 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14576 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11616) );
  NAND4_X1 U14577 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11620) );
  NAND2_X1 U14578 ( .A1(n11620), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11627) );
  AOI22_X1 U14579 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14580 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14581 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11621) );
  NAND4_X1 U14582 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n11625) );
  NAND2_X1 U14583 ( .A1(n11625), .A2(n16617), .ZN(n11626) );
  NAND2_X2 U14584 ( .A1(n11627), .A2(n11626), .ZN(n11723) );
  INV_X1 U14585 ( .A(n12200), .ZN(n11641) );
  AOI22_X1 U14586 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14587 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14588 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14589 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U14590 ( .A1(n11632), .A2(n16617), .ZN(n11640) );
  AOI22_X1 U14591 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14592 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14593 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11635) );
  NAND2_X1 U14594 ( .A1(n11641), .A2(n19547), .ZN(n12199) );
  INV_X1 U14595 ( .A(n11723), .ZN(n11642) );
  NAND2_X1 U14596 ( .A1(n11642), .A2(n11725), .ZN(n11727) );
  AOI22_X1 U14597 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14598 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14599 ( .A1(n11709), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9858), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14600 ( .A1(n11866), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11643) );
  NAND4_X1 U14601 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11647) );
  AOI22_X1 U14602 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11704), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14603 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14604 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11649) );
  NAND4_X1 U14605 ( .A1(n11651), .A2(n11650), .A3(n11649), .A4(n11648), .ZN(
        n11652) );
  NAND2_X1 U14606 ( .A1(n11652), .A2(n16617), .ZN(n11653) );
  AOI21_X1 U14607 ( .B1(n12204), .B2(n11727), .A(n11655), .ZN(n11656) );
  NAND2_X1 U14608 ( .A1(n12199), .A2(n11656), .ZN(n12725) );
  AOI22_X1 U14609 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14610 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11657) );
  AND2_X1 U14611 ( .A1(n11657), .A2(n16617), .ZN(n11659) );
  AOI22_X1 U14612 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11658) );
  NAND4_X1 U14613 ( .A1(n11661), .A2(n11660), .A3(n11659), .A4(n11658), .ZN(
        n11668) );
  AOI22_X1 U14614 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11665) );
  NAND3_X1 U14615 ( .A1(n10385), .A2(n11666), .A3(n11665), .ZN(n11667) );
  NAND2_X1 U14616 ( .A1(n12725), .A2(n12727), .ZN(n11683) );
  AOI22_X1 U14617 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14618 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14619 ( .A1(n11709), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9858), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14620 ( .A1(n11866), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14621 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  NAND2_X1 U14622 ( .A1(n11673), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11680) );
  AOI22_X1 U14623 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14624 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14625 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14626 ( .A1(n11866), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9858), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11674) );
  NAND4_X1 U14627 ( .A1(n11677), .A2(n11676), .A3(n11675), .A4(n11674), .ZN(
        n11678) );
  NAND3_X1 U14628 ( .A1(n11683), .A2(n14199), .A3(n11682), .ZN(n11696) );
  AOI22_X1 U14629 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14630 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14631 ( .A1(n11703), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14632 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11684) );
  NAND4_X1 U14633 ( .A1(n11687), .A2(n11686), .A3(n11685), .A4(n11684), .ZN(
        n11688) );
  NAND2_X1 U14634 ( .A1(n11688), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11695) );
  AOI22_X1 U14635 ( .A1(n9858), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14636 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14637 ( .A1(n11709), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14638 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U14639 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11693) );
  NAND2_X1 U14640 ( .A1(n11693), .A2(n16617), .ZN(n11694) );
  INV_X2 U14641 ( .A(n11886), .ZN(n11852) );
  NAND2_X1 U14642 ( .A1(n12737), .A2(n12734), .ZN(n13622) );
  NAND2_X1 U14643 ( .A1(n11696), .A2(n13622), .ZN(n11739) );
  AOI22_X1 U14644 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11866), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14645 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14646 ( .A1(n11709), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11703), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14647 ( .A1(n9857), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11697) );
  NAND4_X1 U14648 ( .A1(n11700), .A2(n11699), .A3(n11698), .A4(n11697), .ZN(
        n11701) );
  NAND2_X1 U14649 ( .A1(n11701), .A2(n16617), .ZN(n11715) );
  AOI22_X1 U14650 ( .A1(n11861), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11705), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11706) );
  NAND3_X1 U14651 ( .A1(n11708), .A2(n11707), .A3(n11706), .ZN(n11713) );
  AOI22_X1 U14652 ( .A1(n11710), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11711) );
  NAND2_X1 U14653 ( .A1(n11715), .A2(n11714), .ZN(n11724) );
  INV_X2 U14654 ( .A(n11724), .ZN(n12730) );
  NAND2_X1 U14655 ( .A1(n11717), .A2(n11720), .ZN(n12179) );
  NAND2_X1 U14656 ( .A1(n12179), .A2(n12730), .ZN(n12464) );
  NAND2_X1 U14657 ( .A1(n12464), .A2(n14199), .ZN(n11718) );
  INV_X1 U14658 ( .A(n13220), .ZN(n12181) );
  NAND2_X1 U14659 ( .A1(n11718), .A2(n12181), .ZN(n11722) );
  INV_X1 U14660 ( .A(n11725), .ZN(n11719) );
  NAND2_X1 U14661 ( .A1(n11719), .A2(n12202), .ZN(n13626) );
  AND2_X2 U14662 ( .A1(n11721), .A2(n11720), .ZN(n11759) );
  INV_X1 U14663 ( .A(n11759), .ZN(n12194) );
  NAND2_X1 U14664 ( .A1(n11722), .A2(n12194), .ZN(n11738) );
  BUF_X2 U14665 ( .A(n11724), .Z(n11733) );
  NAND2_X1 U14666 ( .A1(n11727), .A2(n12727), .ZN(n11728) );
  NAND2_X1 U14667 ( .A1(n11729), .A2(n11728), .ZN(n11749) );
  INV_X1 U14668 ( .A(n11730), .ZN(n11731) );
  NAND2_X1 U14669 ( .A1(n11749), .A2(n11731), .ZN(n11735) );
  NAND2_X1 U14670 ( .A1(n11735), .A2(n11734), .ZN(n11736) );
  NAND2_X1 U14671 ( .A1(n11737), .A2(n11736), .ZN(n12733) );
  NAND3_X1 U14672 ( .A1(n11739), .A2(n11738), .A3(n12733), .ZN(n11772) );
  AND2_X2 U14673 ( .A1(n11772), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11783) );
  NAND2_X1 U14674 ( .A1(n11759), .A2(n14199), .ZN(n11740) );
  NAND2_X1 U14675 ( .A1(n12196), .A2(n11740), .ZN(n12462) );
  INV_X1 U14676 ( .A(n12462), .ZN(n11744) );
  INV_X1 U14677 ( .A(n12148), .ZN(n12735) );
  NAND2_X1 U14678 ( .A1(n12735), .A2(n11743), .ZN(n11754) );
  NAND2_X1 U14679 ( .A1(n11744), .A2(n11754), .ZN(n12456) );
  AOI21_X2 U14680 ( .B1(n11783), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11748), .ZN(n11764) );
  NAND2_X1 U14681 ( .A1(n11852), .A2(n12226), .ZN(n12472) );
  INV_X1 U14682 ( .A(n11749), .ZN(n11750) );
  INV_X1 U14683 ( .A(n12458), .ZN(n11753) );
  NAND2_X1 U14684 ( .A1(n11753), .A2(n11752), .ZN(n11776) );
  OAI211_X1 U14685 ( .C1(n12181), .C2(n12194), .A(n12196), .B(n11754), .ZN(
        n11755) );
  NAND2_X1 U14686 ( .A1(n11755), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11756) );
  NAND2_X1 U14687 ( .A1(n11789), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11761) );
  NAND2_X1 U14688 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11760) );
  OAI211_X1 U14689 ( .C1(n11801), .C2(n15193), .A(n11761), .B(n11760), .ZN(
        n11762) );
  AOI21_X1 U14690 ( .B1(n11787), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11762), .ZN(n11763) );
  NAND2_X1 U14691 ( .A1(n11764), .A2(n11763), .ZN(n11782) );
  INV_X1 U14692 ( .A(n11814), .ZN(n11781) );
  INV_X1 U14693 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U14694 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11766) );
  AND2_X1 U14695 ( .A1(n16651), .A2(n11766), .ZN(n11768) );
  NAND2_X1 U14696 ( .A1(n11789), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11767) );
  OAI211_X1 U14697 ( .C1(n11801), .C2(n11769), .A(n11768), .B(n11767), .ZN(
        n11770) );
  AOI21_X1 U14698 ( .B1(n11787), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11770), .ZN(n11771) );
  BUF_X1 U14699 ( .A(n11772), .Z(n11775) );
  NAND2_X1 U14700 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n11773) );
  NAND2_X1 U14701 ( .A1(n11801), .A2(n11773), .ZN(n11774) );
  INV_X1 U14702 ( .A(n11776), .ZN(n11778) );
  NOR2_X1 U14703 ( .A1(n16651), .A2(n20233), .ZN(n11777) );
  NOR2_X1 U14704 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  NAND2_X2 U14705 ( .A1(n11781), .A2(n11811), .ZN(n11816) );
  OAI21_X1 U14706 ( .B1(n21487), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15818), 
        .ZN(n11785) );
  INV_X1 U14707 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11792) );
  NAND2_X1 U14708 ( .A1(n11789), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11791) );
  NAND2_X1 U14709 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11790) );
  OAI211_X1 U14710 ( .C1(n11801), .C2(n11792), .A(n11791), .B(n11790), .ZN(
        n11793) );
  AOI21_X1 U14711 ( .B1(n12389), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11793), .ZN(n11795) );
  NAND2_X1 U14712 ( .A1(n11794), .A2(n11795), .ZN(n11799) );
  INV_X1 U14713 ( .A(n11794), .ZN(n11797) );
  INV_X1 U14714 ( .A(n11795), .ZN(n11796) );
  NAND2_X1 U14715 ( .A1(n11797), .A2(n11796), .ZN(n11798) );
  OAI22_X1 U14716 ( .A1(n11800), .A2(n16617), .B1(n16651), .B2(n20209), .ZN(
        n11807) );
  NAND2_X1 U14717 ( .A1(n12389), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11805) );
  AOI22_X1 U14718 ( .A1(n11789), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11803) );
  NAND2_X1 U14719 ( .A1(n12379), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11802) );
  NAND2_X1 U14720 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  OR2_X1 U14721 ( .A1(n11807), .A2(n11806), .ZN(n12376) );
  NAND2_X1 U14722 ( .A1(n11807), .A2(n11806), .ZN(n11808) );
  XNOR2_X2 U14723 ( .A(n12375), .B(n12378), .ZN(n13288) );
  XNOR2_X2 U14724 ( .A(n11815), .B(n11820), .ZN(n15836) );
  AOI22_X1 U14725 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12015), .B1(
        n20022), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11838) );
  INV_X1 U14726 ( .A(n11817), .ZN(n11818) );
  NOR2_X1 U14727 ( .A1(n11816), .A2(n11818), .ZN(n11827) );
  INV_X1 U14728 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11819) );
  AND2_X1 U14729 ( .A1(n11820), .A2(n19365), .ZN(n11829) );
  INV_X1 U14730 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12588) );
  NOR2_X1 U14731 ( .A1(n12017), .A2(n12588), .ZN(n11821) );
  NOR2_X1 U14732 ( .A1(n11822), .A2(n11821), .ZN(n11837) );
  NAND2_X1 U14733 ( .A1(n11844), .A2(n15197), .ZN(n11903) );
  INV_X1 U14734 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11823) );
  OR2_X1 U14735 ( .A1(n11903), .A2(n11823), .ZN(n11835) );
  INV_X1 U14736 ( .A(n11827), .ZN(n11824) );
  OR2_X1 U14737 ( .A1(n14338), .A2(n11824), .ZN(n11825) );
  NAND2_X1 U14738 ( .A1(n14338), .A2(n11829), .ZN(n11826) );
  NAND2_X1 U14739 ( .A1(n14338), .A2(n11827), .ZN(n11828) );
  INV_X1 U14740 ( .A(n12007), .ZN(n19775) );
  INV_X1 U14741 ( .A(n11829), .ZN(n11830) );
  OR2_X1 U14742 ( .A1(n14338), .A2(n11830), .ZN(n11831) );
  AOI22_X1 U14743 ( .A1(n19775), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n19579), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11833) );
  NAND3_X1 U14744 ( .A1(n11838), .A2(n11837), .A3(n11836), .ZN(n11854) );
  INV_X1 U14745 ( .A(n11839), .ZN(n11846) );
  NOR2_X1 U14746 ( .A1(n14338), .A2(n15197), .ZN(n11847) );
  NAND2_X1 U14747 ( .A1(n11846), .A2(n11847), .ZN(n19623) );
  INV_X1 U14748 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13506) );
  NOR2_X1 U14749 ( .A1(n14338), .A2(n15836), .ZN(n11845) );
  INV_X1 U14750 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11869) );
  OAI22_X1 U14751 ( .A1(n19623), .A2(n13506), .B1(n19824), .B2(n11869), .ZN(
        n11843) );
  INV_X1 U14752 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12598) );
  INV_X1 U14753 ( .A(n19977), .ZN(n12003) );
  INV_X1 U14754 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11841) );
  OAI22_X1 U14755 ( .A1(n12598), .A2(n12003), .B1(n14262), .B2(n11841), .ZN(
        n11842) );
  NOR2_X1 U14756 ( .A1(n11843), .A2(n11842), .ZN(n11851) );
  INV_X1 U14757 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19545) );
  INV_X1 U14758 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13513) );
  OAI22_X1 U14759 ( .A1(n11899), .A2(n19545), .B1(n12016), .B2(n13513), .ZN(
        n11849) );
  AOI21_X1 U14760 ( .B1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n19736), .A(
        n11849), .ZN(n11850) );
  NAND2_X1 U14761 ( .A1(n11851), .A2(n11850), .ZN(n11853) );
  NOR2_X1 U14762 ( .A1(n15839), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11857) );
  AOI22_X1 U14763 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11913), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11865) );
  NOR2_X1 U14764 ( .A1(n15815), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11859) );
  AND2_X2 U14765 ( .A1(n13409), .A2(n11859), .ZN(n13305) );
  AOI22_X1 U14766 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12109), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11864) );
  INV_X1 U14767 ( .A(n11710), .ZN(n11860) );
  NAND2_X1 U14768 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11863) );
  NAND2_X1 U14769 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11862) );
  NAND4_X1 U14770 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11871) );
  INV_X2 U14771 ( .A(n13482), .ZN(n11872) );
  NAND2_X4 U14772 ( .A1(n11872), .A2(n16617), .ZN(n13447) );
  NAND2_X1 U14773 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11868) );
  INV_X2 U14774 ( .A(n13600), .ZN(n13591) );
  NAND2_X1 U14775 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11867) );
  OAI211_X1 U14776 ( .C1(n13447), .C2(n11869), .A(n11868), .B(n11867), .ZN(
        n11870) );
  NOR2_X1 U14777 ( .A1(n11871), .A2(n11870), .ZN(n11881) );
  NAND2_X1 U14778 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11876) );
  INV_X1 U14779 ( .A(n11709), .ZN(n13408) );
  NAND2_X1 U14780 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11875) );
  AND2_X2 U14781 ( .A1(n13608), .A2(n16617), .ZN(n13428) );
  NAND2_X1 U14782 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11874) );
  AND2_X2 U14783 ( .A1(n11872), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13429) );
  NAND2_X1 U14784 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11873) );
  NAND2_X1 U14785 ( .A1(n11704), .A2(n16617), .ZN(n12612) );
  INV_X1 U14786 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11879) );
  NAND2_X1 U14787 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11878) );
  NAND3_X1 U14788 ( .A1(n16615), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12190) );
  NAND2_X1 U14789 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11877) );
  OAI211_X1 U14790 ( .C1(n12612), .C2(n11879), .A(n11878), .B(n11877), .ZN(
        n11880) );
  INV_X1 U14791 ( .A(n12497), .ZN(n11882) );
  INV_X1 U14792 ( .A(n19824), .ZN(n11885) );
  NAND2_X1 U14793 ( .A1(n19708), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11888) );
  NAND2_X1 U14794 ( .A1(n19579), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11887) );
  NAND4_X1 U14795 ( .A1(n11889), .A2(n14211), .A3(n11888), .A4(n11887), .ZN(
        n11898) );
  NAND2_X1 U14796 ( .A1(n19977), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11894) );
  INV_X1 U14797 ( .A(n14262), .ZN(n11892) );
  NAND2_X1 U14798 ( .A1(n11892), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11893) );
  NAND4_X1 U14799 ( .A1(n11896), .A2(n11895), .A3(n11894), .A4(n11893), .ZN(
        n11897) );
  NOR2_X1 U14800 ( .A1(n11898), .A2(n11897), .ZN(n11907) );
  INV_X1 U14801 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13459) );
  INV_X1 U14802 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13466) );
  OAI22_X1 U14803 ( .A1(n19623), .A2(n13459), .B1(n12016), .B2(n13466), .ZN(
        n11902) );
  INV_X1 U14804 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14252) );
  INV_X1 U14805 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11900) );
  OAI22_X1 U14806 ( .A1(n11899), .A2(n14252), .B1(n19911), .B2(n11900), .ZN(
        n11901) );
  NOR2_X1 U14807 ( .A1(n11902), .A2(n11901), .ZN(n11906) );
  AOI22_X1 U14808 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19671), .B1(
        n19736), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14809 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12015), .B1(
        n20022), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11904) );
  NAND4_X1 U14810 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11964) );
  AOI22_X1 U14811 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12595), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U14812 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13444), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14813 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13429), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11910) );
  INV_X1 U14814 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14235) );
  INV_X1 U14815 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13316) );
  OAI22_X1 U14816 ( .A1(n13371), .A2(n14235), .B1(n12690), .B2(n13316), .ZN(
        n11908) );
  INV_X1 U14817 ( .A(n11908), .ZN(n11909) );
  NAND4_X1 U14818 ( .A1(n11912), .A2(n11911), .A3(n11910), .A4(n11909), .ZN(
        n11921) );
  AOI22_X1 U14819 ( .A1(n11913), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U14820 ( .A1(n12109), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11918) );
  INV_X1 U14821 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n19886) );
  INV_X1 U14822 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13413) );
  OAI22_X1 U14823 ( .A1(n13375), .A2(n19886), .B1(n12612), .B2(n13413), .ZN(
        n11915) );
  INV_X1 U14824 ( .A(n11915), .ZN(n11917) );
  AOI22_X1 U14825 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13438), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11916) );
  NAND4_X1 U14826 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11920) );
  OR2_X1 U14827 ( .A1(n13763), .A2(n14211), .ZN(n11970) );
  INV_X1 U14828 ( .A(n11970), .ZN(n11942) );
  AOI22_X1 U14829 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11913), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14830 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12109), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U14831 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U14832 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11922) );
  NAND4_X1 U14833 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11930) );
  NAND2_X1 U14834 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11928) );
  NAND2_X1 U14835 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11927) );
  NAND2_X1 U14836 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11926) );
  NAND3_X1 U14837 ( .A1(n11928), .A2(n11927), .A3(n11926), .ZN(n11929) );
  NOR2_X1 U14838 ( .A1(n11930), .A2(n11929), .ZN(n11941) );
  NAND2_X1 U14839 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U14840 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U14841 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11932) );
  NAND2_X1 U14842 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11931) );
  NAND4_X1 U14843 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11939) );
  INV_X1 U14844 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11937) );
  NAND2_X1 U14845 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11936) );
  NAND2_X1 U14846 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11935) );
  OAI211_X1 U14847 ( .C1(n12612), .C2(n11937), .A(n11936), .B(n11935), .ZN(
        n11938) );
  NOR2_X1 U14848 ( .A1(n11939), .A2(n11938), .ZN(n11940) );
  INV_X1 U14849 ( .A(n12482), .ZN(n12221) );
  NAND2_X1 U14850 ( .A1(n11942), .A2(n12221), .ZN(n11969) );
  NAND2_X1 U14851 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11946) );
  NAND2_X1 U14852 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11945) );
  NAND2_X1 U14853 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11944) );
  NAND2_X1 U14854 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11943) );
  NAND4_X1 U14855 ( .A1(n11946), .A2(n11945), .A3(n11944), .A4(n11943), .ZN(
        n11951) );
  INV_X1 U14856 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11949) );
  NAND2_X1 U14857 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11948) );
  NAND2_X1 U14858 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11947) );
  OAI211_X1 U14859 ( .C1(n13447), .C2(n11949), .A(n11948), .B(n11947), .ZN(
        n11950) );
  NOR2_X1 U14860 ( .A1(n11951), .A2(n11950), .ZN(n11962) );
  AOI22_X1 U14861 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11913), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U14862 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12109), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11954) );
  NAND2_X1 U14863 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11953) );
  NAND2_X1 U14864 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11952) );
  NAND4_X1 U14865 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n11960) );
  INV_X1 U14866 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11958) );
  NAND2_X1 U14867 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11957) );
  NAND2_X1 U14868 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11956) );
  OAI211_X1 U14869 ( .C1(n12612), .C2(n11958), .A(n11957), .B(n11956), .ZN(
        n11959) );
  NOR2_X1 U14870 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  NAND2_X1 U14871 ( .A1(n11969), .A2(n12489), .ZN(n11963) );
  XOR2_X1 U14872 ( .A(n12489), .B(n11969), .Z(n13797) );
  NAND2_X1 U14873 ( .A1(n11970), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13762) );
  XNOR2_X1 U14874 ( .A(n13763), .B(n12482), .ZN(n11971) );
  NOR2_X1 U14875 ( .A1(n13762), .A2(n11971), .ZN(n11972) );
  INV_X1 U14876 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15833) );
  XNOR2_X1 U14877 ( .A(n13762), .B(n11971), .ZN(n13820) );
  NOR2_X1 U14878 ( .A1(n15833), .A2(n13820), .ZN(n13819) );
  NOR2_X1 U14879 ( .A1(n11972), .A2(n13819), .ZN(n11973) );
  XOR2_X1 U14880 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11973), .Z(
        n13796) );
  NOR2_X1 U14881 ( .A1(n13797), .A2(n13796), .ZN(n13795) );
  INV_X1 U14882 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19537) );
  NOR2_X1 U14883 ( .A1(n11973), .A2(n19537), .ZN(n11974) );
  OR2_X1 U14884 ( .A1(n13795), .A2(n11974), .ZN(n11975) );
  INV_X1 U14885 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16611) );
  XNOR2_X1 U14886 ( .A(n11975), .B(n16611), .ZN(n16556) );
  NAND2_X1 U14887 ( .A1(n11975), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11976) );
  NAND2_X1 U14888 ( .A1(n16555), .A2(n11976), .ZN(n11998) );
  AOI22_X1 U14889 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11913), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U14890 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12109), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11979) );
  NAND2_X1 U14891 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11978) );
  NAND2_X1 U14892 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11977) );
  AND4_X1 U14893 ( .A1(n11980), .A2(n11979), .A3(n11978), .A4(n11977), .ZN(
        n11995) );
  NAND2_X1 U14894 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U14895 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11983) );
  NAND2_X1 U14896 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11982) );
  NAND2_X1 U14897 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11981) );
  AND4_X1 U14898 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n11994) );
  INV_X1 U14899 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12611) );
  NAND2_X1 U14900 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11986) );
  NAND2_X1 U14901 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11985) );
  OAI211_X1 U14902 ( .C1(n13447), .C2(n12611), .A(n11986), .B(n11985), .ZN(
        n11987) );
  INV_X1 U14903 ( .A(n11987), .ZN(n11993) );
  INV_X1 U14904 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11990) );
  NAND2_X1 U14905 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11989) );
  NAND2_X1 U14906 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11988) );
  OAI211_X1 U14907 ( .C1(n11990), .C2(n12690), .A(n11989), .B(n11988), .ZN(
        n11991) );
  INV_X1 U14908 ( .A(n11991), .ZN(n11992) );
  NAND4_X1 U14909 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n12173) );
  INV_X1 U14910 ( .A(n12173), .ZN(n12502) );
  NAND2_X1 U14911 ( .A1(n11996), .A2(n12502), .ZN(n11997) );
  NAND2_X1 U14912 ( .A1(n12049), .A2(n11997), .ZN(n11999) );
  XNOR2_X1 U14913 ( .A(n11998), .B(n11999), .ZN(n19489) );
  INV_X1 U14914 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19502) );
  INV_X1 U14915 ( .A(n11998), .ZN(n12000) );
  NAND2_X1 U14916 ( .A1(n12000), .A2(n11999), .ZN(n12001) );
  INV_X1 U14917 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13555) );
  INV_X1 U14918 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12031) );
  OAI22_X1 U14919 ( .A1(n19623), .A2(n13555), .B1(n19824), .B2(n12031), .ZN(
        n12002) );
  AOI21_X1 U14920 ( .B1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B2(n19671), .A(
        n12002), .ZN(n12024) );
  INV_X1 U14921 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12645) );
  INV_X1 U14922 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12004) );
  OAI22_X1 U14923 ( .A1(n12645), .A2(n12003), .B1(n19911), .B2(n12004), .ZN(
        n12005) );
  INV_X1 U14924 ( .A(n12005), .ZN(n12014) );
  INV_X1 U14925 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12009) );
  INV_X1 U14926 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12008) );
  OAI22_X1 U14927 ( .A1(n12009), .A2(n12006), .B1(n12007), .B2(n12008), .ZN(
        n12010) );
  INV_X1 U14928 ( .A(n12010), .ZN(n12012) );
  AOI22_X1 U14929 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19579), .B1(
        n14202), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U14930 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19736), .B1(
        n12015), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12022) );
  INV_X1 U14931 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13900) );
  INV_X1 U14932 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13562) );
  OAI22_X1 U14933 ( .A1(n11899), .A2(n13900), .B1(n12016), .B2(n13562), .ZN(
        n12020) );
  INV_X1 U14934 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12636) );
  INV_X1 U14935 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12018) );
  OAI22_X1 U14936 ( .A1(n12636), .A2(n12017), .B1(n14262), .B2(n12018), .ZN(
        n12019) );
  NOR2_X1 U14937 ( .A1(n12020), .A2(n12019), .ZN(n12021) );
  NAND4_X1 U14938 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12046) );
  AOI22_X1 U14939 ( .A1(n11913), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U14940 ( .A1(n12109), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12027) );
  NAND2_X1 U14941 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12026) );
  NAND2_X1 U14942 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12025) );
  NAND4_X1 U14943 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12033) );
  NAND2_X1 U14944 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12030) );
  NAND2_X1 U14945 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12029) );
  OAI211_X1 U14946 ( .C1(n12031), .C2(n13447), .A(n12030), .B(n12029), .ZN(
        n12032) );
  NOR2_X1 U14947 ( .A1(n12033), .A2(n12032), .ZN(n12044) );
  NAND2_X1 U14948 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12037) );
  NAND2_X1 U14949 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12036) );
  NAND2_X1 U14950 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12035) );
  NAND2_X1 U14951 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12034) );
  NAND4_X1 U14952 ( .A1(n12037), .A2(n12036), .A3(n12035), .A4(n12034), .ZN(
        n12042) );
  INV_X1 U14953 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12040) );
  NAND2_X1 U14954 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12039) );
  NAND2_X1 U14955 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12038) );
  OAI211_X1 U14956 ( .C1(n12040), .C2(n12690), .A(n12039), .B(n12038), .ZN(
        n12041) );
  NOR2_X1 U14957 ( .A1(n12042), .A2(n12041), .ZN(n12043) );
  NAND2_X1 U14958 ( .A1(n11852), .A2(n12506), .ZN(n12045) );
  XNOR2_X1 U14959 ( .A(n12049), .B(n12050), .ZN(n12219) );
  INV_X1 U14960 ( .A(n12219), .ZN(n12047) );
  INV_X1 U14961 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14403) );
  INV_X1 U14962 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12052) );
  INV_X1 U14963 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12081) );
  OAI22_X1 U14964 ( .A1(n19623), .A2(n12052), .B1(n19824), .B2(n12081), .ZN(
        n12053) );
  AOI21_X1 U14965 ( .B1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n19671), .A(
        n12053), .ZN(n12070) );
  INV_X1 U14966 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12658) );
  INV_X1 U14967 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12054) );
  OAI22_X1 U14968 ( .A1(n12658), .A2(n12003), .B1(n14262), .B2(n12054), .ZN(
        n12055) );
  INV_X1 U14969 ( .A(n12055), .ZN(n12062) );
  NAND2_X1 U14970 ( .A1(n20022), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12061) );
  AOI22_X1 U14971 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19579), .B1(
        n14202), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12060) );
  INV_X1 U14972 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12057) );
  INV_X1 U14973 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12056) );
  OAI22_X1 U14974 ( .A1(n12057), .A2(n12006), .B1(n12007), .B2(n12056), .ZN(
        n12058) );
  INV_X1 U14975 ( .A(n12058), .ZN(n12059) );
  AOI22_X1 U14976 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19736), .B1(
        n12015), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12068) );
  INV_X1 U14977 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19565) );
  INV_X1 U14978 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13579) );
  OAI22_X1 U14979 ( .A1(n11899), .A2(n19565), .B1(n12016), .B2(n13579), .ZN(
        n12066) );
  INV_X1 U14980 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12064) );
  INV_X1 U14981 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12063) );
  OAI22_X1 U14982 ( .A1(n12064), .A2(n12017), .B1(n19911), .B2(n12063), .ZN(
        n12065) );
  NOR2_X1 U14983 ( .A1(n12066), .A2(n12065), .ZN(n12067) );
  NAND4_X1 U14984 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12093) );
  AOI22_X1 U14985 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11913), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U14986 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12109), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12073) );
  NAND2_X1 U14987 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12072) );
  NAND2_X1 U14988 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12071) );
  NAND2_X1 U14989 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12078) );
  NAND2_X1 U14990 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12077) );
  NAND2_X1 U14991 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12076) );
  NAND2_X1 U14992 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12075) );
  NAND2_X1 U14993 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12080) );
  NAND2_X1 U14994 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12079) );
  OAI211_X1 U14995 ( .C1(n13447), .C2(n12081), .A(n12080), .B(n12079), .ZN(
        n12082) );
  INV_X1 U14996 ( .A(n12082), .ZN(n12088) );
  INV_X1 U14997 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12085) );
  NAND2_X1 U14998 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12084) );
  NAND2_X1 U14999 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12083) );
  OAI211_X1 U15000 ( .C1(n12690), .C2(n12085), .A(n12084), .B(n12083), .ZN(
        n12086) );
  INV_X1 U15001 ( .A(n12086), .ZN(n12087) );
  NAND4_X1 U15002 ( .A1(n12090), .A2(n12089), .A3(n12088), .A4(n12087), .ZN(
        n12511) );
  INV_X1 U15003 ( .A(n12511), .ZN(n12091) );
  NAND2_X1 U15004 ( .A1(n12091), .A2(n11852), .ZN(n12092) );
  INV_X1 U15005 ( .A(n12250), .ZN(n12097) );
  INV_X1 U15006 ( .A(n12101), .ZN(n12095) );
  INV_X1 U15007 ( .A(n14398), .ZN(n12096) );
  NAND2_X1 U15008 ( .A1(n12098), .A2(n12250), .ZN(n12099) );
  INV_X1 U15009 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16596) );
  INV_X1 U15010 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12689) );
  INV_X1 U15011 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12681) );
  OAI22_X1 U15012 ( .A1(n12689), .A2(n12515), .B1(n13371), .B2(n12681), .ZN(
        n12105) );
  INV_X1 U15013 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13596) );
  INV_X1 U15014 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12103) );
  OAI22_X1 U15015 ( .A1(n13596), .A2(n13375), .B1(n13447), .B2(n12103), .ZN(
        n12104) );
  NOR2_X1 U15016 ( .A1(n12105), .A2(n12104), .ZN(n12121) );
  INV_X1 U15017 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13601) );
  NAND2_X1 U15018 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12107) );
  NAND2_X1 U15019 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12106) );
  OAI211_X1 U15020 ( .C1(n12612), .C2(n13601), .A(n12107), .B(n12106), .ZN(
        n12108) );
  INV_X1 U15021 ( .A(n12108), .ZN(n12120) );
  AOI22_X1 U15022 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11914), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15023 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11913), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12112) );
  NAND2_X1 U15024 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12111) );
  NAND2_X1 U15025 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12110) );
  INV_X1 U15026 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12116) );
  NAND2_X1 U15027 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12115) );
  NAND2_X1 U15028 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12114) );
  OAI211_X1 U15029 ( .C1(n12690), .C2(n12116), .A(n12115), .B(n12114), .ZN(
        n12117) );
  INV_X1 U15030 ( .A(n12117), .ZN(n12118) );
  XNOR2_X1 U15031 ( .A(n12124), .B(n12787), .ZN(n15546) );
  NAND2_X1 U15032 ( .A1(n12122), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12123) );
  NAND2_X1 U15033 ( .A1(n12126), .A2(n12787), .ZN(n12125) );
  NAND3_X1 U15034 ( .A1(n12126), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n12787), .ZN(n12127) );
  AND2_X1 U15035 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15734) );
  INV_X1 U15036 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16517) );
  INV_X1 U15037 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15783) );
  NOR2_X1 U15038 ( .A1(n16517), .A2(n15783), .ZN(n15782) );
  AND2_X1 U15039 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15782), .ZN(
        n15727) );
  NAND3_X1 U15040 ( .A1(n15734), .A2(n15727), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16564) );
  AND2_X1 U15041 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15510) );
  NAND2_X1 U15042 ( .A1(n15510), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12129) );
  NOR2_X1 U15043 ( .A1(n16564), .A2(n12129), .ZN(n15680) );
  INV_X1 U15044 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15678) );
  INV_X1 U15045 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15669) );
  INV_X1 U15046 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15645) );
  NAND2_X1 U15047 ( .A1(n12130), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15472) );
  INV_X1 U15048 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15636) );
  INV_X1 U15049 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15617) );
  INV_X1 U15050 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15596) );
  INV_X1 U15051 ( .A(n12815), .ZN(n12132) );
  INV_X1 U15052 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12779) );
  NOR2_X2 U15053 ( .A1(n12815), .A2(n12779), .ZN(n15410) );
  INV_X1 U15054 ( .A(n15410), .ZN(n12131) );
  OAI21_X1 U15055 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n12132), .A(
        n12131), .ZN(n15424) );
  NAND2_X1 U15056 ( .A1(n21540), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12134) );
  NAND2_X1 U15057 ( .A1(n15839), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12133) );
  NAND2_X1 U15058 ( .A1(n12134), .A2(n12133), .ZN(n12151) );
  NAND2_X1 U15059 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20233), .ZN(
        n12150) );
  NAND2_X1 U15060 ( .A1(n12135), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12136) );
  NAND2_X1 U15061 ( .A1(n12138), .A2(n12136), .ZN(n12146) );
  INV_X1 U15062 ( .A(n12146), .ZN(n12137) );
  NAND2_X1 U15063 ( .A1(n12147), .A2(n12137), .ZN(n12139) );
  INV_X1 U15064 ( .A(n12145), .ZN(n12140) );
  NOR2_X1 U15065 ( .A1(n21356), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12142) );
  NAND3_X1 U15066 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12143), .A3(
        n15989), .ZN(n12174) );
  XNOR2_X1 U15067 ( .A(n12145), .B(n12144), .ZN(n12175) );
  XNOR2_X1 U15068 ( .A(n12147), .B(n12146), .ZN(n12183) );
  AOI21_X1 U15069 ( .B1(n16637), .B2(n14211), .A(n12183), .ZN(n12158) );
  AND2_X1 U15070 ( .A1(n12362), .A2(n12183), .ZN(n12169) );
  INV_X1 U15071 ( .A(n12183), .ZN(n12156) );
  OAI21_X1 U15072 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20233), .A(
        n12150), .ZN(n12234) );
  OAI21_X1 U15073 ( .B1(n12234), .B2(n12151), .A(n13214), .ZN(n12155) );
  INV_X1 U15074 ( .A(n12234), .ZN(n12167) );
  NAND2_X1 U15075 ( .A1(n12151), .A2(n12150), .ZN(n12168) );
  NAND2_X1 U15076 ( .A1(n12152), .A2(n12168), .ZN(n12184) );
  INV_X1 U15077 ( .A(n12184), .ZN(n12153) );
  OAI211_X1 U15078 ( .C1(n14211), .C2(n12167), .A(n16637), .B(n12153), .ZN(
        n12154) );
  OAI211_X1 U15079 ( .C1(n16632), .C2(n12156), .A(n12155), .B(n12154), .ZN(
        n12157) );
  OAI211_X1 U15080 ( .C1(n12158), .C2(n12169), .A(n12182), .B(n12157), .ZN(
        n12159) );
  OAI21_X1 U15081 ( .B1(n12182), .B2(n12362), .A(n12159), .ZN(n12160) );
  OR2_X1 U15082 ( .A1(n12186), .A2(n12160), .ZN(n12161) );
  MUX2_X1 U15083 ( .A(n12161), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n16656), .Z(n12163) );
  AND2_X1 U15084 ( .A1(n14199), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13785) );
  NAND2_X1 U15085 ( .A1(n12186), .A2(n13785), .ZN(n12162) );
  NAND2_X1 U15086 ( .A1(n16642), .A2(n14211), .ZN(n13783) );
  INV_X1 U15087 ( .A(n12163), .ZN(n12164) );
  NAND2_X1 U15088 ( .A1(n13783), .A2(n12164), .ZN(n12165) );
  OAI21_X1 U15089 ( .B1(n16637), .B2(n16642), .A(n12165), .ZN(n12166) );
  NAND2_X1 U15090 ( .A1(n12166), .A2(n12204), .ZN(n12216) );
  AND2_X1 U15091 ( .A1(n12168), .A2(n12167), .ZN(n12176) );
  INV_X1 U15092 ( .A(n12169), .ZN(n12172) );
  NAND2_X1 U15093 ( .A1(n12170), .A2(n13214), .ZN(n12171) );
  NAND2_X1 U15094 ( .A1(n12172), .A2(n12171), .ZN(n12220) );
  MUX2_X1 U15095 ( .A(n12174), .B(n12173), .S(n13214), .Z(n12228) );
  OAI211_X1 U15096 ( .C1(n12176), .C2(n12220), .A(n12228), .B(n12225), .ZN(
        n12177) );
  INV_X1 U15097 ( .A(n12177), .ZN(n12178) );
  OR2_X1 U15098 ( .A1(n12178), .A2(n12186), .ZN(n20240) );
  OR2_X1 U15099 ( .A1(n12180), .A2(n12181), .ZN(n12218) );
  INV_X1 U15100 ( .A(n12180), .ZN(n12192) );
  NAND2_X1 U15101 ( .A1(n12183), .A2(n12182), .ZN(n12188) );
  NOR2_X1 U15102 ( .A1(n12184), .A2(n12188), .ZN(n12185) );
  OR2_X1 U15103 ( .A1(n12186), .A2(n12185), .ZN(n16638) );
  INV_X1 U15104 ( .A(n16638), .ZN(n12187) );
  OAI21_X1 U15105 ( .B1(n12234), .B2(n12188), .A(n12187), .ZN(n12189) );
  INV_X1 U15106 ( .A(n12189), .ZN(n12191) );
  NAND2_X1 U15107 ( .A1(n15989), .A2(n12190), .ZN(n15986) );
  INV_X1 U15108 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19174) );
  OAI21_X1 U15109 ( .B1(n13444), .B2(n15986), .A(n19174), .ZN(n16650) );
  MUX2_X1 U15110 ( .A(n12191), .B(n16650), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20236) );
  NAND3_X1 U15111 ( .A1(n12192), .A2(n14211), .A3(n20236), .ZN(n12193) );
  INV_X1 U15112 ( .A(n12194), .ZN(n16654) );
  NOR2_X1 U15113 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20121) );
  AOI211_X1 U15114 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n20121), .ZN(n20114) );
  NAND2_X1 U15115 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20108) );
  NAND2_X1 U15116 ( .A1(n20114), .A2(n20108), .ZN(n15820) );
  INV_X1 U15117 ( .A(n15820), .ZN(n16629) );
  NAND2_X1 U15118 ( .A1(n16654), .A2(n16629), .ZN(n12195) );
  OR2_X1 U15119 ( .A1(n16638), .A2(n12195), .ZN(n12210) );
  AND2_X1 U15120 ( .A1(n11727), .A2(n12204), .ZN(n12198) );
  OAI21_X1 U15121 ( .B1(n12198), .B2(n11733), .A(n12197), .ZN(n12208) );
  CLKBUF_X3 U15122 ( .A(n12202), .Z(n19570) );
  NAND2_X1 U15123 ( .A1(n12201), .A2(n19570), .ZN(n12203) );
  NAND2_X1 U15124 ( .A1(n12203), .A2(n13220), .ZN(n12726) );
  NAND2_X1 U15125 ( .A1(n11852), .A2(n12204), .ZN(n12747) );
  NAND2_X1 U15126 ( .A1(n12747), .A2(n16637), .ZN(n12205) );
  NAND3_X1 U15127 ( .A1(n12205), .A2(n12727), .A3(n19570), .ZN(n12206) );
  NAND2_X1 U15128 ( .A1(n12206), .A2(n12730), .ZN(n12207) );
  NAND4_X1 U15129 ( .A1(n12208), .A2(n12199), .A3(n12726), .A4(n12207), .ZN(
        n12748) );
  INV_X1 U15130 ( .A(n12748), .ZN(n12209) );
  NAND2_X1 U15131 ( .A1(n12210), .A2(n12209), .ZN(n15823) );
  MUX2_X1 U15132 ( .A(n16654), .B(n11733), .S(n11852), .Z(n12211) );
  NAND2_X1 U15133 ( .A1(n12211), .A2(n20108), .ZN(n12212) );
  NOR2_X1 U15134 ( .A1(n16638), .A2(n12212), .ZN(n12213) );
  NOR3_X1 U15135 ( .A1(n12791), .A2(n15823), .A3(n12213), .ZN(n12215) );
  INV_X1 U15136 ( .A(n13783), .ZN(n15822) );
  NAND3_X1 U15137 ( .A1(n15822), .A2(n11733), .A3(n16629), .ZN(n12214) );
  NAND3_X1 U15138 ( .A1(n12216), .A2(n12215), .A3(n12214), .ZN(n12217) );
  NOR2_X1 U15139 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16656), .ZN(n13216) );
  INV_X1 U15140 ( .A(n12218), .ZN(n20239) );
  NAND2_X1 U15141 ( .A1(n12219), .A2(n12320), .ZN(n12229) );
  NAND2_X1 U15142 ( .A1(n12221), .A2(n19552), .ZN(n12223) );
  NOR2_X1 U15143 ( .A1(n19552), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12235) );
  INV_X1 U15144 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n15193) );
  NAND2_X1 U15145 ( .A1(n12235), .A2(n15193), .ZN(n12222) );
  NAND2_X1 U15146 ( .A1(n12223), .A2(n12222), .ZN(n12241) );
  NAND2_X1 U15147 ( .A1(n12242), .A2(n12241), .ZN(n12240) );
  INV_X1 U15148 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12382) );
  MUX2_X1 U15149 ( .A(n12228), .B(n12382), .S(n12227), .Z(n12246) );
  MUX2_X1 U15150 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12506), .S(n19552), .Z(
        n12251) );
  XNOR2_X1 U15151 ( .A(n12252), .B(n12251), .ZN(n19350) );
  INV_X1 U15152 ( .A(n12247), .ZN(n12232) );
  NAND2_X1 U15153 ( .A1(n12230), .A2(n12240), .ZN(n12231) );
  NAND2_X1 U15154 ( .A1(n12232), .A2(n12231), .ZN(n15183) );
  MUX2_X1 U15155 ( .A(n12234), .B(n13763), .S(n13214), .Z(n12236) );
  AOI21_X1 U15156 ( .B1(n12236), .B2(n19552), .A(n12235), .ZN(n19366) );
  NAND2_X1 U15157 ( .A1(n19366), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13824) );
  NAND2_X1 U15158 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12237) );
  NOR2_X1 U15159 ( .A1(n19552), .A2(n12237), .ZN(n12238) );
  OR2_X1 U15160 ( .A1(n12241), .A2(n12238), .ZN(n15191) );
  NOR2_X1 U15161 ( .A1(n13824), .A2(n15191), .ZN(n12239) );
  NAND2_X1 U15162 ( .A1(n13824), .A2(n15191), .ZN(n13823) );
  OAI21_X1 U15163 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12239), .A(
        n13823), .ZN(n13801) );
  OAI21_X1 U15164 ( .B1(n12242), .B2(n12241), .A(n12240), .ZN(n14336) );
  XNOR2_X1 U15165 ( .A(n14336), .B(n19537), .ZN(n13800) );
  OR2_X1 U15166 ( .A1(n13801), .A2(n13800), .ZN(n19525) );
  INV_X1 U15167 ( .A(n14336), .ZN(n12243) );
  NAND2_X1 U15168 ( .A1(n12243), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12244) );
  NAND2_X1 U15169 ( .A1(n19525), .A2(n12244), .ZN(n16553) );
  INV_X1 U15170 ( .A(n16553), .ZN(n12245) );
  OAI21_X1 U15171 ( .B1(n12247), .B2(n12246), .A(n12252), .ZN(n14285) );
  XNOR2_X1 U15172 ( .A(n14285), .B(n19502), .ZN(n19491) );
  NAND2_X1 U15173 ( .A1(n12248), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12249) );
  NAND2_X1 U15174 ( .A1(n12250), .A2(n12320), .ZN(n12253) );
  INV_X1 U15175 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12388) );
  MUX2_X1 U15176 ( .A(n12388), .B(n12511), .S(n19552), .Z(n12257) );
  XNOR2_X1 U15177 ( .A(n12258), .B(n12257), .ZN(n19337) );
  NAND2_X1 U15178 ( .A1(n12253), .A2(n19337), .ZN(n12254) );
  INV_X1 U15179 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14431) );
  XNOR2_X1 U15180 ( .A(n12254), .B(n14431), .ZN(n14424) );
  NAND2_X1 U15181 ( .A1(n14423), .A2(n14424), .ZN(n12256) );
  NAND2_X1 U15182 ( .A1(n12254), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12255) );
  INV_X1 U15183 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12392) );
  MUX2_X1 U15184 ( .A(n12392), .B(n12787), .S(n19552), .Z(n12261) );
  NAND2_X1 U15185 ( .A1(n12227), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12259) );
  OR2_X1 U15186 ( .A1(n12270), .A2(n12259), .ZN(n12260) );
  NAND2_X1 U15187 ( .A1(n12269), .A2(n12260), .ZN(n14300) );
  NOR2_X1 U15188 ( .A1(n14300), .A2(n12320), .ZN(n12264) );
  AND2_X1 U15189 ( .A1(n12264), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16532) );
  NOR2_X1 U15190 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  OR2_X1 U15191 ( .A1(n12270), .A2(n12263), .ZN(n19327) );
  NOR2_X1 U15192 ( .A1(n19327), .A2(n16596), .ZN(n16528) );
  INV_X1 U15193 ( .A(n12264), .ZN(n12266) );
  INV_X1 U15194 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12265) );
  NAND2_X1 U15195 ( .A1(n12266), .A2(n12265), .ZN(n16530) );
  NAND2_X1 U15196 ( .A1(n19327), .A2(n16596), .ZN(n16529) );
  AND2_X1 U15197 ( .A1(n16530), .A2(n16529), .ZN(n12267) );
  NAND2_X1 U15198 ( .A1(n12227), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12268) );
  XNOR2_X1 U15199 ( .A(n12269), .B(n12268), .ZN(n19317) );
  NAND2_X1 U15200 ( .A1(n19317), .A2(n12787), .ZN(n12276) );
  INV_X1 U15201 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15725) );
  AND2_X1 U15202 ( .A1(n12276), .A2(n15725), .ZN(n13653) );
  NAND2_X2 U15203 ( .A1(n12270), .A2(n19552), .ZN(n12357) );
  NAND3_X1 U15204 ( .A1(n12272), .A2(n12227), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n12271) );
  OAI211_X1 U15205 ( .C1(n12272), .C2(P2_EBX_REG_10__SCAN_IN), .A(n12357), .B(
        n12271), .ZN(n19304) );
  OAI21_X1 U15206 ( .B1(n19304), .B2(n12320), .A(n16517), .ZN(n16512) );
  INV_X1 U15207 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n14159) );
  AND2_X1 U15208 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n9892), .ZN(n12273) );
  NAND2_X1 U15209 ( .A1(n12227), .A2(n12273), .ZN(n15171) );
  NAND2_X1 U15210 ( .A1(n15171), .A2(n12787), .ZN(n12274) );
  OR2_X1 U15211 ( .A1(n12280), .A2(n12274), .ZN(n12277) );
  AND2_X1 U15212 ( .A1(n12277), .A2(n15783), .ZN(n15775) );
  NAND2_X1 U15213 ( .A1(n12787), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12275) );
  OR2_X1 U15214 ( .A1(n19304), .A2(n12275), .ZN(n16511) );
  OR2_X1 U15215 ( .A1(n12276), .A2(n15725), .ZN(n13652) );
  NAND2_X1 U15216 ( .A1(n16511), .A2(n13652), .ZN(n15772) );
  NOR2_X1 U15217 ( .A1(n12277), .A2(n15783), .ZN(n15776) );
  NOR2_X1 U15218 ( .A1(n15772), .A2(n15776), .ZN(n12278) );
  NAND2_X1 U15219 ( .A1(n12227), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12279) );
  NAND3_X1 U15220 ( .A1(n12227), .A2(P2_EBX_REG_12__SCAN_IN), .A3(n12281), 
        .ZN(n12282) );
  NAND2_X1 U15221 ( .A1(n12299), .A2(n12282), .ZN(n19297) );
  INV_X1 U15222 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15756) );
  NOR2_X1 U15223 ( .A1(n12283), .A2(n15756), .ZN(n15764) );
  INV_X1 U15224 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12404) );
  NOR2_X1 U15225 ( .A1(n19552), .A2(n12404), .ZN(n12298) );
  INV_X1 U15226 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12408) );
  NAND2_X1 U15227 ( .A1(n12227), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12304) );
  NAND2_X1 U15228 ( .A1(n12227), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12287) );
  INV_X1 U15229 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n19222) );
  NOR2_X1 U15230 ( .A1(n19552), .A2(n19222), .ZN(n12308) );
  INV_X1 U15231 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12425) );
  NOR2_X1 U15232 ( .A1(n19552), .A2(n12425), .ZN(n12306) );
  INV_X1 U15233 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n12428) );
  INV_X1 U15234 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n19197) );
  NOR2_X1 U15235 ( .A1(n19552), .A2(n19197), .ZN(n12284) );
  AND2_X1 U15236 ( .A1(n12315), .A2(n12284), .ZN(n12285) );
  NOR2_X1 U15237 ( .A1(n12332), .A2(n12285), .ZN(n19202) );
  INV_X1 U15238 ( .A(n19202), .ZN(n12286) );
  OAI21_X1 U15239 ( .B1(n12286), .B2(n12320), .A(n15645), .ZN(n15467) );
  OR2_X1 U15240 ( .A1(n12288), .A2(n12287), .ZN(n12289) );
  AND2_X1 U15241 ( .A1(n12309), .A2(n12289), .ZN(n19234) );
  NAND2_X1 U15242 ( .A1(n19234), .A2(n12787), .ZN(n12291) );
  INV_X1 U15243 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12290) );
  NAND2_X1 U15244 ( .A1(n12291), .A2(n12290), .ZN(n15504) );
  NAND3_X1 U15245 ( .A1(n12292), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n12227), 
        .ZN(n12293) );
  NAND3_X1 U15246 ( .A1(n12294), .A2(n12357), .A3(n12293), .ZN(n19251) );
  INV_X1 U15247 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15712) );
  OAI21_X1 U15248 ( .B1(n19251), .B2(n12320), .A(n15712), .ZN(n12296) );
  NAND2_X1 U15249 ( .A1(n12787), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12295) );
  XNOR2_X1 U15250 ( .A(n12301), .B(n9969), .ZN(n19272) );
  NAND2_X1 U15251 ( .A1(n19272), .A2(n12787), .ZN(n12297) );
  INV_X1 U15252 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15737) );
  NAND2_X1 U15253 ( .A1(n12297), .A2(n15737), .ZN(n15718) );
  NAND2_X1 U15254 ( .A1(n12299), .A2(n12298), .ZN(n12300) );
  NAND2_X1 U15255 ( .A1(n12301), .A2(n12300), .ZN(n19285) );
  NOR2_X1 U15256 ( .A1(n19285), .A2(n12320), .ZN(n12323) );
  INV_X1 U15257 ( .A(n12323), .ZN(n12303) );
  INV_X1 U15258 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U15259 ( .A1(n12303), .A2(n12302), .ZN(n15714) );
  AND2_X1 U15260 ( .A1(n15718), .A2(n15714), .ZN(n15459) );
  XNOR2_X1 U15261 ( .A(n9920), .B(n12304), .ZN(n12321) );
  INV_X1 U15262 ( .A(n12321), .ZN(n19263) );
  NAND2_X1 U15263 ( .A1(n19263), .A2(n12787), .ZN(n12305) );
  INV_X1 U15264 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16570) );
  NAND2_X1 U15265 ( .A1(n12305), .A2(n16570), .ZN(n15527) );
  AND4_X1 U15266 ( .A1(n15504), .A2(n15462), .A3(n15459), .A4(n15527), .ZN(
        n12317) );
  XNOR2_X1 U15267 ( .A(n12311), .B(n10311), .ZN(n19209) );
  NAND2_X1 U15268 ( .A1(n19209), .A2(n12787), .ZN(n12307) );
  NAND2_X1 U15269 ( .A1(n12307), .A2(n15669), .ZN(n15491) );
  NAND2_X1 U15270 ( .A1(n12309), .A2(n12308), .ZN(n12310) );
  NAND2_X1 U15271 ( .A1(n12311), .A2(n12310), .ZN(n19223) );
  OR2_X1 U15272 ( .A1(n19223), .A2(n12320), .ZN(n12312) );
  NAND2_X1 U15273 ( .A1(n12312), .A2(n15678), .ZN(n15675) );
  AND2_X1 U15274 ( .A1(n15491), .A2(n15675), .ZN(n15464) );
  NAND2_X1 U15275 ( .A1(n12227), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12314) );
  MUX2_X1 U15276 ( .A(n12314), .B(n12227), .S(n12313), .Z(n12316) );
  NAND2_X1 U15277 ( .A1(n12316), .A2(n12315), .ZN(n15163) );
  INV_X1 U15278 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U15279 ( .A1(n12328), .A2(n15655), .ZN(n15479) );
  NAND4_X1 U15280 ( .A1(n15467), .A2(n12317), .A3(n15464), .A4(n15479), .ZN(
        n12331) );
  AND2_X1 U15281 ( .A1(n12787), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12318) );
  NAND2_X1 U15282 ( .A1(n19202), .A2(n12318), .ZN(n15466) );
  AND2_X1 U15283 ( .A1(n12787), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12319) );
  NAND2_X1 U15284 ( .A1(n19234), .A2(n12319), .ZN(n15503) );
  NAND2_X1 U15285 ( .A1(n15503), .A2(n15505), .ZN(n15463) );
  AND2_X1 U15286 ( .A1(n12787), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12322) );
  NAND2_X1 U15287 ( .A1(n19272), .A2(n12322), .ZN(n15717) );
  NAND2_X1 U15288 ( .A1(n12323), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15536) );
  NAND3_X1 U15289 ( .A1(n15526), .A2(n15717), .A3(n15536), .ZN(n12324) );
  NOR2_X1 U15290 ( .A1(n15463), .A2(n12324), .ZN(n12327) );
  AND2_X1 U15291 ( .A1(n12787), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12325) );
  NAND2_X1 U15292 ( .A1(n19209), .A2(n12325), .ZN(n15490) );
  NAND2_X1 U15293 ( .A1(n12787), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12326) );
  NAND4_X1 U15294 ( .A1(n15466), .A2(n12327), .A3(n15490), .A4(n15674), .ZN(
        n12329) );
  NOR2_X1 U15295 ( .A1(n12328), .A2(n15655), .ZN(n15481) );
  NOR2_X1 U15296 ( .A1(n12329), .A2(n15481), .ZN(n12330) );
  NAND2_X1 U15297 ( .A1(n12227), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12333) );
  INV_X1 U15298 ( .A(n12333), .ZN(n12334) );
  NAND2_X1 U15299 ( .A1(n9912), .A2(n12334), .ZN(n12335) );
  NAND2_X1 U15300 ( .A1(n12339), .A2(n12335), .ZN(n16000) );
  NOR2_X1 U15301 ( .A1(n12336), .A2(n15636), .ZN(n15624) );
  INV_X1 U15302 ( .A(n15624), .ZN(n12337) );
  INV_X1 U15303 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12438) );
  NOR2_X1 U15304 ( .A1(n19552), .A2(n12438), .ZN(n12338) );
  NAND2_X1 U15305 ( .A1(n12339), .A2(n12338), .ZN(n12340) );
  AND2_X1 U15306 ( .A1(n12345), .A2(n12340), .ZN(n16455) );
  NAND2_X1 U15307 ( .A1(n16455), .A2(n12787), .ZN(n12341) );
  XNOR2_X1 U15308 ( .A(n12341), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15455) );
  INV_X1 U15309 ( .A(n16455), .ZN(n12342) );
  INV_X1 U15310 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12750) );
  NAND2_X1 U15311 ( .A1(n12227), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12343) );
  MUX2_X1 U15312 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n12343), .S(n12345), .Z(
        n12344) );
  NAND2_X1 U15313 ( .A1(n12344), .A2(n12357), .ZN(n16437) );
  NOR2_X1 U15314 ( .A1(n16437), .A2(n12320), .ZN(n15445) );
  INV_X1 U15315 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15238) );
  NOR2_X1 U15316 ( .A1(n12349), .A2(n15238), .ZN(n12346) );
  NAND2_X1 U15317 ( .A1(n12227), .A2(n12346), .ZN(n12347) );
  NAND2_X1 U15318 ( .A1(n12357), .A2(n12347), .ZN(n12348) );
  AOI21_X1 U15319 ( .B1(n12349), .B2(n15238), .A(n12348), .ZN(n16425) );
  AOI21_X1 U15320 ( .B1(n16425), .B2(n12787), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15435) );
  NAND2_X1 U15321 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n12350), .ZN(n12351) );
  INV_X1 U15322 ( .A(n12359), .ZN(n12358) );
  OAI21_X1 U15323 ( .B1(n19552), .B2(n12351), .A(n12358), .ZN(n12352) );
  INV_X1 U15324 ( .A(n12352), .ZN(n12353) );
  NAND2_X1 U15325 ( .A1(n12357), .A2(n12353), .ZN(n16413) );
  XNOR2_X1 U15326 ( .A(n12355), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15428) );
  INV_X1 U15327 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21537) );
  INV_X1 U15328 ( .A(n16425), .ZN(n12354) );
  OAI21_X1 U15329 ( .B1(n12355), .B2(n21537), .A(n15426), .ZN(n12778) );
  INV_X1 U15330 ( .A(n12778), .ZN(n12356) );
  NAND2_X1 U15331 ( .A1(n12227), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12360) );
  OR2_X1 U15332 ( .A1(n12360), .A2(n12359), .ZN(n12361) );
  NAND2_X1 U15333 ( .A1(n12774), .A2(n12361), .ZN(n16401) );
  NOR2_X1 U15334 ( .A1(n12180), .A2(n12362), .ZN(n20237) );
  NAND2_X1 U15335 ( .A1(n12363), .A2(n12779), .ZN(n15416) );
  NAND3_X1 U15336 ( .A1(n15417), .A2(n19526), .A3(n15416), .ZN(n12772) );
  NAND2_X1 U15337 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12369) );
  INV_X1 U15338 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12366) );
  NAND2_X1 U15339 ( .A1(n12844), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12365) );
  NAND2_X1 U15340 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12364) );
  OAI211_X1 U15341 ( .C1(n12453), .C2(n12366), .A(n12365), .B(n12364), .ZN(
        n12367) );
  INV_X1 U15342 ( .A(n12367), .ZN(n12368) );
  NAND2_X1 U15343 ( .A1(n12369), .A2(n12368), .ZN(n14167) );
  NAND2_X1 U15344 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12374) );
  INV_X1 U15345 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n14295) );
  NAND2_X1 U15346 ( .A1(n12844), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12371) );
  NAND2_X1 U15347 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12370) );
  OAI211_X1 U15348 ( .C1(n12453), .C2(n14295), .A(n12371), .B(n12370), .ZN(
        n12372) );
  INV_X1 U15349 ( .A(n12372), .ZN(n12373) );
  INV_X1 U15350 ( .A(n12376), .ZN(n12377) );
  NAND2_X1 U15351 ( .A1(n12389), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12381) );
  AOI22_X1 U15352 ( .A1(n12844), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12380) );
  OAI211_X1 U15353 ( .C1(n12382), .C2(n12453), .A(n12381), .B(n12380), .ZN(
        n13916) );
  NAND2_X1 U15354 ( .A1(n13917), .A2(n13916), .ZN(n13918) );
  INV_X1 U15355 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19352) );
  NAND2_X1 U15356 ( .A1(n12844), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12384) );
  NAND2_X1 U15357 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12383) );
  OAI211_X1 U15358 ( .C1(n12453), .C2(n19352), .A(n12384), .B(n12383), .ZN(
        n12385) );
  AOI21_X1 U15359 ( .B1(n12389), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12385), .ZN(n13885) );
  NAND2_X1 U15360 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12387) );
  AOI22_X1 U15361 ( .A1(n12844), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12386) );
  OAI211_X1 U15362 ( .C1(n12388), .C2(n12453), .A(n12387), .B(n12386), .ZN(
        n13904) );
  NAND2_X1 U15363 ( .A1(n12844), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12391) );
  NAND2_X1 U15364 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12390) );
  OAI211_X1 U15365 ( .C1(n12453), .C2(n12392), .A(n12391), .B(n12390), .ZN(
        n12393) );
  AOI21_X1 U15366 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n12393), .ZN(n13936) );
  INV_X1 U15367 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12396) );
  NAND2_X1 U15368 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12395) );
  AOI22_X1 U15369 ( .A1(n12844), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12394) );
  OAI211_X1 U15370 ( .C1(n12396), .C2(n12453), .A(n12395), .B(n12394), .ZN(
        n13656) );
  NAND2_X1 U15371 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12398) );
  AOI22_X1 U15372 ( .A1(n12844), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12397) );
  OAI211_X1 U15373 ( .C1(n10305), .C2(n12453), .A(n12398), .B(n12397), .ZN(
        n14092) );
  NAND2_X1 U15374 ( .A1(n12844), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12400) );
  NAND2_X1 U15375 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12399) );
  OAI211_X1 U15376 ( .C1(n12453), .C2(n14159), .A(n12400), .B(n12399), .ZN(
        n12401) );
  AOI21_X1 U15377 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12401), .ZN(n14155) );
  NAND2_X1 U15378 ( .A1(n12844), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12403) );
  NAND2_X1 U15379 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12402) );
  OAI211_X1 U15380 ( .C1(n12453), .C2(n12404), .A(n12403), .B(n12402), .ZN(
        n12405) );
  AOI21_X1 U15381 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12405), .ZN(n14255) );
  NAND2_X1 U15382 ( .A1(n12844), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12407) );
  NAND2_X1 U15383 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12406) );
  OAI211_X1 U15384 ( .C1(n12453), .C2(n12408), .A(n12407), .B(n12406), .ZN(
        n12409) );
  AOI21_X1 U15385 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n12409), .ZN(n14377) );
  INV_X1 U15386 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U15387 ( .A1(n12844), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12411) );
  NAND2_X1 U15388 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12410) );
  OAI211_X1 U15389 ( .C1(n12453), .C2(n12412), .A(n12411), .B(n12410), .ZN(
        n12413) );
  AOI21_X1 U15390 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12413), .ZN(n14374) );
  INV_X1 U15391 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n19250) );
  NAND2_X1 U15392 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12415) );
  AOI22_X1 U15393 ( .A1(n12844), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n12414) );
  OAI211_X1 U15394 ( .C1(n12453), .C2(n19250), .A(n12415), .B(n12414), .ZN(
        n14388) );
  INV_X1 U15395 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12418) );
  NAND2_X1 U15396 ( .A1(n12844), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U15397 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12416) );
  OAI211_X1 U15398 ( .C1(n12453), .C2(n12418), .A(n12417), .B(n12416), .ZN(
        n12419) );
  AOI21_X1 U15399 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12419), .ZN(n14456) );
  NAND2_X1 U15400 ( .A1(n12844), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12421) );
  NAND2_X1 U15401 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12420) );
  OAI211_X1 U15402 ( .C1(n12453), .C2(n19222), .A(n12421), .B(n12420), .ZN(
        n12422) );
  AOI21_X1 U15403 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12422), .ZN(n15290) );
  NAND2_X1 U15404 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12424) );
  AOI22_X1 U15405 ( .A1(n12844), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n12423) );
  OAI211_X1 U15406 ( .C1(n12453), .C2(n12425), .A(n12424), .B(n12423), .ZN(
        n15284) );
  NAND2_X1 U15407 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12427) );
  AOI22_X1 U15408 ( .A1(n12844), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12426) );
  OAI211_X1 U15409 ( .C1(n12453), .C2(n12428), .A(n12427), .B(n12426), .ZN(
        n15153) );
  NAND2_X1 U15410 ( .A1(n12844), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12430) );
  NAND2_X1 U15411 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12429) );
  OAI211_X1 U15412 ( .C1(n12453), .C2(n19197), .A(n12430), .B(n12429), .ZN(
        n12431) );
  AOI21_X1 U15413 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12431), .ZN(n15270) );
  INV_X1 U15414 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12434) );
  NAND2_X1 U15415 ( .A1(n12844), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12433) );
  NAND2_X1 U15416 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12432) );
  OAI211_X1 U15417 ( .C1(n12453), .C2(n12434), .A(n12433), .B(n12432), .ZN(
        n12435) );
  AOI21_X1 U15418 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12435), .ZN(n15258) );
  NAND2_X1 U15419 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12437) );
  AOI22_X1 U15420 ( .A1(n12844), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12436) );
  OAI211_X1 U15421 ( .C1(n12453), .C2(n12438), .A(n12437), .B(n12436), .ZN(
        n15255) );
  INV_X1 U15422 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n12441) );
  NAND2_X1 U15423 ( .A1(n12844), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12440) );
  NAND2_X1 U15424 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12439) );
  OAI211_X1 U15425 ( .C1(n12453), .C2(n12441), .A(n12440), .B(n12439), .ZN(
        n12442) );
  AOI21_X1 U15426 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12442), .ZN(n15246) );
  NAND2_X1 U15427 ( .A1(n12844), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12444) );
  NAND2_X1 U15428 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12443) );
  OAI211_X1 U15429 ( .C1(n12453), .C2(n15238), .A(n12444), .B(n12443), .ZN(
        n12445) );
  AOI21_X1 U15430 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12445), .ZN(n15236) );
  INV_X1 U15431 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12448) );
  NAND2_X1 U15432 ( .A1(n12844), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12447) );
  NAND2_X1 U15433 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12446) );
  OAI211_X1 U15434 ( .C1(n12453), .C2(n12448), .A(n12447), .B(n12446), .ZN(
        n12449) );
  AOI21_X1 U15435 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12449), .ZN(n15225) );
  INV_X1 U15436 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12452) );
  NAND2_X1 U15437 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12451) );
  AOI22_X1 U15438 ( .A1(n12844), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12450) );
  OAI211_X1 U15439 ( .C1(n12453), .C2(n12452), .A(n12451), .B(n12450), .ZN(
        n12454) );
  NOR2_X1 U15440 ( .A1(n15226), .A2(n12454), .ZN(n12455) );
  OR2_X1 U15441 ( .A1(n15137), .A2(n12455), .ZN(n16403) );
  NAND2_X1 U15442 ( .A1(n12457), .A2(n9859), .ZN(n12460) );
  OR2_X1 U15443 ( .A1(n15813), .A2(n12459), .ZN(n15844) );
  NAND2_X1 U15444 ( .A1(n12460), .A2(n15844), .ZN(n12461) );
  AND2_X1 U15445 ( .A1(n12463), .A2(n14211), .ZN(n12466) );
  OR2_X1 U15446 ( .A1(n12464), .A2(n11852), .ZN(n12465) );
  NOR2_X1 U15447 ( .A1(n12465), .A2(n15813), .ZN(n16639) );
  OR2_X1 U15448 ( .A1(n12466), .A2(n16639), .ZN(n12467) );
  NOR2_X1 U15449 ( .A1(n14211), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12468) );
  INV_X1 U15450 ( .A(n12698), .ZN(n12512) );
  INV_X1 U15451 ( .A(n11727), .ZN(n13625) );
  INV_X1 U15452 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n16669) );
  NAND2_X1 U15453 ( .A1(n13625), .A2(n9860), .ZN(n12488) );
  INV_X1 U15454 ( .A(n12481), .ZN(n12469) );
  OAI21_X1 U15455 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n16669), .A(
        n12469), .ZN(n12470) );
  INV_X1 U15456 ( .A(n12472), .ZN(n12473) );
  INV_X1 U15457 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19188) );
  NAND2_X1 U15458 ( .A1(n12719), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12478) );
  INV_X1 U15459 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12475) );
  NAND2_X1 U15460 ( .A1(n14211), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12474) );
  OAI211_X1 U15461 ( .C1(n19570), .C2(n12475), .A(n12474), .B(n16669), .ZN(
        n12476) );
  INV_X1 U15462 ( .A(n12476), .ZN(n12477) );
  NAND2_X1 U15463 ( .A1(n12478), .A2(n12477), .ZN(n13806) );
  NAND2_X1 U15464 ( .A1(n12719), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12480) );
  INV_X2 U15465 ( .A(n9907), .ZN(n12821) );
  AOI22_X1 U15466 ( .A1(n12821), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n9861), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U15467 ( .A1(n12480), .A2(n12479), .ZN(n12485) );
  AOI22_X1 U15468 ( .A1(n11727), .A2(n12481), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12484) );
  OR2_X1 U15469 ( .A1(n12698), .A2(n12482), .ZN(n12483) );
  NAND2_X1 U15470 ( .A1(n12484), .A2(n12483), .ZN(n13984) );
  NAND2_X1 U15471 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12487) );
  OAI211_X1 U15472 ( .C1(n12698), .C2(n12489), .A(n12488), .B(n12487), .ZN(
        n12494) );
  XNOR2_X1 U15473 ( .A(n12495), .B(n12494), .ZN(n13981) );
  INV_X1 U15474 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20133) );
  NAND2_X1 U15475 ( .A1(n12719), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15476 ( .A1(n12821), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12491), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12492) );
  NAND2_X1 U15477 ( .A1(n12493), .A2(n12492), .ZN(n13980) );
  NOR2_X1 U15478 ( .A1(n13981), .A2(n13980), .ZN(n13982) );
  NOR2_X1 U15479 ( .A1(n12495), .A2(n12494), .ZN(n12496) );
  NAND2_X1 U15480 ( .A1(n12719), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15481 ( .A1(n12491), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12500) );
  OR2_X1 U15482 ( .A1(n12698), .A2(n12497), .ZN(n12499) );
  NAND2_X1 U15483 ( .A1(n12821), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12498) );
  NAND4_X1 U15484 ( .A1(n12501), .A2(n12500), .A3(n12499), .A4(n12498), .ZN(
        n15180) );
  NAND2_X1 U15485 ( .A1(n12719), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U15486 ( .A1(n12821), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12491), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12504) );
  OR2_X1 U15487 ( .A1(n12698), .A2(n12502), .ZN(n12503) );
  INV_X1 U15488 ( .A(n12506), .ZN(n12507) );
  AOI22_X1 U15489 ( .A1(n12719), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n12512), 
        .B2(n12507), .ZN(n12509) );
  AOI22_X1 U15490 ( .A1(n12821), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12491), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12508) );
  NAND2_X1 U15491 ( .A1(n12509), .A2(n12508), .ZN(n14408) );
  INV_X1 U15492 ( .A(n14407), .ZN(n12510) );
  AOI21_X1 U15493 ( .B1(n12512), .B2(n12511), .A(n12510), .ZN(n14430) );
  AOI222_X1 U15494 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n12719), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(P2_EAX_REG_6__SCAN_IN), 
        .C2(n12821), .ZN(n14429) );
  OAI22_X2 U15495 ( .A1(n14430), .A2(n14429), .B1(n12320), .B2(n12698), .ZN(
        n15795) );
  INV_X1 U15496 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19470) );
  INV_X1 U15497 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20143) );
  OAI222_X1 U15498 ( .A1(n16596), .A2(n12513), .B1(n9907), .B2(n19470), .C1(
        n12490), .C2(n20143), .ZN(n15794) );
  NAND2_X1 U15499 ( .A1(n12719), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U15500 ( .A1(n12821), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12491), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12535) );
  INV_X1 U15501 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12514) );
  INV_X1 U15502 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13314) );
  OAI22_X1 U15503 ( .A1(n12515), .A2(n12514), .B1(n13375), .B2(n13314), .ZN(
        n12518) );
  INV_X1 U15504 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12516) );
  OAI22_X1 U15505 ( .A1(n13371), .A2(n19886), .B1(n12690), .B2(n12516), .ZN(
        n12517) );
  NOR2_X1 U15506 ( .A1(n12518), .A2(n12517), .ZN(n12532) );
  INV_X1 U15507 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12521) );
  NAND2_X1 U15508 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12520) );
  NAND2_X1 U15509 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12519) );
  OAI211_X1 U15510 ( .C1(n12521), .C2(n12612), .A(n12520), .B(n12519), .ZN(
        n12522) );
  INV_X1 U15511 ( .A(n12522), .ZN(n12531) );
  AOI22_X1 U15512 ( .A1(n11914), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12526) );
  AOI22_X1 U15513 ( .A1(n11913), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12525) );
  NAND2_X1 U15514 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12524) );
  NAND2_X1 U15515 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12523) );
  NAND2_X1 U15516 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12528) );
  NAND2_X1 U15517 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12527) );
  OAI211_X1 U15518 ( .C1(n14235), .C2(n13447), .A(n12528), .B(n12527), .ZN(
        n12529) );
  INV_X1 U15519 ( .A(n12529), .ZN(n12530) );
  NAND4_X1 U15520 ( .A1(n12532), .A2(n12531), .A3(n10384), .A4(n12530), .ZN(
        n13970) );
  INV_X1 U15521 ( .A(n13970), .ZN(n12533) );
  OR2_X1 U15522 ( .A1(n12698), .A2(n12533), .ZN(n12534) );
  AOI22_X1 U15523 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11913), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U15524 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13305), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12539) );
  NAND2_X1 U15525 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12538) );
  NAND2_X1 U15526 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12537) );
  NAND4_X1 U15527 ( .A1(n12540), .A2(n12539), .A3(n12538), .A4(n12537), .ZN(
        n12545) );
  INV_X1 U15528 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12543) );
  NAND2_X1 U15529 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12542) );
  NAND2_X1 U15530 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12541) );
  OAI211_X1 U15531 ( .C1(n13447), .C2(n12543), .A(n12542), .B(n12541), .ZN(
        n12544) );
  NOR2_X1 U15532 ( .A1(n12545), .A2(n12544), .ZN(n12556) );
  NAND2_X1 U15533 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12549) );
  NAND2_X1 U15534 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12548) );
  NAND2_X1 U15535 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12547) );
  NAND2_X1 U15536 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12546) );
  NAND4_X1 U15537 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12554) );
  INV_X1 U15538 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12552) );
  NAND2_X1 U15539 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12551) );
  NAND2_X1 U15540 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12550) );
  OAI211_X1 U15541 ( .C1(n12690), .C2(n12552), .A(n12551), .B(n12550), .ZN(
        n12553) );
  NOR2_X1 U15542 ( .A1(n12554), .A2(n12553), .ZN(n12555) );
  NAND2_X1 U15543 ( .A1(n12719), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15544 ( .A1(n12821), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12491), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12557) );
  OAI211_X1 U15545 ( .C1(n14028), .C2(n12698), .A(n12558), .B(n12557), .ZN(
        n13658) );
  NAND2_X1 U15546 ( .A1(n12719), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15547 ( .A1(n12821), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15548 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11913), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U15549 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12109), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12561) );
  NAND2_X1 U15550 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12560) );
  NAND2_X1 U15551 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12559) );
  NAND4_X1 U15552 ( .A1(n12562), .A2(n12561), .A3(n12560), .A4(n12559), .ZN(
        n12567) );
  INV_X1 U15553 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12565) );
  NAND2_X1 U15554 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12564) );
  NAND2_X1 U15555 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12563) );
  OAI211_X1 U15556 ( .C1(n13447), .C2(n12565), .A(n12564), .B(n12563), .ZN(
        n12566) );
  NOR2_X1 U15557 ( .A1(n12567), .A2(n12566), .ZN(n12578) );
  NAND2_X1 U15558 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12571) );
  NAND2_X1 U15559 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12570) );
  NAND2_X1 U15560 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12569) );
  NAND2_X1 U15561 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12568) );
  NAND4_X1 U15562 ( .A1(n12571), .A2(n12570), .A3(n12569), .A4(n12568), .ZN(
        n12576) );
  INV_X1 U15563 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U15564 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12573) );
  NAND2_X1 U15565 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12572) );
  OAI211_X1 U15566 ( .C1(n13374), .C2(n12574), .A(n12573), .B(n12572), .ZN(
        n12575) );
  NOR2_X1 U15567 ( .A1(n12576), .A2(n12575), .ZN(n12577) );
  OR2_X1 U15568 ( .A1(n12698), .A2(n14088), .ZN(n12579) );
  AOI22_X1 U15569 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11913), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15570 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13305), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12584) );
  NAND2_X1 U15571 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12583) );
  NAND2_X1 U15572 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12582) );
  NAND4_X1 U15573 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n12590) );
  NAND2_X1 U15574 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12587) );
  NAND2_X1 U15575 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12586) );
  OAI211_X1 U15576 ( .C1(n13447), .C2(n12588), .A(n12587), .B(n12586), .ZN(
        n12589) );
  NOR2_X1 U15577 ( .A1(n12590), .A2(n12589), .ZN(n12602) );
  NAND2_X1 U15578 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12594) );
  NAND2_X1 U15579 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12593) );
  NAND2_X1 U15580 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12592) );
  NAND2_X1 U15581 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12591) );
  NAND4_X1 U15582 ( .A1(n12594), .A2(n12593), .A3(n12592), .A4(n12591), .ZN(
        n12600) );
  NAND2_X1 U15583 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12597) );
  NAND2_X1 U15584 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12596) );
  OAI211_X1 U15585 ( .C1(n12690), .C2(n12598), .A(n12597), .B(n12596), .ZN(
        n12599) );
  NOR2_X1 U15586 ( .A1(n12600), .A2(n12599), .ZN(n12601) );
  NAND2_X1 U15587 ( .A1(n12719), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15588 ( .A1(n12821), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12603) );
  OAI211_X1 U15589 ( .C1(n14152), .C2(n12698), .A(n12604), .B(n12603), .ZN(
        n15168) );
  NAND2_X1 U15590 ( .A1(n12719), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15591 ( .A1(n12821), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12628) );
  INV_X1 U15592 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12605) );
  INV_X1 U15593 ( .A(n13428), .ZN(n13372) );
  INV_X1 U15594 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13370) );
  OAI22_X1 U15595 ( .A1(n12605), .A2(n13372), .B1(n13375), .B2(n13370), .ZN(
        n12608) );
  INV_X1 U15596 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13536) );
  INV_X1 U15597 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12606) );
  OAI22_X1 U15598 ( .A1(n13536), .A2(n13371), .B1(n12690), .B2(n12606), .ZN(
        n12607) );
  NOR2_X1 U15599 ( .A1(n12608), .A2(n12607), .ZN(n12625) );
  NAND2_X1 U15600 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12610) );
  NAND2_X1 U15601 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12609) );
  OAI211_X1 U15602 ( .C1(n12612), .C2(n12611), .A(n12610), .B(n12609), .ZN(
        n12613) );
  INV_X1 U15603 ( .A(n12613), .ZN(n12624) );
  AOI22_X1 U15604 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11914), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15605 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11913), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12616) );
  NAND2_X1 U15606 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12615) );
  NAND2_X1 U15607 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12614) );
  AND4_X1 U15608 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n12623) );
  INV_X1 U15609 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12620) );
  NAND2_X1 U15610 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12619) );
  NAND2_X1 U15611 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12618) );
  OAI211_X1 U15612 ( .C1(n13374), .C2(n12620), .A(n12619), .B(n12618), .ZN(
        n12621) );
  INV_X1 U15613 ( .A(n12621), .ZN(n12622) );
  NAND4_X1 U15614 ( .A1(n12625), .A2(n12624), .A3(n12623), .A4(n12622), .ZN(
        n14170) );
  INV_X1 U15615 ( .A(n14170), .ZN(n12626) );
  OR2_X1 U15616 ( .A1(n12698), .A2(n12626), .ZN(n12627) );
  NOR2_X2 U15617 ( .A1(n15761), .A2(n15760), .ZN(n15744) );
  AOI22_X1 U15618 ( .A1(n11913), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15619 ( .A1(n12109), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12632) );
  NAND2_X1 U15620 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12631) );
  NAND2_X1 U15621 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12630) );
  NAND4_X1 U15622 ( .A1(n12633), .A2(n12632), .A3(n12631), .A4(n12630), .ZN(
        n12638) );
  NAND2_X1 U15623 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12635) );
  NAND2_X1 U15624 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12634) );
  OAI211_X1 U15625 ( .C1(n12636), .C2(n13447), .A(n12635), .B(n12634), .ZN(
        n12637) );
  NOR2_X1 U15626 ( .A1(n12638), .A2(n12637), .ZN(n12649) );
  NAND2_X1 U15627 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12642) );
  NAND2_X1 U15628 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12641) );
  NAND2_X1 U15629 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12640) );
  NAND2_X1 U15630 ( .A1(n13429), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12639) );
  NAND4_X1 U15631 ( .A1(n12642), .A2(n12641), .A3(n12640), .A4(n12639), .ZN(
        n12647) );
  NAND2_X1 U15632 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12644) );
  NAND2_X1 U15633 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12643) );
  OAI211_X1 U15634 ( .C1(n12645), .C2(n12690), .A(n12644), .B(n12643), .ZN(
        n12646) );
  NOR2_X1 U15635 ( .A1(n12647), .A2(n12646), .ZN(n12648) );
  NAND2_X1 U15636 ( .A1(n12719), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U15637 ( .A1(n12821), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12650) );
  OAI211_X1 U15638 ( .C1(n14253), .C2(n12698), .A(n12651), .B(n12650), .ZN(
        n15745) );
  NAND2_X1 U15639 ( .A1(n15744), .A2(n15745), .ZN(n15729) );
  AOI22_X1 U15640 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11913), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15641 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12109), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U15642 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12653) );
  NAND2_X1 U15643 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12652) );
  NAND4_X1 U15644 ( .A1(n12655), .A2(n12654), .A3(n12653), .A4(n12652), .ZN(
        n12660) );
  NAND2_X1 U15645 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12657) );
  NAND2_X1 U15646 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12656) );
  OAI211_X1 U15647 ( .C1(n12690), .C2(n12658), .A(n12657), .B(n12656), .ZN(
        n12659) );
  NOR2_X1 U15648 ( .A1(n12660), .A2(n12659), .ZN(n12672) );
  NAND2_X1 U15649 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12665) );
  NAND2_X1 U15650 ( .A1(n13427), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12664) );
  NAND2_X1 U15651 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12663) );
  NAND2_X1 U15652 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12662) );
  NAND4_X1 U15653 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12670) );
  INV_X1 U15654 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U15655 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12667) );
  NAND2_X1 U15656 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12666) );
  OAI211_X1 U15657 ( .C1(n13374), .C2(n12668), .A(n12667), .B(n12666), .ZN(
        n12669) );
  NOR2_X1 U15658 ( .A1(n12670), .A2(n12669), .ZN(n12671) );
  AOI22_X1 U15659 ( .A1(n12821), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12673) );
  OAI21_X1 U15660 ( .B1(n14382), .B2(n12698), .A(n12673), .ZN(n12674) );
  AOI21_X1 U15661 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n12719), .A(n12674), 
        .ZN(n15731) );
  INV_X1 U15662 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12675) );
  OAI22_X1 U15663 ( .A1(n12675), .A2(n13372), .B1(n13371), .B2(n13596), .ZN(
        n12678) );
  INV_X1 U15664 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12676) );
  INV_X1 U15665 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13599) );
  OAI22_X1 U15666 ( .A1(n12676), .A2(n13375), .B1(n13374), .B2(n13599), .ZN(
        n12677) );
  NOR2_X1 U15667 ( .A1(n12678), .A2(n12677), .ZN(n12695) );
  NAND2_X1 U15668 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12680) );
  NAND2_X1 U15669 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12679) );
  OAI211_X1 U15670 ( .C1(n13447), .C2(n12681), .A(n12680), .B(n12679), .ZN(
        n12682) );
  INV_X1 U15671 ( .A(n12682), .ZN(n12694) );
  AOI22_X1 U15672 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11914), .B1(
        n11913), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15673 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13305), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U15674 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12684) );
  NAND2_X1 U15675 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12683) );
  AND4_X1 U15676 ( .A1(n12686), .A2(n12685), .A3(n12684), .A4(n12683), .ZN(
        n12693) );
  NAND2_X1 U15677 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12688) );
  NAND2_X1 U15678 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12687) );
  OAI211_X1 U15679 ( .C1(n12690), .C2(n12689), .A(n12688), .B(n12687), .ZN(
        n12691) );
  INV_X1 U15680 ( .A(n12691), .ZN(n12692) );
  NAND4_X1 U15681 ( .A1(n12695), .A2(n12694), .A3(n12693), .A4(n12692), .ZN(
        n14373) );
  INV_X1 U15682 ( .A(n14373), .ZN(n12699) );
  NAND2_X1 U15683 ( .A1(n12719), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U15684 ( .A1(n12821), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12696) );
  OAI211_X1 U15685 ( .C1(n12699), .C2(n12698), .A(n12697), .B(n12696), .ZN(
        n16565) );
  NAND2_X1 U15686 ( .A1(n15730), .A2(n16565), .ZN(n16566) );
  NAND2_X1 U15687 ( .A1(n12719), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15688 ( .A1(n12821), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12700) );
  NAND2_X1 U15689 ( .A1(n12701), .A2(n12700), .ZN(n15382) );
  NAND2_X1 U15690 ( .A1(n12719), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15691 ( .A1(n12821), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12702) );
  AOI222_X1 U15692 ( .A1(n12719), .A2(P2_REIP_REG_18__SCAN_IN), .B1(n12821), 
        .B2(P2_EAX_REG_18__SCAN_IN), .C1(n12491), .C2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15683) );
  NOR2_X2 U15693 ( .A1(n15682), .A2(n15683), .ZN(n15681) );
  NAND2_X1 U15694 ( .A1(n12719), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15695 ( .A1(n12821), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U15696 ( .A1(n12705), .A2(n12704), .ZN(n15364) );
  AND2_X2 U15697 ( .A1(n15681), .A2(n15364), .ZN(n15366) );
  NAND2_X1 U15698 ( .A1(n12719), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15699 ( .A1(n12821), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12706) );
  NAND2_X1 U15700 ( .A1(n12707), .A2(n12706), .ZN(n15156) );
  NAND2_X1 U15701 ( .A1(n12719), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15702 ( .A1(n12821), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12708) );
  NAND2_X1 U15703 ( .A1(n12709), .A2(n12708), .ZN(n15353) );
  AND2_X2 U15704 ( .A1(n15155), .A2(n15353), .ZN(n15627) );
  NAND2_X1 U15705 ( .A1(n12719), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15706 ( .A1(n12821), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U15707 ( .A1(n12711), .A2(n12710), .ZN(n15628) );
  NAND2_X1 U15708 ( .A1(n12719), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U15709 ( .A1(n12821), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12712) );
  AND2_X1 U15710 ( .A1(n12713), .A2(n12712), .ZN(n15343) );
  NAND2_X1 U15711 ( .A1(n12719), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U15712 ( .A1(n12821), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12714) );
  AND2_X1 U15713 ( .A1(n12715), .A2(n12714), .ZN(n15335) );
  INV_X1 U15714 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20177) );
  AOI22_X1 U15715 ( .A1(n12821), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12716) );
  OAI21_X1 U15716 ( .B1(n12490), .B2(n20177), .A(n12716), .ZN(n15328) );
  NAND2_X1 U15717 ( .A1(n12719), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15718 ( .A1(n12821), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12717) );
  AND2_X1 U15719 ( .A1(n12718), .A2(n12717), .ZN(n15320) );
  NAND2_X1 U15720 ( .A1(n12719), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15721 ( .A1(n12821), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12720) );
  AND2_X1 U15722 ( .A1(n12721), .A2(n12720), .ZN(n12722) );
  AND2_X1 U15723 ( .A1(n9909), .A2(n12722), .ZN(n12723) );
  NOR2_X1 U15724 ( .A1(n12819), .A2(n12723), .ZN(n16404) );
  AND2_X2 U15725 ( .A1(n11745), .A2(n20206), .ZN(n19247) );
  NAND2_X1 U15726 ( .A1(n19247), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15418) );
  INV_X1 U15727 ( .A(n15418), .ZN(n12724) );
  AOI21_X1 U15728 ( .B1(n19517), .B2(n16404), .A(n12724), .ZN(n12753) );
  NAND2_X1 U15729 ( .A1(n12725), .A2(n14211), .ZN(n15814) );
  NAND2_X1 U15730 ( .A1(n15814), .A2(n12726), .ZN(n12728) );
  NAND2_X1 U15731 ( .A1(n12728), .A2(n12727), .ZN(n12741) );
  OAI22_X1 U15732 ( .A1(n12729), .A2(n19547), .B1(n12730), .B2(n16637), .ZN(
        n12731) );
  INV_X1 U15733 ( .A(n12731), .ZN(n12732) );
  AND2_X1 U15734 ( .A1(n12733), .A2(n12732), .ZN(n12740) );
  INV_X1 U15735 ( .A(n12734), .ZN(n12742) );
  NAND2_X1 U15736 ( .A1(n13622), .A2(n12735), .ZN(n12736) );
  OAI211_X1 U15737 ( .C1(n12742), .C2(n12737), .A(n12736), .B(n12729), .ZN(
        n12738) );
  NAND2_X1 U15738 ( .A1(n12738), .A2(n13621), .ZN(n12739) );
  AND3_X1 U15739 ( .A1(n12741), .A2(n12740), .A3(n12739), .ZN(n15851) );
  NAND2_X1 U15740 ( .A1(n15851), .A2(n12744), .ZN(n12745) );
  NAND2_X1 U15741 ( .A1(n12755), .A2(n12745), .ZN(n19512) );
  INV_X1 U15742 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15817) );
  NOR2_X1 U15743 ( .A1(n15833), .A2(n15817), .ZN(n19519) );
  NAND2_X1 U15744 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19519), .ZN(
        n12746) );
  OR2_X1 U15745 ( .A1(n19512), .A2(n12746), .ZN(n12749) );
  NAND2_X1 U15746 ( .A1(n12755), .A2(n13620), .ZN(n19523) );
  NAND2_X1 U15747 ( .A1(n12749), .A2(n19523), .ZN(n14401) );
  INV_X1 U15748 ( .A(n19519), .ZN(n19515) );
  NAND2_X1 U15749 ( .A1(n19537), .A2(n19515), .ZN(n19522) );
  NOR2_X1 U15750 ( .A1(n14403), .A2(n19502), .ZN(n14432) );
  NAND3_X1 U15751 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n14432), .ZN(n15792) );
  INV_X1 U15752 ( .A(n15792), .ZN(n14433) );
  AND4_X1 U15753 ( .A1(n19522), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n14433), .ZN(n12756) );
  AND2_X1 U15754 ( .A1(n15680), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12758) );
  NAND2_X1 U15755 ( .A1(n15781), .A2(n12758), .ZN(n15663) );
  NAND2_X1 U15756 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12760) );
  NOR2_X1 U15757 ( .A1(n15663), .A2(n12760), .ZN(n12762) );
  NAND2_X1 U15758 ( .A1(n12762), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15632) );
  NOR2_X1 U15759 ( .A1(n15601), .A2(n12750), .ZN(n15597) );
  NAND2_X1 U15760 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12765) );
  INV_X1 U15761 ( .A(n12765), .ZN(n12751) );
  NAND2_X1 U15762 ( .A1(n15597), .A2(n12751), .ZN(n15566) );
  OR2_X1 U15763 ( .A1(n15566), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12752) );
  OAI211_X1 U15764 ( .C1(n16403), .C2(n19534), .A(n12753), .B(n12752), .ZN(
        n12770) );
  AND2_X1 U15765 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19519), .ZN(
        n12754) );
  OR2_X1 U15766 ( .A1(n19512), .A2(n12754), .ZN(n19518) );
  INV_X1 U15767 ( .A(n19247), .ZN(n19233) );
  OR2_X1 U15768 ( .A1(n12755), .A2(n19247), .ZN(n19513) );
  AND2_X1 U15769 ( .A1(n19518), .A2(n19513), .ZN(n14399) );
  OR2_X1 U15770 ( .A1(n15726), .A2(n12756), .ZN(n12757) );
  NAND2_X1 U15771 ( .A1(n15780), .A2(n12758), .ZN(n12759) );
  NAND2_X1 U15772 ( .A1(n12759), .A2(n12766), .ZN(n15688) );
  INV_X1 U15773 ( .A(n12760), .ZN(n15654) );
  OR2_X1 U15774 ( .A1(n15779), .A2(n15654), .ZN(n12761) );
  AND2_X1 U15775 ( .A1(n15688), .A2(n12761), .ZN(n15646) );
  NAND2_X1 U15776 ( .A1(n12762), .A2(n15645), .ZN(n15643) );
  AND2_X1 U15777 ( .A1(n15646), .A2(n15643), .ZN(n15637) );
  NOR2_X1 U15778 ( .A1(n15617), .A2(n15636), .ZN(n15612) );
  OAI21_X1 U15779 ( .B1(n15726), .B2(n15612), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12763) );
  INV_X1 U15780 ( .A(n12763), .ZN(n12764) );
  NAND2_X1 U15781 ( .A1(n15637), .A2(n12764), .ZN(n15602) );
  NAND2_X1 U15782 ( .A1(n15602), .A2(n12766), .ZN(n15591) );
  NAND2_X1 U15783 ( .A1(n12766), .A2(n12765), .ZN(n12767) );
  NAND2_X1 U15784 ( .A1(n15591), .A2(n12767), .ZN(n15576) );
  INV_X1 U15785 ( .A(n15576), .ZN(n12768) );
  NOR2_X1 U15786 ( .A1(n12768), .A2(n12779), .ZN(n12769) );
  NOR2_X1 U15787 ( .A1(n12770), .A2(n12769), .ZN(n12771) );
  NAND2_X1 U15788 ( .A1(n10388), .A2(n10389), .ZN(P2_U3019) );
  INV_X1 U15789 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12794) );
  NOR2_X1 U15790 ( .A1(n19552), .A2(n12794), .ZN(n12773) );
  NAND2_X1 U15791 ( .A1(n12774), .A2(n12773), .ZN(n12775) );
  NAND2_X1 U15792 ( .A1(n12784), .A2(n12775), .ZN(n15141) );
  OAI22_X1 U15793 ( .A1(n15408), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15405), .ZN(n12776) );
  INV_X1 U15794 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15409) );
  NAND2_X1 U15795 ( .A1(n15409), .A2(n12779), .ZN(n15567) );
  INV_X1 U15796 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12798) );
  NOR2_X1 U15797 ( .A1(n19552), .A2(n12798), .ZN(n12783) );
  AOI21_X1 U15798 ( .B1(n16388), .B2(n12787), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15397) );
  INV_X1 U15799 ( .A(n16388), .ZN(n12782) );
  INV_X1 U15800 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15558) );
  NOR3_X1 U15801 ( .A1(n12782), .A2(n12320), .A3(n15558), .ZN(n15398) );
  NOR2_X1 U15802 ( .A1(n12835), .A2(n15398), .ZN(n12790) );
  NAND2_X1 U15803 ( .A1(n12227), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12785) );
  INV_X1 U15804 ( .A(n13231), .ZN(n12786) );
  INV_X1 U15805 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12870) );
  INV_X1 U15806 ( .A(n12834), .ZN(n12788) );
  NOR2_X1 U15807 ( .A1(n12788), .A2(n12832), .ZN(n12789) );
  XNOR2_X1 U15808 ( .A(n12790), .B(n12789), .ZN(n12830) );
  AND2_X1 U15809 ( .A1(n14199), .A2(n16665), .ZN(n13221) );
  NAND2_X1 U15810 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12793) );
  AOI22_X1 U15811 ( .A1(n12844), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12792) );
  OAI211_X1 U15812 ( .C1(n12453), .C2(n12794), .A(n12793), .B(n12792), .ZN(
        n15136) );
  NAND2_X1 U15813 ( .A1(n12795), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12797) );
  AOI22_X1 U15814 ( .A1(n12844), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12796) );
  OAI211_X1 U15815 ( .C1(n12453), .C2(n12798), .A(n12797), .B(n12796), .ZN(
        n15204) );
  INV_X1 U15816 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U15817 ( .A1(n12844), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12800) );
  NAND2_X1 U15818 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12799) );
  OAI211_X1 U15819 ( .C1(n12453), .C2(n12801), .A(n12800), .B(n12799), .ZN(
        n12802) );
  AOI21_X1 U15820 ( .B1(n12795), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12802), .ZN(n12803) );
  NAND2_X1 U15821 ( .A1(n15207), .A2(n12803), .ZN(n12804) );
  NAND2_X1 U15822 ( .A1(n9939), .A2(n12804), .ZN(n14545) );
  NOR2_X1 U15823 ( .A1(n15818), .A2(n19913), .ZN(n16649) );
  INV_X1 U15824 ( .A(n16649), .ZN(n13671) );
  OAI211_X1 U15825 ( .C1(P2_STATE2_REG_1__SCAN_IN), .C2(
        P2_STATE2_REG_2__SCAN_IN), .A(n13671), .B(n16656), .ZN(n12805) );
  INV_X1 U15826 ( .A(n14195), .ZN(n19494) );
  NAND2_X1 U15827 ( .A1(n15818), .A2(n19873), .ZN(n20200) );
  INV_X1 U15828 ( .A(n20200), .ZN(n15855) );
  OR2_X1 U15829 ( .A1(n20206), .A2(n15855), .ZN(n20225) );
  NAND2_X1 U15830 ( .A1(n20225), .A2(n16656), .ZN(n12806) );
  INV_X1 U15831 ( .A(n13287), .ZN(n12808) );
  INV_X1 U15832 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20197) );
  NAND2_X1 U15833 ( .A1(n20197), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U15834 ( .A1(n12808), .A2(n12807), .ZN(n13765) );
  INV_X1 U15835 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15497) );
  INV_X1 U15836 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n19196) );
  INV_X1 U15837 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15439) );
  INV_X1 U15838 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16400) );
  INV_X1 U15839 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13180) );
  INV_X1 U15840 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12810) );
  XNOR2_X1 U15841 ( .A(n12849), .B(n12810), .ZN(n16382) );
  INV_X1 U15842 ( .A(n16382), .ZN(n12812) );
  NAND2_X1 U15843 ( .A1(n19247), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12826) );
  OAI21_X1 U15844 ( .B1(n16561), .B2(n12810), .A(n12826), .ZN(n12811) );
  AOI21_X1 U15845 ( .B1(n16550), .B2(n12812), .A(n12811), .ZN(n12813) );
  OAI21_X1 U15846 ( .B1(n14545), .B2(n14195), .A(n12813), .ZN(n12814) );
  AOI21_X1 U15847 ( .B1(n12830), .B2(n19493), .A(n12814), .ZN(n12817) );
  NAND3_X1 U15848 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15557) );
  XNOR2_X1 U15849 ( .A(n15394), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12829) );
  NAND2_X1 U15850 ( .A1(n12817), .A2(n12816), .ZN(P2_U2984) );
  INV_X1 U15851 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20182) );
  AOI22_X1 U15852 ( .A1(n12821), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12818) );
  OAI21_X1 U15853 ( .B1(n12490), .B2(n20182), .A(n12818), .ZN(n15142) );
  AND2_X2 U15854 ( .A1(n12819), .A2(n15142), .ZN(n15301) );
  INV_X1 U15855 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n21456) );
  AOI22_X1 U15856 ( .A1(n12821), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12820) );
  OAI21_X1 U15857 ( .B1(n12490), .B2(n21456), .A(n12820), .ZN(n15300) );
  NAND2_X1 U15858 ( .A1(n12719), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U15859 ( .A1(n12821), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12491), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12822) );
  AND2_X1 U15860 ( .A1(n12823), .A2(n12822), .ZN(n12824) );
  OR2_X2 U15861 ( .A1(n15303), .A2(n12824), .ZN(n12867) );
  NAND2_X1 U15862 ( .A1(n15303), .A2(n12824), .ZN(n12825) );
  INV_X1 U15863 ( .A(n12826), .ZN(n12828) );
  NOR3_X1 U15864 ( .A1(n15566), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15557), .ZN(n12827) );
  INV_X1 U15865 ( .A(n15726), .ZN(n15809) );
  AOI21_X1 U15866 ( .B1(n15809), .B2(n15557), .A(n15576), .ZN(n12864) );
  NAND2_X1 U15867 ( .A1(n9938), .A2(n12831), .ZN(P2_U3016) );
  INV_X1 U15868 ( .A(n12836), .ZN(n12839) );
  NOR2_X1 U15869 ( .A1(n12837), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12838) );
  MUX2_X1 U15870 ( .A(n12839), .B(n12838), .S(n12227), .Z(n16378) );
  NAND2_X1 U15871 ( .A1(n16378), .A2(n12787), .ZN(n12840) );
  XNOR2_X1 U15872 ( .A(n12841), .B(n10386), .ZN(n12860) );
  NAND2_X1 U15873 ( .A1(n12860), .A2(n19493), .ZN(n12859) );
  NAND2_X1 U15874 ( .A1(n15394), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12843) );
  AOI22_X1 U15876 ( .A1(n12844), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12846) );
  NAND2_X1 U15877 ( .A1(n12379), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12845) );
  OAI211_X1 U15878 ( .C1(n11788), .C2(n12842), .A(n12846), .B(n12845), .ZN(
        n12848) );
  NAND2_X1 U15879 ( .A1(n16380), .A2(n19494), .ZN(n12856) );
  INV_X1 U15880 ( .A(n12849), .ZN(n12850) );
  NAND2_X1 U15881 ( .A1(n12850), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12852) );
  INV_X1 U15882 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12851) );
  NAND2_X1 U15883 ( .A1(n19247), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12868) );
  NAND2_X1 U15884 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12853) );
  OAI211_X1 U15885 ( .C1(n19499), .C2(n13179), .A(n12868), .B(n12853), .ZN(
        n12854) );
  INV_X1 U15886 ( .A(n12854), .ZN(n12855) );
  INV_X1 U15887 ( .A(n12857), .ZN(n12858) );
  NAND2_X1 U15888 ( .A1(n12859), .A2(n12858), .ZN(P2_U2983) );
  NAND2_X1 U15889 ( .A1(n12860), .A2(n19526), .ZN(n12879) );
  INV_X1 U15890 ( .A(n12861), .ZN(n12863) );
  NAND2_X1 U15891 ( .A1(n12863), .A2(n12862), .ZN(n12878) );
  INV_X1 U15892 ( .A(n16380), .ZN(n12875) );
  OAI21_X1 U15893 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15726), .A(
        n12864), .ZN(n12865) );
  INV_X1 U15894 ( .A(n12865), .ZN(n12872) );
  AOI222_X1 U15895 ( .A1(n12719), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12821), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12491), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12866) );
  OAI21_X1 U15896 ( .B1(n16379), .B2(n16603), .A(n12868), .ZN(n12869) );
  INV_X1 U15897 ( .A(n12869), .ZN(n12871) );
  INV_X1 U15898 ( .A(n12873), .ZN(n12874) );
  OAI21_X1 U15899 ( .B1(n12875), .B2(n19534), .A(n12874), .ZN(n12876) );
  NAND3_X1 U15900 ( .A1(n12879), .A2(n12878), .A3(n12877), .ZN(P2_U3015) );
  AOI22_X1 U15901 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12884) );
  NOR2_X1 U15902 ( .A1(n17182), .A2(n12880), .ZN(n12917) );
  NOR2_X1 U15903 ( .A1(n12885), .A2(n12880), .ZN(n12926) );
  INV_X2 U15904 ( .A(n17370), .ZN(n15953) );
  AOI22_X1 U15905 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12883) );
  INV_X2 U15906 ( .A(n17220), .ZN(n17450) );
  AOI22_X1 U15907 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17450), .ZN(n12882) );
  BUF_X4 U15908 ( .A(n9821), .Z(n17472) );
  AOI22_X1 U15909 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12881) );
  NAND4_X1 U15910 ( .A1(n12884), .A2(n12883), .A3(n12882), .A4(n12881), .ZN(
        n12894) );
  AOI22_X1 U15911 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17458), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12892) );
  AOI22_X1 U15912 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15918), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12891) );
  INV_X2 U15913 ( .A(n17435), .ZN(n17460) );
  AOI22_X1 U15914 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U15915 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12889) );
  NAND4_X1 U15916 ( .A1(n12892), .A2(n12891), .A3(n12890), .A4(n12889), .ZN(
        n12893) );
  AOI22_X1 U15917 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U15918 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12897) );
  AOI22_X1 U15919 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U15920 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12895) );
  NAND4_X1 U15921 ( .A1(n12898), .A2(n12897), .A3(n12896), .A4(n12895), .ZN(
        n12904) );
  AOI22_X1 U15922 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U15923 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U15924 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12900) );
  INV_X2 U15925 ( .A(n9917), .ZN(n17417) );
  AOI22_X1 U15926 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12899) );
  NAND4_X1 U15927 ( .A1(n12902), .A2(n12901), .A3(n12900), .A4(n12899), .ZN(
        n12903) );
  AOI22_X1 U15928 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U15929 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U15930 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U15931 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12905) );
  NAND4_X1 U15932 ( .A1(n12908), .A2(n12907), .A3(n12906), .A4(n12905), .ZN(
        n12914) );
  AOI22_X1 U15933 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12912) );
  INV_X2 U15934 ( .A(n17370), .ZN(n17471) );
  AOI22_X1 U15935 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U15936 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U15937 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12909) );
  NAND4_X1 U15938 ( .A1(n12912), .A2(n12911), .A3(n12910), .A4(n12909), .ZN(
        n12913) );
  INV_X2 U15939 ( .A(n15920), .ZN(n17480) );
  AOI22_X1 U15940 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12924) );
  AOI22_X1 U15941 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12923) );
  INV_X1 U15942 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17518) );
  AOI22_X1 U15943 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U15944 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12917), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U15945 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U15946 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U15947 ( .A1(n12922), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12932) );
  INV_X2 U15948 ( .A(n13062), .ZN(n17386) );
  AOI22_X1 U15949 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12931) );
  INV_X1 U15950 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n21467) );
  AOI22_X1 U15951 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U15952 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U15953 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12926), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U15954 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U15955 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U15956 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12942) );
  INV_X4 U15957 ( .A(n12956), .ZN(n17457) );
  AOI22_X1 U15958 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12941) );
  INV_X1 U15959 ( .A(n17370), .ZN(n13090) );
  INV_X1 U15960 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U15961 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12933) );
  OAI21_X1 U15962 ( .B1(n9911), .B2(n17300), .A(n12933), .ZN(n12939) );
  AOI22_X1 U15963 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17458), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U15964 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U15965 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U15966 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12934) );
  NAND4_X1 U15967 ( .A1(n12937), .A2(n12936), .A3(n12935), .A4(n12934), .ZN(
        n12938) );
  AOI211_X1 U15968 ( .C1(n13090), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n12939), .B(n12938), .ZN(n12940) );
  NAND3_X1 U15969 ( .A1(n12942), .A2(n12941), .A3(n12940), .ZN(n17659) );
  NAND2_X1 U15970 ( .A1(n12954), .A2(n17659), .ZN(n12975) );
  AOI22_X1 U15971 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U15972 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12952) );
  AOI22_X1 U15973 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12943) );
  OAI21_X1 U15974 ( .B1(n12956), .B2(n21366), .A(n12943), .ZN(n12950) );
  AOI22_X1 U15975 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U15976 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12947) );
  INV_X1 U15977 ( .A(n12944), .ZN(n17459) );
  AOI22_X1 U15978 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U15979 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12945) );
  NAND4_X1 U15980 ( .A1(n12948), .A2(n12947), .A3(n12946), .A4(n12945), .ZN(
        n12949) );
  AOI211_X1 U15981 ( .C1(n15908), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12950), .B(n12949), .ZN(n12951) );
  NAND3_X1 U15982 ( .A1(n12953), .A2(n12952), .A3(n12951), .ZN(n18089) );
  INV_X1 U15983 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16684) );
  INV_X1 U15984 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21488) );
  INV_X1 U15985 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17926) );
  INV_X1 U15986 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21522) );
  NAND2_X1 U15987 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18250) );
  NOR2_X1 U15988 ( .A1(n21522), .A2(n18250), .ZN(n18171) );
  NAND2_X1 U15989 ( .A1(n18171), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17861) );
  NOR2_X1 U15990 ( .A1(n17926), .A2(n17861), .ZN(n17858) );
  AND2_X1 U15991 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17858), .ZN(
        n12995) );
  INV_X1 U15992 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18303) );
  INV_X1 U15993 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18343) );
  INV_X1 U15994 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18327) );
  INV_X1 U15995 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18296) );
  NOR3_X1 U15996 ( .A1(n18343), .A2(n18327), .A3(n18296), .ZN(n13250) );
  NAND2_X1 U15997 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12973), .ZN(
        n12974) );
  INV_X1 U15998 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18446) );
  XOR2_X1 U15999 ( .A(n12955), .B(n13136), .Z(n18129) );
  INV_X1 U16000 ( .A(n12969), .ZN(n17681) );
  NAND2_X1 U16001 ( .A1(n17681), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12968) );
  AOI22_X1 U16002 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9823), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12961) );
  AOI22_X1 U16003 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12960) );
  AOI22_X1 U16004 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U16005 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12958) );
  NAND4_X1 U16006 ( .A1(n12961), .A2(n12960), .A3(n12959), .A4(n12958), .ZN(
        n12967) );
  AOI22_X1 U16007 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U16008 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U16009 ( .A1(n12922), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16010 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12962) );
  NAND4_X1 U16011 ( .A1(n12965), .A2(n12964), .A3(n12963), .A4(n12962), .ZN(
        n12966) );
  NOR2_X2 U16012 ( .A1(n12967), .A2(n12966), .ZN(n18163) );
  INV_X1 U16013 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19125) );
  NOR2_X1 U16014 ( .A1(n18163), .A2(n19125), .ZN(n18162) );
  NAND2_X1 U16015 ( .A1(n18155), .A2(n18162), .ZN(n18154) );
  NAND2_X1 U16016 ( .A1(n12968), .A2(n18154), .ZN(n18147) );
  INV_X1 U16017 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18457) );
  XNOR2_X1 U16018 ( .A(n12970), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18148) );
  NAND2_X1 U16019 ( .A1(n18147), .A2(n18148), .ZN(n18146) );
  OR2_X1 U16020 ( .A1(n18457), .A2(n12970), .ZN(n12971) );
  NAND2_X1 U16021 ( .A1(n18146), .A2(n12971), .ZN(n18130) );
  NAND2_X1 U16022 ( .A1(n18129), .A2(n18130), .ZN(n18128) );
  NOR2_X1 U16023 ( .A1(n18129), .A2(n18130), .ZN(n12972) );
  XOR2_X1 U16024 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12973), .Z(
        n18121) );
  NAND2_X1 U16025 ( .A1(n18118), .A2(n18121), .ZN(n18119) );
  XOR2_X1 U16026 ( .A(n12975), .B(n17655), .Z(n12977) );
  NAND2_X1 U16027 ( .A1(n12977), .A2(n12976), .ZN(n12978) );
  XOR2_X1 U16028 ( .A(n12979), .B(n18089), .Z(n12980) );
  XOR2_X1 U16029 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12980), .Z(
        n18096) );
  NAND2_X1 U16030 ( .A1(n12980), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12981) );
  AOI21_X1 U16031 ( .B1(n17649), .B2(n12982), .A(n18068), .ZN(n12984) );
  NAND2_X1 U16032 ( .A1(n12984), .A2(n17961), .ZN(n12985) );
  NAND2_X1 U16033 ( .A1(n12987), .A2(n18360), .ZN(n18067) );
  NAND2_X1 U16034 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18366) );
  INV_X1 U16035 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18026) );
  NOR2_X1 U16036 ( .A1(n18366), .A2(n18026), .ZN(n18337) );
  INV_X1 U16037 ( .A(n18337), .ZN(n18008) );
  NOR2_X1 U16038 ( .A1(n21466), .A2(n18008), .ZN(n18321) );
  INV_X1 U16039 ( .A(n12993), .ZN(n17949) );
  NOR2_X1 U16040 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18039) );
  INV_X1 U16041 ( .A(n18039), .ZN(n12989) );
  NOR2_X2 U16042 ( .A1(n18043), .A2(n12989), .ZN(n18014) );
  NAND2_X1 U16043 ( .A1(n18014), .A2(n18026), .ZN(n18007) );
  NOR2_X2 U16044 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18007), .ZN(
        n17971) );
  NAND3_X1 U16045 ( .A1(n17971), .A2(n21466), .A3(n18327), .ZN(n12990) );
  NAND2_X1 U16046 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18280) );
  INV_X1 U16047 ( .A(n18280), .ZN(n17924) );
  NAND2_X1 U16048 ( .A1(n17924), .A2(n12995), .ZN(n17853) );
  NAND2_X1 U16049 ( .A1(n18030), .A2(n17926), .ZN(n17925) );
  NOR2_X1 U16050 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17925), .ZN(
        n12991) );
  INV_X1 U16051 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18228) );
  NAND2_X1 U16052 ( .A1(n12991), .A2(n18228), .ZN(n17887) );
  INV_X1 U16053 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18213) );
  INV_X1 U16054 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18244) );
  NAND3_X1 U16055 ( .A1(n17880), .A2(n18213), .A3(n18244), .ZN(n12992) );
  OAI21_X1 U16056 ( .B1(n12993), .B2(n17853), .A(n12992), .ZN(n12994) );
  INV_X1 U16057 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17856) );
  NAND2_X1 U16058 ( .A1(n17924), .A2(n17949), .ZN(n17886) );
  NAND3_X1 U16059 ( .A1(n12995), .A2(n17851), .A3(n17857), .ZN(n12996) );
  INV_X1 U16060 ( .A(n12996), .ZN(n17840) );
  NAND2_X1 U16061 ( .A1(n18030), .A2(n17851), .ZN(n17839) );
  NAND2_X1 U16062 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18174) );
  OR2_X1 U16063 ( .A1(n12996), .A2(n18174), .ZN(n12997) );
  NAND2_X1 U16064 ( .A1(n16684), .A2(n13001), .ZN(n13002) );
  OR2_X1 U16065 ( .A1(n13002), .A2(n18068), .ZN(n16055) );
  NOR2_X1 U16066 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16055), .ZN(
        n12999) );
  MUX2_X1 U16067 ( .A(n18068), .B(n12999), .S(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(n13006) );
  NAND2_X1 U16068 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n13000), .ZN(
        n17806) );
  INV_X1 U16069 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17792) );
  NAND2_X1 U16070 ( .A1(n18068), .A2(n17792), .ZN(n16698) );
  INV_X1 U16071 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16056) );
  NOR2_X1 U16072 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16056), .ZN(
        n13258) );
  AOI21_X1 U16073 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n18030), .ZN(n13005) );
  NOR2_X1 U16074 ( .A1(n18068), .A2(n13003), .ZN(n13004) );
  AOI22_X1 U16075 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13010) );
  AOI22_X1 U16076 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13009) );
  AOI22_X1 U16077 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U16078 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13007) );
  NAND4_X1 U16079 ( .A1(n13010), .A2(n13009), .A3(n13008), .A4(n13007), .ZN(
        n13016) );
  INV_X2 U16080 ( .A(n9911), .ZN(n17479) );
  AOI22_X1 U16081 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U16082 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17458), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U16083 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U16084 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13011) );
  NAND4_X1 U16085 ( .A1(n13014), .A2(n13013), .A3(n13012), .A4(n13011), .ZN(
        n13015) );
  NAND2_X1 U16086 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18968), .ZN(
        n13127) );
  OAI21_X1 U16087 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18968), .A(
        n13127), .ZN(n13130) );
  AOI22_X1 U16088 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18969), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19121), .ZN(n13126) );
  OAI22_X1 U16089 ( .A1(n13017), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13028) );
  INV_X1 U16090 ( .A(n13127), .ZN(n13018) );
  OAI22_X1 U16091 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18502), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13021), .ZN(n13023) );
  NOR2_X1 U16092 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18502), .ZN(
        n13022) );
  NAND2_X1 U16093 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13021), .ZN(
        n13024) );
  AOI22_X1 U16094 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13023), .B1(
        n13022), .B2(n13024), .ZN(n13027) );
  NAND2_X1 U16095 ( .A1(n13126), .A2(n13027), .ZN(n13030) );
  AOI21_X1 U16096 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13024), .A(
        n13023), .ZN(n13025) );
  NAND2_X1 U16097 ( .A1(n13029), .A2(n13028), .ZN(n13026) );
  OAI211_X1 U16098 ( .C1(n13029), .C2(n13028), .A(n13027), .B(n13026), .ZN(
        n13131) );
  OAI211_X1 U16099 ( .C1(n13130), .C2(n13030), .A(n13128), .B(n13131), .ZN(
        n18946) );
  AOI22_X1 U16100 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U16101 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U16102 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U16103 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13031) );
  NAND4_X1 U16104 ( .A1(n13034), .A2(n13033), .A3(n13032), .A4(n13031), .ZN(
        n13040) );
  AOI22_X1 U16105 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13038) );
  AOI22_X1 U16106 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U16107 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U16108 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13035) );
  NAND4_X1 U16109 ( .A1(n13038), .A2(n13037), .A3(n13036), .A4(n13035), .ZN(
        n13039) );
  AOI22_X1 U16110 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13044) );
  AOI22_X1 U16111 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U16112 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16113 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13041) );
  NAND4_X1 U16114 ( .A1(n13044), .A2(n13043), .A3(n13042), .A4(n13041), .ZN(
        n13050) );
  AOI22_X1 U16115 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U16116 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U16117 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U16118 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13045) );
  NAND4_X1 U16119 ( .A1(n13048), .A2(n13047), .A3(n13046), .A4(n13045), .ZN(
        n13049) );
  AOI22_X1 U16120 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17450), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16121 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17433), .ZN(n13053) );
  AOI22_X1 U16122 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U16123 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17472), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13051) );
  NAND4_X1 U16124 ( .A1(n13054), .A2(n13053), .A3(n13052), .A4(n13051), .ZN(
        n13060) );
  AOI22_X1 U16125 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n9823), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17456), .ZN(n13058) );
  AOI22_X1 U16126 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U16127 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n15918), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U16128 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17457), .ZN(n13055) );
  NAND4_X1 U16129 ( .A1(n13058), .A2(n13057), .A3(n13056), .A4(n13055), .ZN(
        n13059) );
  AOI22_X1 U16130 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16131 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13070) );
  INV_X1 U16132 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15907) );
  AOI22_X1 U16133 ( .A1(n12922), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13061) );
  OAI21_X1 U16134 ( .B1(n13062), .B2(n15907), .A(n13061), .ZN(n13068) );
  AOI22_X1 U16135 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16136 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U16137 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16138 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13063) );
  NAND4_X1 U16139 ( .A1(n13066), .A2(n13065), .A3(n13064), .A4(n13063), .ZN(
        n13067) );
  NAND2_X1 U16140 ( .A1(n18545), .A2(n18508), .ZN(n13110) );
  INV_X1 U16141 ( .A(n13110), .ZN(n13114) );
  AOI22_X1 U16142 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U16143 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17458), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13074) );
  AOI22_X1 U16144 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U16145 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13072) );
  NAND4_X1 U16146 ( .A1(n13075), .A2(n13074), .A3(n13073), .A4(n13072), .ZN(
        n13079) );
  AOI22_X1 U16147 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13078) );
  AOI22_X1 U16148 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U16149 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13090), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U16150 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U16151 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13082) );
  AOI22_X1 U16152 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13081) );
  AOI22_X1 U16153 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13080) );
  NAND4_X1 U16154 ( .A1(n13083), .A2(n13082), .A3(n13081), .A4(n13080), .ZN(
        n13089) );
  AOI22_X1 U16155 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16156 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U16157 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U16158 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17458), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13084) );
  NAND4_X1 U16159 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13088) );
  NAND2_X1 U16160 ( .A1(n18531), .A2(n18535), .ZN(n13103) );
  INV_X1 U16161 ( .A(n13103), .ZN(n13240) );
  NAND4_X1 U16162 ( .A1(n18521), .A2(n13117), .A3(n13114), .A4(n13240), .ZN(
        n18949) );
  AOI22_X1 U16163 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13090), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16164 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16165 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16166 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13091) );
  NAND4_X1 U16167 ( .A1(n13094), .A2(n13093), .A3(n13092), .A4(n13091), .ZN(
        n13100) );
  AOI22_X1 U16168 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U16169 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17458), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U16170 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U16171 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9823), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13095) );
  NAND4_X1 U16172 ( .A1(n13098), .A2(n13097), .A3(n13096), .A4(n13095), .ZN(
        n13099) );
  NAND2_X1 U16173 ( .A1(n18516), .A2(n13124), .ZN(n13102) );
  AOI21_X1 U16174 ( .B1(n18545), .B2(n13103), .A(n13117), .ZN(n13101) );
  AOI21_X1 U16175 ( .B1(n13103), .B2(n13102), .A(n13101), .ZN(n13112) );
  INV_X1 U16176 ( .A(n13117), .ZN(n18528) );
  NAND2_X1 U16177 ( .A1(n17526), .A2(n18528), .ZN(n18953) );
  INV_X1 U16178 ( .A(n13115), .ZN(n13113) );
  AND2_X1 U16179 ( .A1(n18953), .A2(n13113), .ZN(n13106) );
  NOR2_X2 U16180 ( .A1(n18535), .A2(n17533), .ZN(n18964) );
  NAND2_X1 U16181 ( .A1(n19152), .A2(n17683), .ZN(n13119) );
  INV_X1 U16182 ( .A(n13119), .ZN(n13104) );
  OAI21_X1 U16183 ( .B1(n17612), .B2(n18964), .A(n13104), .ZN(n13241) );
  OAI211_X1 U16184 ( .C1(n18531), .C2(n13106), .A(n13241), .B(n18516), .ZN(
        n13105) );
  INV_X1 U16185 ( .A(n13105), .ZN(n13108) );
  OAI211_X1 U16186 ( .C1(n18964), .C2(n18508), .A(n18516), .B(n13106), .ZN(
        n13107) );
  OAI21_X1 U16187 ( .B1(n13108), .B2(n18521), .A(n13107), .ZN(n13109) );
  AOI21_X1 U16188 ( .B1(n18521), .B2(n13110), .A(n13109), .ZN(n13111) );
  NAND2_X1 U16189 ( .A1(n13112), .A2(n13111), .ZN(n13122) );
  NAND2_X1 U16190 ( .A1(n18516), .A2(n18521), .ZN(n18952) );
  NOR2_X1 U16191 ( .A1(n17612), .A2(n18521), .ZN(n13121) );
  NAND2_X1 U16192 ( .A1(n18516), .A2(n13121), .ZN(n13120) );
  NOR3_X1 U16193 ( .A1(n18964), .A2(n13115), .A3(n13120), .ZN(n13116) );
  NOR2_X1 U16194 ( .A1(n18516), .A2(n18949), .ZN(n13243) );
  NOR2_X2 U16195 ( .A1(n13118), .A2(n13243), .ZN(n16813) );
  NOR2_X2 U16196 ( .A1(n15972), .A2(n15971), .ZN(n18975) );
  INV_X2 U16197 ( .A(n18975), .ZN(n18967) );
  NAND2_X1 U16198 ( .A1(n13124), .A2(n13119), .ZN(n19163) );
  NOR3_X1 U16199 ( .A1(n17533), .A2(n13120), .A3(n18953), .ZN(n15979) );
  NOR2_X1 U16200 ( .A1(n19152), .A2(n13121), .ZN(n13123) );
  AOI21_X1 U16201 ( .B1(n13123), .B2(n18938), .A(n13122), .ZN(n18951) );
  OAI21_X2 U16202 ( .B1(n18952), .B2(n15971), .A(n18951), .ZN(n18965) );
  OAI21_X1 U16203 ( .B1(n15979), .B2(n13125), .A(n13124), .ZN(n13236) );
  XOR2_X1 U16204 ( .A(n13127), .B(n13126), .Z(n13129) );
  OAI21_X1 U16205 ( .B1(n13131), .B2(n13130), .A(n18941), .ZN(n13132) );
  INV_X1 U16206 ( .A(n13132), .ZN(n18943) );
  NAND2_X1 U16207 ( .A1(n18516), .A2(n18511), .ZN(n13238) );
  NOR2_X1 U16208 ( .A1(n17526), .A2(n13238), .ZN(n13237) );
  NAND2_X1 U16209 ( .A1(n18943), .A2(n13237), .ZN(n13245) );
  OAI22_X2 U16210 ( .A1(n18946), .A2(n18227), .B1(n13236), .B2(n13245), .ZN(
        n18947) );
  NAND2_X1 U16211 ( .A1(n13249), .A2(n18069), .ZN(n13178) );
  INV_X1 U16212 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18170) );
  NOR2_X1 U16213 ( .A1(n18170), .A2(n17792), .ZN(n16682) );
  NAND2_X1 U16214 ( .A1(n16682), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16058) );
  INV_X1 U16215 ( .A(n17853), .ZN(n18196) );
  NAND3_X1 U16216 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18196), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18187) );
  INV_X1 U16217 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18186) );
  NOR2_X1 U16218 ( .A1(n18187), .A2(n18186), .ZN(n13254) );
  INV_X1 U16219 ( .A(n13254), .ZN(n18169) );
  NOR2_X1 U16220 ( .A1(n17681), .A2(n18163), .ZN(n13138) );
  NOR2_X1 U16221 ( .A1(n13138), .A2(n17668), .ZN(n13137) );
  NOR2_X1 U16222 ( .A1(n13136), .A2(n13137), .ZN(n13135) );
  NAND2_X1 U16223 ( .A1(n13135), .A2(n17659), .ZN(n13134) );
  NOR2_X1 U16224 ( .A1(n17655), .A2(n13134), .ZN(n18088) );
  NAND2_X1 U16225 ( .A1(n18088), .A2(n18089), .ZN(n13133) );
  NOR2_X1 U16226 ( .A1(n17649), .A2(n13133), .ZN(n13155) );
  INV_X1 U16227 ( .A(n17649), .ZN(n16703) );
  XNOR2_X1 U16228 ( .A(n16703), .B(n13133), .ZN(n13152) );
  XOR2_X1 U16229 ( .A(n17655), .B(n13134), .Z(n13147) );
  AND2_X1 U16230 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13147), .ZN(
        n13148) );
  XOR2_X1 U16231 ( .A(n17659), .B(n13135), .Z(n13145) );
  AND2_X1 U16232 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13145), .ZN(
        n13146) );
  INV_X1 U16233 ( .A(n13136), .ZN(n17664) );
  XOR2_X1 U16234 ( .A(n17664), .B(n13137), .Z(n13143) );
  NOR2_X1 U16235 ( .A1(n18446), .A2(n13143), .ZN(n13144) );
  XOR2_X1 U16236 ( .A(n17668), .B(n13138), .Z(n13141) );
  NOR2_X1 U16237 ( .A1(n13141), .A2(n18457), .ZN(n13142) );
  NOR2_X1 U16238 ( .A1(n17681), .A2(n19125), .ZN(n13140) );
  NAND3_X1 U16239 ( .A1(n18163), .A2(n17681), .A3(n19125), .ZN(n13139) );
  OAI221_X1 U16240 ( .B1(n13140), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18163), .C2(n17681), .A(n13139), .ZN(n18144) );
  XOR2_X1 U16241 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13141), .Z(
        n18143) );
  NOR2_X1 U16242 ( .A1(n18144), .A2(n18143), .ZN(n18142) );
  NOR2_X1 U16243 ( .A1(n13142), .A2(n18142), .ZN(n18134) );
  XOR2_X1 U16244 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13143), .Z(
        n18133) );
  NOR2_X1 U16245 ( .A1(n18134), .A2(n18133), .ZN(n18132) );
  NOR2_X1 U16246 ( .A1(n13144), .A2(n18132), .ZN(n18116) );
  INV_X1 U16247 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18444) );
  XOR2_X1 U16248 ( .A(n18444), .B(n13145), .Z(n18115) );
  NOR2_X1 U16249 ( .A1(n18116), .A2(n18115), .ZN(n18114) );
  NOR2_X1 U16250 ( .A1(n13146), .A2(n18114), .ZN(n18105) );
  XNOR2_X1 U16251 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n13147), .ZN(
        n18104) );
  INV_X1 U16252 ( .A(n18088), .ZN(n18086) );
  XOR2_X1 U16253 ( .A(n18089), .B(n18086), .Z(n13149) );
  INV_X1 U16254 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18418) );
  AOI222_X1 U16255 ( .A1(n18087), .A2(n13149), .B1(n18087), .B2(n18418), .C1(
        n13149), .C2(n18418), .ZN(n13151) );
  NOR2_X1 U16256 ( .A1(n13152), .A2(n13151), .ZN(n18075) );
  INV_X1 U16257 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18411) );
  NOR2_X1 U16258 ( .A1(n18075), .A2(n18411), .ZN(n13150) );
  NAND2_X1 U16259 ( .A1(n13155), .A2(n13150), .ZN(n13156) );
  INV_X1 U16260 ( .A(n13150), .ZN(n13154) );
  AND2_X1 U16261 ( .A1(n13152), .A2(n13151), .ZN(n18076) );
  AOI21_X1 U16262 ( .B1(n13155), .B2(n13154), .A(n18076), .ZN(n13153) );
  OAI21_X1 U16263 ( .B1(n13155), .B2(n13154), .A(n13153), .ZN(n18059) );
  NAND2_X1 U16264 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18059), .ZN(
        n18058) );
  NAND2_X1 U16265 ( .A1(n13156), .A2(n18058), .ZN(n18023) );
  NOR2_X1 U16266 ( .A1(n18169), .A2(n18306), .ZN(n18177) );
  INV_X1 U16267 ( .A(n18177), .ZN(n13157) );
  NAND2_X1 U16268 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16683), .ZN(
        n13158) );
  XOR2_X1 U16269 ( .A(n13003), .B(n13158), .Z(n13262) );
  INV_X1 U16270 ( .A(n13262), .ZN(n13160) );
  NOR2_X2 U16271 ( .A1(n18511), .A2(n16814), .ZN(n18157) );
  NOR2_X1 U16272 ( .A1(n13160), .A2(n13159), .ZN(n13176) );
  INV_X1 U16273 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19005) );
  OAI21_X1 U16274 ( .B1(n19109), .B2(n19005), .A(n19102), .ZN(n15966) );
  INV_X1 U16275 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19151) );
  INV_X1 U16276 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16857) );
  INV_X1 U16277 ( .A(n18019), .ZN(n16968) );
  NAND3_X1 U16278 ( .A1(n17989), .A2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17974) );
  NAND3_X1 U16279 ( .A1(n17874), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17819) );
  INV_X1 U16280 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16842) );
  INV_X1 U16281 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17812) );
  INV_X1 U16282 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16882) );
  NOR2_X1 U16283 ( .A1(n17812), .A2(n16882), .ZN(n13163) );
  INV_X1 U16284 ( .A(n13163), .ZN(n17801) );
  XOR2_X2 U16285 ( .A(n16857), .B(n13161), .Z(n17157) );
  INV_X1 U16286 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19088) );
  NOR2_X1 U16287 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19124) );
  INV_X1 U16288 ( .A(n19124), .ZN(n17198) );
  NOR2_X1 U16289 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n17198), .ZN(n19165) );
  NAND2_X2 U16290 ( .A1(n19165), .A2(n19099), .ZN(n18484) );
  NOR2_X1 U16291 ( .A1(n19088), .A2(n18484), .ZN(n13255) );
  INV_X1 U16292 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16673) );
  INV_X1 U16293 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21330) );
  NAND2_X1 U16294 ( .A1(n19099), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18165) );
  INV_X1 U16295 ( .A(n18165), .ZN(n17986) );
  NAND3_X1 U16296 ( .A1(n19005), .A2(n19102), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18847) );
  OAI21_X2 U16297 ( .B1(n21330), .B2(n17898), .A(n18540), .ZN(n17988) );
  NAND2_X1 U16298 ( .A1(n13162), .A2(n17988), .ZN(n16672) );
  NOR2_X1 U16299 ( .A1(n16673), .A2(n16672), .ZN(n13168) );
  NOR2_X1 U16300 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17898), .ZN(
        n16690) );
  NOR2_X1 U16301 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16672), .ZN(
        n13166) );
  NOR2_X1 U16302 ( .A1(n21330), .A2(n17786), .ZN(n16843) );
  NAND2_X1 U16303 ( .A1(n16843), .A2(n13163), .ZN(n16689) );
  INV_X1 U16304 ( .A(n16689), .ZN(n16840) );
  NAND2_X1 U16305 ( .A1(n18883), .A2(n13164), .ZN(n13165) );
  OAI211_X1 U16306 ( .C1(n16840), .C2(n18165), .A(n18164), .B(n13165), .ZN(
        n16691) );
  NOR3_X1 U16307 ( .A1(n16690), .A2(n13166), .A3(n16691), .ZN(n16671) );
  INV_X1 U16308 ( .A(n16671), .ZN(n13167) );
  MUX2_X1 U16309 ( .A(n13168), .B(n13167), .S(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n13169) );
  AOI211_X1 U16310 ( .C1(n18006), .C2(n17157), .A(n13255), .B(n13169), .ZN(
        n13174) );
  NAND2_X1 U16311 ( .A1(n18341), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17979) );
  INV_X1 U16312 ( .A(n17979), .ZN(n13170) );
  NOR2_X1 U16313 ( .A1(n18327), .A2(n18296), .ZN(n13251) );
  NOR2_X1 U16314 ( .A1(n18305), .A2(n18169), .ZN(n17791) );
  INV_X1 U16315 ( .A(n17791), .ZN(n18179) );
  NAND2_X1 U16316 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16681), .ZN(
        n13171) );
  XNOR2_X1 U16317 ( .A(n13003), .B(n13171), .ZN(n13260) );
  INV_X1 U16318 ( .A(n13260), .ZN(n13172) );
  NOR2_X2 U16319 ( .A1(n16703), .A2(n18168), .ZN(n18070) );
  NAND2_X1 U16320 ( .A1(n13172), .A2(n18070), .ZN(n13173) );
  NAND2_X1 U16321 ( .A1(n13174), .A2(n13173), .ZN(n13175) );
  NAND2_X1 U16322 ( .A1(n13178), .A2(n13177), .ZN(P3_U2799) );
  AND2_X1 U16323 ( .A1(n13206), .A2(n13180), .ZN(n13181) );
  OR2_X1 U16324 ( .A1(n13181), .A2(n13208), .ZN(n15412) );
  OR2_X1 U16325 ( .A1(n13183), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13184) );
  NAND2_X1 U16326 ( .A1(n13182), .A2(n13184), .ZN(n16420) );
  INV_X1 U16327 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16450) );
  AOI21_X1 U16328 ( .B1(n16450), .B2(n13203), .A(n13204), .ZN(n13185) );
  INV_X1 U16329 ( .A(n13185), .ZN(n16458) );
  AOI21_X1 U16330 ( .B1(n19196), .B2(n13202), .A(n9967), .ZN(n15475) );
  INV_X1 U16331 ( .A(n15475), .ZN(n19205) );
  AOI21_X1 U16332 ( .B1(n10160), .B2(n15497), .A(n13186), .ZN(n15499) );
  INV_X1 U16333 ( .A(n15499), .ZN(n19217) );
  AOI21_X1 U16334 ( .B1(n15530), .B2(n13197), .A(n13199), .ZN(n19262) );
  AOI21_X1 U16335 ( .B1(n15541), .B2(n13195), .A(n13198), .ZN(n15539) );
  AOI21_X1 U16336 ( .B1(n16508), .B2(n13194), .A(n13196), .ZN(n16501) );
  AOI21_X1 U16337 ( .B1(n16527), .B2(n13192), .A(n13187), .ZN(n19315) );
  AOI21_X1 U16338 ( .B1(n15550), .B2(n13191), .A(n13193), .ZN(n19325) );
  AOI21_X1 U16339 ( .B1(n16548), .B2(n13189), .A(n9881), .ZN(n19359) );
  AOI21_X1 U16340 ( .B1(n16562), .B2(n13188), .A(n13190), .ZN(n16549) );
  OAI22_X1 U16341 ( .A1(n16656), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19384) );
  INV_X1 U16342 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15192) );
  OAI22_X1 U16343 ( .A1(n16656), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15192), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15200) );
  AND2_X1 U16344 ( .A1(n19384), .A2(n15200), .ZN(n14330) );
  OAI21_X1 U16345 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n13188), .ZN(n14331) );
  NAND2_X1 U16346 ( .A1(n14330), .A2(n14331), .ZN(n15177) );
  NOR2_X1 U16347 ( .A1(n16549), .A2(n15177), .ZN(n14276) );
  OAI21_X1 U16348 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13190), .A(
        n13189), .ZN(n19498) );
  NAND2_X1 U16349 ( .A1(n14276), .A2(n19498), .ZN(n19357) );
  NOR2_X1 U16350 ( .A1(n19359), .A2(n19357), .ZN(n19339) );
  OAI21_X1 U16351 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9881), .A(
        n13191), .ZN(n19341) );
  NAND2_X1 U16352 ( .A1(n19339), .A2(n19341), .ZN(n19324) );
  NOR2_X1 U16353 ( .A1(n19325), .A2(n19324), .ZN(n14289) );
  OAI21_X1 U16354 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13193), .A(
        n13192), .ZN(n16540) );
  NAND2_X1 U16355 ( .A1(n14289), .A2(n16540), .ZN(n19314) );
  NOR2_X1 U16356 ( .A1(n19315), .A2(n19314), .ZN(n19307) );
  OAI21_X1 U16357 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13187), .A(
        n13194), .ZN(n19308) );
  NAND2_X1 U16358 ( .A1(n19307), .A2(n19308), .ZN(n15164) );
  NOR2_X1 U16359 ( .A1(n16501), .A2(n15164), .ZN(n19294) );
  OAI21_X1 U16360 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13196), .A(
        n13195), .ZN(n19300) );
  NAND2_X1 U16361 ( .A1(n19294), .A2(n19300), .ZN(n19287) );
  NOR2_X1 U16362 ( .A1(n15539), .A2(n19287), .ZN(n19270) );
  OAI21_X1 U16363 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13198), .A(
        n13197), .ZN(n19271) );
  AOI21_X1 U16364 ( .B1(n19262), .B2(n10150), .A(n19261), .ZN(n19257) );
  OAI21_X1 U16365 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13199), .A(
        n9971), .ZN(n19256) );
  NAND2_X1 U16366 ( .A1(n19257), .A2(n19256), .ZN(n19255) );
  NAND2_X1 U16367 ( .A1(n19255), .A2(n9877), .ZN(n19242) );
  AOI21_X1 U16368 ( .B1(n19235), .B2(n9971), .A(n13201), .ZN(n13200) );
  INV_X1 U16369 ( .A(n13200), .ZN(n19243) );
  NAND2_X1 U16370 ( .A1(n19242), .A2(n19243), .ZN(n19241) );
  NAND2_X1 U16371 ( .A1(n9877), .A2(n19241), .ZN(n19228) );
  OAI21_X1 U16372 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13201), .A(
        n10160), .ZN(n19229) );
  NAND2_X1 U16373 ( .A1(n19228), .A2(n19229), .ZN(n19227) );
  NAND2_X1 U16374 ( .A1(n9875), .A2(n19227), .ZN(n19216) );
  NAND2_X1 U16375 ( .A1(n19217), .A2(n19216), .ZN(n19215) );
  NAND2_X1 U16376 ( .A1(n19215), .A2(n9876), .ZN(n15152) );
  OAI21_X1 U16377 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n13186), .A(
        n13202), .ZN(n15485) );
  NAND2_X1 U16378 ( .A1(n15152), .A2(n15485), .ZN(n15151) );
  NAND2_X1 U16379 ( .A1(n9877), .A2(n15151), .ZN(n19204) );
  NAND2_X1 U16380 ( .A1(n19205), .A2(n19204), .ZN(n19203) );
  NAND2_X1 U16381 ( .A1(n19203), .A2(n9876), .ZN(n16005) );
  OAI21_X1 U16382 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n9967), .A(
        n13203), .ZN(n16488) );
  NAND2_X1 U16383 ( .A1(n16005), .A2(n16488), .ZN(n16004) );
  NAND2_X1 U16384 ( .A1(n9876), .A2(n16004), .ZN(n16457) );
  NAND2_X1 U16385 ( .A1(n16458), .A2(n16457), .ZN(n16456) );
  NAND2_X1 U16386 ( .A1(n16456), .A2(n9876), .ZN(n16444) );
  OAI21_X1 U16387 ( .B1(n13204), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n13205), .ZN(n16445) );
  NAND2_X1 U16388 ( .A1(n16444), .A2(n16445), .ZN(n16443) );
  AOI21_X1 U16389 ( .B1(n15439), .B2(n13205), .A(n13183), .ZN(n15442) );
  INV_X1 U16390 ( .A(n15442), .ZN(n16432) );
  NAND2_X1 U16391 ( .A1(n16431), .A2(n16432), .ZN(n16430) );
  NAND2_X1 U16392 ( .A1(n9876), .A2(n16430), .ZN(n16419) );
  NAND2_X1 U16393 ( .A1(n16420), .A2(n16419), .ZN(n16418) );
  INV_X1 U16394 ( .A(n13206), .ZN(n13207) );
  AOI21_X1 U16395 ( .B1(n16400), .B2(n13182), .A(n13207), .ZN(n15421) );
  INV_X1 U16396 ( .A(n15421), .ZN(n16408) );
  NAND2_X1 U16397 ( .A1(n16407), .A2(n16408), .ZN(n16406) );
  NAND2_X1 U16398 ( .A1(n9876), .A2(n16406), .ZN(n15140) );
  NAND2_X1 U16399 ( .A1(n15412), .A2(n15140), .ZN(n15139) );
  NAND2_X1 U16400 ( .A1(n15139), .A2(n9875), .ZN(n16394) );
  OAI21_X1 U16401 ( .B1(n13208), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n12849), .ZN(n16395) );
  NAND2_X1 U16402 ( .A1(n16394), .A2(n16395), .ZN(n16393) );
  NAND2_X1 U16403 ( .A1(n9876), .A2(n16393), .ZN(n16381) );
  INV_X2 U16404 ( .A(n19334), .ZN(n20102) );
  NAND2_X1 U16405 ( .A1(n16382), .A2(n16381), .ZN(n13209) );
  OAI211_X1 U16406 ( .C1(n16381), .C2(n16382), .A(n20102), .B(n13209), .ZN(
        n13235) );
  NAND2_X1 U16407 ( .A1(n12463), .A2(n16665), .ZN(n13210) );
  INV_X1 U16408 ( .A(n20108), .ZN(n20124) );
  NOR2_X1 U16409 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20124), .ZN(n13223) );
  AND2_X1 U16410 ( .A1(n13214), .A2(n13223), .ZN(n13211) );
  INV_X1 U16411 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13212) );
  NOR2_X1 U16412 ( .A1(n13223), .A2(n13212), .ZN(n13213) );
  NAND2_X1 U16413 ( .A1(n13214), .A2(n13213), .ZN(n13215) );
  NOR2_X2 U16414 ( .A1(n13219), .A2(n13215), .ZN(n19367) );
  NOR2_X1 U16415 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19873), .ZN(n19768) );
  NAND2_X1 U16416 ( .A1(n13216), .A2(n19768), .ZN(n16666) );
  NAND2_X1 U16417 ( .A1(n16666), .A2(n19334), .ZN(n13217) );
  NOR2_X1 U16418 ( .A1(n19247), .A2(n13217), .ZN(n13218) );
  NOR2_X2 U16419 ( .A1(n19873), .A2(n19369), .ZN(n19356) );
  NOR2_X1 U16420 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n15820), .ZN(n13224) );
  AND2_X1 U16421 ( .A1(n13220), .A2(n13224), .ZN(n16653) );
  NAND2_X1 U16422 ( .A1(n13640), .A2(n19275), .ZN(n13229) );
  NAND2_X1 U16423 ( .A1(n16654), .A2(n13221), .ZN(n13222) );
  OAI21_X1 U16424 ( .B1(P2_EBX_REG_31__SCAN_IN), .B2(n13223), .A(n14211), .ZN(
        n13226) );
  INV_X1 U16425 ( .A(n13224), .ZN(n13225) );
  NAND2_X1 U16426 ( .A1(n13226), .A2(n13225), .ZN(n13227) );
  NOR2_X2 U16427 ( .A1(n13680), .A2(n13227), .ZN(n19368) );
  AOI22_X1 U16428 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19368), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19369), .ZN(n13228) );
  OAI211_X1 U16429 ( .C1(n12810), .C2(n19378), .A(n13229), .B(n13228), .ZN(
        n13230) );
  AOI21_X1 U16430 ( .B1(n13231), .B2(n19367), .A(n13230), .ZN(n13232) );
  NAND2_X1 U16431 ( .A1(n13235), .A2(n13234), .ZN(P2_U2825) );
  INV_X1 U16432 ( .A(n13236), .ZN(n13242) );
  NAND2_X1 U16433 ( .A1(n13242), .A2(n13237), .ZN(n18942) );
  NAND2_X1 U16434 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19153) );
  NOR2_X1 U16435 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n19017) );
  NOR2_X1 U16436 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19017), .ZN(n19026) );
  INV_X1 U16437 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21390) );
  NOR2_X1 U16438 ( .A1(n19034), .A2(n19161), .ZN(n19027) );
  NAND2_X1 U16439 ( .A1(n19026), .A2(n19090), .ZN(n19150) );
  OAI211_X1 U16440 ( .C1(n18516), .C2(n18511), .A(n13238), .B(n19150), .ZN(
        n13239) );
  NAND2_X1 U16441 ( .A1(n19153), .A2(n13239), .ZN(n16810) );
  AOI211_X1 U16442 ( .C1(n18516), .C2(n18531), .A(n16811), .B(n16810), .ZN(
        n13248) );
  AOI21_X1 U16443 ( .B1(n18516), .B2(n13240), .A(n18528), .ZN(n13246) );
  OAI21_X1 U16444 ( .B1(n13243), .B2(n13242), .A(n13241), .ZN(n13244) );
  INV_X1 U16445 ( .A(n13244), .ZN(n15975) );
  OAI211_X1 U16446 ( .C1(n13246), .C2(n18946), .A(n15975), .B(n13245), .ZN(
        n13247) );
  NOR3_X2 U16447 ( .A1(n17649), .A2(n18942), .A3(n18490), .ZN(n18404) );
  NAND2_X1 U16448 ( .A1(n13249), .A2(n18404), .ZN(n13264) );
  NAND2_X1 U16449 ( .A1(n9866), .A2(n18473), .ZN(n18422) );
  NOR2_X1 U16450 ( .A1(n18942), .A2(n18490), .ZN(n18487) );
  NOR2_X1 U16451 ( .A1(n16703), .A2(n18482), .ZN(n18405) );
  INV_X1 U16452 ( .A(n18405), .ZN(n18335) );
  NOR2_X1 U16453 ( .A1(n18169), .A2(n18490), .ZN(n16710) );
  AND3_X1 U16454 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18419) );
  AND2_X1 U16455 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18419), .ZN(
        n18392) );
  NAND3_X1 U16456 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n18392), .ZN(n18336) );
  AOI21_X1 U16457 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18462) );
  NOR2_X1 U16458 ( .A1(n18336), .A2(n18462), .ZN(n18293) );
  AND2_X1 U16459 ( .A1(n18321), .A2(n18293), .ZN(n18322) );
  NAND2_X1 U16460 ( .A1(n13250), .A2(n18322), .ZN(n18234) );
  INV_X1 U16461 ( .A(n18336), .ZN(n18273) );
  NAND2_X1 U16462 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18272) );
  INV_X1 U16463 ( .A(n18272), .ZN(n18437) );
  NAND2_X1 U16464 ( .A1(n18273), .A2(n18437), .ZN(n18320) );
  NOR2_X1 U16465 ( .A1(n17962), .A2(n18343), .ZN(n18274) );
  INV_X1 U16466 ( .A(n18274), .ZN(n17955) );
  NOR2_X1 U16467 ( .A1(n18320), .A2(n17955), .ZN(n18319) );
  NAND2_X1 U16468 ( .A1(n13251), .A2(n18319), .ZN(n18295) );
  AOI21_X1 U16469 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18965), .A(
        n18967), .ZN(n18466) );
  OAI22_X1 U16470 ( .A1(n18981), .A2(n18234), .B1(n18295), .B2(n18466), .ZN(
        n18195) );
  NAND2_X1 U16471 ( .A1(n16710), .A2(n18195), .ZN(n15996) );
  NOR2_X1 U16472 ( .A1(n16058), .A2(n15996), .ZN(n13257) );
  NAND2_X1 U16473 ( .A1(n18393), .A2(n18473), .ZN(n18475) );
  INV_X1 U16474 ( .A(n18475), .ZN(n18438) );
  NAND2_X1 U16475 ( .A1(n18975), .A2(n18956), .ZN(n18396) );
  NOR2_X1 U16476 ( .A1(n18956), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18461) );
  NOR2_X1 U16477 ( .A1(n18461), .A2(n18295), .ZN(n18276) );
  NAND2_X1 U16478 ( .A1(n17924), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18245) );
  NOR3_X1 U16479 ( .A1(n17861), .A2(n18234), .A3(n18245), .ZN(n18193) );
  NAND2_X1 U16480 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18194) );
  NOR2_X1 U16481 ( .A1(n18174), .A2(n18194), .ZN(n13252) );
  AOI21_X1 U16482 ( .B1(n18193), .B2(n13252), .A(n18981), .ZN(n18173) );
  AOI211_X1 U16483 ( .C1(n18965), .C2(n18170), .A(n18173), .B(n18490), .ZN(
        n13253) );
  OAI221_X1 U16484 ( .B1(n18459), .B2(n13254), .C1(n18459), .C2(n18276), .A(
        n13253), .ZN(n15993) );
  AOI22_X1 U16485 ( .A1(n18438), .A2(n16058), .B1(n18484), .B2(n15993), .ZN(
        n16060) );
  AOI221_X1 U16486 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16060), 
        .C1(n18475), .C2(n16060), .A(n13003), .ZN(n13256) );
  AOI211_X1 U16487 ( .C1(n13258), .C2(n13257), .A(n13256), .B(n13255), .ZN(
        n13259) );
  NAND2_X1 U16488 ( .A1(n13264), .A2(n13263), .ZN(P3_U2831) );
  NAND2_X1 U16489 ( .A1(n19557), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13265) );
  NAND2_X1 U16490 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19907) );
  NAND2_X1 U16491 ( .A1(n19907), .A2(n21487), .ZN(n13267) );
  NAND2_X1 U16492 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20012) );
  INV_X1 U16493 ( .A(n20012), .ZN(n13266) );
  AND2_X1 U16494 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13266), .ZN(
        n13289) );
  INV_X1 U16495 ( .A(n13289), .ZN(n13290) );
  AND2_X1 U16496 ( .A1(n13267), .A2(n13290), .ZN(n19673) );
  AOI22_X1 U16497 ( .A1(n13292), .A2(n16615), .B1(n20206), .B2(n19673), .ZN(
        n13273) );
  INV_X1 U16498 ( .A(n13273), .ZN(n13269) );
  INV_X1 U16499 ( .A(n19557), .ZN(n13757) );
  INV_X1 U16500 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14360) );
  INV_X1 U16501 ( .A(n13271), .ZN(n13272) );
  AND2_X1 U16502 ( .A1(n13273), .A2(n13272), .ZN(n13274) );
  NAND2_X1 U16503 ( .A1(n13275), .A2(n13274), .ZN(n13276) );
  NAND2_X1 U16504 ( .A1(n13292), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13278) );
  OAI21_X1 U16505 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19907), .ZN(n19672) );
  INV_X1 U16506 ( .A(n19672), .ZN(n13277) );
  NAND2_X1 U16507 ( .A1(n13277), .A2(n20206), .ZN(n19882) );
  NAND2_X1 U16508 ( .A1(n13278), .A2(n19882), .ZN(n13279) );
  AOI22_X1 U16509 ( .A1(n13292), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20206), .B2(n20233), .ZN(n13280) );
  NAND2_X1 U16510 ( .A1(n13546), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13282) );
  INV_X1 U16511 ( .A(n13282), .ZN(n13283) );
  NOR2_X1 U16512 ( .A1(n15819), .A2(n13283), .ZN(n13284) );
  NAND2_X1 U16513 ( .A1(n13828), .A2(n13829), .ZN(n13286) );
  NAND2_X1 U16514 ( .A1(n13288), .A2(n13287), .ZN(n13294) );
  NAND2_X1 U16515 ( .A1(n13289), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14272) );
  NAND2_X1 U16516 ( .A1(n20209), .A2(n13290), .ZN(n13291) );
  AND3_X1 U16517 ( .A1(n14272), .A2(n20206), .A3(n13291), .ZN(n19944) );
  AOI21_X1 U16518 ( .B1(n13292), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19944), .ZN(n13293) );
  NAND2_X1 U16519 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n14211), .ZN(
        n13295) );
  NOR2_X1 U16520 ( .A1(n13295), .A2(n19557), .ZN(n13296) );
  NOR2_X1 U16521 ( .A1(n13913), .A2(n19545), .ZN(n13893) );
  OAI211_X1 U16522 ( .C1(n13890), .C2(n13297), .A(n13296), .B(n13891), .ZN(
        n13883) );
  INV_X1 U16523 ( .A(n13883), .ZN(n13298) );
  NAND2_X1 U16524 ( .A1(n13298), .A2(n10383), .ZN(n13901) );
  INV_X1 U16525 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13299) );
  NOR2_X2 U16526 ( .A1(n13901), .A2(n13299), .ZN(n13966) );
  NAND2_X1 U16527 ( .A1(n13966), .A2(n13970), .ZN(n13968) );
  INV_X1 U16528 ( .A(n13968), .ZN(n13301) );
  NAND2_X1 U16529 ( .A1(n13301), .A2(n13300), .ZN(n14029) );
  INV_X1 U16530 ( .A(n14029), .ZN(n13303) );
  NAND2_X1 U16531 ( .A1(n13303), .A2(n13302), .ZN(n14089) );
  AND2_X2 U16532 ( .A1(n14368), .A2(n14373), .ZN(n14370) );
  AOI22_X1 U16533 ( .A1(n11913), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U16534 ( .A1(n12109), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13308) );
  NAND2_X1 U16535 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13307) );
  NAND2_X1 U16536 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13306) );
  NAND4_X1 U16537 ( .A1(n13309), .A2(n13308), .A3(n13307), .A4(n13306), .ZN(
        n13313) );
  NAND2_X1 U16538 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13311) );
  NAND2_X1 U16539 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13310) );
  OAI211_X1 U16540 ( .C1(n19886), .C2(n13447), .A(n13311), .B(n13310), .ZN(
        n13312) );
  NOR2_X1 U16541 ( .A1(n13313), .A2(n13312), .ZN(n13322) );
  OAI22_X1 U16542 ( .A1(n13372), .A2(n13413), .B1(n13371), .B2(n13314), .ZN(
        n13318) );
  INV_X1 U16543 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13315) );
  OAI22_X1 U16544 ( .A1(n13375), .A2(n13316), .B1(n13374), .B2(n13315), .ZN(
        n13317) );
  NOR2_X1 U16545 ( .A1(n13318), .A2(n13317), .ZN(n13321) );
  AOI22_X1 U16546 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U16547 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13319) );
  NAND4_X1 U16548 ( .A1(n13322), .A2(n13321), .A3(n13320), .A4(n13319), .ZN(
        n14387) );
  AOI22_X1 U16549 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11914), .B1(
        n11913), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13326) );
  AOI22_X1 U16550 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13305), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13325) );
  NAND2_X1 U16551 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13324) );
  NAND2_X1 U16552 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13323) );
  AND4_X1 U16553 ( .A1(n13326), .A2(n13325), .A3(n13324), .A4(n13323), .ZN(
        n13328) );
  AOI22_X1 U16554 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13444), .B1(
        n13443), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13327) );
  OAI211_X1 U16555 ( .C1(n13466), .C2(n13447), .A(n13328), .B(n13327), .ZN(
        n13334) );
  AOI22_X1 U16556 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13428), .B1(
        n13427), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U16557 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13429), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13331) );
  AOI22_X1 U16558 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n13432), .B1(
        n13431), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13330) );
  NAND2_X1 U16559 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13329) );
  NAND4_X1 U16560 ( .A1(n13332), .A2(n13331), .A3(n13330), .A4(n13329), .ZN(
        n13333) );
  NOR2_X1 U16561 ( .A1(n13334), .A2(n13333), .ZN(n14451) );
  AOI22_X1 U16562 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13428), .B1(
        n13427), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U16563 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13429), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U16564 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n13431), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13336) );
  NAND2_X1 U16565 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13335) );
  NAND4_X1 U16566 ( .A1(n13338), .A2(n13337), .A3(n13336), .A4(n13335), .ZN(
        n13348) );
  AOI22_X1 U16567 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11914), .B1(
        n11913), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U16568 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13305), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13341) );
  NAND2_X1 U16569 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13340) );
  NAND2_X1 U16570 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13339) );
  NAND4_X1 U16571 ( .A1(n13342), .A2(n13341), .A3(n13340), .A4(n13339), .ZN(
        n13346) );
  INV_X1 U16572 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13489) );
  NAND2_X1 U16573 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n13344) );
  NAND2_X1 U16574 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13343) );
  OAI211_X1 U16575 ( .C1(n13447), .C2(n13489), .A(n13344), .B(n13343), .ZN(
        n13345) );
  OR2_X1 U16576 ( .A1(n13346), .A2(n13345), .ZN(n13347) );
  NOR2_X1 U16577 ( .A1(n13348), .A2(n13347), .ZN(n15293) );
  INV_X1 U16578 ( .A(n15293), .ZN(n13349) );
  AOI22_X1 U16579 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11914), .B1(
        n11913), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13353) );
  AOI22_X1 U16580 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13305), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13352) );
  NAND2_X1 U16581 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13351) );
  NAND2_X1 U16582 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13350) );
  AND4_X1 U16583 ( .A1(n13353), .A2(n13352), .A3(n13351), .A4(n13350), .ZN(
        n13355) );
  AOI22_X1 U16584 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n13444), .B1(
        n13443), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13354) );
  OAI211_X1 U16585 ( .C1(n13513), .C2(n13447), .A(n13355), .B(n13354), .ZN(
        n13361) );
  AOI22_X1 U16586 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13428), .B1(
        n13427), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13359) );
  AOI22_X1 U16587 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13429), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13358) );
  AOI22_X1 U16588 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n13432), .B1(
        n13431), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13357) );
  NAND2_X1 U16589 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13356) );
  NAND4_X1 U16590 ( .A1(n13359), .A2(n13358), .A3(n13357), .A4(n13356), .ZN(
        n13360) );
  OR2_X1 U16591 ( .A1(n13361), .A2(n13360), .ZN(n15283) );
  AOI22_X1 U16592 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11914), .B1(
        n11913), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U16593 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13305), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13364) );
  NAND2_X1 U16594 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13363) );
  NAND2_X1 U16595 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13362) );
  NAND4_X1 U16596 ( .A1(n13365), .A2(n13364), .A3(n13363), .A4(n13362), .ZN(
        n13369) );
  NAND2_X1 U16597 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13367) );
  NAND2_X1 U16598 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13366) );
  OAI211_X1 U16599 ( .C1(n13447), .C2(n13536), .A(n13367), .B(n13366), .ZN(
        n13368) );
  NOR2_X1 U16600 ( .A1(n13369), .A2(n13368), .ZN(n13381) );
  INV_X1 U16601 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13373) );
  OAI22_X1 U16602 ( .A1(n13373), .A2(n13372), .B1(n13371), .B2(n13370), .ZN(
        n13377) );
  INV_X1 U16603 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13529) );
  OAI22_X1 U16604 ( .A1(n11990), .A2(n13375), .B1(n13374), .B2(n13529), .ZN(
        n13376) );
  NOR2_X1 U16605 ( .A1(n13377), .A2(n13376), .ZN(n13380) );
  AOI22_X1 U16606 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13432), .B1(
        n13431), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13379) );
  NAND2_X1 U16607 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13378) );
  NAND4_X1 U16608 ( .A1(n13381), .A2(n13380), .A3(n13379), .A4(n13378), .ZN(
        n15276) );
  NAND2_X1 U16609 ( .A1(n15277), .A2(n15276), .ZN(n15267) );
  AOI22_X1 U16610 ( .A1(n11913), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U16611 ( .A1(n12109), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13384) );
  NAND2_X1 U16612 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13383) );
  NAND2_X1 U16613 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13382) );
  AND4_X1 U16614 ( .A1(n13385), .A2(n13384), .A3(n13383), .A4(n13382), .ZN(
        n13387) );
  AOI22_X1 U16615 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13444), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13386) );
  OAI211_X1 U16616 ( .C1(n13447), .C2(n13562), .A(n13387), .B(n13386), .ZN(
        n13393) );
  AOI22_X1 U16617 ( .A1(n13428), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13427), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13391) );
  AOI22_X1 U16618 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13429), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13390) );
  AOI22_X1 U16619 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13389) );
  NAND2_X1 U16620 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13388) );
  NAND4_X1 U16621 ( .A1(n13391), .A2(n13390), .A3(n13389), .A4(n13388), .ZN(
        n13392) );
  NOR2_X1 U16622 ( .A1(n13393), .A2(n13392), .ZN(n15268) );
  NOR2_X2 U16623 ( .A1(n15267), .A2(n15268), .ZN(n15261) );
  AOI22_X1 U16624 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11914), .B1(
        n11913), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13397) );
  AOI22_X1 U16625 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13305), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13396) );
  NAND2_X1 U16626 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n13395) );
  NAND2_X1 U16627 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13394) );
  AND4_X1 U16628 ( .A1(n13397), .A2(n13396), .A3(n13395), .A4(n13394), .ZN(
        n13399) );
  AOI22_X1 U16629 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13444), .B1(
        n13443), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13398) );
  OAI211_X1 U16630 ( .C1(n13579), .C2(n13447), .A(n13399), .B(n13398), .ZN(
        n13405) );
  AOI22_X1 U16631 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13428), .B1(
        n13427), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U16632 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13429), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U16633 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n13432), .B1(
        n13431), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13401) );
  NAND2_X1 U16634 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n13400) );
  NAND4_X1 U16635 ( .A1(n13403), .A2(n13402), .A3(n13401), .A4(n13400), .ZN(
        n13404) );
  NOR2_X1 U16636 ( .A1(n13405), .A2(n13404), .ZN(n15264) );
  INV_X1 U16637 ( .A(n15264), .ZN(n13406) );
  INV_X2 U16638 ( .A(n13407), .ZN(n13608) );
  AOI22_X1 U16639 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U16640 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13606), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U16641 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13416) );
  NAND2_X1 U16642 ( .A1(n13591), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13412) );
  INV_X1 U16643 ( .A(n13409), .ZN(n13411) );
  NAND2_X1 U16644 ( .A1(n16615), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13410) );
  NAND2_X1 U16645 ( .A1(n13411), .A2(n13410), .ZN(n13598) );
  OAI211_X1 U16646 ( .C1(n13602), .C2(n13413), .A(n13412), .B(n13598), .ZN(
        n13414) );
  INV_X1 U16647 ( .A(n13414), .ZN(n13415) );
  NAND4_X1 U16648 ( .A1(n13418), .A2(n13417), .A3(n13416), .A4(n13415), .ZN(
        n13426) );
  AOI22_X1 U16649 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U16650 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13423) );
  AOI22_X1 U16651 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13422) );
  INV_X1 U16652 ( .A(n11704), .ZN(n13597) );
  NAND2_X1 U16653 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13419) );
  INV_X1 U16654 ( .A(n13598), .ZN(n13577) );
  OAI211_X1 U16655 ( .C1(n13597), .C2(n19886), .A(n13419), .B(n13577), .ZN(
        n13420) );
  INV_X1 U16656 ( .A(n13420), .ZN(n13421) );
  NAND4_X1 U16657 ( .A1(n13424), .A2(n13423), .A3(n13422), .A4(n13421), .ZN(
        n13425) );
  NAND2_X1 U16658 ( .A1(n13426), .A2(n13425), .ZN(n13477) );
  NOR2_X1 U16659 ( .A1(n9859), .A2(n13477), .ZN(n13452) );
  AOI22_X1 U16660 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13428), .B1(
        n13427), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13436) );
  AOI22_X1 U16661 ( .A1(n13430), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13429), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U16662 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n13432), .B1(
        n13431), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U16663 ( .A1(n12595), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13433) );
  NAND4_X1 U16664 ( .A1(n13436), .A2(n13435), .A3(n13434), .A4(n13433), .ZN(
        n13451) );
  AOI22_X1 U16665 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11913), .B1(
        n11914), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13442) );
  AOI22_X1 U16666 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13305), .B1(
        n12109), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13441) );
  NAND2_X1 U16667 ( .A1(n13437), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n13440) );
  NAND2_X1 U16668 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13439) );
  NAND4_X1 U16669 ( .A1(n13442), .A2(n13441), .A3(n13440), .A4(n13439), .ZN(
        n13449) );
  NAND2_X1 U16670 ( .A1(n13443), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n13446) );
  NAND2_X1 U16671 ( .A1(n13444), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13445) );
  OAI211_X1 U16672 ( .C1(n13447), .C2(n13596), .A(n13446), .B(n13445), .ZN(
        n13448) );
  OR2_X1 U16673 ( .A1(n13449), .A2(n13448), .ZN(n13450) );
  NOR2_X1 U16674 ( .A1(n13451), .A2(n13450), .ZN(n13455) );
  XNOR2_X1 U16675 ( .A(n13452), .B(n13455), .ZN(n13475) );
  INV_X1 U16676 ( .A(n13477), .ZN(n13456) );
  NAND2_X1 U16677 ( .A1(n11852), .A2(n13456), .ZN(n15253) );
  NAND2_X1 U16678 ( .A1(n13453), .A2(n13475), .ZN(n13454) );
  INV_X1 U16679 ( .A(n13455), .ZN(n13457) );
  AND2_X1 U16680 ( .A1(n13457), .A2(n13456), .ZN(n13474) );
  AOI22_X1 U16681 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13464) );
  AOI22_X1 U16682 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13463) );
  AOI22_X1 U16683 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13462) );
  NAND2_X1 U16684 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13458) );
  OAI211_X1 U16685 ( .C1(n13597), .C2(n13459), .A(n13458), .B(n13598), .ZN(
        n13460) );
  INV_X1 U16686 ( .A(n13460), .ZN(n13461) );
  NAND4_X1 U16687 ( .A1(n13464), .A2(n13463), .A3(n13462), .A4(n13461), .ZN(
        n13473) );
  AOI22_X1 U16688 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U16689 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13470) );
  INV_X1 U16690 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U16691 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U16692 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13465) );
  OAI211_X1 U16693 ( .C1(n13597), .C2(n13466), .A(n13465), .B(n13577), .ZN(
        n13467) );
  INV_X1 U16694 ( .A(n13467), .ZN(n13468) );
  NAND4_X1 U16695 ( .A1(n13471), .A2(n13470), .A3(n13469), .A4(n13468), .ZN(
        n13472) );
  AND2_X1 U16696 ( .A1(n13473), .A2(n13472), .ZN(n13476) );
  NAND2_X1 U16697 ( .A1(n13474), .A2(n13476), .ZN(n13480) );
  OAI211_X1 U16698 ( .C1(n13474), .C2(n13476), .A(n13546), .B(n13480), .ZN(
        n15242) );
  NOR2_X2 U16699 ( .A1(n15240), .A2(n15242), .ZN(n15241) );
  INV_X1 U16700 ( .A(n13475), .ZN(n13478) );
  NAND2_X1 U16701 ( .A1(n11852), .A2(n13476), .ZN(n15245) );
  NOR3_X1 U16702 ( .A1(n13478), .A2(n13477), .A3(n15245), .ZN(n13479) );
  INV_X1 U16703 ( .A(n13480), .ZN(n13497) );
  AOI22_X1 U16704 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U16705 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13486) );
  AOI22_X1 U16706 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13485) );
  INV_X1 U16707 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n19652) );
  NAND2_X1 U16708 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13481) );
  OAI211_X1 U16709 ( .C1(n19652), .C2(n13482), .A(n13481), .B(n13598), .ZN(
        n13483) );
  INV_X1 U16710 ( .A(n13483), .ZN(n13484) );
  NAND4_X1 U16711 ( .A1(n13487), .A2(n13486), .A3(n13485), .A4(n13484), .ZN(
        n13496) );
  AOI22_X1 U16712 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13494) );
  AOI22_X1 U16713 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13606), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13493) );
  AOI22_X1 U16714 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13492) );
  NAND2_X1 U16715 ( .A1(n13591), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13488) );
  OAI211_X1 U16716 ( .C1(n13597), .C2(n13489), .A(n13488), .B(n13577), .ZN(
        n13490) );
  INV_X1 U16717 ( .A(n13490), .ZN(n13491) );
  NAND4_X1 U16718 ( .A1(n13494), .A2(n13493), .A3(n13492), .A4(n13491), .ZN(
        n13495) );
  AND2_X1 U16719 ( .A1(n13496), .A2(n13495), .ZN(n13499) );
  NAND2_X1 U16720 ( .A1(n13497), .A2(n13499), .ZN(n13521) );
  OAI211_X1 U16721 ( .C1(n13497), .C2(n13499), .A(n13546), .B(n13521), .ZN(
        n13502) );
  INV_X1 U16722 ( .A(n13499), .ZN(n13500) );
  NOR2_X1 U16723 ( .A1(n14211), .A2(n13500), .ZN(n15235) );
  INV_X1 U16724 ( .A(n13501), .ZN(n13503) );
  AOI22_X1 U16725 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13511) );
  AOI22_X1 U16726 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13510) );
  AOI22_X1 U16727 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13509) );
  NAND2_X1 U16728 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13505) );
  OAI211_X1 U16729 ( .C1(n13597), .C2(n13506), .A(n13505), .B(n13598), .ZN(
        n13507) );
  INV_X1 U16730 ( .A(n13507), .ZN(n13508) );
  NAND4_X1 U16731 ( .A1(n13511), .A2(n13510), .A3(n13509), .A4(n13508), .ZN(
        n13520) );
  AOI22_X1 U16732 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U16733 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U16734 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13516) );
  NAND2_X1 U16735 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13512) );
  OAI211_X1 U16736 ( .C1(n13597), .C2(n13513), .A(n13512), .B(n13577), .ZN(
        n13514) );
  INV_X1 U16737 ( .A(n13514), .ZN(n13515) );
  NAND4_X1 U16738 ( .A1(n13518), .A2(n13517), .A3(n13516), .A4(n13515), .ZN(
        n13519) );
  NAND2_X1 U16739 ( .A1(n13520), .A2(n13519), .ZN(n13522) );
  AOI21_X1 U16740 ( .B1(n13521), .B2(n13522), .A(n13913), .ZN(n13524) );
  INV_X1 U16741 ( .A(n13521), .ZN(n13523) );
  INV_X1 U16742 ( .A(n13522), .ZN(n13525) );
  NAND2_X1 U16743 ( .A1(n13523), .A2(n13525), .ZN(n13545) );
  NAND2_X1 U16744 ( .A1(n11852), .A2(n13525), .ZN(n15230) );
  NOR2_X2 U16745 ( .A1(n15228), .A2(n15230), .ZN(n15229) );
  NOR2_X2 U16746 ( .A1(n15229), .A2(n13527), .ZN(n13551) );
  INV_X1 U16747 ( .A(n13551), .ZN(n13548) );
  AOI22_X1 U16748 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13534) );
  AOI22_X1 U16749 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13533) );
  AOI22_X1 U16750 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13532) );
  NAND2_X1 U16751 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13528) );
  OAI211_X1 U16752 ( .C1(n13597), .C2(n13529), .A(n13528), .B(n13598), .ZN(
        n13530) );
  INV_X1 U16753 ( .A(n13530), .ZN(n13531) );
  NAND4_X1 U16754 ( .A1(n13534), .A2(n13533), .A3(n13532), .A4(n13531), .ZN(
        n13543) );
  AOI22_X1 U16755 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U16756 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U16757 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U16758 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13535) );
  OAI211_X1 U16759 ( .C1(n13597), .C2(n13536), .A(n13535), .B(n13577), .ZN(
        n13537) );
  INV_X1 U16760 ( .A(n13537), .ZN(n13538) );
  NAND4_X1 U16761 ( .A1(n13541), .A2(n13540), .A3(n13539), .A4(n13538), .ZN(
        n13542) );
  NAND2_X1 U16762 ( .A1(n13543), .A2(n13542), .ZN(n13544) );
  INV_X1 U16763 ( .A(n13544), .ZN(n13553) );
  INV_X1 U16764 ( .A(n13545), .ZN(n13547) );
  OR2_X1 U16765 ( .A1(n13545), .A2(n13544), .ZN(n15214) );
  OAI211_X1 U16766 ( .C1(n13553), .C2(n13547), .A(n15214), .B(n13546), .ZN(
        n13549) );
  NAND2_X2 U16767 ( .A1(n13548), .A2(n13550), .ZN(n15213) );
  INV_X1 U16768 ( .A(n13549), .ZN(n13550) );
  NAND2_X1 U16769 ( .A1(n9859), .A2(n13553), .ZN(n15221) );
  AOI22_X1 U16770 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13560) );
  AOI22_X1 U16771 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13559) );
  AOI22_X1 U16772 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U16773 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13554) );
  OAI211_X1 U16774 ( .C1(n13597), .C2(n13555), .A(n13554), .B(n13598), .ZN(
        n13556) );
  INV_X1 U16775 ( .A(n13556), .ZN(n13557) );
  NAND4_X1 U16776 ( .A1(n13560), .A2(n13559), .A3(n13558), .A4(n13557), .ZN(
        n13569) );
  AOI22_X1 U16777 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U16778 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13566) );
  AOI22_X1 U16779 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13565) );
  NAND2_X1 U16780 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13561) );
  OAI211_X1 U16781 ( .C1(n13597), .C2(n13562), .A(n13561), .B(n13577), .ZN(
        n13563) );
  INV_X1 U16782 ( .A(n13563), .ZN(n13564) );
  NAND4_X1 U16783 ( .A1(n13567), .A2(n13566), .A3(n13565), .A4(n13564), .ZN(
        n13568) );
  AND2_X1 U16784 ( .A1(n13569), .A2(n13568), .ZN(n15215) );
  NAND2_X1 U16785 ( .A1(n14211), .A2(n15215), .ZN(n13570) );
  NOR2_X1 U16786 ( .A1(n15214), .A2(n13570), .ZN(n13588) );
  AOI22_X1 U16787 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13576) );
  AOI22_X1 U16788 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13575) );
  AOI22_X1 U16789 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11704), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13574) );
  INV_X1 U16790 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n19663) );
  NAND2_X1 U16791 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n13571) );
  OAI211_X1 U16792 ( .C1(n19663), .C2(n13482), .A(n13571), .B(n13598), .ZN(
        n13572) );
  INV_X1 U16793 ( .A(n13572), .ZN(n13573) );
  NAND4_X1 U16794 ( .A1(n13576), .A2(n13575), .A3(n13574), .A4(n13573), .ZN(
        n13586) );
  AOI22_X1 U16795 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13584) );
  AOI22_X1 U16796 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13583) );
  AOI22_X1 U16797 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13582) );
  NAND2_X1 U16798 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n13578) );
  OAI211_X1 U16799 ( .C1(n13597), .C2(n13579), .A(n13578), .B(n13577), .ZN(
        n13580) );
  INV_X1 U16800 ( .A(n13580), .ZN(n13581) );
  NAND4_X1 U16801 ( .A1(n13584), .A2(n13583), .A3(n13582), .A4(n13581), .ZN(
        n13585) );
  AND2_X1 U16802 ( .A1(n13586), .A2(n13585), .ZN(n13587) );
  NAND2_X1 U16803 ( .A1(n13588), .A2(n13587), .ZN(n13589) );
  OAI21_X1 U16804 ( .B1(n13588), .B2(n13587), .A(n13589), .ZN(n15210) );
  INV_X1 U16805 ( .A(n13589), .ZN(n13590) );
  AOI22_X1 U16806 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13593) );
  AOI22_X1 U16807 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13592) );
  NAND2_X1 U16808 ( .A1(n13593), .A2(n13592), .ZN(n13615) );
  AOI22_X1 U16809 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11702), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13595) );
  AOI21_X1 U16810 ( .B1(n13606), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n13598), .ZN(n13594) );
  OAI211_X1 U16811 ( .C1(n13597), .C2(n13596), .A(n13595), .B(n13594), .ZN(
        n13614) );
  OAI21_X1 U16812 ( .B1(n13600), .B2(n13599), .A(n13598), .ZN(n13605) );
  INV_X1 U16813 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13603) );
  OAI22_X1 U16814 ( .A1(n13482), .A2(n13603), .B1(n13602), .B2(n13601), .ZN(
        n13604) );
  AOI211_X1 U16815 ( .C1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n11704), .A(
        n13605), .B(n13604), .ZN(n13612) );
  AOI22_X1 U16816 ( .A1(n13607), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13606), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13611) );
  AOI22_X1 U16817 ( .A1(n13609), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13608), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13610) );
  NAND3_X1 U16818 ( .A1(n13612), .A2(n13611), .A3(n13610), .ZN(n13613) );
  OAI21_X1 U16819 ( .B1(n13615), .B2(n13614), .A(n13613), .ZN(n13616) );
  XNOR2_X1 U16820 ( .A(n13617), .B(n13616), .ZN(n14548) );
  AND2_X1 U16821 ( .A1(n12729), .A2(n20108), .ZN(n16630) );
  NAND2_X1 U16822 ( .A1(n12463), .A2(n16630), .ZN(n13618) );
  NOR2_X1 U16823 ( .A1(n16638), .A2(n13618), .ZN(n13619) );
  AOI21_X1 U16824 ( .B1(n16642), .B2(n13620), .A(n13619), .ZN(n15826) );
  NAND4_X1 U16825 ( .A1(n13622), .A2(n13621), .A3(n12735), .A4(n19557), .ZN(
        n13623) );
  NAND2_X1 U16826 ( .A1(n15826), .A2(n13623), .ZN(n13624) );
  INV_X1 U16827 ( .A(n13626), .ZN(n13627) );
  NOR4_X1 U16828 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_14__SCAN_IN), .ZN(n13631) );
  NOR4_X1 U16829 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13630) );
  NOR4_X1 U16830 ( .A1(P2_ADDRESS_REG_9__SCAN_IN), .A2(
        P2_ADDRESS_REG_8__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13629) );
  NOR4_X1 U16831 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P2_ADDRESS_REG_12__SCAN_IN), .A3(P2_ADDRESS_REG_11__SCAN_IN), .A4(
        P2_ADDRESS_REG_10__SCAN_IN), .ZN(n13628) );
  NAND4_X1 U16832 ( .A1(n13631), .A2(n13630), .A3(n13629), .A4(n13628), .ZN(
        n13636) );
  NOR4_X1 U16833 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_5__SCAN_IN), .ZN(n13634) );
  NOR4_X1 U16834 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13633) );
  NOR4_X1 U16835 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13632) );
  INV_X1 U16836 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20136) );
  NAND4_X1 U16837 ( .A1(n13634), .A2(n13633), .A3(n13632), .A4(n20136), .ZN(
        n13635) );
  MUX2_X1 U16838 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n14196), .Z(n19393) );
  INV_X1 U16839 ( .A(n19393), .ZN(n13638) );
  INV_X1 U16840 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13637) );
  OAI22_X1 U16841 ( .A1(n15386), .A2(n13638), .B1(n19415), .B2(n13637), .ZN(
        n13639) );
  AOI21_X1 U16842 ( .B1(n13640), .B2(n19443), .A(n13639), .ZN(n13644) );
  INV_X1 U16843 ( .A(n13641), .ZN(n13642) );
  NAND2_X1 U16844 ( .A1(n19415), .A2(n13642), .ZN(n13991) );
  NOR2_X2 U16845 ( .A1(n13991), .A2(n14196), .ZN(n19385) );
  AOI22_X1 U16846 ( .A1(n19385), .A2(BUF1_REG_30__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n13643) );
  AND2_X1 U16847 ( .A1(n13644), .A2(n13643), .ZN(n13645) );
  OAI21_X1 U16848 ( .B1(n14548), .B2(n19419), .A(n13645), .ZN(P2_U2889) );
  INV_X1 U16849 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20234) );
  NOR2_X1 U16850 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n20234), .ZN(n13647) );
  NOR4_X1 U16851 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_BE_N_REG_3__SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13646) );
  INV_X1 U16852 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n21341) );
  NAND4_X1 U16853 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13647), .A3(n13646), .A4(
        n21341), .ZN(n13650) );
  INV_X1 U16854 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21525) );
  NOR3_X1 U16855 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21525), .ZN(n13649) );
  NOR4_X1 U16856 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13648) );
  NAND4_X1 U16857 ( .A1(n20497), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13649), .A4(
        n13648), .ZN(U214) );
  NOR2_X1 U16858 ( .A1(n13708), .A2(n13650), .ZN(n16716) );
  NAND2_X1 U16859 ( .A1(n16716), .A2(U214), .ZN(U212) );
  NAND2_X1 U16860 ( .A1(n13651), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16516) );
  OAI21_X1 U16861 ( .B1(n13651), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16516), .ZN(n16522) );
  NOR2_X1 U16862 ( .A1(n16522), .A2(n16604), .ZN(n13667) );
  INV_X1 U16863 ( .A(n13652), .ZN(n16509) );
  OR2_X1 U16864 ( .A1(n16509), .A2(n13653), .ZN(n13654) );
  XNOR2_X1 U16865 ( .A(n13655), .B(n13654), .ZN(n16521) );
  NOR2_X1 U16866 ( .A1(n16521), .A2(n16587), .ZN(n13666) );
  NOR2_X1 U16867 ( .A1(n15780), .A2(n15725), .ZN(n13665) );
  NOR2_X1 U16868 ( .A1(n13965), .A2(n13656), .ZN(n13657) );
  NOR2_X1 U16869 ( .A1(n14093), .A2(n13657), .ZN(n16524) );
  INV_X1 U16870 ( .A(n16524), .ZN(n19319) );
  NAND2_X1 U16871 ( .A1(n15781), .A2(n15725), .ZN(n13663) );
  OR2_X1 U16872 ( .A1(n13658), .A2(n14292), .ZN(n13659) );
  NAND2_X1 U16873 ( .A1(n13659), .A2(n16579), .ZN(n19407) );
  INV_X1 U16874 ( .A(n19407), .ZN(n13661) );
  INV_X1 U16875 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20146) );
  NOR2_X1 U16876 ( .A1(n20146), .A2(n19348), .ZN(n13660) );
  AOI21_X1 U16877 ( .B1(n19517), .B2(n13661), .A(n13660), .ZN(n13662) );
  OAI211_X1 U16878 ( .C1(n19534), .C2(n19319), .A(n13663), .B(n13662), .ZN(
        n13664) );
  INV_X1 U16879 ( .A(n16665), .ZN(n20098) );
  OR2_X1 U16880 ( .A1(n12197), .A2(n20098), .ZN(n13782) );
  NOR2_X1 U16881 ( .A1(n16638), .A2(n13782), .ZN(n19381) );
  INV_X1 U16882 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13668) );
  NAND2_X1 U16883 ( .A1(n20206), .A2(n15818), .ZN(n13669) );
  OAI211_X1 U16884 ( .C1(n19381), .C2(n13668), .A(n13680), .B(n13669), .ZN(
        P2_U2814) );
  NOR2_X1 U16885 ( .A1(n19170), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13670)
         );
  INV_X1 U16886 ( .A(n12729), .ZN(n13676) );
  AOI22_X1 U16887 ( .A1(n13670), .A2(n13669), .B1(n13676), .B2(n19170), .ZN(
        P2_U3612) );
  NOR2_X1 U16888 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13671), .ZN(n19485) );
  AOI21_X1 U16889 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n16651), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13672) );
  AOI211_X1 U16890 ( .C1(n19466), .C2(n20108), .A(n13672), .B(n19170), .ZN(
        n13679) );
  INV_X1 U16891 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20120) );
  AOI21_X1 U16892 ( .B1(n15818), .B2(n19913), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n13673) );
  AOI21_X1 U16893 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20108), .A(n13673), 
        .ZN(n13674) );
  NOR2_X1 U16894 ( .A1(n13679), .A2(n13674), .ZN(n13678) );
  OAI21_X1 U16895 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n14211), .A(n20114), 
        .ZN(n13675) );
  NAND3_X1 U16896 ( .A1(n13676), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13675), 
        .ZN(n13677) );
  AOI22_X1 U16897 ( .A1(n13679), .A2(n20120), .B1(n13678), .B2(n13677), .ZN(
        P2_U3610) );
  INV_X1 U16898 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19468) );
  NOR3_X4 U16899 ( .A1(n13680), .A2(n11852), .A3(n20124), .ZN(n13744) );
  MUX2_X1 U16900 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n13708), .Z(n19410) );
  NAND2_X1 U16901 ( .A1(n13744), .A2(n19410), .ZN(n13687) );
  OAI21_X1 U16902 ( .B1(n11852), .B2(n20108), .A(n13681), .ZN(n13710) );
  NAND2_X1 U16903 ( .A1(n13710), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13682) );
  OAI211_X1 U16904 ( .C1(n19468), .C2(n13781), .A(n13687), .B(n13682), .ZN(
        P2_U2975) );
  INV_X1 U16905 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n21305) );
  MUX2_X1 U16906 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n14196), .Z(n19398) );
  NAND2_X1 U16907 ( .A1(n13744), .A2(n19398), .ZN(n13685) );
  NAND2_X1 U16908 ( .A1(n13710), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13683) );
  OAI211_X1 U16909 ( .C1(n21305), .C2(n13781), .A(n13685), .B(n13683), .ZN(
        P2_U2964) );
  INV_X1 U16910 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19459) );
  NAND2_X1 U16911 ( .A1(n13710), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13684) );
  OAI211_X1 U16912 ( .C1(n19459), .C2(n13781), .A(n13685), .B(n13684), .ZN(
        P2_U2979) );
  INV_X1 U16913 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13794) );
  NAND2_X1 U16914 ( .A1(n13710), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13686) );
  OAI211_X1 U16915 ( .C1(n13794), .C2(n13781), .A(n13687), .B(n13686), .ZN(
        P2_U2960) );
  NAND2_X1 U16916 ( .A1(n13744), .A2(n19393), .ZN(n13712) );
  NAND2_X1 U16917 ( .A1(n13710), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13688) );
  OAI211_X1 U16918 ( .C1(n13637), .C2(n13781), .A(n13712), .B(n13688), .ZN(
        P2_U2966) );
  INV_X1 U16919 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19463) );
  MUX2_X1 U16920 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n14196), .Z(n19403) );
  NAND2_X1 U16921 ( .A1(n13744), .A2(n19403), .ZN(n13691) );
  NAND2_X1 U16922 ( .A1(n13710), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13689) );
  OAI211_X1 U16923 ( .C1(n19463), .C2(n13781), .A(n13691), .B(n13689), .ZN(
        P2_U2977) );
  INV_X1 U16924 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13789) );
  NAND2_X1 U16925 ( .A1(n13710), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13690) );
  OAI211_X1 U16926 ( .C1(n13789), .C2(n13781), .A(n13691), .B(n13690), .ZN(
        P2_U2962) );
  INV_X1 U16927 ( .A(n13781), .ZN(n13746) );
  AOI22_X1 U16928 ( .A1(n13746), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13710), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13692) );
  OAI22_X1 U16929 ( .A1(n13708), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14194), .ZN(n19548) );
  INV_X1 U16930 ( .A(n19548), .ZN(n16469) );
  NAND2_X1 U16931 ( .A1(n13744), .A2(n16469), .ZN(n13734) );
  NAND2_X1 U16932 ( .A1(n13692), .A2(n13734), .ZN(P2_U2956) );
  AOI22_X1 U16933 ( .A1(n13746), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13710), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13696) );
  INV_X1 U16934 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14530) );
  OR2_X1 U16935 ( .A1(n13708), .A2(n14530), .ZN(n13694) );
  NAND2_X1 U16936 ( .A1(n14196), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13693) );
  AND2_X1 U16937 ( .A1(n13694), .A2(n13693), .ZN(n19396) );
  INV_X1 U16938 ( .A(n19396), .ZN(n13695) );
  NAND2_X1 U16939 ( .A1(n13744), .A2(n13695), .ZN(n13724) );
  NAND2_X1 U16940 ( .A1(n13696), .A2(n13724), .ZN(P2_U2980) );
  AOI22_X1 U16941 ( .A1(n13746), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13745), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U16942 ( .A1(n14194), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13708), .ZN(n19553) );
  INV_X1 U16943 ( .A(n19553), .ZN(n13697) );
  NAND2_X1 U16944 ( .A1(n13744), .A2(n13697), .ZN(n13732) );
  NAND2_X1 U16945 ( .A1(n13698), .A2(n13732), .ZN(P2_U2957) );
  AOI22_X1 U16946 ( .A1(n13746), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13710), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U16947 ( .A1(n14194), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14196), .ZN(n19451) );
  INV_X1 U16948 ( .A(n19451), .ZN(n13699) );
  NAND2_X1 U16949 ( .A1(n13744), .A2(n13699), .ZN(n13720) );
  NAND2_X1 U16950 ( .A1(n13700), .A2(n13720), .ZN(P2_U2952) );
  AOI22_X1 U16951 ( .A1(n13746), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13745), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U16952 ( .A1(n14194), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13708), .ZN(n19572) );
  INV_X1 U16953 ( .A(n19572), .ZN(n13701) );
  NAND2_X1 U16954 ( .A1(n13744), .A2(n13701), .ZN(n13736) );
  NAND2_X1 U16955 ( .A1(n13702), .A2(n13736), .ZN(P2_U2959) );
  AOI22_X1 U16956 ( .A1(n13746), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13745), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U16957 ( .A1(n14194), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14196), .ZN(n19542) );
  INV_X1 U16958 ( .A(n19542), .ZN(n13703) );
  NAND2_X1 U16959 ( .A1(n13744), .A2(n13703), .ZN(n13730) );
  NAND2_X1 U16960 ( .A1(n13704), .A2(n13730), .ZN(P2_U2955) );
  AOI22_X1 U16961 ( .A1(n13746), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13745), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13706) );
  AOI22_X1 U16962 ( .A1(n14194), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13708), .ZN(n19441) );
  INV_X1 U16963 ( .A(n19441), .ZN(n13705) );
  NAND2_X1 U16964 ( .A1(n13744), .A2(n13705), .ZN(n13722) );
  NAND2_X1 U16965 ( .A1(n13706), .A2(n13722), .ZN(P2_U2953) );
  AOI22_X1 U16966 ( .A1(n13746), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13745), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13707) );
  OAI22_X1 U16967 ( .A1(n13708), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14194), .ZN(n14354) );
  INV_X1 U16968 ( .A(n14354), .ZN(n16476) );
  NAND2_X1 U16969 ( .A1(n13744), .A2(n16476), .ZN(n13713) );
  NAND2_X1 U16970 ( .A1(n13707), .A2(n13713), .ZN(P2_U2954) );
  AOI22_X1 U16971 ( .A1(n13746), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13745), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13709) );
  OAI22_X1 U16972 ( .A1(n13708), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14194), .ZN(n19558) );
  INV_X1 U16973 ( .A(n19558), .ZN(n16462) );
  NAND2_X1 U16974 ( .A1(n13744), .A2(n16462), .ZN(n13738) );
  NAND2_X1 U16975 ( .A1(n13709), .A2(n13738), .ZN(P2_U2958) );
  INV_X1 U16976 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19456) );
  NAND2_X1 U16977 ( .A1(n13745), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13711) );
  OAI211_X1 U16978 ( .C1(n19456), .C2(n13781), .A(n13712), .B(n13711), .ZN(
        P2_U2981) );
  AOI22_X1 U16979 ( .A1(n13746), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13745), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13714) );
  NAND2_X1 U16980 ( .A1(n13714), .A2(n13713), .ZN(P2_U2969) );
  AOI22_X1 U16981 ( .A1(n13746), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13745), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13719) );
  INV_X1 U16982 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13715) );
  OR2_X1 U16983 ( .A1(n14196), .A2(n13715), .ZN(n13717) );
  NAND2_X1 U16984 ( .A1(n14196), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13716) );
  AND2_X1 U16985 ( .A1(n13717), .A2(n13716), .ZN(n19401) );
  INV_X1 U16986 ( .A(n19401), .ZN(n13718) );
  NAND2_X1 U16987 ( .A1(n13744), .A2(n13718), .ZN(n13742) );
  NAND2_X1 U16988 ( .A1(n13719), .A2(n13742), .ZN(P2_U2963) );
  AOI22_X1 U16989 ( .A1(n13746), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n13745), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13721) );
  NAND2_X1 U16990 ( .A1(n13721), .A2(n13720), .ZN(P2_U2967) );
  AOI22_X1 U16991 ( .A1(n13746), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13745), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13723) );
  NAND2_X1 U16992 ( .A1(n13723), .A2(n13722), .ZN(P2_U2968) );
  AOI22_X1 U16993 ( .A1(n13746), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13745), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13725) );
  NAND2_X1 U16994 ( .A1(n13725), .A2(n13724), .ZN(P2_U2965) );
  AOI22_X1 U16995 ( .A1(n13746), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13745), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13729) );
  INV_X1 U16996 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14448) );
  OR2_X1 U16997 ( .A1(n14196), .A2(n14448), .ZN(n13727) );
  NAND2_X1 U16998 ( .A1(n14196), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13726) );
  AND2_X1 U16999 ( .A1(n13727), .A2(n13726), .ZN(n19406) );
  INV_X1 U17000 ( .A(n19406), .ZN(n13728) );
  NAND2_X1 U17001 ( .A1(n13744), .A2(n13728), .ZN(n13740) );
  NAND2_X1 U17002 ( .A1(n13729), .A2(n13740), .ZN(P2_U2961) );
  AOI22_X1 U17003 ( .A1(n13746), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13745), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13731) );
  NAND2_X1 U17004 ( .A1(n13731), .A2(n13730), .ZN(P2_U2970) );
  AOI22_X1 U17005 ( .A1(n13746), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13745), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U17006 ( .A1(n13733), .A2(n13732), .ZN(P2_U2972) );
  AOI22_X1 U17007 ( .A1(n13746), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13745), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13735) );
  NAND2_X1 U17008 ( .A1(n13735), .A2(n13734), .ZN(P2_U2971) );
  AOI22_X1 U17009 ( .A1(n13746), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13745), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13737) );
  NAND2_X1 U17010 ( .A1(n13737), .A2(n13736), .ZN(P2_U2974) );
  AOI22_X1 U17011 ( .A1(n13746), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13745), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13739) );
  NAND2_X1 U17012 ( .A1(n13739), .A2(n13738), .ZN(P2_U2973) );
  AOI22_X1 U17013 ( .A1(n13746), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13745), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13741) );
  NAND2_X1 U17014 ( .A1(n13741), .A2(n13740), .ZN(P2_U2976) );
  AOI22_X1 U17015 ( .A1(n13746), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13745), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13743) );
  NAND2_X1 U17016 ( .A1(n13743), .A2(n13742), .ZN(P2_U2978) );
  INV_X1 U17017 ( .A(n13744), .ZN(n13748) );
  AOI22_X1 U17018 ( .A1(n14194), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14196), .ZN(n19390) );
  AOI22_X1 U17019 ( .A1(n13746), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13745), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n13747) );
  OAI21_X1 U17020 ( .B1(n13748), .B2(n19390), .A(n13747), .ZN(P2_U2982) );
  INV_X1 U17021 ( .A(n16642), .ZN(n13752) );
  NAND2_X1 U17022 ( .A1(n13752), .A2(n16639), .ZN(n15824) );
  NAND2_X1 U17023 ( .A1(n15824), .A2(n12744), .ZN(n13753) );
  INV_X1 U17024 ( .A(n13754), .ZN(n13920) );
  MUX2_X1 U17025 ( .A(n15193), .B(n15197), .S(n13920), .Z(n13755) );
  OAI21_X1 U17026 ( .B1(n19676), .B2(n15289), .A(n13755), .ZN(P2_U2886) );
  INV_X1 U17027 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19541) );
  NAND2_X1 U17028 ( .A1(n14211), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13756) );
  AND4_X1 U17029 ( .A1(n13757), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13756), 
        .A4(n19873), .ZN(n13758) );
  NOR2_X1 U17030 ( .A1(n15273), .A2(n13805), .ZN(n13759) );
  AOI21_X1 U17031 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n15273), .A(n13759), .ZN(
        n13760) );
  OAI21_X1 U17032 ( .B1(n15289), .B2(n20228), .A(n13760), .ZN(P2_U2887) );
  OAI21_X1 U17033 ( .B1(n19366), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13824), .ZN(n13761) );
  INV_X1 U17034 ( .A(n13761), .ZN(n13811) );
  OAI21_X1 U17035 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13763), .A(
        n13762), .ZN(n13808) );
  NAND2_X1 U17036 ( .A1(n19247), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13804) );
  OAI21_X1 U17037 ( .B1(n16543), .B2(n13808), .A(n13804), .ZN(n13764) );
  AOI21_X1 U17038 ( .B1(n19493), .B2(n13811), .A(n13764), .ZN(n13767) );
  OAI21_X1 U17039 ( .B1(n19488), .B2(n13765), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13766) );
  OAI211_X1 U17040 ( .C1(n14195), .C2(n13805), .A(n13767), .B(n13766), .ZN(
        P2_U3014) );
  NOR3_X1 U17041 ( .A1(n14306), .A2(n10210), .A3(n21230), .ZN(n21229) );
  NAND2_X1 U17042 ( .A1(n11420), .A2(n13777), .ZN(n13815) );
  AOI22_X1 U17043 ( .A1(n13815), .A2(n11551), .B1(n16010), .B2(n13768), .ZN(
        n20250) );
  OAI21_X1 U17044 ( .B1(n21229), .B2(n21132), .A(n20250), .ZN(n16028) );
  AND2_X1 U17045 ( .A1(n16028), .A2(n13876), .ZN(n20259) );
  INV_X1 U17046 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13780) );
  INV_X1 U17047 ( .A(n11420), .ZN(n13776) );
  INV_X1 U17048 ( .A(n16010), .ZN(n13769) );
  NAND2_X1 U17049 ( .A1(n13848), .A2(n13769), .ZN(n13775) );
  NAND4_X1 U17050 ( .A1(n13771), .A2(n10542), .A3(n13770), .A4(n20501), .ZN(
        n13772) );
  NAND2_X1 U17051 ( .A1(n13837), .A2(n13772), .ZN(n13773) );
  OAI21_X1 U17052 ( .B1(n16032), .B2(n13773), .A(n16010), .ZN(n13774) );
  OAI211_X1 U17053 ( .C1(n13777), .C2(n13776), .A(n13775), .B(n13774), .ZN(
        n13778) );
  AND2_X1 U17054 ( .A1(n13778), .A2(n20550), .ZN(n16030) );
  NAND2_X1 U17055 ( .A1(n20259), .A2(n16030), .ZN(n13779) );
  OAI21_X1 U17056 ( .B1(n20259), .B2(n13780), .A(n13779), .ZN(P1_U3484) );
  INV_X1 U17057 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15330) );
  OAI21_X1 U17058 ( .B1(n13783), .B2(n13782), .A(n13781), .ZN(n13784) );
  AND2_X1 U17059 ( .A1(n13784), .A2(n20114), .ZN(n19452) );
  NAND2_X1 U17060 ( .A1(n19452), .A2(n13785), .ZN(n13933) );
  AOI22_X1 U17061 ( .A1(n19466), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13786) );
  OAI21_X1 U17062 ( .B1(n15330), .B2(n13933), .A(n13786), .ZN(P2_U2926) );
  AOI22_X1 U17063 ( .A1(n19466), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13787) );
  OAI21_X1 U17064 ( .B1(n21305), .B2(n13933), .A(n13787), .ZN(P2_U2923) );
  AOI22_X1 U17065 ( .A1(n19466), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13788) );
  OAI21_X1 U17066 ( .B1(n13789), .B2(n13933), .A(n13788), .ZN(P2_U2925) );
  INV_X1 U17067 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15314) );
  AOI22_X1 U17068 ( .A1(n19466), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13790) );
  OAI21_X1 U17069 ( .B1(n15314), .B2(n13933), .A(n13790), .ZN(P2_U2924) );
  AOI22_X1 U17070 ( .A1(n19466), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13791) );
  OAI21_X1 U17071 ( .B1(n13637), .B2(n13933), .A(n13791), .ZN(P2_U2921) );
  INV_X1 U17072 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U17073 ( .A1(n19466), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13792) );
  OAI21_X1 U17074 ( .B1(n15304), .B2(n13933), .A(n13792), .ZN(P2_U2922) );
  AOI22_X1 U17075 ( .A1(n19466), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13793) );
  OAI21_X1 U17076 ( .B1(n13794), .B2(n13933), .A(n13793), .ZN(P2_U2927) );
  AOI21_X1 U17077 ( .B1(n13797), .B2(n13796), .A(n13795), .ZN(n19521) );
  AOI22_X1 U17078 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19247), .ZN(n13798) );
  OAI21_X1 U17079 ( .B1(n19499), .B2(n14331), .A(n13798), .ZN(n13799) );
  AOI21_X1 U17080 ( .B1(n19521), .B2(n19495), .A(n13799), .ZN(n13803) );
  NAND2_X1 U17081 ( .A1(n13801), .A2(n13800), .ZN(n19524) );
  NAND3_X1 U17082 ( .A1(n19525), .A2(n19493), .A3(n19524), .ZN(n13802) );
  OAI211_X1 U17083 ( .C1(n19533), .C2(n14195), .A(n13803), .B(n13802), .ZN(
        P2_U3012) );
  OAI21_X1 U17084 ( .B1(n19534), .B2(n13805), .A(n13804), .ZN(n13810) );
  XNOR2_X1 U17085 ( .A(n13807), .B(n13806), .ZN(n19370) );
  OAI22_X1 U17086 ( .A1(n16604), .A2(n13808), .B1(n16603), .B2(n19370), .ZN(
        n13809) );
  AOI211_X1 U17087 ( .C1(n19526), .C2(n13811), .A(n13810), .B(n13809), .ZN(
        n13813) );
  MUX2_X1 U17088 ( .A(n15726), .B(n19513), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13812) );
  NAND2_X1 U17089 ( .A1(n13813), .A2(n13812), .ZN(P2_U3046) );
  NAND2_X1 U17090 ( .A1(n21206), .A2(n16040), .ZN(n20254) );
  INV_X1 U17091 ( .A(n20254), .ZN(n13814) );
  NOR2_X1 U17092 ( .A1(n13814), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13818)
         );
  INV_X1 U17093 ( .A(n11551), .ZN(n13816) );
  OAI21_X1 U17094 ( .B1(n14306), .B2(n11476), .A(n21225), .ZN(n13817) );
  OAI21_X1 U17095 ( .B1(n13818), .B2(n21225), .A(n13817), .ZN(P1_U3487) );
  AOI21_X1 U17096 ( .B1(n15833), .B2(n13820), .A(n13819), .ZN(n15808) );
  NAND2_X1 U17097 ( .A1(n19495), .A2(n15808), .ZN(n13821) );
  NAND2_X1 U17098 ( .A1(n19247), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15805) );
  OAI211_X1 U17099 ( .C1(n16561), .C2(n15192), .A(n13821), .B(n15805), .ZN(
        n13822) );
  AOI21_X1 U17100 ( .B1(n16550), .B2(n15192), .A(n13822), .ZN(n13827) );
  OAI21_X1 U17101 ( .B1(n15191), .B2(n13824), .A(n13823), .ZN(n13825) );
  XOR2_X1 U17102 ( .A(n13825), .B(n15833), .Z(n15804) );
  NAND2_X1 U17103 ( .A1(n15804), .A2(n19493), .ZN(n13826) );
  OAI211_X1 U17104 ( .C1(n15197), .C2(n14195), .A(n13827), .B(n13826), .ZN(
        P2_U3013) );
  INV_X1 U17105 ( .A(n13829), .ZN(n13830) );
  INV_X1 U17106 ( .A(n19677), .ZN(n20212) );
  MUX2_X1 U17107 ( .A(n19533), .B(n11792), .S(n15273), .Z(n13831) );
  OAI21_X1 U17108 ( .B1(n20212), .B2(n15289), .A(n13831), .ZN(P2_U2885) );
  INV_X1 U17109 ( .A(n14066), .ZN(n16366) );
  NAND3_X1 U17110 ( .A1(n13852), .A2(n13834), .A3(n13833), .ZN(n13835) );
  OR3_X1 U17111 ( .A1(n13836), .A2(n16366), .A3(n13835), .ZN(n15128) );
  INV_X1 U17112 ( .A(n15128), .ZN(n13844) );
  INV_X1 U17113 ( .A(n13837), .ZN(n13838) );
  OR2_X1 U17114 ( .A1(n13848), .A2(n13838), .ZN(n14048) );
  XNOR2_X1 U17115 ( .A(n13839), .B(n10394), .ZN(n13845) );
  INV_X1 U17116 ( .A(n13845), .ZN(n13841) );
  INV_X1 U17117 ( .A(n16012), .ZN(n13867) );
  XNOR2_X1 U17118 ( .A(n10394), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13840) );
  AOI22_X1 U17119 ( .A1(n14048), .A2(n13841), .B1(n13867), .B2(n13840), .ZN(
        n13843) );
  NAND3_X1 U17120 ( .A1(n13844), .A2(n14043), .A3(n13845), .ZN(n13842) );
  OAI211_X1 U17121 ( .C1(n13832), .C2(n13844), .A(n13843), .B(n13842), .ZN(
        n14060) );
  NOR2_X1 U17122 ( .A1(n16040), .A2(n20473), .ZN(n15131) );
  OAI22_X1 U17123 ( .A1(n11418), .A2(n14133), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15132) );
  INV_X1 U17124 ( .A(n15132), .ZN(n13846) );
  AOI222_X1 U17125 ( .A1(n14060), .A2(n21189), .B1(n15131), .B2(n13846), .C1(
        n13845), .C2(n21188), .ZN(n13864) );
  INV_X1 U17126 ( .A(n13847), .ZN(n13851) );
  NAND2_X1 U17127 ( .A1(n13848), .A2(n16010), .ZN(n13875) );
  OR2_X1 U17128 ( .A1(n14319), .A2(n20523), .ZN(n13849) );
  AND4_X1 U17129 ( .A1(n13851), .A2(n13875), .A3(n13850), .A4(n13849), .ZN(
        n13858) );
  NAND2_X1 U17130 ( .A1(n16012), .A2(n13852), .ZN(n13855) );
  NOR2_X1 U17131 ( .A1(n16066), .A2(n21132), .ZN(n13854) );
  AOI21_X1 U17132 ( .B1(n13855), .B2(n13854), .A(n13853), .ZN(n13856) );
  OR2_X1 U17133 ( .A1(n13856), .A2(n16010), .ZN(n13857) );
  NAND2_X1 U17134 ( .A1(n16014), .A2(n13876), .ZN(n13861) );
  NAND2_X1 U17135 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16372) );
  INV_X1 U17136 ( .A(n16372), .ZN(n16043) );
  NAND2_X1 U17137 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16043), .ZN(n16376) );
  INV_X1 U17138 ( .A(n16376), .ZN(n13859) );
  NAND2_X1 U17139 ( .A1(n13859), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13860) );
  NAND2_X1 U17140 ( .A1(n13861), .A2(n13860), .ZN(n16365) );
  AND2_X1 U17141 ( .A1(n20500), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13862) );
  OR2_X1 U17142 ( .A1(n16365), .A2(n13862), .ZN(n21192) );
  NAND2_X1 U17143 ( .A1(n13869), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13863) );
  OAI21_X1 U17144 ( .B1(n13864), .B2(n13869), .A(n13863), .ZN(P1_U3472) );
  AOI22_X1 U17145 ( .A1(n21209), .A2(n15128), .B1(n15125), .B2(n10273), .ZN(
        n16011) );
  INV_X1 U17146 ( .A(n16011), .ZN(n13866) );
  OAI22_X1 U17147 ( .A1(n16040), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15129), .ZN(n13865) );
  AOI21_X1 U17148 ( .B1(n13866), .B2(n21189), .A(n13865), .ZN(n13870) );
  AOI21_X1 U17149 ( .B1(n13867), .B2(n21189), .A(n13869), .ZN(n13868) );
  OAI22_X1 U17150 ( .A1(n13870), .A2(n13869), .B1(n13868), .B2(n10273), .ZN(
        P1_U3474) );
  OAI21_X1 U17151 ( .B1(n13872), .B2(n13871), .A(n14021), .ZN(n14536) );
  OR2_X1 U17152 ( .A1(n13873), .A2(n11545), .ZN(n13874) );
  NAND2_X1 U17153 ( .A1(n13875), .A2(n13874), .ZN(n13877) );
  OR2_X1 U17154 ( .A1(n14538), .A2(n10210), .ZN(n13879) );
  AND2_X1 U17155 ( .A1(n13880), .A2(n13879), .ZN(n20478) );
  INV_X1 U17156 ( .A(n20478), .ZN(n13881) );
  AOI22_X1 U17157 ( .A1(n14721), .A2(n13881), .B1(n14720), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13882) );
  OAI21_X1 U17158 ( .B1(n14536), .B2(n14772), .A(n13882), .ZN(P1_U2871) );
  XOR2_X1 U17159 ( .A(n13884), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13889)
         );
  NAND2_X1 U17160 ( .A1(n13885), .A2(n13918), .ZN(n13887) );
  INV_X1 U17161 ( .A(n13903), .ZN(n13886) );
  INV_X1 U17162 ( .A(n19360), .ZN(n14409) );
  MUX2_X1 U17163 ( .A(n14409), .B(n19352), .S(n15273), .Z(n13888) );
  OAI21_X1 U17164 ( .B1(n13889), .B2(n15289), .A(n13888), .ZN(P2_U2882) );
  INV_X1 U17165 ( .A(n13890), .ZN(n13894) );
  NAND2_X1 U17166 ( .A1(n13892), .A2(n13893), .ZN(n13911) );
  NAND2_X1 U17167 ( .A1(n13891), .A2(n13911), .ZN(n13895) );
  NAND2_X1 U17168 ( .A1(n13894), .A2(n13895), .ZN(n13897) );
  INV_X1 U17169 ( .A(n13895), .ZN(n13896) );
  INV_X1 U17170 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n15182) );
  NOR2_X1 U17171 ( .A1(n13920), .A2(n15182), .ZN(n13898) );
  AOI21_X1 U17172 ( .B1(n16601), .B2(n13920), .A(n13898), .ZN(n13899) );
  OAI21_X1 U17173 ( .B1(n20202), .B2(n15289), .A(n13899), .ZN(P2_U2884) );
  NOR2_X1 U17174 ( .A1(n13884), .A2(n13900), .ZN(n13902) );
  OAI211_X1 U17175 ( .C1(n13902), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15294), .B(n13901), .ZN(n13908) );
  OR2_X1 U17176 ( .A1(n13904), .A2(n13903), .ZN(n13905) );
  NAND2_X1 U17177 ( .A1(n13905), .A2(n13935), .ZN(n19342) );
  INV_X1 U17178 ( .A(n19342), .ZN(n13906) );
  NAND2_X1 U17179 ( .A1(n13920), .A2(n13906), .ZN(n13907) );
  OAI211_X1 U17180 ( .C1(n13920), .C2(n12388), .A(n13908), .B(n13907), .ZN(
        P2_U2881) );
  INV_X1 U17181 ( .A(n13909), .ZN(n13915) );
  INV_X1 U17182 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13912) );
  NAND2_X1 U17183 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19557), .ZN(
        n13910) );
  OAI211_X1 U17184 ( .C1(n13913), .C2(n13912), .A(n13911), .B(n13910), .ZN(
        n13914) );
  OAI21_X1 U17185 ( .B1(n13915), .B2(n13914), .A(n13884), .ZN(n19425) );
  OR2_X1 U17186 ( .A1(n13917), .A2(n13916), .ZN(n13919) );
  AND2_X1 U17187 ( .A1(n13919), .A2(n13918), .ZN(n19501) );
  NOR2_X1 U17188 ( .A1(n13920), .A2(n12382), .ZN(n13921) );
  AOI21_X1 U17189 ( .B1(n19501), .B2(n13920), .A(n13921), .ZN(n13922) );
  OAI21_X1 U17190 ( .B1(n19425), .B2(n15289), .A(n13922), .ZN(P2_U2883) );
  INV_X1 U17191 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n15385) );
  AOI22_X1 U17192 ( .A1(n19485), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13923) );
  OAI21_X1 U17193 ( .B1(n15385), .B2(n13933), .A(n13923), .ZN(P2_U2935) );
  INV_X1 U17194 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U17195 ( .A1(n19466), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13924) );
  OAI21_X1 U17196 ( .B1(n13925), .B2(n13933), .A(n13924), .ZN(P2_U2931) );
  INV_X1 U17197 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U17198 ( .A1(n19466), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13926) );
  OAI21_X1 U17199 ( .B1(n13927), .B2(n13933), .A(n13926), .ZN(P2_U2929) );
  INV_X1 U17200 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n21469) );
  AOI22_X1 U17201 ( .A1(n19466), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13928) );
  OAI21_X1 U17202 ( .B1(n21469), .B2(n13933), .A(n13928), .ZN(P2_U2934) );
  INV_X1 U17203 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15356) );
  AOI22_X1 U17204 ( .A1(n19466), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13929) );
  OAI21_X1 U17205 ( .B1(n15356), .B2(n13933), .A(n13929), .ZN(P2_U2930) );
  INV_X1 U17206 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n21317) );
  AOI22_X1 U17207 ( .A1(n19466), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13930) );
  OAI21_X1 U17208 ( .B1(n21317), .B2(n13933), .A(n13930), .ZN(P2_U2932) );
  INV_X1 U17209 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15346) );
  AOI22_X1 U17210 ( .A1(n19466), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13931) );
  OAI21_X1 U17211 ( .B1(n15346), .B2(n13933), .A(n13931), .ZN(P2_U2928) );
  INV_X1 U17212 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13934) );
  AOI22_X1 U17213 ( .A1(n19466), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13932) );
  OAI21_X1 U17214 ( .B1(n13934), .B2(n13933), .A(n13932), .ZN(P2_U2933) );
  XOR2_X1 U17215 ( .A(n13901), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13938)
         );
  AOI21_X1 U17216 ( .B1(n13936), .B2(n13935), .A(n13964), .ZN(n15796) );
  INV_X1 U17217 ( .A(n15796), .ZN(n19330) );
  MUX2_X1 U17218 ( .A(n19330), .B(n12392), .S(n15273), .Z(n13937) );
  OAI21_X1 U17219 ( .B1(n13938), .B2(n15289), .A(n13937), .ZN(P2_U2880) );
  INV_X1 U17220 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13943) );
  NOR2_X1 U17221 ( .A1(n13939), .A2(n16066), .ZN(n16038) );
  INV_X1 U17222 ( .A(n16038), .ZN(n13940) );
  OAI21_X1 U17223 ( .B1(n16012), .B2(n16066), .A(n13940), .ZN(n13941) );
  OR2_X1 U17224 ( .A1(n16372), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20380) );
  INV_X2 U17225 ( .A(n20380), .ZN(n20387) );
  AOI22_X1 U17226 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13942) );
  OAI21_X1 U17227 ( .B1(n13943), .B2(n20365), .A(n13942), .ZN(P1_U2912) );
  AOI22_X1 U17228 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13944) );
  OAI21_X1 U17229 ( .B1(n14789), .B2(n20365), .A(n13944), .ZN(P1_U2910) );
  AOI22_X1 U17230 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13945) );
  OAI21_X1 U17231 ( .B1(n14823), .B2(n20365), .A(n13945), .ZN(P1_U2918) );
  INV_X1 U17232 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13947) );
  AOI22_X1 U17233 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13946) );
  OAI21_X1 U17234 ( .B1(n13947), .B2(n20365), .A(n13946), .ZN(P1_U2911) );
  INV_X1 U17235 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13949) );
  AOI22_X1 U17236 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13948) );
  OAI21_X1 U17237 ( .B1(n13949), .B2(n20365), .A(n13948), .ZN(P1_U2920) );
  INV_X1 U17238 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U17239 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13950) );
  OAI21_X1 U17240 ( .B1(n13951), .B2(n20365), .A(n13950), .ZN(P1_U2919) );
  INV_X1 U17241 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U17242 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13952) );
  OAI21_X1 U17243 ( .B1(n13953), .B2(n20365), .A(n13952), .ZN(P1_U2908) );
  INV_X1 U17244 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U17245 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13954) );
  OAI21_X1 U17246 ( .B1(n13955), .B2(n20365), .A(n13954), .ZN(P1_U2913) );
  INV_X1 U17247 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U17248 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13956) );
  OAI21_X1 U17249 ( .B1(n13957), .B2(n20365), .A(n13956), .ZN(P1_U2917) );
  INV_X1 U17250 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14816) );
  AOI22_X1 U17251 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13958) );
  OAI21_X1 U17252 ( .B1(n14816), .B2(n20365), .A(n13958), .ZN(P1_U2916) );
  INV_X1 U17253 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21493) );
  AOI22_X1 U17254 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13959) );
  OAI21_X1 U17255 ( .B1(n21493), .B2(n20365), .A(n13959), .ZN(P1_U2915) );
  INV_X1 U17256 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U17257 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13960) );
  OAI21_X1 U17258 ( .B1(n13961), .B2(n20365), .A(n13960), .ZN(P1_U2914) );
  INV_X1 U17259 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13963) );
  AOI22_X1 U17260 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13962) );
  OAI21_X1 U17261 ( .B1(n13963), .B2(n20365), .A(n13962), .ZN(P1_U2909) );
  AOI21_X1 U17262 ( .B1(n9982), .B2(n10335), .A(n13965), .ZN(n16537) );
  INV_X1 U17263 ( .A(n16537), .ZN(n16591) );
  OAI211_X1 U17264 ( .C1(n13967), .C2(n13970), .A(n13969), .B(n15294), .ZN(
        n13972) );
  NAND2_X1 U17265 ( .A1(n13754), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13971) );
  OAI211_X1 U17266 ( .C1(n16591), .C2(n13754), .A(n13972), .B(n13971), .ZN(
        P2_U2879) );
  AND2_X1 U17267 ( .A1(n21231), .A2(n21132), .ZN(n13973) );
  OR2_X1 U17268 ( .A1(n20397), .A2(n20517), .ZN(n14097) );
  INV_X1 U17269 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13979) );
  NOR2_X2 U17270 ( .A1(n20397), .A2(n13974), .ZN(n20411) );
  INV_X1 U17271 ( .A(n20411), .ZN(n13978) );
  INV_X1 U17272 ( .A(n20497), .ZN(n20495) );
  INV_X1 U17273 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13975) );
  NOR2_X1 U17274 ( .A1(n20495), .A2(n13975), .ZN(n13976) );
  AOI21_X1 U17275 ( .B1(DATAI_15_), .B2(n20495), .A(n13976), .ZN(n14837) );
  INV_X1 U17276 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13977) );
  OAI222_X1 U17277 ( .A1(n14097), .A2(n13979), .B1(n13978), .B2(n14837), .C1(
        n13977), .C2(n14015), .ZN(P1_U2967) );
  NAND2_X1 U17278 ( .A1(n13981), .A2(n13980), .ZN(n13983) );
  NAND2_X1 U17279 ( .A1(n13983), .A2(n10288), .ZN(n20214) );
  INV_X1 U17280 ( .A(n20214), .ZN(n13994) );
  INV_X1 U17281 ( .A(n19443), .ZN(n15324) );
  XNOR2_X1 U17282 ( .A(n20212), .B(n20214), .ZN(n13989) );
  XNOR2_X1 U17283 ( .A(n13985), .B(n13984), .ZN(n20223) );
  NOR2_X1 U17284 ( .A1(n20221), .A2(n20223), .ZN(n13986) );
  AOI21_X1 U17285 ( .B1(n20223), .B2(n20221), .A(n13986), .ZN(n19437) );
  INV_X1 U17286 ( .A(n19370), .ZN(n19446) );
  NAND2_X1 U17287 ( .A1(n19447), .A2(n19446), .ZN(n19445) );
  NAND2_X1 U17288 ( .A1(n19437), .A2(n19445), .ZN(n19436) );
  INV_X1 U17289 ( .A(n13986), .ZN(n13987) );
  NAND2_X1 U17290 ( .A1(n19436), .A2(n13987), .ZN(n13988) );
  NAND2_X1 U17291 ( .A1(n13988), .A2(n13989), .ZN(n19417) );
  OAI21_X1 U17292 ( .B1(n13989), .B2(n13988), .A(n19417), .ZN(n13990) );
  NAND2_X1 U17293 ( .A1(n13990), .A2(n19444), .ZN(n13993) );
  NAND2_X1 U17294 ( .A1(n15386), .A2(n13991), .ZN(n19409) );
  AOI22_X1 U17295 ( .A1(n19409), .A2(n16476), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19442), .ZN(n13992) );
  OAI211_X1 U17296 ( .C1(n13994), .C2(n15324), .A(n13993), .B(n13992), .ZN(
        P2_U2917) );
  INV_X1 U17297 ( .A(n14097), .ZN(n20393) );
  AOI22_X1 U17298 ( .A1(n20393), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20425), .ZN(n13998) );
  NAND2_X1 U17299 ( .A1(n20495), .A2(DATAI_5_), .ZN(n13996) );
  NAND2_X1 U17300 ( .A1(n20497), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13995) );
  AND2_X1 U17301 ( .A1(n13996), .A2(n13995), .ZN(n20542) );
  INV_X1 U17302 ( .A(n20542), .ZN(n13997) );
  NAND2_X1 U17303 ( .A1(n20411), .A2(n13997), .ZN(n14110) );
  NAND2_X1 U17304 ( .A1(n13998), .A2(n14110), .ZN(P1_U2957) );
  AOI22_X1 U17305 ( .A1(n20393), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20425), .ZN(n14002) );
  NAND2_X1 U17306 ( .A1(n20495), .A2(DATAI_3_), .ZN(n14000) );
  NAND2_X1 U17307 ( .A1(n20497), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13999) );
  AND2_X1 U17308 ( .A1(n14000), .A2(n13999), .ZN(n20531) );
  INV_X1 U17309 ( .A(n20531), .ZN(n14001) );
  NAND2_X1 U17310 ( .A1(n20411), .A2(n14001), .ZN(n14114) );
  NAND2_X1 U17311 ( .A1(n14002), .A2(n14114), .ZN(P1_U2955) );
  AOI22_X1 U17312 ( .A1(n20393), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20425), .ZN(n14006) );
  NAND2_X1 U17313 ( .A1(n20495), .A2(DATAI_4_), .ZN(n14004) );
  NAND2_X1 U17314 ( .A1(n20497), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14003) );
  AND2_X1 U17315 ( .A1(n14004), .A2(n14003), .ZN(n20537) );
  INV_X1 U17316 ( .A(n20537), .ZN(n14005) );
  NAND2_X1 U17317 ( .A1(n20411), .A2(n14005), .ZN(n14108) );
  NAND2_X1 U17318 ( .A1(n14006), .A2(n14108), .ZN(P1_U2956) );
  AOI22_X1 U17319 ( .A1(n20393), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20425), .ZN(n14010) );
  NAND2_X1 U17320 ( .A1(n20495), .A2(DATAI_6_), .ZN(n14008) );
  NAND2_X1 U17321 ( .A1(n20497), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14007) );
  AND2_X1 U17322 ( .A1(n14008), .A2(n14007), .ZN(n20547) );
  INV_X1 U17323 ( .A(n20547), .ZN(n14009) );
  NAND2_X1 U17324 ( .A1(n20411), .A2(n14009), .ZN(n14118) );
  NAND2_X1 U17325 ( .A1(n14010), .A2(n14118), .ZN(P1_U2958) );
  AOI22_X1 U17326 ( .A1(n20393), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20425), .ZN(n14014) );
  NAND2_X1 U17327 ( .A1(n20495), .A2(DATAI_2_), .ZN(n14012) );
  NAND2_X1 U17328 ( .A1(n20497), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14011) );
  AND2_X1 U17329 ( .A1(n14012), .A2(n14011), .ZN(n20526) );
  INV_X1 U17330 ( .A(n20526), .ZN(n14013) );
  NAND2_X1 U17331 ( .A1(n20411), .A2(n14013), .ZN(n14102) );
  NAND2_X1 U17332 ( .A1(n14014), .A2(n14102), .ZN(P1_U2954) );
  INV_X1 U17333 ( .A(n14015), .ZN(n20425) );
  AOI22_X1 U17334 ( .A1(n20393), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20425), .ZN(n14018) );
  INV_X1 U17335 ( .A(DATAI_7_), .ZN(n14017) );
  NAND2_X1 U17336 ( .A1(n20497), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14016) );
  OAI21_X1 U17337 ( .B1(n20497), .B2(n14017), .A(n14016), .ZN(n14802) );
  NAND2_X1 U17338 ( .A1(n20411), .A2(n14802), .ZN(n14104) );
  NAND2_X1 U17339 ( .A1(n14018), .A2(n14104), .ZN(P1_U2959) );
  INV_X1 U17340 ( .A(n14019), .ZN(n14020) );
  AOI21_X1 U17341 ( .B1(n14022), .B2(n14021), .A(n14020), .ZN(n14130) );
  INV_X1 U17342 ( .A(n14130), .ZN(n14708) );
  NAND2_X1 U17343 ( .A1(n14024), .A2(n14023), .ZN(n14025) );
  NAND2_X1 U17344 ( .A1(n14086), .A2(n14025), .ZN(n20465) );
  INV_X1 U17345 ( .A(n20465), .ZN(n14026) );
  AOI22_X1 U17346 ( .A1(n14721), .A2(n14026), .B1(n14720), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14027) );
  OAI21_X1 U17347 ( .B1(n14708), .B2(n14772), .A(n14027), .ZN(P1_U2870) );
  INV_X1 U17348 ( .A(n13969), .ZN(n14031) );
  OAI211_X1 U17349 ( .C1(n14031), .C2(n13300), .A(n15294), .B(n14030), .ZN(
        n14033) );
  NAND2_X1 U17350 ( .A1(n13920), .A2(n16524), .ZN(n14032) );
  OAI211_X1 U17351 ( .C1(n13920), .C2(n12396), .A(n14033), .B(n14032), .ZN(
        P2_U2878) );
  AND2_X1 U17352 ( .A1(n10549), .A2(n14035), .ZN(n14034) );
  NAND2_X2 U17353 ( .A1(n14836), .A2(n14034), .ZN(n14839) );
  NAND2_X1 U17354 ( .A1(n14836), .A2(n10545), .ZN(n14831) );
  NAND2_X1 U17355 ( .A1(n20495), .A2(DATAI_1_), .ZN(n14038) );
  NAND2_X1 U17356 ( .A1(n20497), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14037) );
  AND2_X1 U17357 ( .A1(n14038), .A2(n14037), .ZN(n20520) );
  OAI222_X1 U17358 ( .A1(n14536), .A2(n14839), .B1(n14838), .B2(n20520), .C1(
        n14836), .C2(n10664), .ZN(P1_U2903) );
  NAND2_X1 U17359 ( .A1(n14039), .A2(n15128), .ZN(n14057) );
  INV_X1 U17360 ( .A(n9862), .ZN(n14042) );
  NAND2_X1 U17361 ( .A1(n13839), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14040) );
  NAND2_X1 U17362 ( .A1(n14040), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14041) );
  NAND2_X1 U17363 ( .A1(n14042), .A2(n14041), .ZN(n21187) );
  NAND2_X1 U17364 ( .A1(n14043), .A2(n21187), .ZN(n14054) );
  MUX2_X1 U17365 ( .A(n14044), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13839), .Z(n14046) );
  NOR2_X1 U17366 ( .A1(n14046), .A2(n14045), .ZN(n14047) );
  NAND2_X1 U17367 ( .A1(n14048), .A2(n14047), .ZN(n14053) );
  NAND2_X1 U17368 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14050) );
  INV_X1 U17369 ( .A(n14050), .ZN(n14049) );
  MUX2_X1 U17370 ( .A(n14050), .B(n14049), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14051) );
  OR2_X1 U17371 ( .A1(n16012), .A2(n14051), .ZN(n14052) );
  OAI211_X1 U17372 ( .C1(n15128), .C2(n14054), .A(n14053), .B(n14052), .ZN(
        n14055) );
  INV_X1 U17373 ( .A(n14055), .ZN(n14056) );
  NAND2_X1 U17374 ( .A1(n14057), .A2(n14056), .ZN(n21190) );
  MUX2_X1 U17375 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21190), .S(
        n16014), .Z(n16026) );
  NAND2_X1 U17376 ( .A1(n16026), .A2(n16040), .ZN(n14059) );
  NOR2_X1 U17377 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16040), .ZN(n14071) );
  NAND2_X1 U17378 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14071), .ZN(
        n14058) );
  NAND2_X1 U17379 ( .A1(n14059), .A2(n14058), .ZN(n14063) );
  MUX2_X1 U17380 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14060), .S(
        n16014), .Z(n16019) );
  AOI22_X1 U17381 ( .A1(n14071), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16019), .B2(n16040), .ZN(n14061) );
  INV_X1 U17382 ( .A(n14061), .ZN(n14062) );
  NAND2_X1 U17383 ( .A1(n14063), .A2(n14062), .ZN(n16033) );
  OR2_X1 U17384 ( .A1(n16033), .A2(n14064), .ZN(n16045) );
  INV_X1 U17385 ( .A(n20665), .ZN(n20929) );
  XNOR2_X1 U17386 ( .A(n14065), .B(n14067), .ZN(n20332) );
  OAI21_X1 U17387 ( .B1(n20332), .B2(n14066), .A(n16014), .ZN(n14070) );
  INV_X1 U17388 ( .A(n16014), .ZN(n14068) );
  AOI21_X1 U17389 ( .B1(n14068), .B2(n14067), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n14069) );
  NAND2_X1 U17390 ( .A1(n14070), .A2(n14069), .ZN(n14073) );
  NAND2_X1 U17391 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n14071), .ZN(
        n14072) );
  NAND2_X1 U17392 ( .A1(n14073), .A2(n14072), .ZN(n16042) );
  NOR2_X1 U17393 ( .A1(n16042), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n14074) );
  AOI21_X1 U17394 ( .B1(n16045), .B2(n14074), .A(n16376), .ZN(n14075) );
  NOR2_X1 U17395 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21235) );
  INV_X1 U17396 ( .A(n20670), .ZN(n20505) );
  NOR3_X1 U17397 ( .A1(n9870), .A2(n21194), .A3(n20927), .ZN(n20563) );
  INV_X1 U17398 ( .A(n9870), .ZN(n14078) );
  NAND2_X1 U17399 ( .A1(n21206), .A2(n20927), .ZN(n21199) );
  NAND2_X1 U17400 ( .A1(n20931), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21208) );
  INV_X1 U17401 ( .A(n21208), .ZN(n21197) );
  OAI22_X1 U17402 ( .A1(n14078), .A2(n21199), .B1(n14077), .B2(n21197), .ZN(
        n14079) );
  OAI21_X1 U17403 ( .B1(n20563), .B2(n14079), .A(n21212), .ZN(n14080) );
  OAI21_X1 U17404 ( .B1(n21212), .B2(n20850), .A(n14080), .ZN(P1_U3477) );
  OAI222_X1 U17405 ( .A1(n14708), .A2(n14839), .B1(n20526), .B2(n14838), .C1(
        n14836), .C2(n10658), .ZN(P1_U2902) );
  OAI21_X1 U17406 ( .B1(n14081), .B2(n14083), .A(n14082), .ZN(n14148) );
  INV_X1 U17407 ( .A(n14163), .ZN(n14084) );
  AOI21_X1 U17408 ( .B1(n14086), .B2(n14085), .A(n14084), .ZN(n20453) );
  AOI22_X1 U17409 ( .A1(n20453), .A2(n14721), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14720), .ZN(n14087) );
  OAI21_X1 U17410 ( .B1(n14148), .B2(n14772), .A(n14087), .ZN(P1_U2869) );
  OAI222_X1 U17411 ( .A1(n14148), .A2(n14839), .B1(n20531), .B2(n14838), .C1(
        n14836), .C2(n10709), .ZN(P1_U2901) );
  INV_X1 U17412 ( .A(n14030), .ZN(n14091) );
  OAI211_X1 U17413 ( .C1(n14091), .C2(n13302), .A(n15294), .B(n14090), .ZN(
        n14096) );
  OR2_X1 U17414 ( .A1(n14093), .A2(n14092), .ZN(n14094) );
  AND2_X1 U17415 ( .A1(n14094), .A2(n14154), .ZN(n19310) );
  NAND2_X1 U17416 ( .A1(n13920), .A2(n19310), .ZN(n14095) );
  OAI211_X1 U17417 ( .C1(n13920), .C2(n10305), .A(n14096), .B(n14095), .ZN(
        P2_U2877) );
  AOI22_X1 U17418 ( .A1(n20426), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20425), .ZN(n14101) );
  NAND2_X1 U17419 ( .A1(n20495), .A2(DATAI_0_), .ZN(n14099) );
  NAND2_X1 U17420 ( .A1(n20497), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14098) );
  AND2_X1 U17421 ( .A1(n14099), .A2(n14098), .ZN(n20510) );
  INV_X1 U17422 ( .A(n20510), .ZN(n14100) );
  NAND2_X1 U17423 ( .A1(n20411), .A2(n14100), .ZN(n14112) );
  NAND2_X1 U17424 ( .A1(n14101), .A2(n14112), .ZN(P1_U2952) );
  AOI22_X1 U17425 ( .A1(n20426), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20425), .ZN(n14103) );
  NAND2_X1 U17426 ( .A1(n14103), .A2(n14102), .ZN(P1_U2939) );
  AOI22_X1 U17427 ( .A1(n20426), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20425), .ZN(n14105) );
  NAND2_X1 U17428 ( .A1(n14105), .A2(n14104), .ZN(P1_U2944) );
  AOI22_X1 U17429 ( .A1(n20426), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20425), .ZN(n14107) );
  INV_X1 U17430 ( .A(n20520), .ZN(n14106) );
  NAND2_X1 U17431 ( .A1(n20411), .A2(n14106), .ZN(n14116) );
  NAND2_X1 U17432 ( .A1(n14107), .A2(n14116), .ZN(P1_U2953) );
  AOI22_X1 U17433 ( .A1(n20426), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20425), .ZN(n14109) );
  NAND2_X1 U17434 ( .A1(n14109), .A2(n14108), .ZN(P1_U2941) );
  AOI22_X1 U17435 ( .A1(n20426), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20425), .ZN(n14111) );
  NAND2_X1 U17436 ( .A1(n14111), .A2(n14110), .ZN(P1_U2942) );
  AOI22_X1 U17437 ( .A1(n20426), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20425), .ZN(n14113) );
  NAND2_X1 U17438 ( .A1(n14113), .A2(n14112), .ZN(P1_U2937) );
  AOI22_X1 U17439 ( .A1(n20426), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20425), .ZN(n14115) );
  NAND2_X1 U17440 ( .A1(n14115), .A2(n14114), .ZN(P1_U2940) );
  AOI22_X1 U17441 ( .A1(n20426), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20425), .ZN(n14117) );
  NAND2_X1 U17442 ( .A1(n14117), .A2(n14116), .ZN(P1_U2938) );
  AOI22_X1 U17443 ( .A1(n20426), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20425), .ZN(n14119) );
  NAND2_X1 U17444 ( .A1(n14119), .A2(n14118), .ZN(P1_U2943) );
  XNOR2_X1 U17445 ( .A(n14121), .B(n14122), .ZN(n20459) );
  NOR2_X1 U17446 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16040), .ZN(n21228) );
  NAND2_X1 U17447 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21228), .ZN(n16370) );
  INV_X1 U17448 ( .A(n16370), .ZN(n14123) );
  NAND2_X1 U17449 ( .A1(n21194), .A2(n14124), .ZN(n21226) );
  NAND2_X1 U17450 ( .A1(n21226), .A2(n20500), .ZN(n14125) );
  NAND2_X1 U17451 ( .A1(n20500), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21119) );
  NAND2_X1 U17452 ( .A1(n20927), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14126) );
  AND2_X1 U17453 ( .A1(n21119), .A2(n14126), .ZN(n20433) );
  INV_X1 U17454 ( .A(n20433), .ZN(n14127) );
  AOI22_X1 U17455 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14128) );
  OAI21_X1 U17456 ( .B1(n14701), .B2(n16219), .A(n14128), .ZN(n14129) );
  AOI21_X1 U17457 ( .B1(n14130), .B2(n16214), .A(n14129), .ZN(n14131) );
  OAI21_X1 U17458 ( .B1(n20258), .B2(n20459), .A(n14131), .ZN(P1_U2997) );
  XNOR2_X1 U17459 ( .A(n9833), .B(n14133), .ZN(n20482) );
  NAND2_X1 U17460 ( .A1(n20482), .A2(n20435), .ZN(n14137) );
  INV_X1 U17461 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20273) );
  OR2_X1 U17462 ( .A1(n20447), .A2(n20273), .ZN(n20477) );
  OAI21_X1 U17463 ( .B1(n20432), .B2(n14135), .A(n20477), .ZN(n14134) );
  AOI21_X1 U17464 ( .B1(n16189), .B2(n14135), .A(n14134), .ZN(n14136) );
  OAI211_X1 U17465 ( .C1(n14536), .C2(n20496), .A(n14137), .B(n14136), .ZN(
        P1_U2998) );
  OR2_X1 U17466 ( .A1(n14138), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14140) );
  AND2_X1 U17467 ( .A1(n14140), .A2(n14139), .ZN(n20485) );
  INV_X1 U17468 ( .A(n20485), .ZN(n14145) );
  OAI21_X1 U17469 ( .B1(n14143), .B2(n14142), .A(n14141), .ZN(n20438) );
  OAI222_X1 U17470 ( .A1(n14145), .A2(n14768), .B1(n14144), .B2(n14770), .C1(
        n20438), .C2(n14767), .ZN(P1_U2872) );
  XNOR2_X1 U17471 ( .A(n14147), .B(n14146), .ZN(n20450) );
  INV_X1 U17472 ( .A(n14148), .ZN(n20358) );
  AOI22_X1 U17473 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14149) );
  OAI21_X1 U17474 ( .B1(n20348), .B2(n16219), .A(n14149), .ZN(n14150) );
  AOI21_X1 U17475 ( .B1(n20358), .B2(n16214), .A(n14150), .ZN(n14151) );
  OAI21_X1 U17476 ( .B1(n20450), .B2(n20258), .A(n14151), .ZN(P1_U2996) );
  AOI211_X1 U17477 ( .C1(n14152), .C2(n14090), .A(n15289), .B(n9904), .ZN(
        n14153) );
  INV_X1 U17478 ( .A(n14153), .ZN(n14158) );
  NAND2_X1 U17479 ( .A1(n14155), .A2(n14154), .ZN(n14156) );
  AND2_X1 U17480 ( .A1(n14156), .A2(n10349), .ZN(n16505) );
  INV_X1 U17481 ( .A(n16505), .ZN(n15786) );
  OR2_X1 U17482 ( .A1(n15273), .A2(n15786), .ZN(n14157) );
  OAI211_X1 U17483 ( .C1(n13920), .C2(n14159), .A(n14158), .B(n14157), .ZN(
        P2_U2876) );
  INV_X1 U17484 ( .A(n14160), .ZN(n14161) );
  AOI21_X1 U17485 ( .B1(n14162), .B2(n14082), .A(n14161), .ZN(n14178) );
  INV_X1 U17486 ( .A(n14178), .ZN(n20336) );
  INV_X1 U17487 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20382) );
  OAI222_X1 U17488 ( .A1(n20336), .A2(n14839), .B1(n20537), .B2(n14838), .C1(
        n14836), .C2(n20382), .ZN(P1_U2900) );
  AOI21_X1 U17489 ( .B1(n14164), .B2(n14163), .A(n14184), .ZN(n20444) );
  INV_X1 U17490 ( .A(n20444), .ZN(n14165) );
  OAI222_X1 U17491 ( .A1(n14165), .A2(n14768), .B1(n14770), .B2(n11463), .C1(
        n20336), .C2(n14767), .ZN(P1_U2868) );
  OR2_X1 U17492 ( .A1(n14167), .A2(n14166), .ZN(n14168) );
  AND2_X1 U17493 ( .A1(n14256), .A2(n14168), .ZN(n19299) );
  INV_X1 U17494 ( .A(n19299), .ZN(n15762) );
  OAI211_X1 U17495 ( .C1(n9904), .C2(n14170), .A(n14169), .B(n15294), .ZN(
        n14172) );
  NAND2_X1 U17496 ( .A1(n13754), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14171) );
  OAI211_X1 U17497 ( .C1(n15762), .C2(n15273), .A(n14172), .B(n14171), .ZN(
        P2_U2875) );
  XNOR2_X1 U17498 ( .A(n14174), .B(n14173), .ZN(n20440) );
  INV_X1 U17499 ( .A(n14175), .ZN(n20334) );
  INV_X1 U17500 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21140) );
  NOR2_X1 U17501 ( .A1(n20447), .A2(n21140), .ZN(n20443) );
  AOI21_X1 U17502 ( .B1(n16209), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20443), .ZN(n14176) );
  OAI21_X1 U17503 ( .B1(n20334), .B2(n16219), .A(n14176), .ZN(n14177) );
  AOI21_X1 U17504 ( .B1(n14178), .B2(n16214), .A(n14177), .ZN(n14179) );
  OAI21_X1 U17505 ( .B1(n20258), .B2(n20440), .A(n14179), .ZN(P1_U2995) );
  AND2_X1 U17506 ( .A1(n14181), .A2(n14160), .ZN(n14182) );
  OR2_X1 U17507 ( .A1(n14180), .A2(n14182), .ZN(n20322) );
  OAI21_X1 U17508 ( .B1(n14184), .B2(n14183), .A(n14221), .ZN(n14185) );
  INV_X1 U17509 ( .A(n14185), .ZN(n20321) );
  AOI22_X1 U17510 ( .A1(n20321), .A2(n14721), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14720), .ZN(n14186) );
  OAI21_X1 U17511 ( .B1(n20322), .B2(n14772), .A(n14186), .ZN(P1_U2867) );
  OAI222_X1 U17512 ( .A1(n20322), .A2(n14839), .B1(n20542), .B2(n14838), .C1(
        n14187), .C2(n14836), .ZN(P1_U2899) );
  OAI222_X1 U17513 ( .A1(n20438), .A2(n14839), .B1(n14838), .B2(n20510), .C1(
        n14836), .C2(n10672), .ZN(P1_U2904) );
  NAND2_X1 U17514 ( .A1(n19704), .A2(n20199), .ZN(n14188) );
  NAND2_X1 U17515 ( .A1(n14188), .A2(n20206), .ZN(n14205) );
  NAND2_X1 U17516 ( .A1(n20209), .A2(n21487), .ZN(n19620) );
  INV_X1 U17517 ( .A(n19620), .ZN(n19618) );
  NAND2_X1 U17518 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19618), .ZN(
        n14204) );
  INV_X1 U17519 ( .A(n14204), .ZN(n14189) );
  OR2_X1 U17520 ( .A1(n14205), .A2(n14189), .ZN(n14193) );
  NAND2_X1 U17521 ( .A1(n14202), .A2(n19873), .ZN(n14191) );
  NOR2_X1 U17522 ( .A1(n19907), .A2(n19620), .ZN(n19665) );
  NOR2_X1 U17523 ( .A1(n19665), .A2(n20206), .ZN(n14190) );
  AOI21_X1 U17524 ( .B1(n14191), .B2(n14190), .A(n19981), .ZN(n14192) );
  NAND2_X1 U17525 ( .A1(n14193), .A2(n14192), .ZN(n19667) );
  INV_X1 U17526 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14209) );
  AOI22_X1 U17527 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19567), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19568), .ZN(n20028) );
  INV_X1 U17528 ( .A(n20028), .ZN(n19883) );
  INV_X1 U17529 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16742) );
  INV_X1 U17530 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n14197) );
  OAI22_X2 U17531 ( .A1(n16742), .A2(n19561), .B1(n14197), .B2(n19559), .ZN(
        n20014) );
  INV_X1 U17532 ( .A(n20014), .ZN(n14232) );
  INV_X1 U17533 ( .A(n19780), .ZN(n14198) );
  INV_X1 U17534 ( .A(n19665), .ZN(n14200) );
  NAND2_X1 U17535 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20020), .ZN(n19546) );
  NAND2_X1 U17536 ( .A1(n14199), .A2(n19569), .ZN(n19771) );
  OAI22_X1 U17537 ( .A1(n14232), .A2(n19697), .B1(n14200), .B2(n19771), .ZN(
        n14201) );
  AOI21_X1 U17538 ( .B1(n19659), .B2(n19883), .A(n14201), .ZN(n14208) );
  OAI21_X1 U17539 ( .B1(n14202), .B2(n19665), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14203) );
  OAI21_X1 U17540 ( .B1(n14205), .B2(n14204), .A(n14203), .ZN(n19666) );
  NAND2_X1 U17541 ( .A1(n19666), .A2(n14206), .ZN(n14207) );
  OAI211_X1 U17542 ( .C1(n19664), .C2(n14209), .A(n14208), .B(n14207), .ZN(
        P2_U3072) );
  INV_X1 U17543 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14215) );
  INV_X1 U17544 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18513) );
  INV_X1 U17545 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16728) );
  OAI22_X2 U17546 ( .A1(n18513), .A2(n19559), .B1(n16728), .B2(n19561), .ZN(
        n20053) );
  INV_X1 U17547 ( .A(n20053), .ZN(n14249) );
  AOI22_X2 U17548 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19568), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19567), .ZN(n20031) );
  INV_X1 U17549 ( .A(n20031), .ZN(n20052) );
  AOI22_X1 U17550 ( .A1(n20052), .A2(n19700), .B1(n20051), .B2(n19665), .ZN(
        n14212) );
  OAI21_X1 U17551 ( .B1(n14249), .B2(n19670), .A(n14212), .ZN(n14213) );
  AOI21_X1 U17552 ( .B1(n14210), .B2(n19666), .A(n14213), .ZN(n14214) );
  OAI21_X1 U17553 ( .B1(n19664), .B2(n14215), .A(n14214), .ZN(P2_U3073) );
  OR2_X1 U17554 ( .A1(n14180), .A2(n14217), .ZN(n14218) );
  AND2_X1 U17555 ( .A1(n14216), .A2(n14218), .ZN(n20308) );
  INV_X1 U17556 ( .A(n20308), .ZN(n14223) );
  INV_X1 U17557 ( .A(n14219), .ZN(n14220) );
  XNOR2_X1 U17558 ( .A(n14221), .B(n14220), .ZN(n20306) );
  AOI22_X1 U17559 ( .A1(n20306), .A2(n14721), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14720), .ZN(n14222) );
  OAI21_X1 U17560 ( .B1(n14223), .B2(n14772), .A(n14222), .ZN(P1_U2866) );
  OAI222_X1 U17561 ( .A1(n14223), .A2(n14839), .B1(n20547), .B2(n14838), .C1(
        n14836), .C2(n10773), .ZN(P1_U2898) );
  NOR2_X1 U17562 ( .A1(n20202), .A2(n20197), .ZN(n19984) );
  INV_X1 U17563 ( .A(n19984), .ZN(n14224) );
  INV_X1 U17564 ( .A(n19583), .ZN(n19589) );
  OAI21_X1 U17565 ( .B1(n14224), .B2(n19589), .A(n20206), .ZN(n14230) );
  NAND2_X1 U17566 ( .A1(n21487), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19912) );
  INV_X1 U17567 ( .A(n19912), .ZN(n19908) );
  NAND2_X1 U17568 ( .A1(n19908), .A2(n21540), .ZN(n19822) );
  INV_X1 U17569 ( .A(n19822), .ZN(n14227) );
  NAND2_X1 U17570 ( .A1(n21540), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19577) );
  NOR2_X1 U17571 ( .A1(n19577), .A2(n19912), .ZN(n19872) );
  INV_X1 U17572 ( .A(n19872), .ZN(n14225) );
  INV_X1 U17573 ( .A(n20206), .ZN(n20198) );
  OAI211_X1 U17574 ( .C1(n12017), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n14225), 
        .B(n20198), .ZN(n14226) );
  OAI211_X1 U17575 ( .C1(n14230), .C2(n14227), .A(n20020), .B(n14226), .ZN(
        n19867) );
  INV_X1 U17576 ( .A(n19867), .ZN(n14236) );
  OAI21_X1 U17577 ( .B1(n14228), .B2(n19872), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14229) );
  OAI21_X1 U17578 ( .B1(n14230), .B2(n19822), .A(n14229), .ZN(n19866) );
  INV_X1 U17579 ( .A(n19771), .ZN(n20013) );
  AOI22_X1 U17580 ( .A1(n19883), .A2(n19857), .B1(n20013), .B2(n19872), .ZN(
        n14231) );
  OAI21_X1 U17581 ( .B1(n14232), .B2(n19900), .A(n14231), .ZN(n14233) );
  AOI21_X1 U17582 ( .B1(n19866), .B2(n14206), .A(n14233), .ZN(n14234) );
  OAI21_X1 U17583 ( .B1(n14236), .B2(n14235), .A(n14234), .ZN(P2_U3120) );
  NAND2_X1 U17584 ( .A1(n19583), .A2(n19675), .ZN(n19617) );
  OAI21_X1 U17585 ( .B1(n20092), .B2(n19605), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14237) );
  NAND2_X1 U17586 ( .A1(n14237), .A2(n20206), .ZN(n14247) );
  NAND2_X1 U17587 ( .A1(n19618), .A2(n21540), .ZN(n19585) );
  NOR2_X1 U17588 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19585), .ZN(
        n19571) );
  INV_X1 U17589 ( .A(n19571), .ZN(n14238) );
  NAND2_X1 U17590 ( .A1(n14272), .A2(n14238), .ZN(n14243) );
  OR2_X1 U17591 ( .A1(n14247), .A2(n14243), .ZN(n14242) );
  OR2_X1 U17592 ( .A1(n11899), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14240) );
  NOR2_X1 U17593 ( .A1(n20206), .A2(n19571), .ZN(n14239) );
  AOI21_X1 U17594 ( .B1(n14240), .B2(n14239), .A(n19981), .ZN(n14241) );
  NAND2_X1 U17595 ( .A1(n14242), .A2(n14241), .ZN(n19574) );
  INV_X1 U17596 ( .A(n14243), .ZN(n14246) );
  INV_X1 U17597 ( .A(n11899), .ZN(n14244) );
  OAI21_X1 U17598 ( .B1(n14244), .B2(n19571), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14245) );
  INV_X1 U17599 ( .A(n20092), .ZN(n14357) );
  AOI22_X1 U17600 ( .A1(n20052), .A2(n19605), .B1(n20051), .B2(n19571), .ZN(
        n14248) );
  OAI21_X1 U17601 ( .B1(n14249), .B2(n14357), .A(n14248), .ZN(n14250) );
  AOI21_X1 U17602 ( .B1(n19573), .B2(n14210), .A(n14250), .ZN(n14251) );
  OAI21_X1 U17603 ( .B1(n19566), .B2(n14252), .A(n14251), .ZN(P2_U3049) );
  INV_X1 U17604 ( .A(n14169), .ZN(n14254) );
  OAI211_X1 U17605 ( .C1(n14254), .C2(n10361), .A(n15294), .B(n9941), .ZN(
        n14259) );
  NAND2_X1 U17606 ( .A1(n14256), .A2(n14255), .ZN(n14257) );
  AND2_X1 U17607 ( .A1(n14378), .A2(n14257), .ZN(n19283) );
  INV_X1 U17608 ( .A(n19283), .ZN(n15747) );
  OR2_X1 U17609 ( .A1(n15273), .A2(n15747), .ZN(n14258) );
  OAI211_X1 U17610 ( .C1(n13920), .C2(n12404), .A(n14259), .B(n14258), .ZN(
        P2_U2874) );
  NAND2_X1 U17611 ( .A1(n19984), .A2(n14269), .ZN(n14260) );
  OR2_X1 U17612 ( .A1(n20209), .A2(n20012), .ZN(n14266) );
  NAND2_X1 U17613 ( .A1(n14260), .A2(n14266), .ZN(n14265) );
  INV_X1 U17614 ( .A(n14272), .ZN(n20088) );
  AND2_X1 U17615 ( .A1(n14272), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14261) );
  NAND2_X1 U17616 ( .A1(n14262), .A2(n14261), .ZN(n14268) );
  OAI211_X1 U17617 ( .C1(n20088), .C2(n19873), .A(n14268), .B(n20020), .ZN(
        n14263) );
  INV_X1 U17618 ( .A(n14263), .ZN(n14264) );
  NAND2_X1 U17619 ( .A1(n14265), .A2(n14264), .ZN(n20093) );
  INV_X1 U17620 ( .A(n20093), .ZN(n20058) );
  INV_X1 U17621 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14275) );
  INV_X1 U17622 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19913) );
  OAI21_X1 U17623 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n14266), .A(n19913), 
        .ZN(n14267) );
  AND2_X1 U17624 ( .A1(n14268), .A2(n14267), .ZN(n20090) );
  AOI22_X1 U17625 ( .A1(n20092), .A2(n20014), .B1(n20054), .B2(n19883), .ZN(
        n14271) );
  OAI21_X1 U17626 ( .B1(n19771), .B2(n14272), .A(n14271), .ZN(n14273) );
  AOI21_X1 U17627 ( .B1(n20090), .B2(n14206), .A(n14273), .ZN(n14274) );
  OAI21_X1 U17628 ( .B1(n20058), .B2(n14275), .A(n14274), .ZN(P2_U3168) );
  INV_X1 U17629 ( .A(n19381), .ZN(n15179) );
  INV_X1 U17630 ( .A(n19498), .ZN(n14279) );
  NOR2_X1 U17631 ( .A1(n9878), .A2(n14276), .ZN(n14278) );
  AOI21_X1 U17632 ( .B1(n14279), .B2(n14278), .A(n19334), .ZN(n14277) );
  OAI21_X1 U17633 ( .B1(n14279), .B2(n14278), .A(n14277), .ZN(n14288) );
  AOI21_X1 U17634 ( .B1(n14281), .B2(n14280), .A(n9972), .ZN(n19504) );
  AOI22_X1 U17635 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19356), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19369), .ZN(n14282) );
  OAI211_X1 U17636 ( .C1(n19353), .C2(n12382), .A(n14282), .B(n19348), .ZN(
        n14283) );
  AOI21_X1 U17637 ( .B1(n19275), .B2(n19504), .A(n14283), .ZN(n14284) );
  OAI21_X1 U17638 ( .B1(n14285), .B2(n19351), .A(n14284), .ZN(n14286) );
  AOI21_X1 U17639 ( .B1(n19501), .B2(n19364), .A(n14286), .ZN(n14287) );
  OAI211_X1 U17640 ( .C1(n19425), .C2(n15179), .A(n14288), .B(n14287), .ZN(
        P2_U2851) );
  NOR2_X1 U17641 ( .A1(n9824), .A2(n14289), .ZN(n14290) );
  XNOR2_X1 U17642 ( .A(n14290), .B(n16540), .ZN(n14291) );
  NAND2_X1 U17643 ( .A1(n14291), .A2(n20102), .ZN(n14299) );
  AOI21_X1 U17644 ( .B1(n14293), .B2(n15793), .A(n14292), .ZN(n19408) );
  AOI22_X1 U17645 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19356), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19369), .ZN(n14294) );
  OAI211_X1 U17646 ( .C1(n19353), .C2(n14295), .A(n14294), .B(n19348), .ZN(
        n14297) );
  NOR2_X1 U17647 ( .A1(n16591), .A2(n19343), .ZN(n14296) );
  AOI211_X1 U17648 ( .C1(n19275), .C2(n19408), .A(n14297), .B(n14296), .ZN(
        n14298) );
  OAI211_X1 U17649 ( .C1(n19351), .C2(n14300), .A(n14299), .B(n14298), .ZN(
        P2_U2847) );
  NAND2_X1 U17650 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21235), .ZN(n16046) );
  NAND2_X1 U17651 ( .A1(n9819), .A2(n21228), .ZN(n14301) );
  OAI211_X1 U17652 ( .C1(n16046), .C2(n20500), .A(n20447), .B(n14301), .ZN(
        n14302) );
  INV_X1 U17653 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14853) );
  XNOR2_X1 U17654 ( .A(n14304), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14843) );
  NOR2_X1 U17655 ( .A1(n14843), .A2(n16040), .ZN(n14305) );
  NAND2_X1 U17656 ( .A1(n21225), .A2(n14306), .ZN(n14307) );
  NAND2_X1 U17657 ( .A1(n20294), .A2(n14307), .ZN(n20357) );
  INV_X1 U17658 ( .A(n20357), .ZN(n20335) );
  AND2_X1 U17659 ( .A1(n21224), .A2(n20927), .ZN(n16037) );
  NAND2_X1 U17660 ( .A1(n14308), .A2(n16037), .ZN(n14311) );
  NOR2_X1 U17661 ( .A1(n14311), .A2(n14309), .ZN(n14310) );
  INV_X1 U17662 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14323) );
  INV_X1 U17663 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14709) );
  OR2_X1 U17664 ( .A1(n11545), .A2(n14709), .ZN(n14313) );
  AND3_X1 U17665 ( .A1(n14313), .A2(n20501), .A3(n14311), .ZN(n14312) );
  NOR2_X1 U17666 ( .A1(n14313), .A2(n16037), .ZN(n14314) );
  NAND2_X1 U17667 ( .A1(n20345), .A2(n20485), .ZN(n14317) );
  AND2_X1 U17668 ( .A1(n14843), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14315) );
  OAI21_X1 U17669 ( .B1(n20351), .B2(n20350), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14316) );
  OAI211_X1 U17670 ( .C1(n20330), .C2(n14144), .A(n14317), .B(n14316), .ZN(
        n14318) );
  INV_X1 U17671 ( .A(n14318), .ZN(n14322) );
  INV_X1 U17672 ( .A(n14319), .ZN(n14320) );
  AND2_X1 U17673 ( .A1(n21225), .A2(n14320), .ZN(n20347) );
  NAND2_X1 U17674 ( .A1(n21209), .A2(n20347), .ZN(n14321) );
  OAI211_X1 U17675 ( .C1(n14558), .C2(n14323), .A(n14322), .B(n14321), .ZN(
        n14324) );
  INV_X1 U17676 ( .A(n14324), .ZN(n14325) );
  OAI21_X1 U17677 ( .B1(n20438), .B2(n20335), .A(n14325), .ZN(P1_U2840) );
  NAND2_X1 U17678 ( .A1(n14216), .A2(n14327), .ZN(n14328) );
  AND2_X1 U17679 ( .A1(n14326), .A2(n14328), .ZN(n16205) );
  INV_X1 U17680 ( .A(n16205), .ZN(n14329) );
  INV_X1 U17681 ( .A(n14802), .ZN(n20556) );
  OAI222_X1 U17682 ( .A1(n14329), .A2(n14839), .B1(n20556), .B2(n14838), .C1(
        n14836), .C2(n10783), .ZN(P1_U2897) );
  NOR2_X1 U17683 ( .A1(n9878), .A2(n14330), .ZN(n15199) );
  XNOR2_X1 U17684 ( .A(n15199), .B(n14331), .ZN(n14332) );
  NAND2_X1 U17685 ( .A1(n14332), .A2(n20102), .ZN(n14340) );
  NAND2_X1 U17686 ( .A1(n20214), .A2(n19275), .ZN(n14335) );
  OAI22_X1 U17687 ( .A1(n11792), .A2(n19353), .B1(n20133), .B2(n19349), .ZN(
        n14333) );
  AOI21_X1 U17688 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19356), .A(
        n14333), .ZN(n14334) );
  OAI211_X1 U17689 ( .C1(n19351), .C2(n14336), .A(n14335), .B(n14334), .ZN(
        n14337) );
  AOI21_X1 U17690 ( .B1(n14338), .B2(n19364), .A(n14337), .ZN(n14339) );
  OAI211_X1 U17691 ( .C1(n15179), .C2(n20212), .A(n14340), .B(n14339), .ZN(
        P2_U2853) );
  AND2_X1 U17692 ( .A1(n14342), .A2(n14341), .ZN(n14343) );
  OR2_X1 U17693 ( .A1(n14343), .A2(n14365), .ZN(n16345) );
  INV_X1 U17694 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14344) );
  OAI22_X1 U17695 ( .A1(n16345), .A2(n14768), .B1(n14344), .B2(n14770), .ZN(
        n14345) );
  AOI21_X1 U17696 ( .B1(n16205), .B2(n14511), .A(n14345), .ZN(n14346) );
  INV_X1 U17697 ( .A(n14346), .ZN(P1_U2865) );
  INV_X1 U17698 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n16344) );
  NAND2_X1 U17699 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n14347) );
  NAND2_X1 U17700 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20346) );
  NOR3_X1 U17701 ( .A1(n20273), .A2(n21140), .A3(n20346), .ZN(n14469) );
  NAND2_X1 U17702 ( .A1(n14469), .A2(n16076), .ZN(n20323) );
  OAI21_X1 U17703 ( .B1(n14347), .B2(n20323), .A(n20324), .ZN(n20314) );
  NAND2_X1 U17704 ( .A1(n20351), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14348) );
  OAI211_X1 U17705 ( .C1(n20333), .C2(n16208), .A(n20447), .B(n14348), .ZN(
        n14351) );
  INV_X1 U17706 ( .A(n14676), .ZN(n16078) );
  NAND2_X1 U17707 ( .A1(n16078), .A2(n14469), .ZN(n20318) );
  NAND3_X1 U17708 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n16344), .ZN(n14349) );
  OAI22_X1 U17709 ( .A1(n20301), .A2(n16345), .B1(n20318), .B2(n14349), .ZN(
        n14350) );
  AOI211_X1 U17710 ( .C1(n20344), .C2(P1_EBX_REG_7__SCAN_IN), .A(n14351), .B(
        n14350), .ZN(n14353) );
  NAND2_X1 U17711 ( .A1(n16205), .A2(n20307), .ZN(n14352) );
  OAI211_X1 U17712 ( .C1(n16344), .C2(n20314), .A(n14353), .B(n14352), .ZN(
        P1_U2833) );
  INV_X1 U17713 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16726) );
  INV_X1 U17714 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n21500) );
  INV_X1 U17715 ( .A(n20033), .ZN(n20063) );
  AOI22_X1 U17716 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19568), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19567), .ZN(n20036) );
  INV_X1 U17717 ( .A(n20036), .ZN(n20060) );
  AOI22_X1 U17718 ( .A1(n20060), .A2(n19605), .B1(n20059), .B2(n19571), .ZN(
        n14356) );
  OAI21_X1 U17719 ( .B1(n20063), .B2(n14357), .A(n14356), .ZN(n14358) );
  AOI21_X1 U17720 ( .B1(n19573), .B2(n14355), .A(n14358), .ZN(n14359) );
  OAI21_X1 U17721 ( .B1(n19566), .B2(n14360), .A(n14359), .ZN(P2_U3050) );
  OAI21_X1 U17722 ( .B1(n10805), .B2(n10379), .A(n14361), .ZN(n20295) );
  INV_X1 U17723 ( .A(DATAI_8_), .ZN(n14362) );
  INV_X1 U17724 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16753) );
  MUX2_X1 U17725 ( .A(n14362), .B(n16753), .S(n20497), .Z(n20390) );
  INV_X1 U17726 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14363) );
  OAI222_X1 U17727 ( .A1(n20295), .A2(n14839), .B1(n20390), .B2(n14838), .C1(
        n14363), .C2(n14836), .ZN(P1_U2896) );
  INV_X1 U17728 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14367) );
  OR2_X1 U17729 ( .A1(n14365), .A2(n14364), .ZN(n14366) );
  NAND2_X1 U17730 ( .A1(n14419), .A2(n14366), .ZN(n20300) );
  OAI222_X1 U17731 ( .A1(n20295), .A2(n14772), .B1(n14770), .B2(n14367), .C1(
        n20300), .C2(n14768), .ZN(P1_U2864) );
  INV_X1 U17732 ( .A(n14371), .ZN(n14372) );
  OAI211_X1 U17733 ( .C1(n14369), .C2(n14373), .A(n14372), .B(n15294), .ZN(
        n14376) );
  AOI21_X1 U17734 ( .B1(n14374), .B2(n14380), .A(n14389), .ZN(n16573) );
  NAND2_X1 U17735 ( .A1(n16573), .A2(n13920), .ZN(n14375) );
  OAI211_X1 U17736 ( .C1(n13920), .C2(n12412), .A(n14376), .B(n14375), .ZN(
        P2_U2872) );
  NAND2_X1 U17737 ( .A1(n14378), .A2(n14377), .ZN(n14379) );
  AND2_X1 U17738 ( .A1(n14380), .A2(n14379), .ZN(n19276) );
  INV_X1 U17739 ( .A(n19276), .ZN(n14381) );
  NOR2_X1 U17740 ( .A1(n14381), .A2(n15273), .ZN(n14384) );
  AOI211_X1 U17741 ( .C1(n14382), .C2(n9941), .A(n15289), .B(n14369), .ZN(
        n14383) );
  AOI211_X1 U17742 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n13754), .A(n14384), .B(
        n14383), .ZN(n14385) );
  INV_X1 U17743 ( .A(n14385), .ZN(P2_U2873) );
  OAI21_X1 U17744 ( .B1(n14371), .B2(n14387), .A(n14386), .ZN(n15393) );
  OAI21_X1 U17745 ( .B1(n14389), .B2(n14388), .A(n14455), .ZN(n15514) );
  NOR2_X1 U17746 ( .A1(n15514), .A2(n15273), .ZN(n14390) );
  AOI21_X1 U17747 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n13754), .A(n14390), .ZN(
        n14391) );
  OAI21_X1 U17748 ( .B1(n15393), .B2(n15289), .A(n14391), .ZN(P2_U2871) );
  XNOR2_X1 U17749 ( .A(n14393), .B(n14392), .ZN(n16542) );
  OAI21_X1 U17750 ( .B1(n14397), .B2(n14395), .A(n14394), .ZN(n14396) );
  OAI21_X1 U17751 ( .B1(n14398), .B2(n14397), .A(n14396), .ZN(n16544) );
  INV_X1 U17752 ( .A(n16544), .ZN(n14412) );
  OAI21_X1 U17753 ( .B1(n19523), .B2(n19522), .A(n14399), .ZN(n14400) );
  INV_X1 U17754 ( .A(n14400), .ZN(n16610) );
  OAI21_X1 U17755 ( .B1(n15726), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n16610), .ZN(n19505) );
  NAND2_X1 U17756 ( .A1(n14401), .A2(n19522), .ZN(n16612) );
  NOR2_X1 U17757 ( .A1(n16611), .A2(n16612), .ZN(n19503) );
  INV_X1 U17758 ( .A(n19503), .ZN(n14402) );
  AOI211_X1 U17759 ( .C1(n14403), .C2(n19502), .A(n14432), .B(n14402), .ZN(
        n14405) );
  INV_X1 U17760 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20139) );
  NOR2_X1 U17761 ( .A1(n20139), .A2(n19348), .ZN(n14404) );
  AOI211_X1 U17762 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n19505), .A(
        n14405), .B(n14404), .ZN(n14406) );
  INV_X1 U17763 ( .A(n14406), .ZN(n14411) );
  OAI21_X1 U17764 ( .B1(n9972), .B2(n14408), .A(n14407), .ZN(n19422) );
  OAI22_X1 U17765 ( .A1(n19422), .A2(n16603), .B1(n19534), .B2(n14409), .ZN(
        n14410) );
  AOI211_X1 U17766 ( .C1(n14412), .C2(n12862), .A(n14411), .B(n14410), .ZN(
        n14413) );
  OAI21_X1 U17767 ( .B1(n16587), .B2(n16542), .A(n14413), .ZN(P2_U3041) );
  AND2_X1 U17768 ( .A1(n14361), .A2(n14414), .ZN(n14416) );
  OR2_X1 U17769 ( .A1(n14416), .A2(n14415), .ZN(n20283) );
  INV_X1 U17770 ( .A(n14462), .ZN(n14417) );
  AOI21_X1 U17771 ( .B1(n14419), .B2(n14418), .A(n14417), .ZN(n20282) );
  AOI22_X1 U17772 ( .A1(n20282), .A2(n14721), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14720), .ZN(n14420) );
  OAI21_X1 U17773 ( .B1(n20283), .B2(n14767), .A(n14420), .ZN(P1_U2863) );
  XNOR2_X1 U17774 ( .A(n14422), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14440) );
  INV_X1 U17775 ( .A(n14424), .ZN(n14425) );
  XNOR2_X1 U17776 ( .A(n14423), .B(n14425), .ZN(n14438) );
  INV_X1 U17777 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20141) );
  OAI22_X1 U17778 ( .A1(n20141), .A2(n19348), .B1(n19499), .B2(n19341), .ZN(
        n14427) );
  INV_X1 U17779 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19336) );
  OAI22_X1 U17780 ( .A1(n14195), .A2(n19342), .B1(n16561), .B2(n19336), .ZN(
        n14426) );
  AOI211_X1 U17781 ( .C1(n14438), .C2(n19493), .A(n14427), .B(n14426), .ZN(
        n14428) );
  OAI21_X1 U17782 ( .B1(n14440), .B2(n16543), .A(n14428), .ZN(P2_U3008) );
  XNOR2_X1 U17783 ( .A(n14430), .B(n14429), .ZN(n19414) );
  NAND3_X1 U17784 ( .A1(n14432), .A2(n19503), .A3(n14431), .ZN(n14436) );
  OAI21_X1 U17785 ( .B1(n15726), .B2(n14433), .A(n16610), .ZN(n16589) );
  OAI22_X1 U17786 ( .A1(n19534), .A2(n19342), .B1(n19233), .B2(n20141), .ZN(
        n14434) );
  AOI21_X1 U17787 ( .B1(n16589), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14434), .ZN(n14435) );
  OAI211_X1 U17788 ( .C1(n19414), .C2(n16603), .A(n14436), .B(n14435), .ZN(
        n14437) );
  AOI21_X1 U17789 ( .B1(n14438), .B2(n19526), .A(n14437), .ZN(n14439) );
  OAI21_X1 U17790 ( .B1(n14440), .B2(n16604), .A(n14439), .ZN(P2_U3040) );
  XNOR2_X1 U17791 ( .A(n14441), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14442) );
  XNOR2_X1 U17792 ( .A(n14443), .B(n14442), .ZN(n16338) );
  NAND2_X1 U17793 ( .A1(n16338), .A2(n20435), .ZN(n14447) );
  INV_X1 U17794 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n14444) );
  OAI22_X1 U17795 ( .A1(n20432), .A2(n20289), .B1(n20447), .B2(n14444), .ZN(
        n14445) );
  AOI21_X1 U17796 ( .B1(n16189), .B2(n20297), .A(n14445), .ZN(n14446) );
  OAI211_X1 U17797 ( .C1(n20496), .C2(n20295), .A(n14447), .B(n14446), .ZN(
        P1_U2991) );
  INV_X1 U17798 ( .A(DATAI_9_), .ZN(n14449) );
  MUX2_X1 U17799 ( .A(n14449), .B(n14448), .S(n20497), .Z(n20394) );
  INV_X1 U17800 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14450) );
  OAI222_X1 U17801 ( .A1(n20283), .A2(n14839), .B1(n20394), .B2(n14838), .C1(
        n14450), .C2(n14836), .ZN(P1_U2895) );
  INV_X1 U17802 ( .A(n14386), .ZN(n14453) );
  INV_X1 U17803 ( .A(n14451), .ZN(n14452) );
  OAI21_X1 U17804 ( .B1(n14453), .B2(n14452), .A(n9949), .ZN(n15380) );
  NAND2_X1 U17805 ( .A1(n13754), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14458) );
  INV_X1 U17806 ( .A(n15291), .ZN(n14454) );
  AOI21_X1 U17807 ( .B1(n14456), .B2(n14455), .A(n14454), .ZN(n19240) );
  NAND2_X1 U17808 ( .A1(n19240), .A2(n13920), .ZN(n14457) );
  OAI211_X1 U17809 ( .C1(n15380), .C2(n15289), .A(n14458), .B(n14457), .ZN(
        P2_U2870) );
  NOR2_X1 U17810 ( .A1(n14415), .A2(n14459), .ZN(n14460) );
  OR2_X1 U17811 ( .A1(n9922), .A2(n14460), .ZN(n15010) );
  AND2_X1 U17812 ( .A1(n14462), .A2(n14461), .ZN(n14463) );
  OR2_X1 U17813 ( .A1(n14463), .A2(n14484), .ZN(n16321) );
  OAI22_X1 U17814 ( .A1(n16321), .A2(n14768), .B1(n14464), .B2(n14770), .ZN(
        n14465) );
  INV_X1 U17815 ( .A(n14465), .ZN(n14466) );
  OAI21_X1 U17816 ( .B1(n15010), .B2(n14767), .A(n14466), .ZN(P1_U2862) );
  INV_X1 U17817 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20288) );
  NAND3_X1 U17818 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n20290) );
  NOR2_X1 U17819 ( .A1(n14444), .A2(n20290), .ZN(n14468) );
  NAND2_X1 U17820 ( .A1(n14469), .A2(n14468), .ZN(n14553) );
  NOR3_X1 U17821 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20288), .A3(n20279), 
        .ZN(n14467) );
  AOI211_X1 U17822 ( .C1(n20351), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20487), .B(n14467), .ZN(n14474) );
  INV_X1 U17823 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21150) );
  NOR2_X1 U17824 ( .A1(n21150), .A2(n20288), .ZN(n16155) );
  NAND3_X1 U17825 ( .A1(n14469), .A2(n14468), .A3(n16076), .ZN(n20276) );
  INV_X1 U17826 ( .A(n20276), .ZN(n14524) );
  AOI21_X1 U17827 ( .B1(n16155), .B2(n14524), .A(n14558), .ZN(n16161) );
  INV_X1 U17828 ( .A(n14470), .ZN(n15007) );
  AOI22_X1 U17829 ( .A1(n20344), .A2(P1_EBX_REG_10__SCAN_IN), .B1(n15007), 
        .B2(n20350), .ZN(n14471) );
  OAI21_X1 U17830 ( .B1(n16321), .B2(n20301), .A(n14471), .ZN(n14472) );
  AOI21_X1 U17831 ( .B1(n16161), .B2(P1_REIP_REG_10__SCAN_IN), .A(n14472), 
        .ZN(n14473) );
  OAI211_X1 U17832 ( .C1(n15010), .C2(n20294), .A(n14474), .B(n14473), .ZN(
        P1_U2830) );
  INV_X1 U17833 ( .A(DATAI_10_), .ZN(n14475) );
  INV_X1 U17834 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16750) );
  MUX2_X1 U17835 ( .A(n14475), .B(n16750), .S(n20497), .Z(n20398) );
  INV_X1 U17836 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14476) );
  OAI222_X1 U17837 ( .A1(n15010), .A2(n14839), .B1(n20398), .B2(n14838), .C1(
        n14476), .C2(n14836), .ZN(P1_U2894) );
  XNOR2_X1 U17838 ( .A(n15002), .B(n16332), .ZN(n14477) );
  XNOR2_X1 U17839 ( .A(n14478), .B(n14477), .ZN(n16327) );
  OAI22_X1 U17840 ( .A1(n20432), .A2(n20277), .B1(n20447), .B2(n20288), .ZN(
        n14480) );
  NOR2_X1 U17841 ( .A1(n20283), .A2(n20496), .ZN(n14479) );
  AOI211_X1 U17842 ( .C1(n16189), .C2(n20284), .A(n14480), .B(n14479), .ZN(
        n14481) );
  OAI21_X1 U17843 ( .B1(n20258), .B2(n16327), .A(n14481), .ZN(P1_U2990) );
  OAI21_X1 U17844 ( .B1(n9922), .B2(n14483), .A(n14482), .ZN(n14493) );
  XNOR2_X1 U17845 ( .A(n14493), .B(n14491), .ZN(n16198) );
  INV_X1 U17846 ( .A(n16198), .ZN(n14490) );
  AOI21_X1 U17847 ( .B1(n9984), .B2(n10105), .A(n14497), .ZN(n16307) );
  AOI22_X1 U17848 ( .A1(n16307), .A2(n14721), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14720), .ZN(n14485) );
  OAI21_X1 U17849 ( .B1(n14490), .B2(n14767), .A(n14485), .ZN(P1_U2861) );
  INV_X1 U17850 ( .A(n14838), .ZN(n14488) );
  INV_X1 U17851 ( .A(DATAI_11_), .ZN(n14487) );
  NAND2_X1 U17852 ( .A1(n20497), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14486) );
  OAI21_X1 U17853 ( .B1(n20497), .B2(n14487), .A(n14486), .ZN(n20401) );
  AOI22_X1 U17854 ( .A1(n14488), .A2(n20401), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14801), .ZN(n14489) );
  OAI21_X1 U17855 ( .B1(n14490), .B2(n14839), .A(n14489), .ZN(P1_U2893) );
  INV_X1 U17856 ( .A(n14491), .ZN(n14492) );
  OAI21_X1 U17857 ( .B1(n14493), .B2(n14492), .A(n14482), .ZN(n14515) );
  XNOR2_X1 U17858 ( .A(n14515), .B(n14514), .ZN(n16193) );
  INV_X1 U17859 ( .A(DATAI_12_), .ZN(n14494) );
  INV_X1 U17860 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16747) );
  MUX2_X1 U17861 ( .A(n14494), .B(n16747), .S(n20497), .Z(n20403) );
  INV_X1 U17862 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14495) );
  OAI222_X1 U17863 ( .A1(n16193), .A2(n14839), .B1(n20403), .B2(n14838), .C1(
        n14495), .C2(n14836), .ZN(P1_U2892) );
  INV_X1 U17864 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14499) );
  OR2_X1 U17865 ( .A1(n14497), .A2(n14496), .ZN(n14498) );
  NAND2_X1 U17866 ( .A1(n14519), .A2(n14498), .ZN(n16300) );
  OAI222_X1 U17867 ( .A1(n16193), .A2(n14772), .B1(n14770), .B2(n14499), .C1(
        n16300), .C2(n14768), .ZN(P1_U2860) );
  NAND2_X1 U17868 ( .A1(n14501), .A2(n14502), .ZN(n14503) );
  AND2_X1 U17869 ( .A1(n14500), .A2(n14503), .ZN(n16142) );
  INV_X1 U17870 ( .A(n16142), .ZN(n14507) );
  INV_X1 U17871 ( .A(DATAI_14_), .ZN(n14505) );
  INV_X1 U17872 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14504) );
  MUX2_X1 U17873 ( .A(n14505), .B(n14504), .S(n20497), .Z(n20409) );
  INV_X1 U17874 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14506) );
  OAI222_X1 U17875 ( .A1(n14507), .A2(n14839), .B1(n20409), .B2(n14838), .C1(
        n14506), .C2(n14836), .ZN(P1_U2890) );
  AND2_X1 U17876 ( .A1(n14521), .A2(n14508), .ZN(n14509) );
  OR2_X1 U17877 ( .A1(n14509), .A2(n14687), .ZN(n16277) );
  OAI22_X1 U17878 ( .A1(n16277), .A2(n14768), .B1(n21404), .B2(n14770), .ZN(
        n14510) );
  AOI21_X1 U17879 ( .B1(n16142), .B2(n14511), .A(n14510), .ZN(n14512) );
  INV_X1 U17880 ( .A(n14512), .ZN(P1_U2858) );
  AOI21_X1 U17881 ( .B1(n14515), .B2(n14514), .A(n14513), .ZN(n14517) );
  INV_X1 U17882 ( .A(n14501), .ZN(n14516) );
  INV_X1 U17883 ( .A(n14996), .ZN(n14533) );
  NAND2_X1 U17884 ( .A1(n14519), .A2(n14518), .ZN(n14520) );
  AND2_X1 U17885 ( .A1(n14521), .A2(n14520), .ZN(n16279) );
  AOI22_X1 U17886 ( .A1(n16279), .A2(n14721), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14720), .ZN(n14522) );
  OAI21_X1 U17887 ( .B1(n14533), .B2(n14767), .A(n14522), .ZN(P1_U2859) );
  INV_X1 U17888 ( .A(n14523), .ZN(n14994) );
  NAND2_X1 U17889 ( .A1(n14996), .A2(n20307), .ZN(n14529) );
  INV_X1 U17890 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21152) );
  NAND3_X1 U17891 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .ZN(n16150) );
  NOR2_X1 U17892 ( .A1(n21152), .A2(n16150), .ZN(n14552) );
  AOI21_X1 U17893 ( .B1(n14552), .B2(n14524), .A(n14558), .ZN(n16152) );
  NOR3_X1 U17894 ( .A1(n21152), .A2(n16150), .A3(n20279), .ZN(n16138) );
  INV_X1 U17895 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n16284) );
  AOI22_X1 U17896 ( .A1(n16279), .A2(n20345), .B1(n20344), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14525) );
  OAI211_X1 U17897 ( .C1(n20342), .C2(n14526), .A(n14525), .B(n20447), .ZN(
        n14527) );
  AOI221_X1 U17898 ( .B1(n16152), .B2(P1_REIP_REG_13__SCAN_IN), .C1(n16138), 
        .C2(n16284), .A(n14527), .ZN(n14528) );
  OAI211_X1 U17899 ( .C1(n14994), .C2(n20333), .A(n14529), .B(n14528), .ZN(
        P1_U2827) );
  INV_X1 U17900 ( .A(DATAI_13_), .ZN(n14531) );
  MUX2_X1 U17901 ( .A(n14531), .B(n14530), .S(n20497), .Z(n20406) );
  INV_X1 U17902 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14532) );
  OAI222_X1 U17903 ( .A1(n14533), .A2(n14839), .B1(n20406), .B2(n14838), .C1(
        n14532), .C2(n14836), .ZN(P1_U2891) );
  NOR2_X1 U17904 ( .A1(n19109), .A2(n19099), .ZN(n19012) );
  NAND2_X1 U17905 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19012), .ZN(n19101) );
  AOI21_X1 U17906 ( .B1(n18957), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15982) );
  AND2_X1 U17907 ( .A1(n9911), .A2(n15982), .ZN(n18494) );
  INV_X1 U17908 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16815) );
  OAI221_X1 U17909 ( .B1(n19101), .B2(n18494), .C1(n19101), .C2(n16815), .A(
        n18541), .ZN(n18501) );
  INV_X1 U17910 ( .A(n18501), .ZN(n18496) );
  INV_X1 U17911 ( .A(n15966), .ZN(n19148) );
  NOR2_X1 U17912 ( .A1(n19109), .A2(n19151), .ZN(n19013) );
  INV_X1 U17913 ( .A(n19013), .ZN(n17984) );
  AOI22_X1 U17914 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n19148), .B2(n17984), .ZN(n15969) );
  NOR2_X1 U17915 ( .A1(n18496), .A2(n15969), .ZN(n14535) );
  INV_X1 U17916 ( .A(n18847), .ZN(n18795) );
  NAND2_X1 U17917 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18968), .ZN(n18549) );
  NAND2_X1 U17918 ( .A1(n18549), .A2(n18501), .ZN(n15967) );
  OR2_X1 U17919 ( .A1(n18795), .A2(n15967), .ZN(n14534) );
  MUX2_X1 U17920 ( .A(n14535), .B(n14534), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17921 ( .A(n20347), .ZN(n20331) );
  INV_X1 U17922 ( .A(n14536), .ZN(n14537) );
  NAND2_X1 U17923 ( .A1(n14537), .A2(n20357), .ZN(n14544) );
  NAND2_X1 U17924 ( .A1(n20345), .A2(n14538), .ZN(n14540) );
  INV_X1 U17925 ( .A(n16076), .ZN(n14698) );
  AOI22_X1 U17926 ( .A1(n20351), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14698), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14539) );
  OAI211_X1 U17927 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20333), .A(
        n14540), .B(n14539), .ZN(n14542) );
  OAI22_X1 U17928 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n14676), .B1(n20330), 
        .B2(n11450), .ZN(n14541) );
  NOR2_X1 U17929 ( .A1(n14542), .A2(n14541), .ZN(n14543) );
  OAI211_X1 U17930 ( .C1(n20331), .C2(n14077), .A(n14544), .B(n14543), .ZN(
        P1_U2839) );
  NOR2_X1 U17931 ( .A1(n14545), .A2(n15273), .ZN(n14546) );
  AOI21_X1 U17932 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15273), .A(n14546), .ZN(
        n14547) );
  OAI21_X1 U17933 ( .B1(n14548), .B2(n15289), .A(n14547), .ZN(P2_U2857) );
  NAND2_X1 U17934 ( .A1(n14549), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14551)
         );
  NAND3_X1 U17935 ( .A1(n14551), .A2(n14550), .A3(n20254), .ZN(P1_U2801) );
  NAND2_X1 U17936 ( .A1(n14845), .A2(n20307), .ZN(n14565) );
  AND2_X1 U17937 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14557) );
  INV_X1 U17938 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14872) );
  INV_X1 U17939 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14885) );
  INV_X1 U17940 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n16091) );
  NAND2_X1 U17941 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14694) );
  INV_X1 U17942 ( .A(n14694), .ZN(n14691) );
  INV_X1 U17943 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21158) );
  INV_X1 U17944 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n14695) );
  NOR2_X1 U17945 ( .A1(n21158), .A2(n14695), .ZN(n16120) );
  NAND4_X1 U17946 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14552), .A3(n14691), 
        .A4(n16120), .ZN(n14673) );
  NOR2_X1 U17947 ( .A1(n14553), .A2(n14673), .ZN(n14675) );
  NAND4_X1 U17948 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14675), .A3(
        P1_REIP_REG_19__SCAN_IN), .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n16087) );
  NOR2_X1 U17949 ( .A1(n16091), .A2(n16087), .ZN(n14636) );
  AND2_X1 U17950 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n14636), .ZN(n14554) );
  NAND4_X1 U17951 ( .A1(n14554), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .A4(P1_REIP_REG_23__SCAN_IN), .ZN(n14560) );
  INV_X1 U17952 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14896) );
  NOR2_X1 U17953 ( .A1(n14560), .A2(n14896), .ZN(n14555) );
  NAND2_X1 U17954 ( .A1(n16076), .A2(n14555), .ZN(n14612) );
  OR3_X1 U17955 ( .A1(n14872), .A2(n14885), .A3(n14612), .ZN(n14556) );
  NAND2_X1 U17956 ( .A1(n20324), .A2(n14556), .ZN(n14596) );
  OAI21_X1 U17957 ( .B1(n14558), .B2(n14557), .A(n14596), .ZN(n14572) );
  INV_X1 U17958 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14559) );
  OAI22_X1 U17959 ( .A1(n14559), .A2(n20342), .B1(n20330), .B2(n14709), .ZN(
        n14563) );
  NOR2_X1 U17960 ( .A1(n14676), .A2(n14560), .ZN(n14627) );
  NAND3_X1 U17961 ( .A1(n14627), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_26__SCAN_IN), .ZN(n14599) );
  NOR2_X1 U17962 ( .A1(n14599), .A2(n14872), .ZN(n14586) );
  INV_X1 U17963 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14561) );
  AND4_X1 U17964 ( .A1(n14586), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .A4(n14561), .ZN(n14562) );
  AOI211_X1 U17965 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14572), .A(n14563), 
        .B(n14562), .ZN(n14564) );
  OAI211_X1 U17966 ( .C1(n14710), .C2(n20301), .A(n14565), .B(n14564), .ZN(
        P1_U2809) );
  XOR2_X1 U17967 ( .A(n14566), .B(n14580), .Z(n14855) );
  INV_X1 U17968 ( .A(n14855), .ZN(n14776) );
  NAND2_X1 U17969 ( .A1(n14587), .A2(n11476), .ZN(n14569) );
  OR2_X1 U17970 ( .A1(n14602), .A2(n14567), .ZN(n14568) );
  NAND2_X1 U17971 ( .A1(n14569), .A2(n14568), .ZN(n14571) );
  XNOR2_X1 U17972 ( .A(n14571), .B(n14570), .ZN(n15013) );
  AOI21_X1 U17973 ( .B1(n14586), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14576) );
  INV_X1 U17974 ( .A(n14572), .ZN(n14575) );
  AOI22_X1 U17975 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20351), .B1(
        n20350), .B2(n14851), .ZN(n14574) );
  NAND2_X1 U17976 ( .A1(n20344), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14573) );
  OAI211_X1 U17977 ( .C1(n14576), .C2(n14575), .A(n14574), .B(n14573), .ZN(
        n14577) );
  AOI21_X1 U17978 ( .B1(n15013), .B2(n20345), .A(n14577), .ZN(n14578) );
  OAI21_X1 U17979 ( .B1(n14776), .B2(n20294), .A(n14578), .ZN(P1_U2810) );
  AOI21_X1 U17980 ( .B1(n14581), .B2(n14579), .A(n14580), .ZN(n14863) );
  INV_X1 U17981 ( .A(n14863), .ZN(n14781) );
  INV_X1 U17982 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U17983 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20351), .B1(
        n20350), .B2(n14859), .ZN(n14583) );
  NAND2_X1 U17984 ( .A1(n20344), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14582) );
  OAI211_X1 U17985 ( .C1(n14596), .C2(n14585), .A(n14583), .B(n14582), .ZN(
        n14584) );
  AOI21_X1 U17986 ( .B1(n14586), .B2(n14585), .A(n14584), .ZN(n14591) );
  INV_X1 U17987 ( .A(n14587), .ZN(n14588) );
  AOI21_X1 U17988 ( .B1(n14589), .B2(n14602), .A(n14588), .ZN(n15022) );
  NAND2_X1 U17989 ( .A1(n15022), .A2(n20345), .ZN(n14590) );
  OAI211_X1 U17990 ( .C1(n14781), .C2(n20294), .A(n14591), .B(n14590), .ZN(
        P1_U2811) );
  INV_X1 U17991 ( .A(n14579), .ZN(n14594) );
  INV_X1 U17992 ( .A(n14871), .ZN(n14785) );
  INV_X1 U17993 ( .A(n14596), .ZN(n14605) );
  AOI22_X1 U17994 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20351), .B1(
        n20350), .B2(n14875), .ZN(n14598) );
  NAND2_X1 U17995 ( .A1(n20344), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14597) );
  OAI211_X1 U17996 ( .C1(n14599), .C2(P1_REIP_REG_28__SCAN_IN), .A(n14598), 
        .B(n14597), .ZN(n14604) );
  OR2_X1 U17997 ( .A1(n14611), .A2(n14600), .ZN(n14601) );
  NAND2_X1 U17998 ( .A1(n14602), .A2(n14601), .ZN(n15033) );
  NOR2_X1 U17999 ( .A1(n15033), .A2(n20301), .ZN(n14603) );
  AOI211_X1 U18000 ( .C1(n14605), .C2(P1_REIP_REG_28__SCAN_IN), .A(n14604), 
        .B(n14603), .ZN(n14606) );
  OAI21_X1 U18001 ( .B1(n14785), .B2(n20294), .A(n14606), .ZN(P1_U2812) );
  OAI21_X1 U18002 ( .B1(n14607), .B2(n14608), .A(n14593), .ZN(n14883) );
  AND2_X1 U18003 ( .A1(n14624), .A2(n14609), .ZN(n14610) );
  OR2_X1 U18004 ( .A1(n14611), .A2(n14610), .ZN(n14714) );
  INV_X1 U18005 ( .A(n14714), .ZN(n15041) );
  NAND2_X1 U18006 ( .A1(n20324), .A2(n14612), .ZN(n14625) );
  OAI22_X1 U18007 ( .A1(n14886), .A2(n20342), .B1(n20333), .B2(n14884), .ZN(
        n14613) );
  AOI21_X1 U18008 ( .B1(n20344), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14613), .ZN(
        n14615) );
  NAND3_X1 U18009 ( .A1(n14627), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n14885), 
        .ZN(n14614) );
  OAI211_X1 U18010 ( .C1(n14625), .C2(n14885), .A(n14615), .B(n14614), .ZN(
        n14616) );
  AOI21_X1 U18011 ( .B1(n15041), .B2(n20345), .A(n14616), .ZN(n14617) );
  OAI21_X1 U18012 ( .B1(n14883), .B2(n20294), .A(n14617), .ZN(P1_U2813) );
  INV_X1 U18013 ( .A(n14618), .ZN(n14619) );
  INV_X1 U18014 ( .A(n14607), .ZN(n14620) );
  OR2_X1 U18015 ( .A1(n14640), .A2(n14622), .ZN(n14623) );
  NAND2_X1 U18016 ( .A1(n14624), .A2(n14623), .ZN(n15051) );
  INV_X1 U18017 ( .A(n15051), .ZN(n14631) );
  INV_X1 U18018 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14716) );
  INV_X1 U18019 ( .A(n14625), .ZN(n14626) );
  OAI21_X1 U18020 ( .B1(n14627), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14626), 
        .ZN(n14629) );
  AOI22_X1 U18021 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20351), .B1(
        n20350), .B2(n14900), .ZN(n14628) );
  OAI211_X1 U18022 ( .C1(n14716), .C2(n20330), .A(n14629), .B(n14628), .ZN(
        n14630) );
  AOI21_X1 U18023 ( .B1(n14631), .B2(n20345), .A(n14630), .ZN(n14632) );
  OAI21_X1 U18024 ( .B1(n14898), .B2(n20294), .A(n14632), .ZN(P1_U2814) );
  INV_X1 U18025 ( .A(n14633), .ZN(n14634) );
  AOI21_X1 U18026 ( .B1(n9974), .B2(n14634), .A(n14619), .ZN(n14910) );
  INV_X1 U18027 ( .A(n14910), .ZN(n14796) );
  AND2_X1 U18028 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14654) );
  NAND3_X1 U18029 ( .A1(n16076), .A2(n14636), .A3(n14654), .ZN(n14635) );
  NAND2_X1 U18030 ( .A1(n20324), .A2(n14635), .ZN(n14668) );
  OAI21_X1 U18031 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n14676), .A(n14668), 
        .ZN(n14645) );
  INV_X1 U18032 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14906) );
  NAND4_X1 U18033 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .A4(n14906), .ZN(n14639) );
  NAND2_X1 U18034 ( .A1(n16078), .A2(n14636), .ZN(n16080) );
  OAI22_X1 U18035 ( .A1(n14907), .A2(n20342), .B1(n20333), .B2(n14905), .ZN(
        n14637) );
  AOI21_X1 U18036 ( .B1(n20344), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14637), .ZN(
        n14638) );
  OAI21_X1 U18037 ( .B1(n14639), .B2(n16080), .A(n14638), .ZN(n14644) );
  INV_X1 U18038 ( .A(n14640), .ZN(n14641) );
  OAI21_X1 U18039 ( .B1(n14642), .B2(n14651), .A(n14641), .ZN(n15058) );
  NOR2_X1 U18040 ( .A1(n15058), .A2(n20301), .ZN(n14643) );
  AOI211_X1 U18041 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14645), .A(n14644), 
        .B(n14643), .ZN(n14646) );
  OAI21_X1 U18042 ( .B1(n14796), .B2(n20294), .A(n14646), .ZN(P1_U2815) );
  AOI21_X1 U18043 ( .B1(n14648), .B2(n14647), .A(n14633), .ZN(n14920) );
  INV_X1 U18044 ( .A(n14920), .ZN(n14800) );
  AND2_X1 U18045 ( .A1(n14662), .A2(n14649), .ZN(n14650) );
  NOR2_X1 U18046 ( .A1(n14651), .A2(n14650), .ZN(n14718) );
  INV_X1 U18047 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21169) );
  INV_X1 U18048 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14918) );
  INV_X1 U18049 ( .A(n14916), .ZN(n14652) );
  OAI22_X1 U18050 ( .A1(n14918), .A2(n20342), .B1(n20333), .B2(n14652), .ZN(
        n14653) );
  AOI21_X1 U18051 ( .B1(n20344), .B2(P1_EBX_REG_24__SCAN_IN), .A(n14653), .ZN(
        n14656) );
  INV_X1 U18052 ( .A(n16080), .ZN(n14665) );
  NAND3_X1 U18053 ( .A1(n14665), .A2(n14654), .A3(n21169), .ZN(n14655) );
  OAI211_X1 U18054 ( .C1(n14668), .C2(n21169), .A(n14656), .B(n14655), .ZN(
        n14657) );
  AOI21_X1 U18055 ( .B1(n14718), .B2(n20345), .A(n14657), .ZN(n14658) );
  OAI21_X1 U18056 ( .B1(n14800), .B2(n20294), .A(n14658), .ZN(P1_U2816) );
  AOI21_X1 U18057 ( .B1(n14661), .B2(n14660), .A(n10193), .ZN(n14929) );
  INV_X1 U18058 ( .A(n14929), .ZN(n14808) );
  INV_X1 U18059 ( .A(n14662), .ZN(n14663) );
  AOI21_X1 U18060 ( .B1(n14728), .B2(n14664), .A(n14663), .ZN(n15080) );
  AOI21_X1 U18061 ( .B1(n14665), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n14669) );
  OAI22_X1 U18062 ( .A1(n14926), .A2(n20342), .B1(n20333), .B2(n14924), .ZN(
        n14666) );
  AOI21_X1 U18063 ( .B1(n20344), .B2(P1_EBX_REG_23__SCAN_IN), .A(n14666), .ZN(
        n14667) );
  OAI21_X1 U18064 ( .B1(n14669), .B2(n14668), .A(n14667), .ZN(n14670) );
  AOI21_X1 U18065 ( .B1(n15080), .B2(n20345), .A(n14670), .ZN(n14671) );
  OAI21_X1 U18066 ( .B1(n14808), .B2(n20294), .A(n14671), .ZN(P1_U2817) );
  OAI21_X1 U18067 ( .B1(n9883), .B2(n10378), .A(n14672), .ZN(n14961) );
  NOR2_X1 U18068 ( .A1(n14673), .A2(n20279), .ZN(n16112) );
  INV_X1 U18069 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21160) );
  INV_X1 U18070 ( .A(n14674), .ZN(n14745) );
  XNOR2_X1 U18071 ( .A(n9908), .B(n14745), .ZN(n16245) );
  OAI21_X1 U18072 ( .B1(n14676), .B2(n14675), .A(n16076), .ZN(n16119) );
  OAI21_X1 U18073 ( .B1(n20342), .B2(n14956), .A(n20447), .ZN(n14678) );
  NOR2_X1 U18074 ( .A1(n20330), .A2(n14750), .ZN(n14677) );
  AOI211_X1 U18075 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n16119), .A(n14678), 
        .B(n14677), .ZN(n14680) );
  NAND2_X1 U18076 ( .A1(n14958), .A2(n20350), .ZN(n14679) );
  OAI211_X1 U18077 ( .C1(n16245), .C2(n20301), .A(n14680), .B(n14679), .ZN(
        n14681) );
  AOI21_X1 U18078 ( .B1(n16112), .B2(n21160), .A(n14681), .ZN(n14682) );
  OAI21_X1 U18079 ( .B1(n14961), .B2(n20294), .A(n14682), .ZN(P1_U2822) );
  INV_X1 U18080 ( .A(n14683), .ZN(n14684) );
  AOI21_X1 U18081 ( .B1(n14685), .B2(n14500), .A(n14684), .ZN(n16182) );
  INV_X1 U18082 ( .A(n16182), .ZN(n14840) );
  NOR2_X1 U18083 ( .A1(n14687), .A2(n14686), .ZN(n14688) );
  OR2_X1 U18084 ( .A1(n14762), .A2(n14688), .ZN(n14769) );
  INV_X1 U18085 ( .A(n14769), .ZN(n15117) );
  AOI22_X1 U18086 ( .A1(n15117), .A2(n20345), .B1(n20344), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14689) );
  OAI211_X1 U18087 ( .C1(n20342), .C2(n14690), .A(n14689), .B(n20447), .ZN(
        n14693) );
  AND2_X1 U18088 ( .A1(n14691), .A2(n16138), .ZN(n16135) );
  NAND2_X1 U18089 ( .A1(n16135), .A2(n14695), .ZN(n16125) );
  INV_X1 U18090 ( .A(n16125), .ZN(n14692) );
  AOI211_X1 U18091 ( .C1(n16181), .C2(n20350), .A(n14693), .B(n14692), .ZN(
        n14697) );
  AOI21_X1 U18092 ( .B1(n14694), .B2(n20324), .A(n16152), .ZN(n16146) );
  OR2_X1 U18093 ( .A1(n16146), .A2(n14695), .ZN(n14696) );
  OAI211_X1 U18094 ( .C1(n14840), .C2(n20294), .A(n14697), .B(n14696), .ZN(
        P1_U2825) );
  INV_X1 U18095 ( .A(n13832), .ZN(n20507) );
  OAI21_X1 U18096 ( .B1(n14698), .B2(n20273), .A(n20324), .ZN(n20361) );
  INV_X1 U18097 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n14699) );
  NOR2_X1 U18098 ( .A1(n20361), .A2(n14699), .ZN(n14706) );
  NAND2_X1 U18099 ( .A1(n16078), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20354) );
  INV_X1 U18100 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14700) );
  OAI22_X1 U18101 ( .A1(n14701), .A2(n20333), .B1(n20342), .B2(n14700), .ZN(
        n14703) );
  NOR2_X1 U18102 ( .A1(n20301), .A2(n20465), .ZN(n14702) );
  AOI211_X1 U18103 ( .C1(n20344), .C2(P1_EBX_REG_2__SCAN_IN), .A(n14703), .B(
        n14702), .ZN(n14704) );
  OAI21_X1 U18104 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n20354), .A(n14704), .ZN(
        n14705) );
  AOI211_X1 U18105 ( .C1(n20347), .C2(n20507), .A(n14706), .B(n14705), .ZN(
        n14707) );
  OAI21_X1 U18106 ( .B1(n14708), .B2(n20335), .A(n14707), .ZN(P1_U2838) );
  OAI22_X1 U18107 ( .A1(n14710), .A2(n14768), .B1(n14770), .B2(n14709), .ZN(
        P1_U2841) );
  AOI22_X1 U18108 ( .A1(n15013), .A2(n14721), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14720), .ZN(n14711) );
  OAI21_X1 U18109 ( .B1(n14776), .B2(n14767), .A(n14711), .ZN(P1_U2842) );
  AOI22_X1 U18110 ( .A1(n15022), .A2(n14721), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14720), .ZN(n14712) );
  OAI21_X1 U18111 ( .B1(n14781), .B2(n14767), .A(n14712), .ZN(P1_U2843) );
  INV_X1 U18112 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14713) );
  OAI222_X1 U18113 ( .A1(n14767), .A2(n14785), .B1(n14713), .B2(n14770), .C1(
        n15033), .C2(n14768), .ZN(P1_U2844) );
  INV_X1 U18114 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14715) );
  OAI222_X1 U18115 ( .A1(n14767), .A2(n14883), .B1(n14715), .B2(n14770), .C1(
        n14714), .C2(n14768), .ZN(P1_U2845) );
  OAI222_X1 U18116 ( .A1(n14767), .A2(n14898), .B1(n14716), .B2(n14770), .C1(
        n15051), .C2(n14768), .ZN(P1_U2846) );
  INV_X1 U18117 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14717) );
  OAI222_X1 U18118 ( .A1(n14767), .A2(n14796), .B1(n14717), .B2(n14770), .C1(
        n15058), .C2(n14768), .ZN(P1_U2847) );
  INV_X1 U18119 ( .A(n14718), .ZN(n15069) );
  OAI222_X1 U18120 ( .A1(n14767), .A2(n14800), .B1(n14719), .B2(n14770), .C1(
        n15069), .C2(n14768), .ZN(P1_U2848) );
  AOI22_X1 U18121 ( .A1(n15080), .A2(n14721), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14720), .ZN(n14722) );
  OAI21_X1 U18122 ( .B1(n14808), .B2(n14772), .A(n14722), .ZN(P1_U2849) );
  NAND2_X1 U18123 ( .A1(n14723), .A2(n14724), .ZN(n14725) );
  AND2_X1 U18124 ( .A1(n14660), .A2(n14725), .ZN(n16084) );
  INV_X1 U18125 ( .A(n16084), .ZN(n14812) );
  OR2_X1 U18126 ( .A1(n14735), .A2(n14726), .ZN(n14727) );
  NAND2_X1 U18127 ( .A1(n14728), .A2(n14727), .ZN(n16233) );
  OAI22_X1 U18128 ( .A1(n16233), .A2(n14768), .B1(n16079), .B2(n14770), .ZN(
        n14729) );
  INV_X1 U18129 ( .A(n14729), .ZN(n14730) );
  OAI21_X1 U18130 ( .B1(n14812), .B2(n14772), .A(n14730), .ZN(P1_U2850) );
  OAI21_X1 U18131 ( .B1(n14731), .B2(n14732), .A(n14723), .ZN(n14944) );
  INV_X1 U18132 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14737) );
  INV_X1 U18133 ( .A(n14746), .ZN(n14734) );
  AOI21_X1 U18134 ( .B1(n14734), .B2(n14741), .A(n14733), .ZN(n14736) );
  OR2_X1 U18135 ( .A1(n14736), .A2(n14735), .ZN(n16093) );
  OAI222_X1 U18136 ( .A1(n14767), .A2(n14944), .B1(n14737), .B2(n14770), .C1(
        n16093), .C2(n14768), .ZN(P1_U2851) );
  INV_X1 U18137 ( .A(n14731), .ZN(n14739) );
  OAI21_X1 U18138 ( .B1(n14740), .B2(n14738), .A(n14739), .ZN(n16102) );
  INV_X1 U18139 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14742) );
  XNOR2_X1 U18140 ( .A(n14746), .B(n14741), .ZN(n16104) );
  INV_X1 U18141 ( .A(n16104), .ZN(n15105) );
  OAI222_X1 U18142 ( .A1(n14767), .A2(n16102), .B1(n14742), .B2(n14770), .C1(
        n14768), .C2(n15105), .ZN(P1_U2852) );
  INV_X1 U18143 ( .A(n14743), .ZN(n14744) );
  OAI21_X1 U18144 ( .B1(n9908), .B2(n14745), .A(n14744), .ZN(n14747) );
  NAND2_X1 U18145 ( .A1(n14747), .A2(n14746), .ZN(n16243) );
  AND2_X1 U18146 ( .A1(n14672), .A2(n14748), .ZN(n14749) );
  OR2_X1 U18147 ( .A1(n14749), .A2(n14738), .ZN(n16108) );
  OAI222_X1 U18148 ( .A1(n16243), .A2(n14768), .B1(n14770), .B2(n11510), .C1(
        n16108), .C2(n14767), .ZN(P1_U2853) );
  OAI22_X1 U18149 ( .A1(n16245), .A2(n14768), .B1(n14750), .B2(n14770), .ZN(
        n14751) );
  INV_X1 U18150 ( .A(n14751), .ZN(n14752) );
  OAI21_X1 U18151 ( .B1(n14961), .B2(n14772), .A(n14752), .ZN(P1_U2854) );
  INV_X1 U18152 ( .A(n14753), .ZN(n14755) );
  AOI21_X1 U18153 ( .B1(n14755), .B2(n10213), .A(n9883), .ZN(n16178) );
  INV_X1 U18154 ( .A(n16178), .ZN(n14830) );
  INV_X1 U18155 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14758) );
  NAND2_X1 U18156 ( .A1(n9952), .A2(n14756), .ZN(n14757) );
  NAND2_X1 U18157 ( .A1(n9908), .A2(n14757), .ZN(n16254) );
  OAI222_X1 U18158 ( .A1(n14830), .A2(n14772), .B1(n14758), .B2(n14770), .C1(
        n16254), .C2(n14768), .ZN(P1_U2855) );
  AND2_X1 U18159 ( .A1(n14683), .A2(n14759), .ZN(n14760) );
  OR2_X1 U18160 ( .A1(n14760), .A2(n14754), .ZN(n16133) );
  OR2_X1 U18161 ( .A1(n14762), .A2(n14761), .ZN(n14763) );
  NAND2_X1 U18162 ( .A1(n9952), .A2(n14763), .ZN(n16261) );
  OAI22_X1 U18163 ( .A1(n16261), .A2(n14768), .B1(n14764), .B2(n14770), .ZN(
        n14765) );
  INV_X1 U18164 ( .A(n14765), .ZN(n14766) );
  OAI21_X1 U18165 ( .B1(n16133), .B2(n14767), .A(n14766), .ZN(P1_U2856) );
  INV_X1 U18166 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14771) );
  OAI222_X1 U18167 ( .A1(n14840), .A2(n14772), .B1(n14771), .B2(n14770), .C1(
        n14769), .C2(n14768), .ZN(P1_U2857) );
  INV_X1 U18168 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n20362) );
  OAI22_X1 U18169 ( .A1(n14831), .A2(n20409), .B1(n20362), .B2(n14836), .ZN(
        n14773) );
  AOI21_X1 U18170 ( .B1(n14833), .B2(BUF1_REG_30__SCAN_IN), .A(n14773), .ZN(
        n14775) );
  NAND2_X1 U18171 ( .A1(n11311), .A2(DATAI_30_), .ZN(n14774) );
  OAI211_X1 U18172 ( .C1(n14776), .C2(n14839), .A(n14775), .B(n14774), .ZN(
        P1_U2874) );
  INV_X1 U18173 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14777) );
  OAI22_X1 U18174 ( .A1(n14831), .A2(n20406), .B1(n14777), .B2(n14836), .ZN(
        n14778) );
  AOI21_X1 U18175 ( .B1(n14833), .B2(BUF1_REG_29__SCAN_IN), .A(n14778), .ZN(
        n14780) );
  NAND2_X1 U18176 ( .A1(n11311), .A2(DATAI_29_), .ZN(n14779) );
  OAI211_X1 U18177 ( .C1(n14781), .C2(n14839), .A(n14780), .B(n14779), .ZN(
        P1_U2875) );
  OAI22_X1 U18178 ( .A1(n14831), .A2(n20403), .B1(n13953), .B2(n14836), .ZN(
        n14782) );
  AOI21_X1 U18179 ( .B1(n14833), .B2(BUF1_REG_28__SCAN_IN), .A(n14782), .ZN(
        n14784) );
  NAND2_X1 U18180 ( .A1(n11311), .A2(DATAI_28_), .ZN(n14783) );
  OAI211_X1 U18181 ( .C1(n14785), .C2(n14839), .A(n14784), .B(n14783), .ZN(
        P1_U2876) );
  INV_X1 U18182 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16724) );
  INV_X1 U18183 ( .A(n14831), .ZN(n14803) );
  AOI22_X1 U18184 ( .A1(n14803), .A2(n20401), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n14801), .ZN(n14786) );
  OAI21_X1 U18185 ( .B1(n16724), .B2(n14805), .A(n14786), .ZN(n14787) );
  AOI21_X1 U18186 ( .B1(n11311), .B2(DATAI_27_), .A(n14787), .ZN(n14788) );
  OAI21_X1 U18187 ( .B1(n14883), .B2(n14839), .A(n14788), .ZN(P1_U2877) );
  INV_X1 U18188 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14789) );
  OAI22_X1 U18189 ( .A1(n14831), .A2(n20398), .B1(n14789), .B2(n14836), .ZN(
        n14790) );
  AOI21_X1 U18190 ( .B1(n14833), .B2(BUF1_REG_26__SCAN_IN), .A(n14790), .ZN(
        n14792) );
  NAND2_X1 U18191 ( .A1(n11311), .A2(DATAI_26_), .ZN(n14791) );
  OAI211_X1 U18192 ( .C1(n14898), .C2(n14839), .A(n14792), .B(n14791), .ZN(
        P1_U2878) );
  OAI22_X1 U18193 ( .A1(n14831), .A2(n20394), .B1(n13947), .B2(n14836), .ZN(
        n14793) );
  AOI21_X1 U18194 ( .B1(n14833), .B2(BUF1_REG_25__SCAN_IN), .A(n14793), .ZN(
        n14795) );
  NAND2_X1 U18195 ( .A1(n11311), .A2(DATAI_25_), .ZN(n14794) );
  OAI211_X1 U18196 ( .C1(n14796), .C2(n14839), .A(n14795), .B(n14794), .ZN(
        P1_U2879) );
  OAI22_X1 U18197 ( .A1(n14831), .A2(n20390), .B1(n13943), .B2(n14836), .ZN(
        n14797) );
  AOI21_X1 U18198 ( .B1(n14833), .B2(BUF1_REG_24__SCAN_IN), .A(n14797), .ZN(
        n14799) );
  NAND2_X1 U18199 ( .A1(n11311), .A2(DATAI_24_), .ZN(n14798) );
  OAI211_X1 U18200 ( .C1(n14800), .C2(n14839), .A(n14799), .B(n14798), .ZN(
        P1_U2880) );
  INV_X1 U18201 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16732) );
  AOI22_X1 U18202 ( .A1(n14803), .A2(n14802), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n14801), .ZN(n14804) );
  OAI21_X1 U18203 ( .B1(n14805), .B2(n16732), .A(n14804), .ZN(n14806) );
  AOI21_X1 U18204 ( .B1(n11311), .B2(DATAI_23_), .A(n14806), .ZN(n14807) );
  OAI21_X1 U18205 ( .B1(n14808), .B2(n14839), .A(n14807), .ZN(P1_U2881) );
  OAI22_X1 U18206 ( .A1(n14831), .A2(n20547), .B1(n13961), .B2(n14836), .ZN(
        n14809) );
  AOI21_X1 U18207 ( .B1(n14833), .B2(BUF1_REG_22__SCAN_IN), .A(n14809), .ZN(
        n14811) );
  NAND2_X1 U18208 ( .A1(n11311), .A2(DATAI_22_), .ZN(n14810) );
  OAI211_X1 U18209 ( .C1(n14812), .C2(n14839), .A(n14811), .B(n14810), .ZN(
        P1_U2882) );
  OAI22_X1 U18210 ( .A1(n14831), .A2(n20542), .B1(n21493), .B2(n14836), .ZN(
        n14813) );
  AOI21_X1 U18211 ( .B1(n14833), .B2(BUF1_REG_21__SCAN_IN), .A(n14813), .ZN(
        n14815) );
  NAND2_X1 U18212 ( .A1(n11311), .A2(DATAI_21_), .ZN(n14814) );
  OAI211_X1 U18213 ( .C1(n14944), .C2(n14839), .A(n14815), .B(n14814), .ZN(
        P1_U2883) );
  OAI22_X1 U18214 ( .A1(n14831), .A2(n20537), .B1(n14816), .B2(n14836), .ZN(
        n14817) );
  AOI21_X1 U18215 ( .B1(n14833), .B2(BUF1_REG_20__SCAN_IN), .A(n14817), .ZN(
        n14819) );
  NAND2_X1 U18216 ( .A1(n11311), .A2(DATAI_20_), .ZN(n14818) );
  OAI211_X1 U18217 ( .C1(n16102), .C2(n14839), .A(n14819), .B(n14818), .ZN(
        P1_U2884) );
  OAI22_X1 U18218 ( .A1(n14831), .A2(n20531), .B1(n13957), .B2(n14836), .ZN(
        n14820) );
  AOI21_X1 U18219 ( .B1(n14833), .B2(BUF1_REG_19__SCAN_IN), .A(n14820), .ZN(
        n14822) );
  NAND2_X1 U18220 ( .A1(n11311), .A2(DATAI_19_), .ZN(n14821) );
  OAI211_X1 U18221 ( .C1(n16108), .C2(n14839), .A(n14822), .B(n14821), .ZN(
        P1_U2885) );
  INV_X1 U18222 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14823) );
  OAI22_X1 U18223 ( .A1(n14831), .A2(n20526), .B1(n14823), .B2(n14836), .ZN(
        n14824) );
  AOI21_X1 U18224 ( .B1(n14833), .B2(BUF1_REG_18__SCAN_IN), .A(n14824), .ZN(
        n14826) );
  NAND2_X1 U18225 ( .A1(n11311), .A2(DATAI_18_), .ZN(n14825) );
  OAI211_X1 U18226 ( .C1(n14961), .C2(n14839), .A(n14826), .B(n14825), .ZN(
        P1_U2886) );
  OAI22_X1 U18227 ( .A1(n14831), .A2(n20520), .B1(n13951), .B2(n14836), .ZN(
        n14827) );
  AOI21_X1 U18228 ( .B1(n14833), .B2(BUF1_REG_17__SCAN_IN), .A(n14827), .ZN(
        n14829) );
  NAND2_X1 U18229 ( .A1(n11311), .A2(DATAI_17_), .ZN(n14828) );
  OAI211_X1 U18230 ( .C1(n14830), .C2(n14839), .A(n14829), .B(n14828), .ZN(
        P1_U2887) );
  OAI22_X1 U18231 ( .A1(n14831), .A2(n20510), .B1(n13949), .B2(n14836), .ZN(
        n14832) );
  AOI21_X1 U18232 ( .B1(n14833), .B2(BUF1_REG_16__SCAN_IN), .A(n14832), .ZN(
        n14835) );
  NAND2_X1 U18233 ( .A1(n11311), .A2(DATAI_16_), .ZN(n14834) );
  OAI211_X1 U18234 ( .C1(n16133), .C2(n14839), .A(n14835), .B(n14834), .ZN(
        P1_U2888) );
  OAI222_X1 U18235 ( .A1(n14840), .A2(n14839), .B1(n14838), .B2(n14837), .C1(
        n14836), .C2(n13979), .ZN(P1_U2889) );
  NAND2_X1 U18236 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14841) );
  OAI211_X1 U18237 ( .C1(n16219), .C2(n14843), .A(n14842), .B(n14841), .ZN(
        n14844) );
  OAI21_X1 U18238 ( .B1(n14847), .B2(n20258), .A(n14846), .ZN(P1_U2968) );
  NAND2_X1 U18239 ( .A1(n14849), .A2(n14848), .ZN(n14850) );
  XNOR2_X1 U18240 ( .A(n14850), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15018) );
  NAND2_X1 U18241 ( .A1(n16189), .A2(n14851), .ZN(n14852) );
  NAND2_X1 U18242 ( .A1(n20487), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15011) );
  OAI211_X1 U18243 ( .C1(n14853), .C2(n20432), .A(n14852), .B(n15011), .ZN(
        n14854) );
  AOI21_X1 U18244 ( .B1(n14855), .B2(n16214), .A(n14854), .ZN(n14856) );
  OAI21_X1 U18245 ( .B1(n15018), .B2(n20258), .A(n14856), .ZN(P1_U2969) );
  NAND2_X1 U18246 ( .A1(n16189), .A2(n14859), .ZN(n14860) );
  NAND2_X1 U18247 ( .A1(n20487), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15019) );
  OAI211_X1 U18248 ( .C1(n14861), .C2(n20432), .A(n14860), .B(n15019), .ZN(
        n14862) );
  AOI21_X1 U18249 ( .B1(n14863), .B2(n16214), .A(n14862), .ZN(n14864) );
  OAI21_X1 U18250 ( .B1(n15026), .B2(n20258), .A(n14864), .ZN(P1_U2970) );
  INV_X1 U18251 ( .A(n9832), .ZN(n14866) );
  NAND2_X1 U18252 ( .A1(n14999), .A2(n15048), .ZN(n14892) );
  NAND2_X1 U18253 ( .A1(n14892), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14865) );
  OAI22_X1 U18254 ( .A1(n14866), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n14865), .B2(n14923), .ZN(n14868) );
  MUX2_X1 U18255 ( .A(n14881), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15002), .Z(n14867) );
  NAND2_X1 U18256 ( .A1(n14868), .A2(n14867), .ZN(n14870) );
  XNOR2_X1 U18257 ( .A(n14870), .B(n14869), .ZN(n15037) );
  NAND2_X1 U18258 ( .A1(n14871), .A2(n16214), .ZN(n14877) );
  NOR2_X1 U18259 ( .A1(n20447), .A2(n14872), .ZN(n15027) );
  NOR2_X1 U18260 ( .A1(n20432), .A2(n14873), .ZN(n14874) );
  AOI211_X1 U18261 ( .C1(n16189), .C2(n14875), .A(n15027), .B(n14874), .ZN(
        n14876) );
  OAI211_X1 U18262 ( .C1(n15037), .C2(n20258), .A(n14877), .B(n14876), .ZN(
        P1_U2971) );
  INV_X1 U18263 ( .A(n14878), .ZN(n14879) );
  MUX2_X1 U18264 ( .A(n14880), .B(n14879), .S(n15002), .Z(n14882) );
  XNOR2_X1 U18265 ( .A(n14882), .B(n14881), .ZN(n15046) );
  INV_X1 U18266 ( .A(n14883), .ZN(n14889) );
  NOR2_X1 U18267 ( .A1(n16219), .A2(n14884), .ZN(n14888) );
  OR2_X1 U18268 ( .A1(n20447), .A2(n14885), .ZN(n15038) );
  OAI21_X1 U18269 ( .B1(n20432), .B2(n14886), .A(n15038), .ZN(n14887) );
  AOI211_X1 U18270 ( .C1(n14889), .C2(n16214), .A(n14888), .B(n14887), .ZN(
        n14890) );
  OAI21_X1 U18271 ( .B1(n20258), .B2(n15046), .A(n14890), .ZN(P1_U2972) );
  OAI211_X1 U18272 ( .C1(n9832), .C2(n14999), .A(n14891), .B(n14892), .ZN(
        n14895) );
  XNOR2_X1 U18273 ( .A(n14895), .B(n14894), .ZN(n15054) );
  INV_X1 U18274 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14897) );
  OR2_X1 U18275 ( .A1(n20447), .A2(n14896), .ZN(n15050) );
  OAI21_X1 U18276 ( .B1(n20432), .B2(n14897), .A(n15050), .ZN(n14899) );
  AND2_X1 U18277 ( .A1(n15002), .A2(n15076), .ZN(n14912) );
  NOR2_X1 U18278 ( .A1(n14923), .A2(n14912), .ZN(n14901) );
  MUX2_X1 U18279 ( .A(n16194), .B(n14901), .S(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n14903) );
  NAND2_X1 U18280 ( .A1(n14902), .A2(n16194), .ZN(n14914) );
  NAND2_X1 U18281 ( .A1(n14903), .A2(n14914), .ZN(n14904) );
  XNOR2_X1 U18282 ( .A(n14904), .B(n15055), .ZN(n15062) );
  NOR2_X1 U18283 ( .A1(n16219), .A2(n14905), .ZN(n14909) );
  OR2_X1 U18284 ( .A1(n20447), .A2(n14906), .ZN(n15057) );
  OAI21_X1 U18285 ( .B1(n20432), .B2(n14907), .A(n15057), .ZN(n14908) );
  AOI211_X1 U18286 ( .C1(n14910), .C2(n16214), .A(n14909), .B(n14908), .ZN(
        n14911) );
  OAI21_X1 U18287 ( .B1(n20258), .B2(n15062), .A(n14911), .ZN(P1_U2974) );
  INV_X1 U18288 ( .A(n14912), .ZN(n14913) );
  NAND3_X1 U18289 ( .A1(n14914), .A2(n14891), .A3(n14913), .ZN(n14915) );
  XNOR2_X1 U18290 ( .A(n14915), .B(n15065), .ZN(n15073) );
  NAND2_X1 U18291 ( .A1(n16189), .A2(n14916), .ZN(n14917) );
  NAND2_X1 U18292 ( .A1(n20487), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15068) );
  OAI211_X1 U18293 ( .C1(n20432), .C2(n14918), .A(n14917), .B(n15068), .ZN(
        n14919) );
  AOI21_X1 U18294 ( .B1(n14920), .B2(n16214), .A(n14919), .ZN(n14921) );
  OAI21_X1 U18295 ( .B1(n20258), .B2(n15073), .A(n14921), .ZN(P1_U2975) );
  XNOR2_X1 U18296 ( .A(n15002), .B(n15076), .ZN(n14922) );
  XNOR2_X1 U18297 ( .A(n14923), .B(n14922), .ZN(n15082) );
  NOR2_X1 U18298 ( .A1(n16219), .A2(n14924), .ZN(n14928) );
  INV_X1 U18299 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14925) );
  OR2_X1 U18300 ( .A1(n20447), .A2(n14925), .ZN(n15074) );
  OAI21_X1 U18301 ( .B1(n20432), .B2(n14926), .A(n15074), .ZN(n14927) );
  AOI211_X1 U18302 ( .C1(n14929), .C2(n16214), .A(n14928), .B(n14927), .ZN(
        n14930) );
  OAI21_X1 U18303 ( .B1(n20258), .B2(n15082), .A(n14930), .ZN(P1_U2976) );
  OAI21_X1 U18304 ( .B1(n14932), .B2(n14999), .A(n14931), .ZN(n14933) );
  XNOR2_X1 U18305 ( .A(n14933), .B(n16224), .ZN(n16228) );
  NAND2_X1 U18306 ( .A1(n16084), .A2(n16214), .ZN(n14938) );
  INV_X1 U18307 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14934) );
  OAI22_X1 U18308 ( .A1(n20432), .A2(n14935), .B1(n20447), .B2(n14934), .ZN(
        n14936) );
  AOI21_X1 U18309 ( .B1(n16189), .B2(n16083), .A(n14936), .ZN(n14937) );
  OAI211_X1 U18310 ( .C1(n16228), .C2(n20258), .A(n14938), .B(n14937), .ZN(
        P1_U2977) );
  OAI21_X1 U18311 ( .B1(n15002), .B2(n16246), .A(n14939), .ZN(n16166) );
  NAND2_X1 U18312 ( .A1(n16194), .A2(n14940), .ZN(n16165) );
  NAND2_X1 U18313 ( .A1(n14999), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16164) );
  OAI22_X1 U18314 ( .A1(n16166), .A2(n16165), .B1(n14939), .B2(n16164), .ZN(
        n14950) );
  NAND2_X1 U18315 ( .A1(n14950), .A2(n14949), .ZN(n14948) );
  INV_X1 U18316 ( .A(n16164), .ZN(n14941) );
  NAND2_X1 U18317 ( .A1(n14941), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14942) );
  OAI22_X1 U18318 ( .A1(n14948), .A2(n15002), .B1(n14939), .B2(n14942), .ZN(
        n14943) );
  XNOR2_X1 U18319 ( .A(n14943), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15092) );
  INV_X1 U18320 ( .A(n14944), .ZN(n16095) );
  NAND2_X1 U18321 ( .A1(n20487), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U18322 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14945) );
  OAI211_X1 U18323 ( .C1(n16219), .C2(n16098), .A(n15088), .B(n14945), .ZN(
        n14946) );
  AOI21_X1 U18324 ( .B1(n16095), .B2(n16214), .A(n14946), .ZN(n14947) );
  OAI21_X1 U18325 ( .B1(n15092), .B2(n20258), .A(n14947), .ZN(P1_U2978) );
  OAI21_X1 U18326 ( .B1(n14950), .B2(n14949), .A(n14948), .ZN(n15093) );
  NAND2_X1 U18327 ( .A1(n15093), .A2(n20435), .ZN(n14953) );
  AND2_X1 U18328 ( .A1(n20487), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15102) );
  INV_X1 U18329 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16107) );
  NOR2_X1 U18330 ( .A1(n20432), .A2(n16107), .ZN(n14951) );
  AOI211_X1 U18331 ( .C1(n16189), .C2(n16099), .A(n15102), .B(n14951), .ZN(
        n14952) );
  OAI211_X1 U18332 ( .C1(n20496), .C2(n16102), .A(n14953), .B(n14952), .ZN(
        P1_U2979) );
  INV_X1 U18333 ( .A(n16244), .ZN(n14955) );
  NAND3_X1 U18334 ( .A1(n14955), .A2(n20435), .A3(n14939), .ZN(n14960) );
  OAI22_X1 U18335 ( .A1(n20432), .A2(n14956), .B1(n20447), .B2(n21160), .ZN(
        n14957) );
  AOI21_X1 U18336 ( .B1(n14958), .B2(n16189), .A(n14957), .ZN(n14959) );
  OAI211_X1 U18337 ( .C1(n20496), .C2(n14961), .A(n14960), .B(n14959), .ZN(
        P1_U2981) );
  NAND2_X1 U18338 ( .A1(n15114), .A2(n16262), .ZN(n16266) );
  NOR2_X1 U18339 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14962) );
  NOR2_X1 U18340 ( .A1(n14999), .A2(n14962), .ZN(n14963) );
  NOR2_X1 U18341 ( .A1(n14976), .A2(n14963), .ZN(n14964) );
  NAND2_X1 U18342 ( .A1(n14965), .A2(n14964), .ZN(n15108) );
  INV_X1 U18343 ( .A(n15107), .ZN(n14966) );
  OR2_X1 U18344 ( .A1(n15108), .A2(n14966), .ZN(n14968) );
  NAND2_X1 U18345 ( .A1(n16266), .A2(n14968), .ZN(n14970) );
  INV_X1 U18346 ( .A(n14967), .ZN(n14969) );
  OAI22_X1 U18347 ( .A1(n14970), .A2(n9950), .B1(n14969), .B2(n14968), .ZN(
        n16265) );
  NAND2_X1 U18348 ( .A1(n16265), .A2(n20435), .ZN(n14974) );
  OAI22_X1 U18349 ( .A1(n20432), .A2(n14971), .B1(n20447), .B2(n21158), .ZN(
        n14972) );
  AOI21_X1 U18350 ( .B1(n16126), .B2(n16189), .A(n14972), .ZN(n14973) );
  OAI211_X1 U18351 ( .C1(n20496), .C2(n16133), .A(n14974), .B(n14973), .ZN(
        P1_U2983) );
  NOR2_X1 U18352 ( .A1(n14988), .A2(n14976), .ZN(n14979) );
  OAI21_X1 U18353 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n14981) );
  XNOR2_X1 U18354 ( .A(n15002), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14980) );
  XNOR2_X1 U18355 ( .A(n14981), .B(n14980), .ZN(n16271) );
  AOI22_X1 U18356 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14982) );
  OAI21_X1 U18357 ( .B1(n16140), .B2(n16219), .A(n14982), .ZN(n14983) );
  AOI21_X1 U18358 ( .B1(n16142), .B2(n16214), .A(n14983), .ZN(n14984) );
  OAI21_X1 U18359 ( .B1(n16271), .B2(n20258), .A(n14984), .ZN(P1_U2985) );
  INV_X1 U18360 ( .A(n14985), .ZN(n14986) );
  AOI21_X1 U18361 ( .B1(n14988), .B2(n14987), .A(n14986), .ZN(n16188) );
  AND2_X1 U18362 ( .A1(n14989), .A2(n14990), .ZN(n16187) );
  NAND2_X1 U18363 ( .A1(n16188), .A2(n16187), .ZN(n16186) );
  NAND2_X1 U18364 ( .A1(n16186), .A2(n14990), .ZN(n14992) );
  XNOR2_X1 U18365 ( .A(n14992), .B(n14991), .ZN(n16278) );
  AOI22_X1 U18366 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14993) );
  OAI21_X1 U18367 ( .B1(n16219), .B2(n14994), .A(n14993), .ZN(n14995) );
  AOI21_X1 U18368 ( .B1(n14996), .B2(n16214), .A(n14995), .ZN(n14997) );
  OAI21_X1 U18369 ( .B1(n16278), .B2(n20258), .A(n14997), .ZN(P1_U2986) );
  NAND2_X1 U18370 ( .A1(n9831), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15001) );
  XNOR2_X1 U18371 ( .A(n14975), .B(n16325), .ZN(n15000) );
  MUX2_X1 U18372 ( .A(n15001), .B(n15000), .S(n14999), .Z(n15004) );
  NOR3_X1 U18373 ( .A1(n9831), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15002), .ZN(n16195) );
  INV_X1 U18374 ( .A(n16195), .ZN(n15003) );
  NAND2_X1 U18375 ( .A1(n15004), .A2(n15003), .ZN(n16323) );
  NAND2_X1 U18376 ( .A1(n16323), .A2(n20435), .ZN(n15009) );
  INV_X1 U18377 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15005) );
  OAI22_X1 U18378 ( .A1(n20432), .A2(n15005), .B1(n20447), .B2(n21150), .ZN(
        n15006) );
  AOI21_X1 U18379 ( .B1(n16189), .B2(n15007), .A(n15006), .ZN(n15008) );
  OAI211_X1 U18380 ( .C1(n20496), .C2(n15010), .A(n15009), .B(n15008), .ZN(
        P1_U2989) );
  INV_X1 U18381 ( .A(n15011), .ZN(n15012) );
  AOI21_X1 U18382 ( .B1(n15013), .B2(n20486), .A(n15012), .ZN(n15017) );
  OAI21_X1 U18383 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15015), .A(
        n15014), .ZN(n15016) );
  OAI211_X1 U18384 ( .C1(n15018), .C2(n20449), .A(n15017), .B(n15016), .ZN(
        P1_U3001) );
  INV_X1 U18385 ( .A(n15019), .ZN(n15021) );
  NOR3_X1 U18386 ( .A1(n15039), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15028), .ZN(n15020) );
  AOI211_X1 U18387 ( .C1(n15022), .C2(n20486), .A(n15021), .B(n15020), .ZN(
        n15025) );
  OR2_X1 U18388 ( .A1(n15023), .A2(n11414), .ZN(n15024) );
  OAI211_X1 U18389 ( .C1(n15026), .C2(n20449), .A(n15025), .B(n15024), .ZN(
        P1_U3002) );
  INV_X1 U18390 ( .A(n15027), .ZN(n15032) );
  INV_X1 U18391 ( .A(n15039), .ZN(n15030) );
  NAND3_X1 U18392 ( .A1(n15030), .A2(n15029), .A3(n15028), .ZN(n15031) );
  OAI211_X1 U18393 ( .C1(n15033), .C2(n20479), .A(n15032), .B(n15031), .ZN(
        n15034) );
  INV_X1 U18394 ( .A(n15034), .ZN(n15036) );
  NAND3_X1 U18395 ( .A1(n15043), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15042), .ZN(n15035) );
  OAI211_X1 U18396 ( .C1(n15037), .C2(n20449), .A(n15036), .B(n15035), .ZN(
        P1_U3003) );
  OAI21_X1 U18397 ( .B1(n15039), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15038), .ZN(n15040) );
  AOI21_X1 U18398 ( .B1(n15041), .B2(n20486), .A(n15040), .ZN(n15045) );
  NAND3_X1 U18399 ( .A1(n15043), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15042), .ZN(n15044) );
  OAI211_X1 U18400 ( .C1(n15046), .C2(n20449), .A(n15045), .B(n15044), .ZN(
        P1_U3004) );
  INV_X1 U18401 ( .A(n15047), .ZN(n15060) );
  OR3_X1 U18402 ( .A1(n15075), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15048), .ZN(n15049) );
  OAI211_X1 U18403 ( .C1(n15051), .C2(n20479), .A(n15050), .B(n15049), .ZN(
        n15052) );
  AOI21_X1 U18404 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15060), .A(
        n15052), .ZN(n15053) );
  OAI21_X1 U18405 ( .B1(n15054), .B2(n20449), .A(n15053), .ZN(P1_U3005) );
  INV_X1 U18406 ( .A(n15075), .ZN(n15066) );
  NAND4_X1 U18407 ( .A1(n15066), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n15055), .ZN(n15056) );
  OAI211_X1 U18408 ( .C1(n15058), .C2(n20479), .A(n15057), .B(n15056), .ZN(
        n15059) );
  AOI21_X1 U18409 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15060), .A(
        n15059), .ZN(n15061) );
  OAI21_X1 U18410 ( .B1(n15062), .B2(n20449), .A(n15061), .ZN(P1_U3006) );
  OAI21_X1 U18411 ( .B1(n15064), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15063), .ZN(n15071) );
  NAND3_X1 U18412 ( .A1(n15066), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15065), .ZN(n15067) );
  OAI211_X1 U18413 ( .C1(n15069), .C2(n20479), .A(n15068), .B(n15067), .ZN(
        n15070) );
  AOI21_X1 U18414 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15071), .A(
        n15070), .ZN(n15072) );
  OAI21_X1 U18415 ( .B1(n15073), .B2(n20449), .A(n15072), .ZN(P1_U3007) );
  OAI21_X1 U18416 ( .B1(n15075), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15074), .ZN(n15079) );
  NOR2_X1 U18417 ( .A1(n15077), .A2(n15076), .ZN(n15078) );
  AOI211_X1 U18418 ( .C1(n20486), .C2(n15080), .A(n15079), .B(n15078), .ZN(
        n15081) );
  OAI21_X1 U18419 ( .B1(n15082), .B2(n20449), .A(n15081), .ZN(P1_U3008) );
  NOR3_X1 U18420 ( .A1(n16282), .A2(n15083), .A3(n20473), .ZN(n15084) );
  NOR2_X1 U18421 ( .A1(n15084), .A2(n16234), .ZN(n16281) );
  NOR2_X1 U18422 ( .A1(n16281), .A2(n16235), .ZN(n15096) );
  NOR2_X1 U18423 ( .A1(n16283), .A2(n15085), .ZN(n15086) );
  OR2_X1 U18424 ( .A1(n15096), .A2(n15086), .ZN(n15094) );
  AND2_X1 U18425 ( .A1(n15094), .A2(n15087), .ZN(n16227) );
  NAND2_X1 U18426 ( .A1(n16227), .A2(n16225), .ZN(n15089) );
  OAI211_X1 U18427 ( .C1(n20479), .C2(n16093), .A(n15089), .B(n15088), .ZN(
        n15090) );
  AOI21_X1 U18428 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n16229), .A(
        n15090), .ZN(n15091) );
  OAI21_X1 U18429 ( .B1(n15092), .B2(n20449), .A(n15091), .ZN(P1_U3010) );
  NAND2_X1 U18430 ( .A1(n15093), .A2(n20489), .ZN(n15104) );
  INV_X1 U18431 ( .A(n15094), .ZN(n15095) );
  NOR3_X1 U18432 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14940), .A3(
        n15095), .ZN(n15101) );
  OAI21_X1 U18433 ( .B1(n15097), .B2(n15096), .A(n14940), .ZN(n15098) );
  INV_X1 U18434 ( .A(n15098), .ZN(n16238) );
  OAI21_X1 U18435 ( .B1(n16239), .B2(n16238), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15099) );
  INV_X1 U18436 ( .A(n15099), .ZN(n15100) );
  NOR3_X1 U18437 ( .A1(n15102), .A2(n15101), .A3(n15100), .ZN(n15103) );
  OAI211_X1 U18438 ( .C1(n15105), .C2(n20479), .A(n15104), .B(n15103), .ZN(
        P1_U3011) );
  NAND2_X1 U18439 ( .A1(n15107), .A2(n15106), .ZN(n15109) );
  XOR2_X1 U18440 ( .A(n15109), .B(n15108), .Z(n16185) );
  NAND2_X1 U18441 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16268), .ZN(
        n15115) );
  OAI21_X1 U18442 ( .B1(n16292), .B2(n15111), .A(n15110), .ZN(n16287) );
  AOI21_X1 U18443 ( .B1(n15112), .B2(n20474), .A(n16287), .ZN(n16263) );
  NAND2_X1 U18444 ( .A1(n20487), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15113) );
  OAI221_X1 U18445 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15115), 
        .C1(n15114), .C2(n16263), .A(n15113), .ZN(n15116) );
  AOI21_X1 U18446 ( .B1(n15117), .B2(n20486), .A(n15116), .ZN(n15118) );
  OAI21_X1 U18447 ( .B1(n16185), .B2(n20449), .A(n15118), .ZN(P1_U3016) );
  NAND2_X1 U18448 ( .A1(n9870), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21068) );
  XNOR2_X1 U18449 ( .A(n15120), .B(n21068), .ZN(n15121) );
  OAI22_X1 U18450 ( .A1(n15121), .A2(n21194), .B1(n13832), .B2(n21197), .ZN(
        n15122) );
  MUX2_X1 U18451 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15122), .S(
        n21212), .Z(P1_U3476) );
  INV_X1 U18452 ( .A(n14077), .ZN(n21016) );
  INV_X1 U18453 ( .A(n14064), .ZN(n15124) );
  INV_X1 U18454 ( .A(n13839), .ZN(n15123) );
  NAND3_X1 U18455 ( .A1(n15125), .A2(n15124), .A3(n15123), .ZN(n15126) );
  OAI21_X1 U18456 ( .B1(n16012), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n15126), .ZN(n15127) );
  AOI21_X1 U18457 ( .B1(n21016), .B2(n15128), .A(n15127), .ZN(n16013) );
  NOR3_X1 U18458 ( .A1(n14064), .A2(n13839), .A3(n15129), .ZN(n15130) );
  AOI21_X1 U18459 ( .B1(n15132), .B2(n15131), .A(n15130), .ZN(n15133) );
  OAI21_X1 U18460 ( .B1(n16013), .B2(n15134), .A(n15133), .ZN(n15135) );
  MUX2_X1 U18461 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15135), .S(
        n21192), .Z(P1_U3473) );
  NOR2_X1 U18462 ( .A1(n15137), .A2(n15136), .ZN(n15138) );
  OAI211_X1 U18463 ( .C1(n15140), .C2(n15412), .A(n20102), .B(n15139), .ZN(
        n15150) );
  INV_X1 U18464 ( .A(n15141), .ZN(n15148) );
  OAI22_X1 U18465 ( .A1(n12794), .A2(n19353), .B1(n20182), .B2(n19349), .ZN(
        n15147) );
  INV_X1 U18466 ( .A(n15142), .ZN(n15144) );
  INV_X1 U18467 ( .A(n12819), .ZN(n15143) );
  AOI21_X1 U18468 ( .B1(n15144), .B2(n15143), .A(n15301), .ZN(n15570) );
  INV_X1 U18469 ( .A(n15570), .ZN(n15145) );
  OAI22_X1 U18470 ( .A1(n15145), .A2(n19371), .B1(n13180), .B2(n19378), .ZN(
        n15146) );
  AOI211_X1 U18471 ( .C1(n15148), .C2(n19367), .A(n15147), .B(n15146), .ZN(
        n15149) );
  OAI211_X1 U18472 ( .C1(n19343), .C2(n15573), .A(n15150), .B(n15149), .ZN(
        P2_U2827) );
  OAI211_X1 U18473 ( .C1(n15485), .C2(n15152), .A(n20102), .B(n15151), .ZN(
        n15162) );
  OR2_X1 U18474 ( .A1(n15286), .A2(n15153), .ZN(n15154) );
  AND2_X1 U18475 ( .A1(n15271), .A2(n15154), .ZN(n15651) );
  NOR2_X1 U18476 ( .A1(n15366), .A2(n15156), .ZN(n15157) );
  OR2_X1 U18477 ( .A1(n15155), .A2(n15157), .ZN(n16470) );
  OAI22_X1 U18478 ( .A1(n19353), .A2(n12428), .B1(n16470), .B2(n19371), .ZN(
        n15160) );
  AOI22_X1 U18479 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19356), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19369), .ZN(n15158) );
  INV_X1 U18480 ( .A(n15158), .ZN(n15159) );
  AOI211_X1 U18481 ( .C1(n15651), .C2(n19364), .A(n15160), .B(n15159), .ZN(
        n15161) );
  OAI211_X1 U18482 ( .C1(n15163), .C2(n19351), .A(n15162), .B(n15161), .ZN(
        P2_U2835) );
  NOR2_X1 U18483 ( .A1(n19334), .A2(n9876), .ZN(n15198) );
  NAND2_X1 U18484 ( .A1(n9875), .A2(n20102), .ZN(n19383) );
  NOR2_X1 U18485 ( .A1(n19294), .A2(n19383), .ZN(n19301) );
  NAND2_X1 U18486 ( .A1(n16501), .A2(n15164), .ZN(n15165) );
  AOI22_X1 U18487 ( .A1(n16501), .A2(n15198), .B1(n19301), .B2(n15165), .ZN(
        n15176) );
  INV_X1 U18488 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20150) );
  OAI22_X1 U18489 ( .A1(n16508), .A2(n19378), .B1(n20150), .B2(n19349), .ZN(
        n15166) );
  AOI211_X1 U18490 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n19368), .A(n19247), .B(
        n15166), .ZN(n15175) );
  OR2_X1 U18491 ( .A1(n15168), .A2(n15167), .ZN(n15169) );
  NAND2_X1 U18492 ( .A1(n15169), .A2(n15761), .ZN(n19402) );
  INV_X1 U18493 ( .A(n19402), .ZN(n15170) );
  AOI22_X1 U18494 ( .A1(n19364), .A2(n16505), .B1(n19275), .B2(n15170), .ZN(
        n15174) );
  INV_X1 U18495 ( .A(n12280), .ZN(n15172) );
  NAND3_X1 U18496 ( .A1(n15172), .A2(n19367), .A3(n15171), .ZN(n15173) );
  NAND4_X1 U18497 ( .A1(n15176), .A2(n15175), .A3(n15174), .A4(n15173), .ZN(
        P2_U2844) );
  NAND2_X1 U18498 ( .A1(n9876), .A2(n15177), .ZN(n15178) );
  XNOR2_X1 U18499 ( .A(n16549), .B(n15178), .ZN(n15189) );
  NOR2_X1 U18500 ( .A1(n20202), .A2(n15179), .ZN(n15188) );
  XNOR2_X1 U18501 ( .A(n15181), .B(n15180), .ZN(n19429) );
  INV_X1 U18502 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20135) );
  OAI22_X1 U18503 ( .A1(n15182), .A2(n19353), .B1(n20135), .B2(n19349), .ZN(
        n15185) );
  OAI22_X1 U18504 ( .A1(n19351), .A2(n15183), .B1(n16562), .B2(n19378), .ZN(
        n15184) );
  AOI211_X1 U18505 ( .C1(n16601), .C2(n19364), .A(n15185), .B(n15184), .ZN(
        n15186) );
  OAI21_X1 U18506 ( .B1(n19429), .B2(n19371), .A(n15186), .ZN(n15187) );
  AOI211_X1 U18507 ( .C1(n15189), .C2(n20102), .A(n15188), .B(n15187), .ZN(
        n15190) );
  INV_X1 U18508 ( .A(n15190), .ZN(P2_U2852) );
  INV_X1 U18509 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20132) );
  OAI22_X1 U18510 ( .A1(n19351), .A2(n15191), .B1(n19349), .B2(n20132), .ZN(
        n15195) );
  OAI22_X1 U18511 ( .A1(n19353), .A2(n15193), .B1(n15192), .B2(n19378), .ZN(
        n15194) );
  AOI211_X1 U18512 ( .C1(n19275), .C2(n20223), .A(n15195), .B(n15194), .ZN(
        n15196) );
  OAI21_X1 U18513 ( .B1(n15197), .B2(n19343), .A(n15196), .ZN(n15202) );
  INV_X1 U18514 ( .A(n15198), .ZN(n19377) );
  OAI21_X1 U18515 ( .B1(n19384), .B2(n15200), .A(n15199), .ZN(n15832) );
  OAI22_X1 U18516 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19377), .B1(
        n15832), .B2(n19334), .ZN(n15201) );
  AOI211_X1 U18517 ( .C1(n20221), .C2(n19381), .A(n15202), .B(n15201), .ZN(
        n15203) );
  INV_X1 U18518 ( .A(n15203), .ZN(P2_U2854) );
  MUX2_X1 U18519 ( .A(n16380), .B(P2_EBX_REG_31__SCAN_IN), .S(n15273), .Z(
        P2_U2856) );
  OR2_X1 U18520 ( .A1(n15205), .A2(n15204), .ZN(n15206) );
  NAND2_X1 U18521 ( .A1(n15207), .A2(n15206), .ZN(n16391) );
  INV_X1 U18522 ( .A(n15208), .ZN(n15299) );
  NAND2_X1 U18523 ( .A1(n15209), .A2(n15210), .ZN(n15298) );
  NAND3_X1 U18524 ( .A1(n15299), .A2(n15294), .A3(n15298), .ZN(n15212) );
  NAND2_X1 U18525 ( .A1(n15273), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15211) );
  OAI211_X1 U18526 ( .C1(n15273), .C2(n16391), .A(n15212), .B(n15211), .ZN(
        P2_U2858) );
  NAND2_X1 U18527 ( .A1(n15213), .A2(n15214), .ZN(n15216) );
  XNOR2_X1 U18528 ( .A(n15216), .B(n15215), .ZN(n15313) );
  NOR2_X1 U18529 ( .A1(n15573), .A2(n13754), .ZN(n15217) );
  AOI21_X1 U18530 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15273), .A(n15217), .ZN(
        n15218) );
  OAI21_X1 U18531 ( .B1(n15313), .B2(n15289), .A(n15218), .ZN(P2_U2859) );
  AOI21_X1 U18532 ( .B1(n15219), .B2(n15221), .A(n15220), .ZN(n15222) );
  INV_X1 U18533 ( .A(n15222), .ZN(n15318) );
  NOR2_X1 U18534 ( .A1(n16403), .A2(n15273), .ZN(n15223) );
  AOI21_X1 U18535 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n13754), .A(n15223), .ZN(
        n15224) );
  OAI21_X1 U18536 ( .B1(n15318), .B2(n15289), .A(n15224), .ZN(P2_U2860) );
  AND2_X1 U18537 ( .A1(n9944), .A2(n15225), .ZN(n15227) );
  OR2_X1 U18538 ( .A1(n15227), .A2(n15226), .ZN(n16416) );
  AOI21_X1 U18539 ( .B1(n15228), .B2(n15230), .A(n15229), .ZN(n15326) );
  NAND2_X1 U18540 ( .A1(n15326), .A2(n15294), .ZN(n15232) );
  NAND2_X1 U18541 ( .A1(n13754), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15231) );
  OAI211_X1 U18542 ( .C1(n16416), .C2(n13754), .A(n15232), .B(n15231), .ZN(
        P2_U2861) );
  OAI21_X1 U18543 ( .B1(n15233), .B2(n15235), .A(n15234), .ZN(n15334) );
  NAND2_X1 U18544 ( .A1(n9893), .A2(n15236), .ZN(n15237) );
  NAND2_X1 U18545 ( .A1(n9944), .A2(n15237), .ZN(n16428) );
  MUX2_X1 U18546 ( .A(n16428), .B(n15238), .S(n15273), .Z(n15239) );
  OAI21_X1 U18547 ( .B1(n15334), .B2(n15289), .A(n15239), .ZN(P2_U2862) );
  CLKBUF_X1 U18548 ( .A(n15240), .Z(n15243) );
  AOI21_X1 U18549 ( .B1(n15243), .B2(n15242), .A(n15241), .ZN(n15244) );
  XOR2_X1 U18550 ( .A(n15245), .B(n15244), .Z(n15342) );
  NAND2_X1 U18551 ( .A1(n9951), .A2(n15246), .ZN(n15247) );
  NAND2_X1 U18552 ( .A1(n9893), .A2(n15247), .ZN(n16441) );
  NOR2_X1 U18553 ( .A1(n16441), .A2(n15273), .ZN(n15248) );
  AOI21_X1 U18554 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n13754), .A(n15248), .ZN(
        n15249) );
  OAI21_X1 U18555 ( .B1(n15342), .B2(n15289), .A(n15249), .ZN(P2_U2863) );
  INV_X1 U18556 ( .A(n15251), .ZN(n15252) );
  AOI21_X1 U18557 ( .B1(n15250), .B2(n15253), .A(n15252), .ZN(n15254) );
  INV_X1 U18558 ( .A(n15254), .ZN(n15352) );
  OR2_X1 U18559 ( .A1(n15259), .A2(n15255), .ZN(n15256) );
  NAND2_X1 U18560 ( .A1(n9951), .A2(n15256), .ZN(n16453) );
  MUX2_X1 U18561 ( .A(n16453), .B(n12438), .S(n15273), .Z(n15257) );
  OAI21_X1 U18562 ( .B1(n15352), .B2(n15289), .A(n15257), .ZN(P2_U2864) );
  AND2_X1 U18563 ( .A1(n9946), .A2(n15258), .ZN(n15260) );
  OR2_X1 U18564 ( .A1(n15260), .A2(n15259), .ZN(n16002) );
  INV_X1 U18565 ( .A(n15261), .ZN(n15263) );
  AOI21_X1 U18566 ( .B1(n15264), .B2(n15263), .A(n13453), .ZN(n16465) );
  NAND2_X1 U18567 ( .A1(n16465), .A2(n15294), .ZN(n15266) );
  NAND2_X1 U18568 ( .A1(n13754), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15265) );
  OAI211_X1 U18569 ( .C1(n16002), .C2(n15273), .A(n15266), .B(n15265), .ZN(
        P2_U2865) );
  INV_X1 U18570 ( .A(n15267), .ZN(n15278) );
  INV_X1 U18571 ( .A(n15268), .ZN(n15269) );
  OAI21_X1 U18572 ( .B1(n15278), .B2(n15269), .A(n15263), .ZN(n15363) );
  NAND2_X1 U18573 ( .A1(n13754), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15275) );
  NAND2_X1 U18574 ( .A1(n15271), .A2(n15270), .ZN(n15272) );
  NAND2_X1 U18575 ( .A1(n9946), .A2(n15272), .ZN(n19200) );
  OR2_X1 U18576 ( .A1(n19200), .A2(n15273), .ZN(n15274) );
  OAI211_X1 U18577 ( .C1(n15363), .C2(n15289), .A(n15275), .B(n15274), .ZN(
        P2_U2866) );
  INV_X1 U18578 ( .A(n15276), .ZN(n15279) );
  INV_X1 U18579 ( .A(n15277), .ZN(n15282) );
  AOI21_X1 U18580 ( .B1(n15279), .B2(n15282), .A(n15278), .ZN(n16472) );
  NAND2_X1 U18581 ( .A1(n16472), .A2(n15294), .ZN(n15281) );
  NAND2_X1 U18582 ( .A1(n15651), .A2(n13920), .ZN(n15280) );
  OAI211_X1 U18583 ( .C1(n13920), .C2(n12428), .A(n15281), .B(n15280), .ZN(
        P2_U2867) );
  OAI21_X1 U18584 ( .B1(n9894), .B2(n15283), .A(n15282), .ZN(n15372) );
  NOR2_X1 U18585 ( .A1(n9940), .A2(n15284), .ZN(n15285) );
  OR2_X1 U18586 ( .A1(n15286), .A2(n15285), .ZN(n19213) );
  NOR2_X1 U18587 ( .A1(n19213), .A2(n15273), .ZN(n15287) );
  AOI21_X1 U18588 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15273), .A(n15287), .ZN(
        n15288) );
  OAI21_X1 U18589 ( .B1(n15372), .B2(n15289), .A(n15288), .ZN(P2_U2868) );
  AND2_X1 U18590 ( .A1(n15291), .A2(n15290), .ZN(n15292) );
  NOR2_X1 U18591 ( .A1(n9940), .A2(n15292), .ZN(n19226) );
  INV_X1 U18592 ( .A(n19226), .ZN(n15297) );
  AOI21_X1 U18593 ( .B1(n15293), .B2(n9949), .A(n9894), .ZN(n16478) );
  NAND2_X1 U18594 ( .A1(n16478), .A2(n15294), .ZN(n15296) );
  NAND2_X1 U18595 ( .A1(n13754), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15295) );
  OAI211_X1 U18596 ( .C1(n15297), .C2(n13754), .A(n15296), .B(n15295), .ZN(
        P2_U2869) );
  NAND3_X1 U18597 ( .A1(n15299), .A2(n19444), .A3(n15298), .ZN(n15308) );
  OR2_X1 U18598 ( .A1(n15301), .A2(n15300), .ZN(n15302) );
  OAI22_X1 U18599 ( .A1(n15386), .A2(n19396), .B1(n19415), .B2(n15304), .ZN(
        n15305) );
  AOI21_X1 U18600 ( .B1(n19443), .B2(n16389), .A(n15305), .ZN(n15307) );
  AOI22_X1 U18601 ( .A1(n19385), .A2(BUF1_REG_29__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15306) );
  NAND3_X1 U18602 ( .A1(n15308), .A2(n15307), .A3(n15306), .ZN(P2_U2890) );
  INV_X1 U18603 ( .A(n19398), .ZN(n15309) );
  OAI22_X1 U18604 ( .A1(n15386), .A2(n15309), .B1(n19415), .B2(n21305), .ZN(
        n15310) );
  AOI21_X1 U18605 ( .B1(n19443), .B2(n15570), .A(n15310), .ZN(n15312) );
  AOI22_X1 U18606 ( .A1(n19385), .A2(BUF1_REG_28__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15311) );
  OAI211_X1 U18607 ( .C1(n15313), .C2(n19419), .A(n15312), .B(n15311), .ZN(
        P2_U2891) );
  OAI22_X1 U18608 ( .A1(n15386), .A2(n19401), .B1(n19415), .B2(n15314), .ZN(
        n15315) );
  AOI21_X1 U18609 ( .B1(n19443), .B2(n16404), .A(n15315), .ZN(n15317) );
  AOI22_X1 U18610 ( .A1(n19385), .A2(BUF1_REG_27__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15316) );
  OAI211_X1 U18611 ( .C1(n15318), .C2(n19419), .A(n15317), .B(n15316), .ZN(
        P2_U2892) );
  NAND2_X1 U18612 ( .A1(n15319), .A2(n15320), .ZN(n15321) );
  NAND2_X1 U18613 ( .A1(n9909), .A2(n15321), .ZN(n16415) );
  AOI22_X1 U18614 ( .A1(n19385), .A2(BUF1_REG_26__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15323) );
  INV_X1 U18615 ( .A(n15386), .ZN(n16477) );
  AOI22_X1 U18616 ( .A1(n16477), .A2(n19403), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19442), .ZN(n15322) );
  OAI211_X1 U18617 ( .C1(n15324), .C2(n16415), .A(n15323), .B(n15322), .ZN(
        n15325) );
  AOI21_X1 U18618 ( .B1(n15326), .B2(n19444), .A(n15325), .ZN(n15327) );
  INV_X1 U18619 ( .A(n15327), .ZN(P2_U2893) );
  OR2_X1 U18620 ( .A1(n15337), .A2(n15328), .ZN(n15329) );
  AND2_X1 U18621 ( .A1(n15319), .A2(n15329), .ZN(n16426) );
  OAI22_X1 U18622 ( .A1(n15386), .A2(n19406), .B1(n19415), .B2(n15330), .ZN(
        n15331) );
  AOI21_X1 U18623 ( .B1(n19443), .B2(n16426), .A(n15331), .ZN(n15333) );
  AOI22_X1 U18624 ( .A1(n19385), .A2(BUF1_REG_25__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15332) );
  OAI211_X1 U18625 ( .C1(n15334), .C2(n19419), .A(n15333), .B(n15332), .ZN(
        P2_U2894) );
  AND2_X1 U18626 ( .A1(n15345), .A2(n15335), .ZN(n15336) );
  NOR2_X1 U18627 ( .A1(n15337), .A2(n15336), .ZN(n16439) );
  INV_X1 U18628 ( .A(n19410), .ZN(n15338) );
  OAI22_X1 U18629 ( .A1(n15386), .A2(n15338), .B1(n19415), .B2(n13794), .ZN(
        n15339) );
  AOI21_X1 U18630 ( .B1(n19443), .B2(n16439), .A(n15339), .ZN(n15341) );
  AOI22_X1 U18631 ( .A1(n19385), .A2(BUF1_REG_24__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15340) );
  OAI211_X1 U18632 ( .C1(n15342), .C2(n19419), .A(n15341), .B(n15340), .ZN(
        P2_U2895) );
  NAND2_X1 U18633 ( .A1(n15630), .A2(n15343), .ZN(n15344) );
  NAND2_X1 U18634 ( .A1(n15345), .A2(n15344), .ZN(n16461) );
  INV_X1 U18635 ( .A(n16461), .ZN(n15350) );
  OAI22_X1 U18636 ( .A1(n15386), .A2(n19572), .B1(n19415), .B2(n15346), .ZN(
        n15349) );
  INV_X1 U18637 ( .A(n19385), .ZN(n15388) );
  INV_X1 U18638 ( .A(n19387), .ZN(n15387) );
  INV_X1 U18639 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15347) );
  OAI22_X1 U18640 ( .A1(n15388), .A2(n16732), .B1(n15387), .B2(n15347), .ZN(
        n15348) );
  AOI211_X1 U18641 ( .C1(n19443), .C2(n15350), .A(n15349), .B(n15348), .ZN(
        n15351) );
  OAI21_X1 U18642 ( .B1(n15352), .B2(n19419), .A(n15351), .ZN(P2_U2896) );
  OR2_X1 U18643 ( .A1(n15155), .A2(n15353), .ZN(n15355) );
  NAND2_X1 U18644 ( .A1(n15355), .A2(n15354), .ZN(n19208) );
  INV_X1 U18645 ( .A(n19208), .ZN(n15361) );
  OAI22_X1 U18646 ( .A1(n15386), .A2(n19553), .B1(n19415), .B2(n15356), .ZN(
        n15360) );
  INV_X1 U18647 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15358) );
  INV_X1 U18648 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15357) );
  OAI22_X1 U18649 ( .A1(n15388), .A2(n15358), .B1(n15387), .B2(n15357), .ZN(
        n15359) );
  AOI211_X1 U18650 ( .C1(n19443), .C2(n15361), .A(n15360), .B(n15359), .ZN(
        n15362) );
  OAI21_X1 U18651 ( .B1(n15363), .B2(n19419), .A(n15362), .ZN(P2_U2898) );
  NOR2_X1 U18652 ( .A1(n15364), .A2(n15681), .ZN(n15365) );
  OR2_X1 U18653 ( .A1(n15366), .A2(n15365), .ZN(n19212) );
  INV_X1 U18654 ( .A(n19212), .ZN(n15370) );
  OAI22_X1 U18655 ( .A1(n15386), .A2(n19542), .B1(n19415), .B2(n21317), .ZN(
        n15369) );
  INV_X1 U18656 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15367) );
  OAI22_X1 U18657 ( .A1(n15388), .A2(n16738), .B1(n15387), .B2(n15367), .ZN(
        n15368) );
  AOI211_X1 U18658 ( .C1(n19443), .C2(n15370), .A(n15369), .B(n15368), .ZN(
        n15371) );
  OAI21_X1 U18659 ( .B1(n15372), .B2(n19419), .A(n15371), .ZN(P2_U2900) );
  NAND2_X1 U18660 ( .A1(n15384), .A2(n15373), .ZN(n15374) );
  NAND2_X1 U18661 ( .A1(n15682), .A2(n15374), .ZN(n15692) );
  INV_X1 U18662 ( .A(n15692), .ZN(n19239) );
  OAI22_X1 U18663 ( .A1(n15386), .A2(n19441), .B1(n19415), .B2(n21469), .ZN(
        n15378) );
  INV_X1 U18664 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n15376) );
  INV_X1 U18665 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15375) );
  OAI22_X1 U18666 ( .A1(n15388), .A2(n15376), .B1(n15387), .B2(n15375), .ZN(
        n15377) );
  AOI211_X1 U18667 ( .C1(n19443), .C2(n19239), .A(n15378), .B(n15377), .ZN(
        n15379) );
  OAI21_X1 U18668 ( .B1(n15380), .B2(n19419), .A(n15379), .ZN(P2_U2902) );
  OR2_X1 U18669 ( .A1(n15382), .A2(n15381), .ZN(n15383) );
  NAND2_X1 U18670 ( .A1(n15384), .A2(n15383), .ZN(n19260) );
  INV_X1 U18671 ( .A(n19260), .ZN(n15391) );
  OAI22_X1 U18672 ( .A1(n15386), .A2(n19451), .B1(n19415), .B2(n15385), .ZN(
        n15390) );
  OAI22_X1 U18673 ( .A1(n15388), .A2(n16742), .B1(n15387), .B2(n14197), .ZN(
        n15389) );
  AOI211_X1 U18674 ( .C1(n19443), .C2(n15391), .A(n15390), .B(n15389), .ZN(
        n15392) );
  OAI21_X1 U18675 ( .B1(n15393), .B2(n19419), .A(n15392), .ZN(P2_U2903) );
  AOI21_X1 U18676 ( .B1(n15410), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15395) );
  OR2_X1 U18677 ( .A1(n15395), .A2(n15394), .ZN(n15565) );
  INV_X1 U18678 ( .A(n15396), .ZN(n15400) );
  OR2_X1 U18679 ( .A1(n15398), .A2(n15397), .ZN(n15399) );
  XNOR2_X1 U18680 ( .A(n15400), .B(n15399), .ZN(n15556) );
  NOR2_X1 U18681 ( .A1(n16391), .A2(n14195), .ZN(n15403) );
  NAND2_X1 U18682 ( .A1(n19247), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15560) );
  NAND2_X1 U18683 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15401) );
  OAI211_X1 U18684 ( .C1(n19499), .C2(n16395), .A(n15560), .B(n15401), .ZN(
        n15402) );
  AOI211_X1 U18685 ( .C1(n15556), .C2(n19493), .A(n15403), .B(n15402), .ZN(
        n15404) );
  OAI21_X1 U18686 ( .B1(n16543), .B2(n15565), .A(n15404), .ZN(P2_U2985) );
  NAND2_X1 U18687 ( .A1(n15406), .A2(n15405), .ZN(n15407) );
  XNOR2_X1 U18688 ( .A(n15410), .B(n15409), .ZN(n15577) );
  NOR2_X1 U18689 ( .A1(n15573), .A2(n14195), .ZN(n15414) );
  NAND2_X1 U18690 ( .A1(n19247), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15572) );
  NAND2_X1 U18691 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15411) );
  OAI211_X1 U18692 ( .C1(n19499), .C2(n15412), .A(n15572), .B(n15411), .ZN(
        n15413) );
  AOI211_X1 U18693 ( .C1(n15577), .C2(n19495), .A(n15414), .B(n15413), .ZN(
        n15415) );
  OAI21_X1 U18694 ( .B1(n15580), .B2(n16541), .A(n15415), .ZN(P2_U2986) );
  NAND3_X1 U18695 ( .A1(n15417), .A2(n19493), .A3(n15416), .ZN(n15423) );
  OAI21_X1 U18696 ( .B1(n16561), .B2(n16400), .A(n15418), .ZN(n15420) );
  NOR2_X1 U18697 ( .A1(n16403), .A2(n14195), .ZN(n15419) );
  AOI211_X1 U18698 ( .C1(n16550), .C2(n15421), .A(n15420), .B(n15419), .ZN(
        n15422) );
  OAI211_X1 U18699 ( .C1(n16543), .C2(n15424), .A(n15423), .B(n15422), .ZN(
        P2_U2987) );
  OAI21_X1 U18700 ( .B1(n15425), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12815), .ZN(n15589) );
  INV_X1 U18701 ( .A(n15426), .ZN(n15434) );
  NOR2_X1 U18702 ( .A1(n15427), .A2(n15434), .ZN(n15429) );
  XNOR2_X1 U18703 ( .A(n15429), .B(n15428), .ZN(n15587) );
  NOR2_X1 U18704 ( .A1(n16416), .A2(n14195), .ZN(n15432) );
  NAND2_X1 U18705 ( .A1(n19247), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15581) );
  NAND2_X1 U18706 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15430) );
  OAI211_X1 U18707 ( .C1(n19499), .C2(n16420), .A(n15581), .B(n15430), .ZN(
        n15431) );
  AOI211_X1 U18708 ( .C1(n15587), .C2(n19493), .A(n15432), .B(n15431), .ZN(
        n15433) );
  OAI21_X1 U18709 ( .B1(n16543), .B2(n15589), .A(n15433), .ZN(P2_U2988) );
  NOR2_X1 U18710 ( .A1(n15435), .A2(n15434), .ZN(n15437) );
  XOR2_X1 U18711 ( .A(n15437), .B(n15436), .Z(n15600) );
  AOI21_X1 U18712 ( .B1(n15596), .B2(n15438), .A(n15425), .ZN(n15590) );
  NAND2_X1 U18713 ( .A1(n15590), .A2(n19495), .ZN(n15444) );
  NAND2_X1 U18714 ( .A1(n19247), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15593) );
  OAI21_X1 U18715 ( .B1(n16561), .B2(n15439), .A(n15593), .ZN(n15441) );
  NOR2_X1 U18716 ( .A1(n16428), .A2(n14195), .ZN(n15440) );
  AOI211_X1 U18717 ( .C1(n16550), .C2(n15442), .A(n15441), .B(n15440), .ZN(
        n15443) );
  OAI211_X1 U18718 ( .C1(n16541), .C2(n15600), .A(n15444), .B(n15443), .ZN(
        P2_U2989) );
  OAI21_X1 U18719 ( .B1(n15452), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15438), .ZN(n15610) );
  XOR2_X1 U18720 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15445), .Z(
        n15446) );
  XNOR2_X1 U18721 ( .A(n15447), .B(n15446), .ZN(n15608) );
  INV_X1 U18722 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20175) );
  NOR2_X1 U18723 ( .A1(n19348), .A2(n20175), .ZN(n15604) );
  NOR2_X1 U18724 ( .A1(n19499), .A2(n16445), .ZN(n15448) );
  AOI211_X1 U18725 ( .C1(n19488), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15604), .B(n15448), .ZN(n15449) );
  OAI21_X1 U18726 ( .B1(n16441), .B2(n14195), .A(n15449), .ZN(n15450) );
  AOI21_X1 U18727 ( .B1(n15608), .B2(n19493), .A(n15450), .ZN(n15451) );
  OAI21_X1 U18728 ( .B1(n15610), .B2(n16543), .A(n15451), .ZN(P2_U2990) );
  INV_X1 U18729 ( .A(n15452), .ZN(n15453) );
  OAI21_X1 U18730 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n10099), .A(
        n15453), .ZN(n15621) );
  XNOR2_X1 U18731 ( .A(n10009), .B(n15455), .ZN(n15619) );
  OAI22_X1 U18732 ( .A1(n16561), .A2(n16450), .B1(n19499), .B2(n16458), .ZN(
        n15457) );
  NAND2_X1 U18733 ( .A1(n19247), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15611) );
  OAI21_X1 U18734 ( .B1(n16453), .B2(n14195), .A(n15611), .ZN(n15456) );
  AOI211_X1 U18735 ( .C1(n15619), .C2(n19493), .A(n15457), .B(n15456), .ZN(
        n15458) );
  OAI21_X1 U18736 ( .B1(n15621), .B2(n16543), .A(n15458), .ZN(P2_U2991) );
  INV_X1 U18737 ( .A(n15459), .ZN(n15460) );
  OAI21_X1 U18738 ( .B1(n15716), .B2(n15460), .A(n15717), .ZN(n15528) );
  INV_X1 U18739 ( .A(n15526), .ZN(n15461) );
  INV_X1 U18740 ( .A(n15462), .ZN(n15521) );
  INV_X1 U18741 ( .A(n15464), .ZN(n15465) );
  AOI21_X1 U18742 ( .B1(n15493), .B2(n15490), .A(n15465), .ZN(n15483) );
  AOI21_X1 U18743 ( .B1(n15483), .B2(n15479), .A(n15481), .ZN(n15469) );
  NAND2_X1 U18744 ( .A1(n15467), .A2(n15466), .ZN(n15468) );
  XNOR2_X1 U18745 ( .A(n15469), .B(n15468), .ZN(n15650) );
  INV_X1 U18746 ( .A(n15472), .ZN(n15473) );
  AOI21_X1 U18747 ( .B1(n15645), .B2(n15471), .A(n15473), .ZN(n15648) );
  NAND2_X1 U18748 ( .A1(n19247), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15640) );
  OAI21_X1 U18749 ( .B1(n16561), .B2(n19196), .A(n15640), .ZN(n15474) );
  AOI21_X1 U18750 ( .B1(n16550), .B2(n15475), .A(n15474), .ZN(n15476) );
  OAI21_X1 U18751 ( .B1(n19200), .B2(n14195), .A(n15476), .ZN(n15477) );
  AOI21_X1 U18752 ( .B1(n15648), .B2(n19495), .A(n15477), .ZN(n15478) );
  OAI21_X1 U18753 ( .B1(n15650), .B2(n16541), .A(n15478), .ZN(P2_U2993) );
  INV_X1 U18754 ( .A(n15479), .ZN(n15480) );
  NOR2_X1 U18755 ( .A1(n15481), .A2(n15480), .ZN(n15482) );
  XNOR2_X1 U18756 ( .A(n15483), .B(n15482), .ZN(n15662) );
  NAND2_X1 U18757 ( .A1(n19247), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15652) );
  NAND2_X1 U18758 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15484) );
  OAI211_X1 U18759 ( .C1(n19499), .C2(n15485), .A(n15652), .B(n15484), .ZN(
        n15488) );
  OAI21_X1 U18760 ( .B1(n15486), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15471), .ZN(n15659) );
  NOR2_X1 U18761 ( .A1(n15659), .A2(n16543), .ZN(n15487) );
  AOI211_X1 U18762 ( .C1(n19494), .C2(n15651), .A(n15488), .B(n15487), .ZN(
        n15489) );
  OAI21_X1 U18763 ( .B1(n15662), .B2(n16541), .A(n15489), .ZN(P2_U2994) );
  NAND2_X1 U18764 ( .A1(n15491), .A2(n15490), .ZN(n15495) );
  INV_X1 U18765 ( .A(n15675), .ZN(n15492) );
  NOR2_X1 U18766 ( .A1(n15493), .A2(n15492), .ZN(n15494) );
  XOR2_X1 U18767 ( .A(n15495), .B(n15494), .Z(n15673) );
  AOI21_X1 U18768 ( .B1(n15669), .B2(n15496), .A(n15486), .ZN(n15671) );
  NAND2_X1 U18769 ( .A1(n19247), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15664) );
  OAI21_X1 U18770 ( .B1(n16561), .B2(n15497), .A(n15664), .ZN(n15498) );
  AOI21_X1 U18771 ( .B1(n15499), .B2(n16550), .A(n15498), .ZN(n15500) );
  OAI21_X1 U18772 ( .B1(n19213), .B2(n14195), .A(n15500), .ZN(n15501) );
  AOI21_X1 U18773 ( .B1(n15671), .B2(n19495), .A(n15501), .ZN(n15502) );
  OAI21_X1 U18774 ( .B1(n15673), .B2(n16541), .A(n15502), .ZN(P2_U2995) );
  NAND2_X1 U18775 ( .A1(n15504), .A2(n15503), .ZN(n15507) );
  NAND2_X1 U18776 ( .A1(n9910), .A2(n15505), .ZN(n15506) );
  XOR2_X1 U18777 ( .A(n15507), .B(n15506), .Z(n15704) );
  INV_X1 U18778 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20162) );
  NOR2_X1 U18779 ( .A1(n20162), .A2(n19348), .ZN(n15509) );
  OAI22_X1 U18780 ( .A1(n16561), .A2(n19235), .B1(n19499), .B2(n19243), .ZN(
        n15508) );
  AOI211_X1 U18781 ( .C1(n19494), .C2(n19240), .A(n15509), .B(n15508), .ZN(
        n15513) );
  INV_X1 U18782 ( .A(n16564), .ZN(n15696) );
  NAND2_X1 U18783 ( .A1(n13651), .A2(n15696), .ZN(n15525) );
  INV_X1 U18784 ( .A(n15510), .ZN(n15693) );
  NOR2_X1 U18785 ( .A1(n15525), .A2(n15693), .ZN(n15698) );
  OAI211_X1 U18786 ( .C1(n15698), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19495), .B(n15511), .ZN(n15512) );
  OAI211_X1 U18787 ( .C1(n15704), .C2(n16541), .A(n15513), .B(n15512), .ZN(
        P2_U2997) );
  INV_X1 U18788 ( .A(n15514), .ZN(n19254) );
  INV_X1 U18789 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15517) );
  INV_X1 U18790 ( .A(n19256), .ZN(n15515) );
  NAND2_X1 U18791 ( .A1(n15515), .A2(n16550), .ZN(n15516) );
  NAND2_X1 U18792 ( .A1(n19247), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15705) );
  OAI211_X1 U18793 ( .C1(n15517), .C2(n16561), .A(n15516), .B(n15705), .ZN(
        n15520) );
  INV_X1 U18794 ( .A(n15525), .ZN(n15722) );
  AOI21_X1 U18795 ( .B1(n15722), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15518) );
  NOR3_X1 U18796 ( .A1(n15518), .A2(n15698), .A3(n16543), .ZN(n15519) );
  AOI211_X1 U18797 ( .C1(n19254), .C2(n19494), .A(n15520), .B(n15519), .ZN(
        n15524) );
  NAND2_X1 U18798 ( .A1(n15522), .A2(n15521), .ZN(n15709) );
  NAND3_X1 U18799 ( .A1(n9910), .A2(n19493), .A3(n15709), .ZN(n15523) );
  NAND2_X1 U18800 ( .A1(n15524), .A2(n15523), .ZN(P2_U2998) );
  XNOR2_X1 U18801 ( .A(n15525), .B(n16570), .ZN(n16572) );
  NAND2_X1 U18802 ( .A1(n15527), .A2(n15526), .ZN(n15529) );
  XOR2_X1 U18803 ( .A(n15529), .B(n15528), .Z(n16577) );
  INV_X1 U18804 ( .A(n16577), .ZN(n15534) );
  INV_X1 U18805 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20158) );
  OAI22_X1 U18806 ( .A1(n16561), .A2(n15530), .B1(n20158), .B2(n19348), .ZN(
        n15533) );
  INV_X1 U18807 ( .A(n16573), .ZN(n19265) );
  INV_X1 U18808 ( .A(n19262), .ZN(n15531) );
  OAI22_X1 U18809 ( .A1(n19265), .A2(n14195), .B1(n19499), .B2(n15531), .ZN(
        n15532) );
  AOI211_X1 U18810 ( .C1(n15534), .C2(n19493), .A(n15533), .B(n15532), .ZN(
        n15535) );
  OAI21_X1 U18811 ( .B1(n16543), .B2(n16572), .A(n15535), .ZN(P2_U2999) );
  NAND2_X1 U18812 ( .A1(n15536), .A2(n15714), .ZN(n15537) );
  XNOR2_X1 U18813 ( .A(n15538), .B(n15537), .ZN(n15752) );
  INV_X1 U18814 ( .A(n15539), .ZN(n19289) );
  INV_X1 U18815 ( .A(n15782), .ZN(n15724) );
  NAND2_X1 U18816 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15753), .ZN(
        n15754) );
  AND2_X1 U18817 ( .A1(n15753), .A2(n15734), .ZN(n15721) );
  AOI21_X1 U18818 ( .B1(n12302), .B2(n15754), .A(n15721), .ZN(n15750) );
  INV_X1 U18819 ( .A(n15750), .ZN(n15540) );
  OAI22_X1 U18820 ( .A1(n19499), .A2(n19289), .B1(n16543), .B2(n15540), .ZN(
        n15543) );
  INV_X1 U18821 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20154) );
  OAI22_X1 U18822 ( .A1(n16561), .A2(n15541), .B1(n20154), .B2(n19348), .ZN(
        n15542) );
  AOI211_X1 U18823 ( .C1(n19494), .C2(n19283), .A(n15543), .B(n15542), .ZN(
        n15544) );
  OAI21_X1 U18824 ( .B1(n15752), .B2(n16541), .A(n15544), .ZN(P2_U3001) );
  XNOR2_X1 U18825 ( .A(n15545), .B(n15546), .ZN(n15803) );
  INV_X1 U18826 ( .A(n16529), .ZN(n15548) );
  NOR2_X1 U18827 ( .A1(n16528), .A2(n15548), .ZN(n15549) );
  XNOR2_X1 U18828 ( .A(n15547), .B(n15549), .ZN(n15799) );
  INV_X1 U18829 ( .A(n15799), .ZN(n15554) );
  OAI22_X1 U18830 ( .A1(n16561), .A2(n15550), .B1(n20143), .B2(n19348), .ZN(
        n15553) );
  INV_X1 U18831 ( .A(n19325), .ZN(n15551) );
  OAI22_X1 U18832 ( .A1(n14195), .A2(n19330), .B1(n19499), .B2(n15551), .ZN(
        n15552) );
  AOI211_X1 U18833 ( .C1(n15554), .C2(n19493), .A(n15553), .B(n15552), .ZN(
        n15555) );
  OAI21_X1 U18834 ( .B1(n15803), .B2(n16543), .A(n15555), .ZN(P2_U3007) );
  NAND2_X1 U18835 ( .A1(n15556), .A2(n19526), .ZN(n15564) );
  NAND2_X1 U18836 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15568) );
  AOI211_X1 U18837 ( .C1(n15568), .C2(n15558), .A(n10326), .B(n15566), .ZN(
        n15562) );
  NAND2_X1 U18838 ( .A1(n19517), .A2(n16389), .ZN(n15559) );
  OAI211_X1 U18839 ( .C1(n16391), .C2(n19534), .A(n15560), .B(n15559), .ZN(
        n15561) );
  AOI211_X1 U18840 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15576), .A(
        n15562), .B(n15561), .ZN(n15563) );
  OAI211_X1 U18841 ( .C1(n15565), .C2(n16604), .A(n15564), .B(n15563), .ZN(
        P2_U3017) );
  INV_X1 U18842 ( .A(n15566), .ZN(n15569) );
  AND3_X1 U18843 ( .A1(n15569), .A2(n15568), .A3(n15567), .ZN(n15575) );
  NAND2_X1 U18844 ( .A1(n19517), .A2(n15570), .ZN(n15571) );
  OAI211_X1 U18845 ( .C1(n15573), .C2(n19534), .A(n15572), .B(n15571), .ZN(
        n15574) );
  AOI211_X1 U18846 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15576), .A(
        n15575), .B(n15574), .ZN(n15579) );
  NAND2_X1 U18847 ( .A1(n15577), .A2(n12862), .ZN(n15578) );
  OAI211_X1 U18848 ( .C1(n15580), .C2(n16587), .A(n15579), .B(n15578), .ZN(
        P2_U3018) );
  XOR2_X1 U18849 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n15584) );
  OAI21_X1 U18850 ( .B1(n16603), .B2(n16415), .A(n15581), .ZN(n15583) );
  NOR2_X1 U18851 ( .A1(n16416), .A2(n19534), .ZN(n15582) );
  AOI211_X1 U18852 ( .C1(n15584), .C2(n15597), .A(n15583), .B(n15582), .ZN(
        n15585) );
  OAI21_X1 U18853 ( .B1(n21537), .B2(n15591), .A(n15585), .ZN(n15586) );
  AOI21_X1 U18854 ( .B1(n15587), .B2(n19526), .A(n15586), .ZN(n15588) );
  OAI21_X1 U18855 ( .B1(n16604), .B2(n15589), .A(n15588), .ZN(P2_U3020) );
  NAND2_X1 U18856 ( .A1(n15590), .A2(n12862), .ZN(n15599) );
  NOR2_X1 U18857 ( .A1(n15591), .A2(n15596), .ZN(n15595) );
  NAND2_X1 U18858 ( .A1(n19517), .A2(n16426), .ZN(n15592) );
  OAI211_X1 U18859 ( .C1(n16428), .C2(n19534), .A(n15593), .B(n15592), .ZN(
        n15594) );
  AOI211_X1 U18860 ( .C1(n15597), .C2(n15596), .A(n15595), .B(n15594), .ZN(
        n15598) );
  OAI211_X1 U18861 ( .C1(n15600), .C2(n16587), .A(n15599), .B(n15598), .ZN(
        P2_U3021) );
  INV_X1 U18862 ( .A(n15601), .ZN(n15603) );
  OAI21_X1 U18863 ( .B1(n15603), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15602), .ZN(n15606) );
  AOI21_X1 U18864 ( .B1(n19517), .B2(n16439), .A(n15604), .ZN(n15605) );
  OAI211_X1 U18865 ( .C1(n16441), .C2(n19534), .A(n15606), .B(n15605), .ZN(
        n15607) );
  AOI21_X1 U18866 ( .B1(n15608), .B2(n19526), .A(n15607), .ZN(n15609) );
  OAI21_X1 U18867 ( .B1(n15610), .B2(n16604), .A(n15609), .ZN(P2_U3022) );
  INV_X1 U18868 ( .A(n16453), .ZN(n15615) );
  OAI21_X1 U18869 ( .B1(n16603), .B2(n16461), .A(n15611), .ZN(n15614) );
  AOI211_X1 U18870 ( .C1(n15617), .C2(n15636), .A(n15612), .B(n15632), .ZN(
        n15613) );
  AOI211_X1 U18871 ( .C1(n15615), .C2(n19500), .A(n15614), .B(n15613), .ZN(
        n15616) );
  OAI21_X1 U18872 ( .B1(n15637), .B2(n15617), .A(n15616), .ZN(n15618) );
  AOI21_X1 U18873 ( .B1(n15619), .B2(n19526), .A(n15618), .ZN(n15620) );
  OAI21_X1 U18874 ( .B1(n15621), .B2(n16604), .A(n15620), .ZN(P2_U3023) );
  NAND2_X1 U18875 ( .A1(n15472), .A2(n15636), .ZN(n15622) );
  NAND2_X1 U18876 ( .A1(n15623), .A2(n15622), .ZN(n16482) );
  OR2_X1 U18877 ( .A1(n15624), .A2(n9960), .ZN(n15625) );
  XNOR2_X1 U18878 ( .A(n15626), .B(n15625), .ZN(n16485) );
  INV_X1 U18879 ( .A(n16002), .ZN(n16484) );
  OR2_X1 U18880 ( .A1(n15628), .A2(n15627), .ZN(n15629) );
  NAND2_X1 U18881 ( .A1(n15630), .A2(n15629), .ZN(n16463) );
  NAND2_X1 U18882 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19247), .ZN(n15631) );
  OAI21_X1 U18883 ( .B1(n16603), .B2(n16463), .A(n15631), .ZN(n15634) );
  NOR2_X1 U18884 ( .A1(n15632), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15633) );
  AOI211_X1 U18885 ( .C1(n16484), .C2(n19500), .A(n15634), .B(n15633), .ZN(
        n15635) );
  OAI21_X1 U18886 ( .B1(n15637), .B2(n15636), .A(n15635), .ZN(n15638) );
  AOI21_X1 U18887 ( .B1(n16485), .B2(n19526), .A(n15638), .ZN(n15639) );
  OAI21_X1 U18888 ( .B1(n16482), .B2(n16604), .A(n15639), .ZN(P2_U3024) );
  INV_X1 U18889 ( .A(n19200), .ZN(n15642) );
  OAI21_X1 U18890 ( .B1(n16603), .B2(n19208), .A(n15640), .ZN(n15641) );
  AOI21_X1 U18891 ( .B1(n15642), .B2(n19500), .A(n15641), .ZN(n15644) );
  OAI211_X1 U18892 ( .C1(n15646), .C2(n15645), .A(n15644), .B(n15643), .ZN(
        n15647) );
  AOI21_X1 U18893 ( .B1(n15648), .B2(n12862), .A(n15647), .ZN(n15649) );
  OAI21_X1 U18894 ( .B1(n15650), .B2(n16587), .A(n15649), .ZN(P2_U3025) );
  INV_X1 U18895 ( .A(n15688), .ZN(n15658) );
  NAND2_X1 U18896 ( .A1(n15651), .A2(n19500), .ZN(n15653) );
  OAI211_X1 U18897 ( .C1(n16603), .C2(n16470), .A(n15653), .B(n15652), .ZN(
        n15657) );
  AOI211_X1 U18898 ( .C1(n15655), .C2(n15669), .A(n15654), .B(n15663), .ZN(
        n15656) );
  AOI211_X1 U18899 ( .C1(n15658), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15657), .B(n15656), .ZN(n15661) );
  OR2_X1 U18900 ( .A1(n15659), .A2(n16604), .ZN(n15660) );
  OAI211_X1 U18901 ( .C1(n15662), .C2(n16587), .A(n15661), .B(n15660), .ZN(
        P2_U3026) );
  INV_X1 U18902 ( .A(n15663), .ZN(n15667) );
  NOR2_X1 U18903 ( .A1(n16603), .A2(n19212), .ZN(n15666) );
  OAI21_X1 U18904 ( .B1(n19213), .B2(n19534), .A(n15664), .ZN(n15665) );
  AOI211_X1 U18905 ( .C1(n15667), .C2(n15669), .A(n15666), .B(n15665), .ZN(
        n15668) );
  OAI21_X1 U18906 ( .B1(n15669), .B2(n15688), .A(n15668), .ZN(n15670) );
  AOI21_X1 U18907 ( .B1(n15671), .B2(n12862), .A(n15670), .ZN(n15672) );
  OAI21_X1 U18908 ( .B1(n15673), .B2(n16587), .A(n15672), .ZN(P2_U3027) );
  NAND2_X1 U18909 ( .A1(n15675), .A2(n15674), .ZN(n15677) );
  XOR2_X1 U18910 ( .A(n15677), .B(n15676), .Z(n16490) );
  INV_X1 U18911 ( .A(n16490), .ZN(n15691) );
  NAND2_X1 U18912 ( .A1(n15511), .A2(n15678), .ZN(n15679) );
  AND2_X1 U18913 ( .A1(n15496), .A2(n15679), .ZN(n16489) );
  AOI21_X1 U18914 ( .B1(n15781), .B2(n15680), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15687) );
  AOI21_X1 U18915 ( .B1(n15683), .B2(n15682), .A(n15681), .ZN(n19225) );
  INV_X1 U18916 ( .A(n19225), .ZN(n15684) );
  INV_X1 U18917 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20164) );
  OAI22_X1 U18918 ( .A1(n16603), .A2(n15684), .B1(n20164), .B2(n19348), .ZN(
        n15685) );
  AOI21_X1 U18919 ( .B1(n19226), .B2(n19500), .A(n15685), .ZN(n15686) );
  OAI21_X1 U18920 ( .B1(n15688), .B2(n15687), .A(n15686), .ZN(n15689) );
  AOI21_X1 U18921 ( .B1(n16489), .B2(n12862), .A(n15689), .ZN(n15690) );
  OAI21_X1 U18922 ( .B1(n15691), .B2(n16587), .A(n15690), .ZN(P2_U3028) );
  OAI22_X1 U18923 ( .A1(n16603), .A2(n15692), .B1(n20162), .B2(n19348), .ZN(
        n15695) );
  AOI22_X1 U18924 ( .A1(n15722), .A2(n12862), .B1(n15696), .B2(n15781), .ZN(
        n15706) );
  NOR3_X1 U18925 ( .A1(n15706), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15693), .ZN(n15694) );
  AOI211_X1 U18926 ( .C1(n19240), .C2(n19500), .A(n15695), .B(n15694), .ZN(
        n15703) );
  INV_X1 U18927 ( .A(n19512), .ZN(n15700) );
  OR2_X1 U18928 ( .A1(n15726), .A2(n15696), .ZN(n15697) );
  NAND2_X1 U18929 ( .A1(n15780), .A2(n15697), .ZN(n16569) );
  AOI21_X1 U18930 ( .B1(n16604), .B2(n19523), .A(n15698), .ZN(n15699) );
  AOI211_X1 U18931 ( .C1(n15700), .C2(n16570), .A(n16569), .B(n15699), .ZN(
        n15713) );
  OAI21_X1 U18932 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15726), .A(
        n15713), .ZN(n15701) );
  NAND2_X1 U18933 ( .A1(n15701), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15702) );
  OAI211_X1 U18934 ( .C1(n15704), .C2(n16587), .A(n15703), .B(n15702), .ZN(
        P2_U3029) );
  OAI21_X1 U18935 ( .B1(n16603), .B2(n19260), .A(n15705), .ZN(n15708) );
  NOR3_X1 U18936 ( .A1(n15706), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16570), .ZN(n15707) );
  AOI211_X1 U18937 ( .C1(n19500), .C2(n19254), .A(n15708), .B(n15707), .ZN(
        n15711) );
  NAND3_X1 U18938 ( .A1(n9910), .A2(n19526), .A3(n15709), .ZN(n15710) );
  OAI211_X1 U18939 ( .C1(n15713), .C2(n15712), .A(n15711), .B(n15710), .ZN(
        P2_U3030) );
  INV_X1 U18940 ( .A(n15714), .ZN(n15715) );
  NOR2_X1 U18941 ( .A1(n15716), .A2(n15715), .ZN(n15720) );
  NAND2_X1 U18942 ( .A1(n15718), .A2(n15717), .ZN(n15719) );
  XNOR2_X1 U18943 ( .A(n15720), .B(n15719), .ZN(n16493) );
  INV_X1 U18944 ( .A(n16493), .ZN(n15741) );
  INV_X1 U18945 ( .A(n15721), .ZN(n15723) );
  AOI21_X1 U18946 ( .B1(n15723), .B2(n15737), .A(n15722), .ZN(n16494) );
  NAND2_X1 U18947 ( .A1(n16494), .A2(n12862), .ZN(n15740) );
  INV_X1 U18948 ( .A(n15734), .ZN(n15728) );
  INV_X1 U18949 ( .A(n15781), .ZN(n16563) );
  NOR3_X1 U18950 ( .A1(n15725), .A2(n15724), .A3(n16563), .ZN(n15759) );
  OAI21_X1 U18951 ( .B1(n15727), .B2(n15726), .A(n15780), .ZN(n15758) );
  AOI21_X1 U18952 ( .B1(n15728), .B2(n15759), .A(n15758), .ZN(n15743) );
  AOI21_X1 U18953 ( .B1(n15731), .B2(n15729), .A(n15730), .ZN(n19392) );
  NAND2_X1 U18954 ( .A1(n19517), .A2(n19392), .ZN(n15736) );
  INV_X1 U18955 ( .A(n15759), .ZN(n15732) );
  NOR2_X1 U18956 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15732), .ZN(
        n15733) );
  AOI22_X1 U18957 ( .A1(n19247), .A2(P2_REIP_REG_14__SCAN_IN), .B1(n15734), 
        .B2(n15733), .ZN(n15735) );
  OAI211_X1 U18958 ( .C1(n15743), .C2(n15737), .A(n15736), .B(n15735), .ZN(
        n15738) );
  AOI21_X1 U18959 ( .B1(n19500), .B2(n19276), .A(n15738), .ZN(n15739) );
  OAI211_X1 U18960 ( .C1(n15741), .C2(n16587), .A(n15740), .B(n15739), .ZN(
        P2_U3032) );
  AOI21_X1 U18961 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15759), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15742) );
  OAI22_X1 U18962 ( .A1(n19233), .A2(n20154), .B1(n15743), .B2(n15742), .ZN(
        n15749) );
  OR2_X1 U18963 ( .A1(n15745), .A2(n15744), .ZN(n15746) );
  NAND2_X1 U18964 ( .A1(n15746), .A2(n15729), .ZN(n19397) );
  OAI22_X1 U18965 ( .A1(n19534), .A2(n15747), .B1(n16603), .B2(n19397), .ZN(
        n15748) );
  AOI211_X1 U18966 ( .C1(n12862), .C2(n15750), .A(n15749), .B(n15748), .ZN(
        n15751) );
  OAI21_X1 U18967 ( .B1(n15752), .B2(n16587), .A(n15751), .ZN(P2_U3033) );
  INV_X1 U18968 ( .A(n15753), .ZN(n15771) );
  INV_X1 U18969 ( .A(n15754), .ZN(n15755) );
  AOI21_X1 U18970 ( .B1(n15771), .B2(n15756), .A(n15755), .ZN(n16497) );
  NAND2_X1 U18971 ( .A1(n16497), .A2(n12862), .ZN(n15770) );
  INV_X1 U18972 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20152) );
  NOR2_X1 U18973 ( .A1(n20152), .A2(n19348), .ZN(n15757) );
  AOI221_X1 U18974 ( .B1(n15759), .B2(n15756), .C1(n15758), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n15757), .ZN(n15769) );
  XNOR2_X1 U18975 ( .A(n15761), .B(n15760), .ZN(n19400) );
  OAI22_X1 U18976 ( .A1(n19534), .A2(n15762), .B1(n16603), .B2(n19400), .ZN(
        n15763) );
  INV_X1 U18977 ( .A(n15763), .ZN(n15768) );
  OR2_X1 U18978 ( .A1(n15764), .A2(n9977), .ZN(n15765) );
  XNOR2_X1 U18979 ( .A(n15766), .B(n15765), .ZN(n16498) );
  NAND2_X1 U18980 ( .A1(n16498), .A2(n19526), .ZN(n15767) );
  NAND4_X1 U18981 ( .A1(n15770), .A2(n15769), .A3(n15768), .A4(n15767), .ZN(
        P2_U3034) );
  NOR2_X1 U18982 ( .A1(n16516), .A2(n16517), .ZN(n16515) );
  OAI21_X1 U18983 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16515), .A(
        n15771), .ZN(n16503) );
  INV_X1 U18984 ( .A(n15772), .ZN(n15773) );
  NAND2_X1 U18985 ( .A1(n15774), .A2(n15773), .ZN(n15778) );
  NOR2_X1 U18986 ( .A1(n15776), .A2(n15775), .ZN(n15777) );
  XNOR2_X1 U18987 ( .A(n15778), .B(n15777), .ZN(n16502) );
  AOI21_X1 U18988 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15780), .A(
        n15779), .ZN(n16583) );
  NOR2_X1 U18989 ( .A1(n20150), .A2(n19348), .ZN(n15785) );
  NAND2_X1 U18990 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15781), .ZN(
        n16580) );
  AOI211_X1 U18991 ( .C1(n16517), .C2(n15783), .A(n15782), .B(n16580), .ZN(
        n15784) );
  AOI211_X1 U18992 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16583), .A(
        n15785), .B(n15784), .ZN(n15789) );
  OAI22_X1 U18993 ( .A1(n19534), .A2(n15786), .B1(n16603), .B2(n19402), .ZN(
        n15787) );
  INV_X1 U18994 ( .A(n15787), .ZN(n15788) );
  OAI211_X1 U18995 ( .C1(n16502), .C2(n16587), .A(n15789), .B(n15788), .ZN(
        n15790) );
  INV_X1 U18996 ( .A(n15790), .ZN(n15791) );
  OAI21_X1 U18997 ( .B1(n16503), .B2(n16604), .A(n15791), .ZN(P2_U3035) );
  NOR2_X1 U18998 ( .A1(n15792), .A2(n16612), .ZN(n16595) );
  OAI21_X1 U18999 ( .B1(n15795), .B2(n15794), .A(n15793), .ZN(n19413) );
  AOI22_X1 U19000 ( .A1(n19500), .A2(n15796), .B1(n19247), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n15798) );
  NAND2_X1 U19001 ( .A1(n16589), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15797) );
  OAI211_X1 U19002 ( .C1(n19413), .C2(n16603), .A(n15798), .B(n15797), .ZN(
        n15801) );
  NOR2_X1 U19003 ( .A1(n15799), .A2(n16587), .ZN(n15800) );
  AOI211_X1 U19004 ( .C1(n16595), .C2(n16596), .A(n15801), .B(n15800), .ZN(
        n15802) );
  OAI21_X1 U19005 ( .B1(n15803), .B2(n16604), .A(n15802), .ZN(P2_U3039) );
  NAND2_X1 U19006 ( .A1(n19526), .A2(n15804), .ZN(n15806) );
  OAI211_X1 U19007 ( .C1(n19513), .C2(n15833), .A(n15806), .B(n15805), .ZN(
        n15807) );
  AOI21_X1 U19008 ( .B1(n15836), .B2(n19500), .A(n15807), .ZN(n15812) );
  AOI22_X1 U19009 ( .A1(n12862), .A2(n15808), .B1(n19517), .B2(n20223), .ZN(
        n15811) );
  OAI211_X1 U19010 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15809), .B(n19515), .ZN(n15810) );
  NAND3_X1 U19011 ( .A1(n15812), .A2(n15811), .A3(n15810), .ZN(P2_U3045) );
  INV_X1 U19012 ( .A(n15851), .ZN(n15870) );
  NAND2_X1 U19013 ( .A1(n15814), .A2(n15813), .ZN(n15838) );
  MUX2_X1 U19014 ( .A(n12457), .B(n15838), .S(n15815), .Z(n15816) );
  AOI21_X1 U19015 ( .B1(n19365), .B2(n15870), .A(n15816), .ZN(n16618) );
  OAI22_X1 U19016 ( .A1(n9876), .A2(n15817), .B1(n19384), .B2(n9824), .ZN(
        n15834) );
  OAI222_X1 U19017 ( .A1(n16660), .A2(n15819), .B1(n20200), .B2(n16618), .C1(
        n15818), .C2(n15834), .ZN(n15831) );
  NOR2_X1 U19018 ( .A1(n12197), .A2(n15820), .ZN(n15821) );
  NAND2_X1 U19019 ( .A1(n15822), .A2(n15821), .ZN(n15827) );
  INV_X1 U19020 ( .A(n15823), .ZN(n15825) );
  NAND4_X1 U19021 ( .A1(n15827), .A2(n15826), .A3(n15825), .A4(n15824), .ZN(
        n16628) );
  NAND2_X1 U19022 ( .A1(n16628), .A2(n16665), .ZN(n15830) );
  NAND2_X1 U19023 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16649), .ZN(n16668) );
  NOR2_X1 U19024 ( .A1(n19174), .A2(n16668), .ZN(n15828) );
  AOI21_X1 U19025 ( .B1(n16656), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n15828), 
        .ZN(n15829) );
  NAND2_X1 U19026 ( .A1(n15830), .A2(n15829), .ZN(n15990) );
  MUX2_X1 U19027 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15831), .S(
        n15990), .Z(P2_U3601) );
  OAI21_X1 U19028 ( .B1(n9876), .B2(n15833), .A(n15832), .ZN(n15854) );
  INV_X1 U19029 ( .A(n15834), .ZN(n15835) );
  NOR2_X1 U19030 ( .A1(n15835), .A2(n15818), .ZN(n15853) );
  INV_X1 U19031 ( .A(n15853), .ZN(n15842) );
  NAND2_X1 U19032 ( .A1(n15836), .A2(n15870), .ZN(n15841) );
  NOR2_X1 U19033 ( .A1(n11858), .A2(n11856), .ZN(n15837) );
  AOI22_X1 U19034 ( .A1(n12457), .A2(n15839), .B1(n15838), .B2(n15837), .ZN(
        n15840) );
  AND2_X1 U19035 ( .A1(n15841), .A2(n15840), .ZN(n16622) );
  OAI222_X1 U19036 ( .A1(n19676), .A2(n16660), .B1(n15854), .B2(n15842), .C1(
        n16622), .C2(n20200), .ZN(n15843) );
  MUX2_X1 U19037 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15843), .S(
        n15990), .Z(P2_U3600) );
  AOI21_X1 U19038 ( .B1(n15844), .B2(n12744), .A(n11872), .ZN(n15860) );
  NOR2_X1 U19039 ( .A1(n11856), .A2(n16615), .ZN(n15859) );
  INV_X1 U19040 ( .A(n15859), .ZN(n15863) );
  NOR2_X1 U19041 ( .A1(n15845), .A2(n15846), .ZN(n15847) );
  AOI22_X1 U19042 ( .A1(n15860), .A2(n15863), .B1(n15847), .B2(n12457), .ZN(
        n15850) );
  INV_X1 U19043 ( .A(n16639), .ZN(n15848) );
  NAND2_X1 U19044 ( .A1(n16641), .A2(n15848), .ZN(n15864) );
  OAI21_X1 U19045 ( .B1(n11872), .B2(n15859), .A(n15864), .ZN(n15849) );
  OAI211_X1 U19046 ( .C1(n19533), .C2(n15851), .A(n15850), .B(n15849), .ZN(
        n16624) );
  INV_X1 U19047 ( .A(n16660), .ZN(n15852) );
  AOI222_X1 U19048 ( .A1(n16624), .A2(n15855), .B1(n15854), .B2(n15853), .C1(
        n15852), .C2(n19677), .ZN(n15858) );
  INV_X1 U19049 ( .A(n15990), .ZN(n15857) );
  NAND2_X1 U19050 ( .A1(n15857), .A2(n16615), .ZN(n15856) );
  OAI21_X1 U19051 ( .B1(n15858), .B2(n15857), .A(n15856), .ZN(P2_U3599) );
  INV_X1 U19052 ( .A(n12457), .ZN(n15862) );
  INV_X1 U19053 ( .A(n15860), .ZN(n15861) );
  OAI211_X1 U19054 ( .C1(n15846), .C2(n15862), .A(n15863), .B(n15861), .ZN(
        n15868) );
  NAND2_X1 U19055 ( .A1(n15864), .A2(n15863), .ZN(n15866) );
  AOI21_X1 U19056 ( .B1(n12457), .B2(n15846), .A(n11872), .ZN(n15865) );
  NAND2_X1 U19057 ( .A1(n15866), .A2(n15865), .ZN(n15867) );
  MUX2_X1 U19058 ( .A(n15868), .B(n15867), .S(n16617), .Z(n15869) );
  AOI21_X1 U19059 ( .B1(n16601), .B2(n15870), .A(n15869), .ZN(n16616) );
  OAI22_X1 U19060 ( .A1(n20202), .A2(n16660), .B1(n16616), .B2(n20200), .ZN(
        n15871) );
  MUX2_X1 U19061 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15871), .S(
        n15990), .Z(P2_U3596) );
  NAND4_X1 U19062 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(P3_EBX_REG_12__SCAN_IN), .ZN(n17337)
         );
  INV_X1 U19063 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17429) );
  INV_X1 U19064 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17085) );
  INV_X1 U19065 ( .A(n18946), .ZN(n15978) );
  NOR2_X1 U19066 ( .A1(n18545), .A2(n18528), .ZN(n15872) );
  INV_X1 U19067 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17512) );
  NAND2_X1 U19068 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17513) );
  NOR2_X1 U19069 ( .A1(n17512), .A2(n17513), .ZN(n17504) );
  NAND4_X1 U19070 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17519), .A4(n17504), .ZN(n17502) );
  NAND4_X1 U19071 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(P3_EBX_REG_5__SCAN_IN), .ZN(n15874) );
  NAND2_X1 U19072 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17431), .ZN(n17428) );
  NAND4_X1 U19073 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .A4(n17411), .ZN(n15875) );
  NAND3_X1 U19074 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n17323), .ZN(n17295) );
  INV_X1 U19075 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16922) );
  INV_X1 U19076 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17258) );
  INV_X1 U19077 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17271) );
  INV_X1 U19078 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17296) );
  NOR4_X1 U19079 ( .A1(n16922), .A2(n17258), .A3(n17271), .A4(n17296), .ZN(
        n17203) );
  NAND2_X1 U19080 ( .A1(n17297), .A2(n17203), .ZN(n17248) );
  NAND3_X1 U19081 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17263), .ZN(n17250) );
  NAND2_X1 U19082 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17243), .ZN(n15952) );
  INV_X1 U19083 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16881) );
  INV_X1 U19084 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17242) );
  NOR2_X1 U19085 ( .A1(n16881), .A2(n17242), .ZN(n17238) );
  NAND2_X1 U19086 ( .A1(n17612), .A2(n17519), .ZN(n17525) );
  INV_X1 U19087 ( .A(n17519), .ZN(n17522) );
  NOR2_X1 U19088 ( .A1(n17523), .A2(n17243), .ZN(n17244) );
  INV_X1 U19089 ( .A(n17244), .ZN(n17252) );
  OAI21_X1 U19090 ( .B1(n17238), .B2(n17525), .A(n17252), .ZN(n17236) );
  AOI22_X1 U19091 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15879) );
  AOI22_X1 U19092 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15878) );
  AOI22_X1 U19093 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15877) );
  AOI22_X1 U19094 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15876) );
  NAND4_X1 U19095 ( .A1(n15879), .A2(n15878), .A3(n15877), .A4(n15876), .ZN(
        n15885) );
  AOI22_X1 U19096 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15883) );
  AOI22_X1 U19097 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15882) );
  AOI22_X1 U19098 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15881) );
  AOI22_X1 U19099 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15880) );
  NAND4_X1 U19100 ( .A1(n15883), .A2(n15882), .A3(n15881), .A4(n15880), .ZN(
        n15884) );
  NOR2_X1 U19101 ( .A1(n15885), .A2(n15884), .ZN(n15950) );
  AOI22_X1 U19102 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15889) );
  AOI22_X1 U19103 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15888) );
  AOI22_X1 U19104 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15887) );
  AOI22_X1 U19105 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15886) );
  NAND4_X1 U19106 ( .A1(n15889), .A2(n15888), .A3(n15887), .A4(n15886), .ZN(
        n15895) );
  AOI22_X1 U19107 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15893) );
  AOI22_X1 U19108 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15892) );
  AOI22_X1 U19109 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15891) );
  AOI22_X1 U19110 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15890) );
  NAND4_X1 U19111 ( .A1(n15893), .A2(n15892), .A3(n15891), .A4(n15890), .ZN(
        n15894) );
  NOR2_X1 U19112 ( .A1(n15895), .A2(n15894), .ZN(n17247) );
  AOI22_X1 U19113 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15899) );
  AOI22_X1 U19114 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15898) );
  AOI22_X1 U19115 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15897) );
  AOI22_X1 U19116 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15896) );
  NAND4_X1 U19117 ( .A1(n15899), .A2(n15898), .A3(n15897), .A4(n15896), .ZN(
        n15905) );
  AOI22_X1 U19118 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15903) );
  AOI22_X1 U19119 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15918), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15902) );
  AOI22_X1 U19120 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15901) );
  AOI22_X1 U19121 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15900) );
  NAND4_X1 U19122 ( .A1(n15903), .A2(n15902), .A3(n15901), .A4(n15900), .ZN(
        n15904) );
  NOR2_X1 U19123 ( .A1(n15905), .A2(n15904), .ZN(n17260) );
  AOI22_X1 U19124 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15917) );
  AOI22_X1 U19125 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15916) );
  AOI22_X1 U19126 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15906) );
  OAI21_X1 U19127 ( .B1(n9915), .B2(n15907), .A(n15906), .ZN(n15914) );
  AOI22_X1 U19128 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15912) );
  AOI22_X1 U19129 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15911) );
  AOI22_X1 U19130 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15910) );
  AOI22_X1 U19131 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15909) );
  NAND4_X1 U19132 ( .A1(n15912), .A2(n15911), .A3(n15910), .A4(n15909), .ZN(
        n15913) );
  AOI211_X1 U19133 ( .C1(n17343), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n15914), .B(n15913), .ZN(n15915) );
  NAND3_X1 U19134 ( .A1(n15917), .A2(n15916), .A3(n15915), .ZN(n17265) );
  AOI22_X1 U19135 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15929) );
  AOI22_X1 U19136 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17479), .ZN(n15928) );
  INV_X1 U19137 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n21409) );
  AOI22_X1 U19138 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17460), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15919) );
  OAI21_X1 U19139 ( .B1(n15920), .B2(n21409), .A(n15919), .ZN(n15926) );
  AOI22_X1 U19140 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15924) );
  AOI22_X1 U19141 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17368), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17457), .ZN(n15923) );
  AOI22_X1 U19142 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17459), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15922) );
  AOI22_X1 U19143 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17450), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17472), .ZN(n15921) );
  NAND4_X1 U19144 ( .A1(n15924), .A2(n15923), .A3(n15922), .A4(n15921), .ZN(
        n15925) );
  AOI211_X1 U19145 ( .C1(n15908), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n15926), .B(n15925), .ZN(n15927) );
  NAND3_X1 U19146 ( .A1(n15929), .A2(n15928), .A3(n15927), .ZN(n17266) );
  NAND2_X1 U19147 ( .A1(n17265), .A2(n17266), .ZN(n17264) );
  NOR2_X1 U19148 ( .A1(n17260), .A2(n17264), .ZN(n17259) );
  AOI22_X1 U19149 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15939) );
  AOI22_X1 U19150 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15938) );
  AOI22_X1 U19151 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15930) );
  OAI21_X1 U19152 ( .B1(n9917), .B2(n21467), .A(n15930), .ZN(n15936) );
  AOI22_X1 U19153 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15934) );
  AOI22_X1 U19154 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15933) );
  AOI22_X1 U19155 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15932) );
  AOI22_X1 U19156 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15931) );
  NAND4_X1 U19157 ( .A1(n15934), .A2(n15933), .A3(n15932), .A4(n15931), .ZN(
        n15935) );
  AOI211_X1 U19158 ( .C1(n15908), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n15936), .B(n15935), .ZN(n15937) );
  NAND3_X1 U19159 ( .A1(n15939), .A2(n15938), .A3(n15937), .ZN(n17255) );
  NAND2_X1 U19160 ( .A1(n17259), .A2(n17255), .ZN(n17254) );
  NOR2_X1 U19161 ( .A1(n17247), .A2(n17254), .ZN(n17246) );
  AOI22_X1 U19162 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15949) );
  AOI22_X1 U19163 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15948) );
  AOI22_X1 U19164 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15940) );
  OAI21_X1 U19165 ( .B1(n10390), .B2(n17300), .A(n15940), .ZN(n15946) );
  AOI22_X1 U19166 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15944) );
  AOI22_X1 U19167 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15943) );
  AOI22_X1 U19168 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15942) );
  AOI22_X1 U19169 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15941) );
  NAND4_X1 U19170 ( .A1(n15944), .A2(n15943), .A3(n15942), .A4(n15941), .ZN(
        n15945) );
  AOI211_X1 U19171 ( .C1(n17458), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n15946), .B(n15945), .ZN(n15947) );
  NAND3_X1 U19172 ( .A1(n15949), .A2(n15948), .A3(n15947), .ZN(n17241) );
  NAND2_X1 U19173 ( .A1(n17246), .A2(n17241), .ZN(n17240) );
  NOR2_X1 U19174 ( .A1(n15950), .A2(n17240), .ZN(n17235) );
  AOI21_X1 U19175 ( .B1(n15950), .B2(n17240), .A(n17235), .ZN(n17543) );
  AOI22_X1 U19176 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17236), .B1(n17543), 
        .B2(n17523), .ZN(n15951) );
  OAI21_X1 U19177 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15952), .A(n15951), .ZN(
        P3_U2675) );
  AOI22_X1 U19178 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15957) );
  AOI22_X1 U19179 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15956) );
  AOI22_X1 U19180 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15955) );
  AOI22_X1 U19181 ( .A1(n17432), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15953), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15954) );
  NAND4_X1 U19182 ( .A1(n15957), .A2(n15956), .A3(n15955), .A4(n15954), .ZN(
        n15963) );
  AOI22_X1 U19183 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15961) );
  AOI22_X1 U19184 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15960) );
  AOI22_X1 U19185 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15959) );
  AOI22_X1 U19186 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17459), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15958) );
  NAND4_X1 U19187 ( .A1(n15961), .A2(n15960), .A3(n15959), .A4(n15958), .ZN(
        n15962) );
  NOR2_X1 U19188 ( .A1(n15963), .A2(n15962), .ZN(n17623) );
  AOI21_X1 U19189 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17411), .A(
        P3_EBX_REG_13__SCAN_IN), .ZN(n15965) );
  INV_X1 U19190 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17396) );
  NAND2_X1 U19191 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17411), .ZN(n15964) );
  OAI21_X1 U19192 ( .B1(n17396), .B2(n15964), .A(n17517), .ZN(n17399) );
  OAI22_X1 U19193 ( .A1(n17623), .A2(n17517), .B1(n15965), .B2(n17399), .ZN(
        P3_U2690) );
  NAND2_X1 U19194 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18679) );
  NOR2_X1 U19195 ( .A1(n15966), .A2(n19013), .ZN(n15968) );
  AOI221_X1 U19196 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18679), .C1(n15968), 
        .C2(n18679), .A(n15967), .ZN(n18500) );
  NOR2_X1 U19197 ( .A1(n15969), .A2(n18969), .ZN(n15970) );
  OAI21_X1 U19198 ( .B1(n15970), .B2(n18795), .A(n18501), .ZN(n18498) );
  AOI22_X1 U19199 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18500), .B1(
        n18498), .B2(n18497), .ZN(P3_U2865) );
  NAND2_X1 U19200 ( .A1(n19099), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18507) );
  INV_X1 U19201 ( .A(n18507), .ZN(n15981) );
  NAND2_X1 U19202 ( .A1(n18941), .A2(n19153), .ZN(n15976) );
  NOR2_X1 U19203 ( .A1(n18511), .A2(n17721), .ZN(n18996) );
  INV_X1 U19204 ( .A(n19150), .ZN(n15973) );
  OAI21_X1 U19205 ( .B1(n15974), .B2(n18996), .A(n15973), .ZN(n17682) );
  OAI21_X1 U19206 ( .B1(n15976), .B2(n17682), .A(n15975), .ZN(n15977) );
  AOI211_X1 U19207 ( .C1(n15979), .C2(n15978), .A(n16071), .B(n15977), .ZN(
        n18983) );
  OAI22_X1 U19208 ( .A1(n18983), .A2(n19149), .B1(n16815), .B2(n19101), .ZN(
        n15980) );
  INV_X1 U19209 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15984) );
  NOR2_X1 U19210 ( .A1(n15982), .A2(n18939), .ZN(n18948) );
  NAND3_X1 U19211 ( .A1(n19126), .A2(n19124), .A3(n18948), .ZN(n15983) );
  OAI21_X1 U19212 ( .B1(n19126), .B2(n15984), .A(n15983), .ZN(P3_U3284) );
  INV_X1 U19213 ( .A(n15985), .ZN(n16634) );
  INV_X1 U19214 ( .A(n15986), .ZN(n16633) );
  NOR4_X1 U19215 ( .A1(n16634), .A2(n16633), .A3(n16632), .A4(n20200), .ZN(
        n15987) );
  NAND2_X1 U19216 ( .A1(n15990), .A2(n15987), .ZN(n15988) );
  OAI21_X1 U19217 ( .B1(n15990), .B2(n15989), .A(n15988), .ZN(P2_U3595) );
  INV_X2 U19218 ( .A(n18484), .ZN(n18479) );
  AOI21_X1 U19219 ( .B1(n16684), .B2(n15992), .A(n15991), .ZN(n16687) );
  AOI22_X1 U19220 ( .A1(n18479), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18404), 
        .B2(n16687), .ZN(n15999) );
  OAI22_X1 U19221 ( .A1(n16683), .A2(n18422), .B1(n16681), .B2(n18335), .ZN(
        n16061) );
  INV_X1 U19222 ( .A(n18375), .ZN(n18342) );
  AOI21_X1 U19223 ( .B1(n18342), .B2(n18170), .A(n15993), .ZN(n16707) );
  OAI22_X1 U19224 ( .A1(n18479), .A2(n16707), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18475), .ZN(n15994) );
  OAI21_X1 U19225 ( .B1(n16061), .B2(n15994), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15998) );
  INV_X1 U19226 ( .A(n18306), .ZN(n17964) );
  NAND3_X1 U19227 ( .A1(n9866), .A2(n17964), .A3(n16710), .ZN(n15995) );
  OAI211_X1 U19228 ( .C1(n18335), .C2(n18179), .A(n15996), .B(n15995), .ZN(
        n16059) );
  NAND3_X1 U19229 ( .A1(n16682), .A2(n16684), .A3(n16059), .ZN(n15997) );
  NAND3_X1 U19230 ( .A1(n15999), .A2(n15998), .A3(n15997), .ZN(P3_U2833) );
  INV_X1 U19231 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20171) );
  OAI22_X1 U19232 ( .A1(n16000), .A2(n19351), .B1(n20171), .B2(n19349), .ZN(
        n16001) );
  INV_X1 U19233 ( .A(n16001), .ZN(n16009) );
  AOI22_X1 U19234 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19368), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19356), .ZN(n16008) );
  OAI22_X1 U19235 ( .A1(n16002), .A2(n19343), .B1(n16463), .B2(n19371), .ZN(
        n16003) );
  INV_X1 U19236 ( .A(n16003), .ZN(n16007) );
  OAI211_X1 U19237 ( .C1(n16488), .C2(n16005), .A(n20102), .B(n16004), .ZN(
        n16006) );
  NAND4_X1 U19238 ( .A1(n16009), .A2(n16008), .A3(n16007), .A4(n16006), .ZN(
        P2_U2833) );
  NOR2_X1 U19239 ( .A1(n16010), .A2(n16046), .ZN(n16053) );
  OAI211_X1 U19240 ( .C1(n10273), .C2(n16012), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16011), .ZN(n16016) );
  INV_X1 U19241 ( .A(n16013), .ZN(n16015) );
  OAI211_X1 U19242 ( .C1(n20850), .C2(n16016), .A(n16015), .B(n16014), .ZN(
        n16018) );
  NAND2_X1 U19243 ( .A1(n20850), .A2(n16016), .ZN(n16017) );
  NAND2_X1 U19244 ( .A1(n16018), .A2(n16017), .ZN(n16020) );
  INV_X1 U19245 ( .A(n16020), .ZN(n16022) );
  AOI21_X1 U19246 ( .B1(n16020), .B2(n20922), .A(n16019), .ZN(n16021) );
  AOI21_X1 U19247 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16022), .A(
        n16021), .ZN(n16027) );
  INV_X1 U19248 ( .A(n16027), .ZN(n16024) );
  INV_X1 U19249 ( .A(n16026), .ZN(n16023) );
  AOI21_X1 U19250 ( .B1(n16024), .B2(n16023), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16025) );
  AOI21_X1 U19251 ( .B1(n16027), .B2(n16026), .A(n16025), .ZN(n16035) );
  INV_X1 U19252 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n16029) );
  AOI21_X1 U19253 ( .B1(n16029), .B2(n13780), .A(n16028), .ZN(n16031) );
  NOR4_X1 U19254 ( .A1(n16042), .A2(n16032), .A3(n16031), .A4(n16030), .ZN(
        n16034) );
  OAI211_X1 U19255 ( .C1(n16035), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n16034), .B(n16033), .ZN(n16048) );
  INV_X1 U19256 ( .A(n16049), .ZN(n21120) );
  NAND3_X1 U19257 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21132), .A3(n20500), 
        .ZN(n16036) );
  AOI22_X1 U19258 ( .A1(n16038), .A2(n16037), .B1(n21120), .B2(n16036), .ZN(
        n16371) );
  INV_X1 U19259 ( .A(n16371), .ZN(n16039) );
  AOI221_X1 U19260 ( .B1(n16040), .B2(n20500), .C1(n16040), .C2(n16048), .A(
        n16039), .ZN(n16041) );
  INV_X1 U19261 ( .A(n16041), .ZN(n16377) );
  NAND2_X1 U19262 ( .A1(n16377), .A2(n20500), .ZN(n16052) );
  INV_X1 U19263 ( .A(n16042), .ZN(n16044) );
  NAND3_X1 U19264 ( .A1(n16045), .A2(n16044), .A3(n16043), .ZN(n21211) );
  OAI211_X1 U19265 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21224), .A(n21211), 
        .B(n16046), .ZN(n16047) );
  AOI21_X1 U19266 ( .B1(n16049), .B2(n16048), .A(n16047), .ZN(n16050) );
  AND2_X1 U19267 ( .A1(n16377), .A2(n16050), .ZN(n16051) );
  OAI22_X1 U19268 ( .A1(n16053), .A2(n16052), .B1(n16051), .B2(n20500), .ZN(
        P1_U3161) );
  NAND2_X1 U19269 ( .A1(n16055), .A2(n16054), .ZN(n16057) );
  XOR2_X1 U19270 ( .A(n16057), .B(n16056), .Z(n16680) );
  NOR2_X1 U19271 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16058), .ZN(
        n16676) );
  AOI22_X1 U19272 ( .A1(n18479), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16676), 
        .B2(n16059), .ZN(n16064) );
  INV_X1 U19273 ( .A(n16060), .ZN(n16062) );
  OAI21_X1 U19274 ( .B1(n16062), .B2(n16061), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16063) );
  OAI211_X1 U19275 ( .C1(n16680), .C2(n18390), .A(n16064), .B(n16063), .ZN(
        P3_U2832) );
  INV_X1 U19276 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21128) );
  INV_X1 U19277 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21452) );
  NOR2_X1 U19278 ( .A1(n21136), .A2(n21452), .ZN(n21131) );
  INV_X1 U19279 ( .A(HOLD), .ZN(n20118) );
  NOR2_X1 U19280 ( .A1(n21128), .A2(n20118), .ZN(n21124) );
  INV_X1 U19281 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21137) );
  OAI22_X1 U19282 ( .A1(n21131), .A2(n21124), .B1(n21137), .B2(n20118), .ZN(
        n16065) );
  OAI211_X1 U19283 ( .C1(n21224), .C2(n21128), .A(n16066), .B(n16065), .ZN(
        P1_U3195) );
  INV_X1 U19284 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16717) );
  NOR2_X1 U19285 ( .A1(n20379), .A2(n16717), .ZN(P1_U2905) );
  NAND2_X1 U19286 ( .A1(n20108), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20099) );
  AND2_X1 U19287 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20217) );
  AOI21_X1 U19288 ( .B1(n16656), .B2(n20217), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16067) );
  OAI21_X1 U19289 ( .B1(n15818), .B2(n20099), .A(n16067), .ZN(n16068) );
  AND2_X1 U19290 ( .A1(n16668), .A2(n16068), .ZN(P2_U3178) );
  OAI221_X1 U19291 ( .B1(n19174), .B2(n16668), .C1(n20236), .C2(n16668), .A(
        n19981), .ZN(n20232) );
  NOR2_X1 U19292 ( .A1(n21356), .A2(n20232), .ZN(P2_U3047) );
  INV_X1 U19293 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21494) );
  NOR3_X1 U19294 ( .A1(n16069), .A2(n17683), .A3(n18511), .ZN(n16070) );
  NOR2_X1 U19295 ( .A1(n18545), .A2(n17674), .ZN(n17677) );
  INV_X1 U19296 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18503) );
  OAI22_X1 U19297 ( .A1(n17673), .A2(n18503), .B1(n17680), .B2(n18163), .ZN(
        n16073) );
  AOI221_X1 U19298 ( .B1(n21494), .B2(n17677), .C1(P3_EAX_REG_0__SCAN_IN), 
        .C2(n17674), .A(n16073), .ZN(n16074) );
  INV_X1 U19299 ( .A(n16074), .ZN(P3_U2735) );
  INV_X1 U19300 ( .A(n16087), .ZN(n16075) );
  NAND2_X1 U19301 ( .A1(n16076), .A2(n16075), .ZN(n16077) );
  NAND2_X1 U19302 ( .A1(n20324), .A2(n16077), .ZN(n16100) );
  NAND2_X1 U19303 ( .A1(n16078), .A2(n16091), .ZN(n16088) );
  AOI21_X1 U19304 ( .B1(n16100), .B2(n16088), .A(n14934), .ZN(n16082) );
  OAI22_X1 U19305 ( .A1(n16080), .A2(P1_REIP_REG_22__SCAN_IN), .B1(n16079), 
        .B2(n20330), .ZN(n16081) );
  AOI211_X1 U19306 ( .C1(n20351), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16082), .B(n16081), .ZN(n16086) );
  AOI22_X1 U19307 ( .A1(n16084), .A2(n20307), .B1(n16083), .B2(n20350), .ZN(
        n16085) );
  OAI211_X1 U19308 ( .C1(n20301), .C2(n16233), .A(n16086), .B(n16085), .ZN(
        P1_U2818) );
  AOI22_X1 U19309 ( .A1(n20344), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20351), .ZN(n16090) );
  OR2_X1 U19310 ( .A1(n16088), .A2(n16087), .ZN(n16089) );
  OAI211_X1 U19311 ( .C1(n16100), .C2(n16091), .A(n16090), .B(n16089), .ZN(
        n16092) );
  INV_X1 U19312 ( .A(n16092), .ZN(n16097) );
  INV_X1 U19313 ( .A(n16093), .ZN(n16094) );
  AOI22_X1 U19314 ( .A1(n16095), .A2(n20307), .B1(n16094), .B2(n20345), .ZN(
        n16096) );
  OAI211_X1 U19315 ( .C1(n16098), .C2(n20333), .A(n16097), .B(n16096), .ZN(
        P1_U2819) );
  AOI22_X1 U19316 ( .A1(n20344), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n20350), 
        .B2(n16099), .ZN(n16106) );
  INV_X1 U19317 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n16110) );
  NOR2_X1 U19318 ( .A1(n16110), .A2(n21160), .ZN(n16109) );
  AOI21_X1 U19319 ( .B1(n16109), .B2(n16112), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n16101) );
  OAI22_X1 U19320 ( .A1(n16102), .A2(n20294), .B1(n16101), .B2(n16100), .ZN(
        n16103) );
  AOI21_X1 U19321 ( .B1(n20345), .B2(n16104), .A(n16103), .ZN(n16105) );
  OAI211_X1 U19322 ( .C1(n16107), .C2(n20342), .A(n16106), .B(n16105), .ZN(
        P1_U2820) );
  INV_X1 U19323 ( .A(n16108), .ZN(n16168) );
  AOI21_X1 U19324 ( .B1(n16110), .B2(n21160), .A(n16109), .ZN(n16111) );
  AOI22_X1 U19325 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n16119), .B1(n16112), 
        .B2(n16111), .ZN(n16115) );
  OAI21_X1 U19326 ( .B1(n20342), .B2(n10975), .A(n20447), .ZN(n16113) );
  AOI21_X1 U19327 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(n20344), .A(n16113), .ZN(
        n16114) );
  OAI211_X1 U19328 ( .C1(n20301), .C2(n16243), .A(n16115), .B(n16114), .ZN(
        n16116) );
  AOI21_X1 U19329 ( .B1(n16168), .B2(n20307), .A(n16116), .ZN(n16117) );
  OAI21_X1 U19330 ( .B1(n16171), .B2(n20333), .A(n16117), .ZN(P1_U2821) );
  AOI22_X1 U19331 ( .A1(n20344), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20351), .ZN(n16124) );
  AOI21_X1 U19332 ( .B1(n20350), .B2(n16177), .A(n20487), .ZN(n16123) );
  INV_X1 U19333 ( .A(n16254), .ZN(n16118) );
  AOI22_X1 U19334 ( .A1(n16178), .A2(n20307), .B1(n20345), .B2(n16118), .ZN(
        n16122) );
  OAI221_X1 U19335 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n16120), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(n16135), .A(n16119), .ZN(n16121) );
  NAND4_X1 U19336 ( .A1(n16124), .A2(n16123), .A3(n16122), .A4(n16121), .ZN(
        P1_U2823) );
  AOI21_X1 U19337 ( .B1(n16146), .B2(n16125), .A(n21158), .ZN(n16131) );
  NAND2_X1 U19338 ( .A1(n16126), .A2(n20350), .ZN(n16129) );
  NAND2_X1 U19339 ( .A1(n20344), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n16128) );
  NAND2_X1 U19340 ( .A1(n20351), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16127) );
  NAND4_X1 U19341 ( .A1(n16129), .A2(n16128), .A3(n20447), .A4(n16127), .ZN(
        n16130) );
  NOR2_X1 U19342 ( .A1(n16131), .A2(n16130), .ZN(n16132) );
  OAI21_X1 U19343 ( .B1(n16133), .B2(n20294), .A(n16132), .ZN(n16134) );
  INV_X1 U19344 ( .A(n16134), .ZN(n16137) );
  NAND3_X1 U19345 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n16135), .A3(n21158), 
        .ZN(n16136) );
  OAI211_X1 U19346 ( .C1(n16261), .C2(n20301), .A(n16137), .B(n16136), .ZN(
        P1_U2824) );
  AOI21_X1 U19347 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n16138), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n16145) );
  OAI22_X1 U19348 ( .A1(n16277), .A2(n20301), .B1(n21404), .B2(n20330), .ZN(
        n16139) );
  AOI211_X1 U19349 ( .C1(n20351), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20487), .B(n16139), .ZN(n16144) );
  INV_X1 U19350 ( .A(n16140), .ZN(n16141) );
  AOI22_X1 U19351 ( .A1(n16142), .A2(n20307), .B1(n16141), .B2(n20350), .ZN(
        n16143) );
  OAI211_X1 U19352 ( .C1(n16146), .C2(n16145), .A(n16144), .B(n16143), .ZN(
        P1_U2826) );
  OAI21_X1 U19353 ( .B1(n20342), .B2(n16147), .A(n20447), .ZN(n16149) );
  NOR2_X1 U19354 ( .A1(n16300), .A2(n20301), .ZN(n16148) );
  AOI211_X1 U19355 ( .C1(n20344), .C2(P1_EBX_REG_12__SCAN_IN), .A(n16149), .B(
        n16148), .ZN(n16154) );
  OAI21_X1 U19356 ( .B1(n16150), .B2(n20279), .A(n21152), .ZN(n16151) );
  AOI22_X1 U19357 ( .A1(n16190), .A2(n20350), .B1(n16152), .B2(n16151), .ZN(
        n16153) );
  OAI211_X1 U19358 ( .C1(n20294), .C2(n16193), .A(n16154), .B(n16153), .ZN(
        P1_U2828) );
  INV_X1 U19359 ( .A(n16155), .ZN(n16156) );
  NOR3_X1 U19360 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n20279), .A3(n16156), 
        .ZN(n16160) );
  INV_X1 U19361 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16158) );
  AOI22_X1 U19362 ( .A1(n16307), .A2(n20345), .B1(n20344), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n16157) );
  OAI211_X1 U19363 ( .C1(n20342), .C2(n16158), .A(n16157), .B(n20447), .ZN(
        n16159) );
  NOR2_X1 U19364 ( .A1(n16160), .A2(n16159), .ZN(n16163) );
  AOI22_X1 U19365 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n16161), .B1(n20307), 
        .B2(n16198), .ZN(n16162) );
  OAI211_X1 U19366 ( .C1(n16201), .C2(n20333), .A(n16163), .B(n16162), .ZN(
        P1_U2829) );
  AOI22_X1 U19367 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16170) );
  NAND2_X1 U19368 ( .A1(n16165), .A2(n16164), .ZN(n16167) );
  XOR2_X1 U19369 ( .A(n16167), .B(n16166), .Z(n16240) );
  AOI22_X1 U19370 ( .A1(n16240), .A2(n20435), .B1(n16214), .B2(n16168), .ZN(
        n16169) );
  OAI211_X1 U19371 ( .C1(n16219), .C2(n16171), .A(n16170), .B(n16169), .ZN(
        P1_U2980) );
  NAND2_X1 U19372 ( .A1(n16173), .A2(n16172), .ZN(n16175) );
  NOR2_X1 U19373 ( .A1(n16175), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16174) );
  MUX2_X1 U19374 ( .A(n16175), .B(n16174), .S(n16194), .Z(n16176) );
  XNOR2_X1 U19375 ( .A(n16176), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16255) );
  AOI22_X1 U19376 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16180) );
  AOI22_X1 U19377 ( .A1(n16178), .A2(n16214), .B1(n16177), .B2(n16189), .ZN(
        n16179) );
  OAI211_X1 U19378 ( .C1(n20258), .C2(n16255), .A(n16180), .B(n16179), .ZN(
        P1_U2982) );
  AOI22_X1 U19379 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16184) );
  AOI22_X1 U19380 ( .A1(n16182), .A2(n16214), .B1(n16189), .B2(n16181), .ZN(
        n16183) );
  OAI211_X1 U19381 ( .C1(n16185), .C2(n20258), .A(n16184), .B(n16183), .ZN(
        P1_U2984) );
  AOI22_X1 U19382 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16192) );
  OAI21_X1 U19383 ( .B1(n16188), .B2(n16187), .A(n16186), .ZN(n16302) );
  AOI22_X1 U19384 ( .A1(n16302), .A2(n20435), .B1(n16190), .B2(n16189), .ZN(
        n16191) );
  OAI211_X1 U19385 ( .C1(n20496), .C2(n16193), .A(n16192), .B(n16191), .ZN(
        P1_U2987) );
  AOI22_X1 U19386 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16200) );
  NOR3_X1 U19387 ( .A1(n14975), .A2(n16194), .A3(n16325), .ZN(n16196) );
  NOR2_X1 U19388 ( .A1(n16196), .A2(n16195), .ZN(n16197) );
  XNOR2_X1 U19389 ( .A(n16197), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16310) );
  AOI22_X1 U19390 ( .A1(n20435), .A2(n16310), .B1(n16214), .B2(n16198), .ZN(
        n16199) );
  OAI211_X1 U19391 ( .C1(n16219), .C2(n16201), .A(n16200), .B(n16199), .ZN(
        P1_U2988) );
  AOI22_X1 U19392 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16207) );
  XNOR2_X1 U19393 ( .A(n16202), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16203) );
  XNOR2_X1 U19394 ( .A(n16204), .B(n16203), .ZN(n16347) );
  AOI22_X1 U19395 ( .A1(n16347), .A2(n20435), .B1(n16214), .B2(n16205), .ZN(
        n16206) );
  OAI211_X1 U19396 ( .C1(n16219), .C2(n16208), .A(n16207), .B(n16206), .ZN(
        P1_U2992) );
  AOI22_X1 U19397 ( .A1(n16209), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20487), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16216) );
  NAND2_X1 U19398 ( .A1(n16211), .A2(n16210), .ZN(n16212) );
  XNOR2_X1 U19399 ( .A(n16213), .B(n16212), .ZN(n16353) );
  AOI22_X1 U19400 ( .A1(n16353), .A2(n20435), .B1(n16214), .B2(n20308), .ZN(
        n16215) );
  OAI211_X1 U19401 ( .C1(n16219), .C2(n20304), .A(n16216), .B(n16215), .ZN(
        P1_U2993) );
  XNOR2_X1 U19402 ( .A(n16218), .B(n16217), .ZN(n16359) );
  OAI222_X1 U19403 ( .A1(n16219), .A2(n20328), .B1(n16359), .B2(n20258), .C1(
        n20496), .C2(n20322), .ZN(n16220) );
  INV_X1 U19404 ( .A(n16220), .ZN(n16222) );
  INV_X1 U19405 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20302) );
  NOR2_X1 U19406 ( .A1(n20447), .A2(n20302), .ZN(n16362) );
  INV_X1 U19407 ( .A(n16362), .ZN(n16221) );
  OAI211_X1 U19408 ( .C1(n20316), .C2(n20432), .A(n16222), .B(n16221), .ZN(
        P1_U2994) );
  AOI21_X1 U19409 ( .B1(n16225), .B2(n16224), .A(n16223), .ZN(n16226) );
  AOI22_X1 U19410 ( .A1(n20487), .A2(P1_REIP_REG_22__SCAN_IN), .B1(n16227), 
        .B2(n16226), .ZN(n16232) );
  INV_X1 U19411 ( .A(n16228), .ZN(n16230) );
  AOI22_X1 U19412 ( .A1(n16230), .A2(n20489), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16229), .ZN(n16231) );
  OAI211_X1 U19413 ( .C1(n20479), .C2(n16233), .A(n16232), .B(n16231), .ZN(
        P1_U3009) );
  INV_X1 U19414 ( .A(n16234), .ZN(n16236) );
  AOI21_X1 U19415 ( .B1(n16282), .B2(n16236), .A(n16235), .ZN(n16237) );
  AOI22_X1 U19416 ( .A1(n20487), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n16238), 
        .B2(n16237), .ZN(n16242) );
  AOI22_X1 U19417 ( .A1(n16240), .A2(n20489), .B1(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16239), .ZN(n16241) );
  OAI211_X1 U19418 ( .C1(n20479), .C2(n16243), .A(n16242), .B(n16241), .ZN(
        P1_U3012) );
  NAND2_X1 U19419 ( .A1(n16246), .A2(n16268), .ZN(n16251) );
  NOR2_X1 U19420 ( .A1(n16244), .A2(n20449), .ZN(n16248) );
  AOI21_X1 U19421 ( .B1(n20474), .B2(n16252), .A(n16287), .ZN(n16260) );
  OAI22_X1 U19422 ( .A1(n16260), .A2(n16246), .B1(n16245), .B2(n20479), .ZN(
        n16247) );
  AOI21_X1 U19423 ( .B1(n16248), .B2(n14939), .A(n16247), .ZN(n16250) );
  NAND2_X1 U19424 ( .A1(n20487), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16249) );
  OAI211_X1 U19425 ( .C1(n16252), .C2(n16251), .A(n16250), .B(n16249), .ZN(
        P1_U3013) );
  AOI21_X1 U19426 ( .B1(n16253), .B2(n16268), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16259) );
  OAI22_X1 U19427 ( .A1(n16255), .A2(n20449), .B1(n20479), .B2(n16254), .ZN(
        n16256) );
  INV_X1 U19428 ( .A(n16256), .ZN(n16258) );
  NAND2_X1 U19429 ( .A1(n20487), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16257) );
  OAI211_X1 U19430 ( .C1(n16260), .C2(n16259), .A(n16258), .B(n16257), .ZN(
        P1_U3014) );
  OAI22_X1 U19431 ( .A1(n16263), .A2(n16262), .B1(n20479), .B2(n16261), .ZN(
        n16264) );
  AOI21_X1 U19432 ( .B1(n16265), .B2(n20489), .A(n16264), .ZN(n16270) );
  NAND2_X1 U19433 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16267) );
  NAND4_X1 U19434 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16268), .A3(
        n16267), .A4(n16266), .ZN(n16269) );
  OAI211_X1 U19435 ( .C1(n21158), .C2(n20447), .A(n16270), .B(n16269), .ZN(
        P1_U3015) );
  AOI22_X1 U19436 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16287), .B1(
        n20487), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16276) );
  INV_X1 U19437 ( .A(n16271), .ZN(n16274) );
  NAND2_X1 U19438 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16299), .ZN(
        n20471) );
  NAND2_X1 U19439 ( .A1(n16333), .A2(n16336), .ZN(n16358) );
  NOR3_X1 U19440 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16290), .A3(
        n16272), .ZN(n16273) );
  AOI21_X1 U19441 ( .B1(n16274), .B2(n20489), .A(n16273), .ZN(n16275) );
  OAI211_X1 U19442 ( .C1(n20479), .C2(n16277), .A(n16276), .B(n16275), .ZN(
        P1_U3017) );
  INV_X1 U19443 ( .A(n16278), .ZN(n16280) );
  AOI22_X1 U19444 ( .A1(n16280), .A2(n20489), .B1(n20486), .B2(n16279), .ZN(
        n16289) );
  OAI21_X1 U19445 ( .B1(n16283), .B2(n16282), .A(n16281), .ZN(n16286) );
  NOR2_X1 U19446 ( .A1(n20447), .A2(n16284), .ZN(n16285) );
  AOI221_X1 U19447 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16287), 
        .C1(n21526), .C2(n16286), .A(n16285), .ZN(n16288) );
  NAND2_X1 U19448 ( .A1(n16289), .A2(n16288), .ZN(P1_U3018) );
  NAND2_X1 U19449 ( .A1(n16291), .A2(n16352), .ZN(n16306) );
  AOI21_X1 U19450 ( .B1(n16334), .B2(n16291), .A(n16333), .ZN(n16297) );
  INV_X1 U19451 ( .A(n16308), .ZN(n16293) );
  AOI21_X1 U19452 ( .B1(n16294), .B2(n16293), .A(n16292), .ZN(n16296) );
  INV_X1 U19453 ( .A(n20457), .ZN(n16295) );
  OAI21_X1 U19454 ( .B1(n16333), .B2(n20460), .A(n16295), .ZN(n16314) );
  NOR3_X1 U19455 ( .A1(n16297), .A2(n16296), .A3(n16314), .ZN(n16313) );
  INV_X1 U19456 ( .A(n16313), .ZN(n16298) );
  AOI21_X1 U19457 ( .B1(n16299), .B2(n21502), .A(n16298), .ZN(n16304) );
  OAI22_X1 U19458 ( .A1(n16300), .A2(n20479), .B1(n21152), .B2(n20447), .ZN(
        n16301) );
  AOI21_X1 U19459 ( .B1(n16302), .B2(n20489), .A(n16301), .ZN(n16303) );
  OAI221_X1 U19460 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16306), 
        .C1(n16305), .C2(n16304), .A(n16303), .ZN(P1_U3019) );
  AOI22_X1 U19461 ( .A1(n20487), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20486), 
        .B2(n16307), .ZN(n16312) );
  NOR2_X1 U19462 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16308), .ZN(
        n16309) );
  AOI22_X1 U19463 ( .A1(n16310), .A2(n20489), .B1(n16309), .B2(n16352), .ZN(
        n16311) );
  OAI211_X1 U19464 ( .C1(n16313), .C2(n21502), .A(n16312), .B(n16311), .ZN(
        P1_U3020) );
  NAND2_X1 U19465 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16315) );
  AOI21_X1 U19466 ( .B1(n16315), .B2(n20458), .A(n16314), .ZN(n20456) );
  NAND2_X1 U19467 ( .A1(n16318), .A2(n20456), .ZN(n16316) );
  OAI22_X1 U19468 ( .A1(n20474), .A2(n20457), .B1(n16317), .B2(n16316), .ZN(
        n16331) );
  NAND2_X1 U19469 ( .A1(n16318), .A2(n16352), .ZN(n16326) );
  AOI221_X1 U19470 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16325), .C2(n16332), .A(
        n16326), .ZN(n16319) );
  AOI21_X1 U19471 ( .B1(n20487), .B2(P1_REIP_REG_10__SCAN_IN), .A(n16319), 
        .ZN(n16320) );
  OAI21_X1 U19472 ( .B1(n16321), .B2(n20479), .A(n16320), .ZN(n16322) );
  AOI21_X1 U19473 ( .B1(n16323), .B2(n20489), .A(n16322), .ZN(n16324) );
  OAI21_X1 U19474 ( .B1(n16325), .B2(n16331), .A(n16324), .ZN(P1_U3021) );
  NOR2_X1 U19475 ( .A1(n20447), .A2(n20288), .ZN(n16329) );
  OAI22_X1 U19476 ( .A1(n16327), .A2(n20449), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16326), .ZN(n16328) );
  AOI211_X1 U19477 ( .C1(n20486), .C2(n20282), .A(n16329), .B(n16328), .ZN(
        n16330) );
  OAI21_X1 U19478 ( .B1(n16332), .B2(n16331), .A(n16330), .ZN(P1_U3022) );
  OR2_X1 U19479 ( .A1(n20439), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16364) );
  OAI21_X1 U19480 ( .B1(n16334), .B2(n16333), .A(n20456), .ZN(n16335) );
  AOI21_X1 U19481 ( .B1(n20439), .B2(n20458), .A(n16335), .ZN(n16360) );
  OAI21_X1 U19482 ( .B1(n16336), .B2(n16364), .A(n16360), .ZN(n16354) );
  AOI21_X1 U19483 ( .B1(n16337), .B2(n20474), .A(n16354), .ZN(n16349) );
  NAND2_X1 U19484 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16352), .ZN(
        n16351) );
  AOI221_X1 U19485 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16343), .C2(n16350), .A(
        n16351), .ZN(n16341) );
  AND2_X1 U19486 ( .A1(n16338), .A2(n20489), .ZN(n16340) );
  OAI22_X1 U19487 ( .A1(n20300), .A2(n20479), .B1(n14444), .B2(n20447), .ZN(
        n16339) );
  NOR3_X1 U19488 ( .A1(n16341), .A2(n16340), .A3(n16339), .ZN(n16342) );
  OAI21_X1 U19489 ( .B1(n16349), .B2(n16343), .A(n16342), .ZN(P1_U3023) );
  OAI22_X1 U19490 ( .A1(n16345), .A2(n20479), .B1(n16344), .B2(n20447), .ZN(
        n16346) );
  AOI21_X1 U19491 ( .B1(n16347), .B2(n20489), .A(n16346), .ZN(n16348) );
  OAI221_X1 U19492 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16351), .C1(
        n16350), .C2(n16349), .A(n16348), .ZN(P1_U3024) );
  INV_X1 U19493 ( .A(n16352), .ZN(n16357) );
  AOI22_X1 U19494 ( .A1(n20487), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20486), 
        .B2(n20306), .ZN(n16356) );
  AOI22_X1 U19495 ( .A1(n16354), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16353), .B2(n20489), .ZN(n16355) );
  OAI211_X1 U19496 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16357), .A(
        n16356), .B(n16355), .ZN(P1_U3025) );
  NAND2_X1 U19497 ( .A1(n20460), .A2(n16358), .ZN(n20448) );
  OAI22_X1 U19498 ( .A1(n16360), .A2(n11360), .B1(n20449), .B2(n16359), .ZN(
        n16361) );
  AOI211_X1 U19499 ( .C1(n20486), .C2(n20321), .A(n16362), .B(n16361), .ZN(
        n16363) );
  OAI21_X1 U19500 ( .B1(n16364), .B2(n20448), .A(n16363), .ZN(P1_U3026) );
  INV_X1 U19501 ( .A(n20332), .ZN(n16367) );
  NAND4_X1 U19502 ( .A1(n16367), .A2(n21189), .A3(n16366), .A4(n16365), .ZN(
        n16368) );
  OAI21_X1 U19503 ( .B1(n21192), .B2(n14067), .A(n16368), .ZN(P1_U3468) );
  NAND2_X1 U19504 ( .A1(n20931), .A2(n21224), .ZN(n16375) );
  NAND4_X1 U19505 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20980), .A4(n21224), .ZN(n16369) );
  AND2_X1 U19506 ( .A1(n16370), .A2(n16369), .ZN(n21121) );
  AOI21_X1 U19507 ( .B1(n21121), .B2(n16372), .A(n16371), .ZN(n16374) );
  AOI21_X1 U19508 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16377), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16373) );
  AOI211_X1 U19509 ( .C1(n21235), .C2(n16375), .A(n16374), .B(n16373), .ZN(
        P1_U3162) );
  OAI221_X1 U19510 ( .B1(n20931), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20931), 
        .C2(n16377), .A(n16376), .ZN(P1_U3466) );
  AOI22_X1 U19511 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n19368), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n19369), .ZN(n16387) );
  AOI22_X1 U19512 ( .A1(n16378), .A2(n19367), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19356), .ZN(n16386) );
  INV_X1 U19513 ( .A(n16379), .ZN(n19386) );
  AOI22_X1 U19514 ( .A1(n16380), .A2(n19364), .B1(n19275), .B2(n19386), .ZN(
        n16385) );
  INV_X1 U19515 ( .A(n19383), .ZN(n16383) );
  NAND3_X1 U19516 ( .A1(n16383), .A2(n16382), .A3(n16381), .ZN(n16384) );
  NAND4_X1 U19517 ( .A1(n16387), .A2(n16386), .A3(n16385), .A4(n16384), .ZN(
        P2_U2824) );
  AOI22_X1 U19518 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19368), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19369), .ZN(n16399) );
  AOI22_X1 U19519 ( .A1(n16388), .A2(n19367), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19356), .ZN(n16398) );
  INV_X1 U19520 ( .A(n16389), .ZN(n16390) );
  OAI22_X1 U19521 ( .A1(n16391), .A2(n19343), .B1(n16390), .B2(n19371), .ZN(
        n16392) );
  INV_X1 U19522 ( .A(n16392), .ZN(n16397) );
  OAI211_X1 U19523 ( .C1(n16395), .C2(n16394), .A(n20102), .B(n16393), .ZN(
        n16396) );
  NAND4_X1 U19524 ( .A1(n16399), .A2(n16398), .A3(n16397), .A4(n16396), .ZN(
        P2_U2826) );
  AOI22_X1 U19525 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19368), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19369), .ZN(n16412) );
  OAI22_X1 U19526 ( .A1(n16401), .A2(n19351), .B1(n16400), .B2(n19378), .ZN(
        n16402) );
  INV_X1 U19527 ( .A(n16402), .ZN(n16411) );
  INV_X1 U19528 ( .A(n16403), .ZN(n16405) );
  AOI22_X1 U19529 ( .A1(n16405), .A2(n19364), .B1(n16404), .B2(n19275), .ZN(
        n16410) );
  OAI211_X1 U19530 ( .C1(n16408), .C2(n16407), .A(n20102), .B(n16406), .ZN(
        n16409) );
  NAND4_X1 U19531 ( .A1(n16412), .A2(n16411), .A3(n16410), .A4(n16409), .ZN(
        P2_U2828) );
  AOI22_X1 U19532 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19368), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19369), .ZN(n16424) );
  OAI22_X1 U19533 ( .A1(n16413), .A2(n19351), .B1(n10159), .B2(n19378), .ZN(
        n16414) );
  INV_X1 U19534 ( .A(n16414), .ZN(n16423) );
  OAI22_X1 U19535 ( .A1(n16416), .A2(n19343), .B1(n16415), .B2(n19371), .ZN(
        n16417) );
  INV_X1 U19536 ( .A(n16417), .ZN(n16422) );
  OAI211_X1 U19537 ( .C1(n16420), .C2(n16419), .A(n20102), .B(n16418), .ZN(
        n16421) );
  NAND4_X1 U19538 ( .A1(n16424), .A2(n16423), .A3(n16422), .A4(n16421), .ZN(
        P2_U2829) );
  AOI22_X1 U19539 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19368), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19369), .ZN(n16436) );
  AOI22_X1 U19540 ( .A1(n16425), .A2(n19367), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19356), .ZN(n16435) );
  INV_X1 U19541 ( .A(n16426), .ZN(n16427) );
  OAI22_X1 U19542 ( .A1(n16428), .A2(n19343), .B1(n16427), .B2(n19371), .ZN(
        n16429) );
  INV_X1 U19543 ( .A(n16429), .ZN(n16434) );
  OAI211_X1 U19544 ( .C1(n16432), .C2(n16431), .A(n20102), .B(n16430), .ZN(
        n16433) );
  NAND4_X1 U19545 ( .A1(n16436), .A2(n16435), .A3(n16434), .A4(n16433), .ZN(
        P2_U2830) );
  AOI22_X1 U19546 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19368), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19369), .ZN(n16449) );
  INV_X1 U19547 ( .A(n16437), .ZN(n16438) );
  AOI22_X1 U19548 ( .A1(n16438), .A2(n19367), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19356), .ZN(n16448) );
  INV_X1 U19549 ( .A(n16439), .ZN(n16440) );
  OAI22_X1 U19550 ( .A1(n16441), .A2(n19343), .B1(n16440), .B2(n19371), .ZN(
        n16442) );
  INV_X1 U19551 ( .A(n16442), .ZN(n16447) );
  OAI211_X1 U19552 ( .C1(n16445), .C2(n16444), .A(n20102), .B(n16443), .ZN(
        n16446) );
  NAND4_X1 U19553 ( .A1(n16449), .A2(n16448), .A3(n16447), .A4(n16446), .ZN(
        P2_U2831) );
  INV_X1 U19554 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20173) );
  OAI22_X1 U19555 ( .A1(n16450), .A2(n19378), .B1(n20173), .B2(n19349), .ZN(
        n16451) );
  AOI21_X1 U19556 ( .B1(n19368), .B2(P2_EBX_REG_23__SCAN_IN), .A(n16451), .ZN(
        n16452) );
  OAI21_X1 U19557 ( .B1(n16453), .B2(n19343), .A(n16452), .ZN(n16454) );
  AOI21_X1 U19558 ( .B1(n16455), .B2(n19367), .A(n16454), .ZN(n16460) );
  OAI211_X1 U19559 ( .C1(n16458), .C2(n16457), .A(n20102), .B(n16456), .ZN(
        n16459) );
  OAI211_X1 U19560 ( .C1(n16461), .C2(n19371), .A(n16460), .B(n16459), .ZN(
        P2_U2832) );
  AOI22_X1 U19561 ( .A1(n16477), .A2(n16462), .B1(n19442), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16468) );
  AOI22_X1 U19562 ( .A1(n19385), .A2(BUF1_REG_22__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16467) );
  INV_X1 U19563 ( .A(n16463), .ZN(n16464) );
  AOI22_X1 U19564 ( .A1(n16465), .A2(n19444), .B1(n19443), .B2(n16464), .ZN(
        n16466) );
  NAND3_X1 U19565 ( .A1(n16468), .A2(n16467), .A3(n16466), .ZN(P2_U2897) );
  AOI22_X1 U19566 ( .A1(n16477), .A2(n16469), .B1(n19442), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19567 ( .A1(n19385), .A2(BUF1_REG_20__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16474) );
  INV_X1 U19568 ( .A(n16470), .ZN(n16471) );
  AOI22_X1 U19569 ( .A1(n16472), .A2(n19444), .B1(n19443), .B2(n16471), .ZN(
        n16473) );
  NAND3_X1 U19570 ( .A1(n16475), .A2(n16474), .A3(n16473), .ZN(P2_U2899) );
  AOI22_X1 U19571 ( .A1(n16477), .A2(n16476), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19442), .ZN(n16481) );
  AOI22_X1 U19572 ( .A1(n19385), .A2(BUF1_REG_18__SCAN_IN), .B1(n19387), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16480) );
  AOI22_X1 U19573 ( .A1(n16478), .A2(n19444), .B1(n19443), .B2(n19225), .ZN(
        n16479) );
  NAND3_X1 U19574 ( .A1(n16481), .A2(n16480), .A3(n16479), .ZN(P2_U2901) );
  AOI22_X1 U19575 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19247), .ZN(n16487) );
  INV_X1 U19576 ( .A(n16482), .ZN(n16483) );
  AOI222_X1 U19577 ( .A1(n16485), .A2(n19493), .B1(n19494), .B2(n16484), .C1(
        n19495), .C2(n16483), .ZN(n16486) );
  OAI211_X1 U19578 ( .C1(n19499), .C2(n16488), .A(n16487), .B(n16486), .ZN(
        P2_U2992) );
  AOI22_X1 U19579 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19247), .ZN(n16492) );
  AOI222_X1 U19580 ( .A1(n16490), .A2(n19493), .B1(n19495), .B2(n16489), .C1(
        n19494), .C2(n19226), .ZN(n16491) );
  OAI211_X1 U19581 ( .C1(n19499), .C2(n19229), .A(n16492), .B(n16491), .ZN(
        P2_U2996) );
  AOI22_X1 U19582 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19247), .ZN(n16496) );
  AOI222_X1 U19583 ( .A1(n16494), .A2(n19495), .B1(n19493), .B2(n16493), .C1(
        n19494), .C2(n19276), .ZN(n16495) );
  OAI211_X1 U19584 ( .C1(n19499), .C2(n19271), .A(n16496), .B(n16495), .ZN(
        P2_U3000) );
  AOI22_X1 U19585 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19247), .ZN(n16500) );
  AOI222_X1 U19586 ( .A1(n16498), .A2(n19493), .B1(n19494), .B2(n19299), .C1(
        n19495), .C2(n16497), .ZN(n16499) );
  OAI211_X1 U19587 ( .C1(n19499), .C2(n19300), .A(n16500), .B(n16499), .ZN(
        P2_U3002) );
  AOI22_X1 U19588 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19247), .B1(n16550), 
        .B2(n16501), .ZN(n16507) );
  OAI22_X1 U19589 ( .A1(n16503), .A2(n16543), .B1(n16502), .B2(n16541), .ZN(
        n16504) );
  AOI21_X1 U19590 ( .B1(n19494), .B2(n16505), .A(n16504), .ZN(n16506) );
  OAI211_X1 U19591 ( .C1(n16561), .C2(n16508), .A(n16507), .B(n16506), .ZN(
        P2_U3003) );
  AOI22_X1 U19592 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19247), .ZN(n16520) );
  NOR2_X1 U19593 ( .A1(n16510), .A2(n16509), .ZN(n16514) );
  NAND2_X1 U19594 ( .A1(n16512), .A2(n16511), .ZN(n16513) );
  XNOR2_X1 U19595 ( .A(n16514), .B(n16513), .ZN(n16588) );
  INV_X1 U19596 ( .A(n16588), .ZN(n16518) );
  AOI21_X1 U19597 ( .B1(n16517), .B2(n16516), .A(n16515), .ZN(n16584) );
  AOI222_X1 U19598 ( .A1(n16518), .A2(n19493), .B1(n19494), .B2(n19310), .C1(
        n19495), .C2(n16584), .ZN(n16519) );
  OAI211_X1 U19599 ( .C1(n19499), .C2(n19308), .A(n16520), .B(n16519), .ZN(
        P2_U3004) );
  AOI22_X1 U19600 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19247), .B1(n16550), 
        .B2(n19315), .ZN(n16526) );
  OAI22_X1 U19601 ( .A1(n16522), .A2(n16543), .B1(n16541), .B2(n16521), .ZN(
        n16523) );
  AOI21_X1 U19602 ( .B1(n19494), .B2(n16524), .A(n16523), .ZN(n16525) );
  OAI211_X1 U19603 ( .C1(n16561), .C2(n16527), .A(n16526), .B(n16525), .ZN(
        P2_U3005) );
  AOI22_X1 U19604 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19247), .ZN(n16539) );
  AOI21_X1 U19605 ( .B1(n15547), .B2(n16529), .A(n16528), .ZN(n16534) );
  INV_X1 U19606 ( .A(n16530), .ZN(n16531) );
  NOR2_X1 U19607 ( .A1(n16532), .A2(n16531), .ZN(n16533) );
  XNOR2_X1 U19608 ( .A(n16534), .B(n16533), .ZN(n16594) );
  XOR2_X1 U19609 ( .A(n16535), .B(n16536), .Z(n16590) );
  AOI222_X1 U19610 ( .A1(n16594), .A2(n19493), .B1(n19494), .B2(n16537), .C1(
        n16590), .C2(n19495), .ZN(n16538) );
  OAI211_X1 U19611 ( .C1(n19499), .C2(n16540), .A(n16539), .B(n16538), .ZN(
        P2_U3006) );
  AOI22_X1 U19612 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19247), .B1(n16550), 
        .B2(n19359), .ZN(n16547) );
  OAI22_X1 U19613 ( .A1(n16544), .A2(n16543), .B1(n16542), .B2(n16541), .ZN(
        n16545) );
  AOI21_X1 U19614 ( .B1(n19494), .B2(n19360), .A(n16545), .ZN(n16546) );
  OAI211_X1 U19615 ( .C1(n16561), .C2(n16548), .A(n16547), .B(n16546), .ZN(
        P2_U3009) );
  AOI22_X1 U19616 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19247), .B1(n16550), 
        .B2(n16549), .ZN(n16560) );
  NAND2_X1 U19617 ( .A1(n16552), .A2(n16551), .ZN(n16554) );
  XNOR2_X1 U19618 ( .A(n16554), .B(n16553), .ZN(n16608) );
  OAI21_X1 U19619 ( .B1(n16557), .B2(n16556), .A(n16555), .ZN(n16605) );
  INV_X1 U19620 ( .A(n16605), .ZN(n16558) );
  AOI222_X1 U19621 ( .A1(n16608), .A2(n19493), .B1(n19495), .B2(n16558), .C1(
        n16601), .C2(n19494), .ZN(n16559) );
  OAI211_X1 U19622 ( .C1(n16562), .C2(n16561), .A(n16560), .B(n16559), .ZN(
        P2_U3011) );
  NOR2_X1 U19623 ( .A1(n16564), .A2(n16563), .ZN(n16571) );
  OR2_X1 U19624 ( .A1(n16565), .A2(n15730), .ZN(n16567) );
  NAND2_X1 U19625 ( .A1(n16567), .A2(n16566), .ZN(n19391) );
  OAI22_X1 U19626 ( .A1(n16603), .A2(n19391), .B1(n20158), .B2(n19348), .ZN(
        n16568) );
  AOI221_X1 U19627 ( .B1(n16571), .B2(n16570), .C1(n16569), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n16568), .ZN(n16576) );
  INV_X1 U19628 ( .A(n16572), .ZN(n16574) );
  AOI22_X1 U19629 ( .A1(n16574), .A2(n12862), .B1(n19500), .B2(n16573), .ZN(
        n16575) );
  OAI211_X1 U19630 ( .C1(n16577), .C2(n16587), .A(n16576), .B(n16575), .ZN(
        P2_U3031) );
  INV_X1 U19631 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20148) );
  NOR2_X1 U19632 ( .A1(n20148), .A2(n19348), .ZN(n16582) );
  XNOR2_X1 U19633 ( .A(n16579), .B(n16578), .ZN(n19405) );
  OAI22_X1 U19634 ( .A1(n16603), .A2(n19405), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16580), .ZN(n16581) );
  AOI211_X1 U19635 ( .C1(n16583), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16582), .B(n16581), .ZN(n16586) );
  AOI22_X1 U19636 ( .A1(n16584), .A2(n12862), .B1(n19500), .B2(n19310), .ZN(
        n16585) );
  OAI211_X1 U19637 ( .C1(n16588), .C2(n16587), .A(n16586), .B(n16585), .ZN(
        P2_U3036) );
  AOI22_X1 U19638 ( .A1(n16589), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19517), .B2(n19408), .ZN(n16600) );
  INV_X1 U19639 ( .A(n16590), .ZN(n16592) );
  OAI22_X1 U19640 ( .A1(n16592), .A2(n16604), .B1(n19534), .B2(n16591), .ZN(
        n16593) );
  AOI21_X1 U19641 ( .B1(n19526), .B2(n16594), .A(n16593), .ZN(n16599) );
  NAND2_X1 U19642 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19247), .ZN(n16598) );
  OAI221_X1 U19643 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n12265), .C2(n16596), .A(
        n16595), .ZN(n16597) );
  NAND4_X1 U19644 ( .A1(n16600), .A2(n16599), .A3(n16598), .A4(n16597), .ZN(
        P2_U3038) );
  AOI22_X1 U19645 ( .A1(n16601), .A2(n19500), .B1(P2_REIP_REG_3__SCAN_IN), 
        .B2(n19247), .ZN(n16602) );
  OAI21_X1 U19646 ( .B1(n19429), .B2(n16603), .A(n16602), .ZN(n16607) );
  NOR2_X1 U19647 ( .A1(n16605), .A2(n16604), .ZN(n16606) );
  AOI211_X1 U19648 ( .C1(n16608), .C2(n19526), .A(n16607), .B(n16606), .ZN(
        n16609) );
  OAI221_X1 U19649 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16612), .C1(
        n16611), .C2(n16610), .A(n16609), .ZN(P2_U3043) );
  NAND2_X1 U19650 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19913), .ZN(n20100) );
  INV_X1 U19651 ( .A(n16624), .ZN(n16613) );
  NAND2_X1 U19652 ( .A1(n16613), .A2(n16628), .ZN(n16614) );
  OAI21_X1 U19653 ( .B1(n16615), .B2(n16628), .A(n16614), .ZN(n16648) );
  MUX2_X1 U19654 ( .A(n16617), .B(n16616), .S(n16628), .Z(n16647) );
  OAI22_X1 U19655 ( .A1(n16648), .A2(n19620), .B1(n16647), .B2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16627) );
  INV_X1 U19656 ( .A(n16618), .ZN(n16619) );
  OAI21_X1 U19657 ( .B1(n16619), .B2(n20233), .A(n21540), .ZN(n16621) );
  OAI21_X1 U19658 ( .B1(n16619), .B2(n19907), .A(n16628), .ZN(n16620) );
  AOI21_X1 U19659 ( .B1(n16622), .B2(n16621), .A(n16620), .ZN(n16623) );
  OAI21_X1 U19660 ( .B1(n16624), .B2(n21487), .A(n16623), .ZN(n16625) );
  AOI21_X1 U19661 ( .B1(n16647), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16625), .ZN(n16626) );
  OAI21_X1 U19662 ( .B1(n16627), .B2(n16626), .A(n21356), .ZN(n16646) );
  INV_X1 U19663 ( .A(n16628), .ZN(n16644) );
  INV_X1 U19664 ( .A(n12463), .ZN(n16631) );
  NOR4_X1 U19665 ( .A1(n16638), .A2(n16631), .A3(n16630), .A4(n16629), .ZN(
        n19172) );
  OAI21_X1 U19666 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n19172), .ZN(n16636) );
  OR3_X1 U19667 ( .A1(n16634), .A2(n16633), .A3(n16632), .ZN(n16635) );
  OAI211_X1 U19668 ( .C1(n16637), .C2(n12180), .A(n16636), .B(n16635), .ZN(
        n16643) );
  AOI22_X1 U19669 ( .A1(n16642), .A2(n16639), .B1(n12463), .B2(n16638), .ZN(
        n16640) );
  OAI21_X1 U19670 ( .B1(n16642), .B2(n16641), .A(n16640), .ZN(n20241) );
  AOI211_X1 U19671 ( .C1(n16644), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16643), .B(n20241), .ZN(n16645) );
  OAI211_X1 U19672 ( .C1(n16648), .C2(n16647), .A(n16646), .B(n16645), .ZN(
        n16664) );
  NAND2_X1 U19673 ( .A1(n16650), .A2(n16649), .ZN(n20226) );
  OAI21_X1 U19674 ( .B1(n16664), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16655) );
  NAND2_X1 U19675 ( .A1(n16651), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16652) );
  AOI21_X1 U19676 ( .B1(n16654), .B2(n16653), .A(n16652), .ZN(n16657) );
  NAND2_X1 U19677 ( .A1(n16655), .A2(n16657), .ZN(n20104) );
  AOI21_X1 U19678 ( .B1(n20226), .B2(n20104), .A(n16656), .ZN(n16663) );
  NAND2_X1 U19679 ( .A1(n15818), .A2(n19913), .ZN(n16659) );
  AOI21_X1 U19680 ( .B1(n16657), .B2(n20124), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16658) );
  OAI21_X1 U19681 ( .B1(n16660), .B2(n16659), .A(n16658), .ZN(n16661) );
  INV_X1 U19682 ( .A(n16661), .ZN(n16662) );
  AOI211_X1 U19683 ( .C1(n16665), .C2(n16664), .A(n16663), .B(n16662), .ZN(
        n16667) );
  OAI211_X1 U19684 ( .C1(n20108), .C2(n20100), .A(n16667), .B(n16666), .ZN(
        P2_U3176) );
  OAI221_X1 U19685 ( .B1(n19873), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n16669), 
        .C2(n20104), .A(n16668), .ZN(P2_U3593) );
  AOI22_X1 U19686 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16688), .B1(
        n16670), .B2(n16673), .ZN(n16860) );
  AOI21_X1 U19687 ( .B1(n16673), .B2(n16672), .A(n16671), .ZN(n16675) );
  INV_X1 U19688 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21437) );
  NOR2_X1 U19689 ( .A1(n18484), .A2(n21437), .ZN(n16674) );
  AOI211_X1 U19690 ( .C1(n18006), .C2(n16860), .A(n16675), .B(n16674), .ZN(
        n16679) );
  OAI22_X1 U19691 ( .A1(n16681), .A2(n18025), .B1(n16683), .B2(n13159), .ZN(
        n16677) );
  OAI22_X1 U19692 ( .A1(n18025), .A2(n18305), .B1(n13159), .B2(n18306), .ZN(
        n17951) );
  NOR3_X1 U19693 ( .A1(n17931), .A2(n18186), .A3(n18187), .ZN(n17814) );
  AOI22_X1 U19694 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16677), .B1(
        n16676), .B2(n17814), .ZN(n16678) );
  OAI211_X1 U19695 ( .C1(n16680), .C2(n18057), .A(n16679), .B(n16678), .ZN(
        P3_U2800) );
  NAND2_X1 U19696 ( .A1(n17791), .A2(n16682), .ZN(n16704) );
  AOI211_X1 U19697 ( .C1(n16684), .C2(n16704), .A(n16681), .B(n18025), .ZN(
        n16686) );
  NAND2_X1 U19698 ( .A1(n16682), .A2(n18177), .ZN(n16705) );
  AOI211_X1 U19699 ( .C1(n16684), .C2(n16705), .A(n16683), .B(n13159), .ZN(
        n16685) );
  AOI211_X1 U19700 ( .C1(n16687), .C2(n18069), .A(n16686), .B(n16685), .ZN(
        n16695) );
  NAND2_X1 U19701 ( .A1(n18479), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16694) );
  AOI21_X1 U19702 ( .B1(n10167), .B2(n16689), .A(n16688), .ZN(n16870) );
  OAI21_X1 U19703 ( .B1(n16690), .B2(n18006), .A(n16870), .ZN(n16693) );
  OAI221_X1 U19704 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18883), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n9983), .A(n16691), .ZN(n16692) );
  NAND4_X1 U19705 ( .A1(n16695), .A2(n16694), .A3(n16693), .A4(n16692), .ZN(
        P3_U2801) );
  AOI21_X1 U19706 ( .B1(n17806), .B2(n18068), .A(n16696), .ZN(n17796) );
  INV_X1 U19707 ( .A(n17796), .ZN(n16697) );
  NOR2_X1 U19708 ( .A1(n16698), .A2(n16697), .ZN(n16700) );
  OAI21_X1 U19709 ( .B1(n18068), .B2(n17792), .A(n16698), .ZN(n16701) );
  NOR3_X1 U19710 ( .A1(n17807), .A2(n18390), .A3(n16701), .ZN(n16699) );
  AOI21_X1 U19711 ( .B1(n16700), .B2(n18487), .A(n16699), .ZN(n16713) );
  INV_X1 U19712 ( .A(n16701), .ZN(n17795) );
  NOR2_X1 U19713 ( .A1(n17796), .A2(n17795), .ZN(n17794) );
  NOR2_X1 U19714 ( .A1(n16703), .A2(n18942), .ZN(n18361) );
  AOI22_X1 U19715 ( .A1(n9866), .A2(n16705), .B1(n18361), .B2(n16704), .ZN(
        n16706) );
  NAND2_X1 U19716 ( .A1(n16707), .A2(n16706), .ZN(n16708) );
  OAI211_X1 U19717 ( .C1(n16709), .C2(n16708), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18484), .ZN(n16712) );
  NAND2_X1 U19718 ( .A1(n18479), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17803) );
  INV_X1 U19719 ( .A(n18361), .ZN(n18340) );
  OAI22_X1 U19720 ( .A1(n18227), .A2(n18306), .B1(n18305), .B2(n18340), .ZN(
        n18275) );
  INV_X1 U19721 ( .A(n18246), .ZN(n18236) );
  NAND4_X1 U19722 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16710), .A3(
        n17792), .A4(n18236), .ZN(n16711) );
  NAND4_X1 U19723 ( .A1(n16713), .A2(n16712), .A3(n17803), .A4(n16711), .ZN(
        P3_U2834) );
  NOR3_X1 U19724 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16715) );
  NOR4_X1 U19725 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16714) );
  NAND4_X1 U19726 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16715), .A3(n16714), .A4(
        U215), .ZN(U213) );
  INV_X1 U19727 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16799) );
  INV_X2 U19728 ( .A(U214), .ZN(n16760) );
  NOR2_X1 U19729 ( .A1(n16760), .A2(n16716), .ZN(n16767) );
  OAI222_X1 U19730 ( .A1(U212), .A2(n16799), .B1(n16764), .B2(n16718), .C1(
        U214), .C2(n16717), .ZN(U216) );
  INV_X1 U19731 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19556) );
  AOI22_X1 U19732 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16759), .ZN(n16719) );
  OAI21_X1 U19733 ( .B1(n19556), .B2(n16764), .A(n16719), .ZN(U217) );
  AOI222_X1 U19734 ( .A1(n16759), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(n16767), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n16760), .C2(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n16720) );
  INV_X1 U19735 ( .A(n16720), .ZN(U218) );
  INV_X1 U19736 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16722) );
  AOI22_X1 U19737 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16759), .ZN(n16721) );
  OAI21_X1 U19738 ( .B1(n16722), .B2(n16764), .A(n16721), .ZN(U219) );
  AOI22_X1 U19739 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16759), .ZN(n16723) );
  OAI21_X1 U19740 ( .B1(n16724), .B2(n16764), .A(n16723), .ZN(U220) );
  AOI22_X1 U19741 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16759), .ZN(n16725) );
  OAI21_X1 U19742 ( .B1(n16726), .B2(n16764), .A(n16725), .ZN(U221) );
  AOI22_X1 U19743 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16759), .ZN(n16727) );
  OAI21_X1 U19744 ( .B1(n16728), .B2(n16764), .A(n16727), .ZN(U222) );
  INV_X1 U19745 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16730) );
  AOI22_X1 U19746 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16759), .ZN(n16729) );
  OAI21_X1 U19747 ( .B1(n16730), .B2(n16764), .A(n16729), .ZN(U223) );
  AOI22_X1 U19748 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16759), .ZN(n16731) );
  OAI21_X1 U19749 ( .B1(n16732), .B2(n16764), .A(n16731), .ZN(U224) );
  INV_X1 U19750 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19562) );
  AOI22_X1 U19751 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16759), .ZN(n16733) );
  OAI21_X1 U19752 ( .B1(n19562), .B2(n16764), .A(n16733), .ZN(U225) );
  AOI22_X1 U19753 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16759), .ZN(n16734) );
  OAI21_X1 U19754 ( .B1(n15358), .B2(n16764), .A(n16734), .ZN(U226) );
  INV_X1 U19755 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16736) );
  AOI22_X1 U19756 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16759), .ZN(n16735) );
  OAI21_X1 U19757 ( .B1(n16736), .B2(n16764), .A(n16735), .ZN(U227) );
  INV_X1 U19758 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16738) );
  AOI22_X1 U19759 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16759), .ZN(n16737) );
  OAI21_X1 U19760 ( .B1(n16738), .B2(n16764), .A(n16737), .ZN(U228) );
  AOI222_X1 U19761 ( .A1(n16759), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n16767), 
        .B2(BUF1_REG_18__SCAN_IN), .C1(n16760), .C2(P1_DATAO_REG_18__SCAN_IN), 
        .ZN(n16739) );
  INV_X1 U19762 ( .A(n16739), .ZN(U229) );
  AOI22_X1 U19763 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16759), .ZN(n16740) );
  OAI21_X1 U19764 ( .B1(n15376), .B2(n16764), .A(n16740), .ZN(U230) );
  AOI22_X1 U19765 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16759), .ZN(n16741) );
  OAI21_X1 U19766 ( .B1(n16742), .B2(n16764), .A(n16741), .ZN(U231) );
  AOI22_X1 U19767 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16759), .ZN(n16743) );
  OAI21_X1 U19768 ( .B1(n13975), .B2(n16764), .A(n16743), .ZN(U232) );
  AOI22_X1 U19769 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16759), .ZN(n16744) );
  OAI21_X1 U19770 ( .B1(n14504), .B2(n16764), .A(n16744), .ZN(U233) );
  AOI22_X1 U19771 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16759), .ZN(n16745) );
  OAI21_X1 U19772 ( .B1(n14530), .B2(n16764), .A(n16745), .ZN(U234) );
  AOI22_X1 U19773 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16759), .ZN(n16746) );
  OAI21_X1 U19774 ( .B1(n16747), .B2(n16764), .A(n16746), .ZN(U235) );
  AOI22_X1 U19775 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16759), .ZN(n16748) );
  OAI21_X1 U19776 ( .B1(n13715), .B2(n16764), .A(n16748), .ZN(U236) );
  AOI22_X1 U19777 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16759), .ZN(n16749) );
  OAI21_X1 U19778 ( .B1(n16750), .B2(n16764), .A(n16749), .ZN(U237) );
  AOI22_X1 U19779 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16759), .ZN(n16751) );
  OAI21_X1 U19780 ( .B1(n14448), .B2(n16764), .A(n16751), .ZN(U238) );
  AOI22_X1 U19781 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16759), .ZN(n16752) );
  OAI21_X1 U19782 ( .B1(n16753), .B2(n16764), .A(n16752), .ZN(U239) );
  INV_X1 U19783 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16755) );
  AOI22_X1 U19784 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16759), .ZN(n16754) );
  OAI21_X1 U19785 ( .B1(n16755), .B2(n16764), .A(n16754), .ZN(U240) );
  INV_X1 U19786 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16757) );
  AOI22_X1 U19787 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16759), .ZN(n16756) );
  OAI21_X1 U19788 ( .B1(n16757), .B2(n16764), .A(n16756), .ZN(U241) );
  INV_X1 U19789 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n21439) );
  AOI22_X1 U19790 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16767), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16759), .ZN(n16758) );
  OAI21_X1 U19791 ( .B1(n21439), .B2(U214), .A(n16758), .ZN(U242) );
  INV_X1 U19792 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16762) );
  AOI22_X1 U19793 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16759), .ZN(n16761) );
  OAI21_X1 U19794 ( .B1(n16762), .B2(n16764), .A(n16761), .ZN(U243) );
  INV_X1 U19795 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n21382) );
  AOI22_X1 U19796 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16760), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16759), .ZN(n16763) );
  OAI21_X1 U19797 ( .B1(n21382), .B2(n16764), .A(n16763), .ZN(U244) );
  INV_X1 U19798 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16771) );
  INV_X1 U19799 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16765) );
  INV_X1 U19800 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n21443) );
  OAI222_X1 U19801 ( .A1(U212), .A2(n16771), .B1(n16764), .B2(n16765), .C1(
        U214), .C2(n21443), .ZN(U245) );
  INV_X1 U19802 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16770) );
  AOI22_X1 U19803 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16767), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16760), .ZN(n16766) );
  OAI21_X1 U19804 ( .B1(n16770), .B2(U212), .A(n16766), .ZN(U246) );
  INV_X1 U19805 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16769) );
  AOI22_X1 U19806 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16767), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16760), .ZN(n16768) );
  OAI21_X1 U19807 ( .B1(n16769), .B2(U212), .A(n16768), .ZN(U247) );
  AOI22_X1 U19808 ( .A1(n16800), .A2(n16769), .B1(n18503), .B2(U215), .ZN(U251) );
  INV_X1 U19809 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18512) );
  AOI22_X1 U19810 ( .A1(n16800), .A2(n16770), .B1(n18512), .B2(U215), .ZN(U252) );
  INV_X1 U19811 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18517) );
  AOI22_X1 U19812 ( .A1(n16800), .A2(n16771), .B1(n18517), .B2(U215), .ZN(U253) );
  OAI22_X1 U19813 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16800), .ZN(n16772) );
  INV_X1 U19814 ( .A(n16772), .ZN(U254) );
  OAI22_X1 U19815 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16785), .ZN(n16773) );
  INV_X1 U19816 ( .A(n16773), .ZN(U255) );
  OAI22_X1 U19817 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16785), .ZN(n16774) );
  INV_X1 U19818 ( .A(n16774), .ZN(U256) );
  OAI22_X1 U19819 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16785), .ZN(n16775) );
  INV_X1 U19820 ( .A(n16775), .ZN(U257) );
  OAI22_X1 U19821 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16785), .ZN(n16776) );
  INV_X1 U19822 ( .A(n16776), .ZN(U258) );
  OAI22_X1 U19823 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16785), .ZN(n16777) );
  INV_X1 U19824 ( .A(n16777), .ZN(U259) );
  OAI22_X1 U19825 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16785), .ZN(n16778) );
  INV_X1 U19826 ( .A(n16778), .ZN(U260) );
  OAI22_X1 U19827 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16785), .ZN(n16779) );
  INV_X1 U19828 ( .A(n16779), .ZN(U261) );
  OAI22_X1 U19829 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16800), .ZN(n16780) );
  INV_X1 U19830 ( .A(n16780), .ZN(U262) );
  OAI22_X1 U19831 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16785), .ZN(n16781) );
  INV_X1 U19832 ( .A(n16781), .ZN(U263) );
  OAI22_X1 U19833 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16800), .ZN(n16782) );
  INV_X1 U19834 ( .A(n16782), .ZN(U264) );
  OAI22_X1 U19835 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16785), .ZN(n16783) );
  INV_X1 U19836 ( .A(n16783), .ZN(U265) );
  OAI22_X1 U19837 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16800), .ZN(n16784) );
  INV_X1 U19838 ( .A(n16784), .ZN(U266) );
  OAI22_X1 U19839 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16785), .ZN(n16786) );
  INV_X1 U19840 ( .A(n16786), .ZN(U267) );
  OAI22_X1 U19841 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16800), .ZN(n16787) );
  INV_X1 U19842 ( .A(n16787), .ZN(U268) );
  INV_X1 U19843 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n21398) );
  INV_X1 U19844 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18518) );
  AOI22_X1 U19845 ( .A1(n16800), .A2(n21398), .B1(n18518), .B2(U215), .ZN(U269) );
  OAI22_X1 U19846 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16800), .ZN(n16788) );
  INV_X1 U19847 ( .A(n16788), .ZN(U270) );
  OAI22_X1 U19848 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16800), .ZN(n16789) );
  INV_X1 U19849 ( .A(n16789), .ZN(U271) );
  OAI22_X1 U19850 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16800), .ZN(n16790) );
  INV_X1 U19851 ( .A(n16790), .ZN(U272) );
  OAI22_X1 U19852 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16800), .ZN(n16791) );
  INV_X1 U19853 ( .A(n16791), .ZN(U273) );
  OAI22_X1 U19854 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16800), .ZN(n16792) );
  INV_X1 U19855 ( .A(n16792), .ZN(U274) );
  OAI22_X1 U19856 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16800), .ZN(n16793) );
  INV_X1 U19857 ( .A(n16793), .ZN(U275) );
  OAI22_X1 U19858 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16800), .ZN(n16794) );
  INV_X1 U19859 ( .A(n16794), .ZN(U276) );
  OAI22_X1 U19860 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16800), .ZN(n16795) );
  INV_X1 U19861 ( .A(n16795), .ZN(U277) );
  OAI22_X1 U19862 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16800), .ZN(n16796) );
  INV_X1 U19863 ( .A(n16796), .ZN(U278) );
  OAI22_X1 U19864 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16800), .ZN(n16797) );
  INV_X1 U19865 ( .A(n16797), .ZN(U279) );
  OAI22_X1 U19866 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16800), .ZN(n16798) );
  INV_X1 U19867 ( .A(n16798), .ZN(U280) );
  INV_X1 U19868 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16801) );
  INV_X1 U19869 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n21395) );
  AOI22_X1 U19870 ( .A1(n16800), .A2(n16801), .B1(n21395), .B2(U215), .ZN(U281) );
  INV_X1 U19871 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18539) );
  AOI22_X1 U19872 ( .A1(n16800), .A2(n16799), .B1(n18539), .B2(U215), .ZN(U282) );
  INV_X1 U19873 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16802) );
  INV_X1 U19874 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n21505) );
  OAI222_X1 U19875 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n16802), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n16801), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n21505), .ZN(n16804) );
  INV_X2 U19876 ( .A(n16805), .ZN(n16803) );
  INV_X1 U19877 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19051) );
  INV_X1 U19878 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20149) );
  AOI22_X1 U19879 ( .A1(n16803), .A2(n19051), .B1(n20149), .B2(n16805), .ZN(
        U347) );
  INV_X1 U19880 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n21503) );
  INV_X1 U19881 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20147) );
  AOI22_X1 U19882 ( .A1(n16803), .A2(n21503), .B1(n20147), .B2(n16805), .ZN(
        U348) );
  INV_X1 U19883 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19047) );
  INV_X1 U19884 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20145) );
  AOI22_X1 U19885 ( .A1(n16803), .A2(n19047), .B1(n20145), .B2(n16805), .ZN(
        U349) );
  INV_X1 U19886 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19046) );
  INV_X1 U19887 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n21517) );
  AOI22_X1 U19888 ( .A1(n16803), .A2(n19046), .B1(n21517), .B2(n16805), .ZN(
        U350) );
  INV_X1 U19889 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19044) );
  INV_X1 U19890 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20142) );
  AOI22_X1 U19891 ( .A1(n16803), .A2(n19044), .B1(n20142), .B2(n16805), .ZN(
        U351) );
  INV_X1 U19892 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19042) );
  INV_X1 U19893 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20140) );
  AOI22_X1 U19894 ( .A1(n16803), .A2(n19042), .B1(n20140), .B2(n16805), .ZN(
        U352) );
  INV_X1 U19895 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19040) );
  INV_X1 U19896 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20138) );
  AOI22_X1 U19897 ( .A1(n16803), .A2(n19040), .B1(n20138), .B2(n16805), .ZN(
        U353) );
  INV_X1 U19898 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19038) );
  AOI22_X1 U19899 ( .A1(n16803), .A2(n19038), .B1(n20136), .B2(n16805), .ZN(
        U354) );
  INV_X1 U19900 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19089) );
  INV_X1 U19901 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20188) );
  AOI22_X1 U19902 ( .A1(n16803), .A2(n19089), .B1(n20188), .B2(n16804), .ZN(
        U355) );
  INV_X1 U19903 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19087) );
  INV_X1 U19904 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20184) );
  AOI22_X1 U19905 ( .A1(n16803), .A2(n19087), .B1(n20184), .B2(n16805), .ZN(
        U356) );
  INV_X1 U19906 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19085) );
  INV_X1 U19907 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20183) );
  AOI22_X1 U19908 ( .A1(n16803), .A2(n19085), .B1(n20183), .B2(n16805), .ZN(
        U357) );
  INV_X1 U19909 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19082) );
  INV_X1 U19910 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20180) );
  AOI22_X1 U19911 ( .A1(n16803), .A2(n19082), .B1(n20180), .B2(n16804), .ZN(
        U358) );
  INV_X1 U19912 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19080) );
  INV_X1 U19913 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20179) );
  AOI22_X1 U19914 ( .A1(n16803), .A2(n19080), .B1(n20179), .B2(n16804), .ZN(
        U359) );
  INV_X1 U19915 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19079) );
  INV_X1 U19916 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n21436) );
  AOI22_X1 U19917 ( .A1(n16803), .A2(n19079), .B1(n21436), .B2(n16804), .ZN(
        U360) );
  INV_X1 U19918 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19077) );
  INV_X1 U19919 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20176) );
  AOI22_X1 U19920 ( .A1(n16803), .A2(n19077), .B1(n20176), .B2(n16804), .ZN(
        U361) );
  INV_X1 U19921 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19074) );
  INV_X1 U19922 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20174) );
  AOI22_X1 U19923 ( .A1(n16803), .A2(n19074), .B1(n20174), .B2(n16804), .ZN(
        U362) );
  INV_X1 U19924 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19073) );
  INV_X1 U19925 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20172) );
  AOI22_X1 U19926 ( .A1(n16803), .A2(n19073), .B1(n20172), .B2(n16805), .ZN(
        U363) );
  INV_X1 U19927 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19070) );
  INV_X1 U19928 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20170) );
  AOI22_X1 U19929 ( .A1(n16803), .A2(n19070), .B1(n20170), .B2(n16805), .ZN(
        U364) );
  INV_X1 U19930 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19036) );
  INV_X1 U19931 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20134) );
  AOI22_X1 U19932 ( .A1(n16803), .A2(n19036), .B1(n20134), .B2(n16805), .ZN(
        U365) );
  INV_X1 U19933 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19069) );
  INV_X1 U19934 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20168) );
  AOI22_X1 U19935 ( .A1(n16803), .A2(n19069), .B1(n20168), .B2(n16805), .ZN(
        U366) );
  INV_X1 U19936 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19067) );
  INV_X1 U19937 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n21378) );
  AOI22_X1 U19938 ( .A1(n16803), .A2(n19067), .B1(n21378), .B2(n16805), .ZN(
        U367) );
  INV_X1 U19939 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19066) );
  INV_X1 U19940 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20165) );
  AOI22_X1 U19941 ( .A1(n16803), .A2(n19066), .B1(n20165), .B2(n16805), .ZN(
        U368) );
  INV_X1 U19942 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19063) );
  INV_X1 U19943 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20163) );
  AOI22_X1 U19944 ( .A1(n16803), .A2(n19063), .B1(n20163), .B2(n16805), .ZN(
        U369) );
  INV_X1 U19945 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n21485) );
  INV_X1 U19946 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20161) );
  AOI22_X1 U19947 ( .A1(n16803), .A2(n21485), .B1(n20161), .B2(n16805), .ZN(
        U370) );
  INV_X1 U19948 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19061) );
  INV_X1 U19949 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20159) );
  AOI22_X1 U19950 ( .A1(n16803), .A2(n19061), .B1(n20159), .B2(n16805), .ZN(
        U371) );
  INV_X1 U19951 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19058) );
  INV_X1 U19952 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20157) );
  AOI22_X1 U19953 ( .A1(n16803), .A2(n19058), .B1(n20157), .B2(n16805), .ZN(
        U372) );
  INV_X1 U19954 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19057) );
  INV_X1 U19955 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20155) );
  AOI22_X1 U19956 ( .A1(n16803), .A2(n19057), .B1(n20155), .B2(n16805), .ZN(
        U373) );
  INV_X1 U19957 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19055) );
  INV_X1 U19958 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20153) );
  AOI22_X1 U19959 ( .A1(n16803), .A2(n19055), .B1(n20153), .B2(n16804), .ZN(
        U374) );
  INV_X1 U19960 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19053) );
  INV_X1 U19961 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20151) );
  AOI22_X1 U19962 ( .A1(n16803), .A2(n19053), .B1(n20151), .B2(n16804), .ZN(
        U375) );
  INV_X1 U19963 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19035) );
  INV_X1 U19964 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20131) );
  AOI22_X1 U19965 ( .A1(n16803), .A2(n19035), .B1(n20131), .B2(n16805), .ZN(
        U376) );
  NOR2_X1 U19966 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21390), .ZN(n19022) );
  NOR2_X1 U19967 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_0__SCAN_IN), 
        .ZN(n19018) );
  AOI21_X1 U19968 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n19022), .A(n19018), 
        .ZN(n19016) );
  INV_X1 U19969 ( .A(n19016), .ZN(n19097) );
  AOI21_X1 U19970 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19097), .ZN(n16806) );
  INV_X1 U19971 ( .A(n16806), .ZN(P3_U2633) );
  NAND2_X1 U19972 ( .A1(n19005), .A2(n19102), .ZN(n16808) );
  INV_X1 U19973 ( .A(n19008), .ZN(n16831) );
  OAI21_X1 U19974 ( .B1(n16813), .B2(n17720), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16807) );
  OAI21_X1 U19975 ( .B1(n16808), .B2(n16831), .A(n16807), .ZN(P3_U2634) );
  INV_X2 U19976 ( .A(n19161), .ZN(n19140) );
  AOI21_X1 U19977 ( .B1(n19034), .B2(n21390), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16809) );
  AOI22_X1 U19978 ( .A1(n19140), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16809), 
        .B2(n19161), .ZN(P3_U2635) );
  OAI21_X1 U19979 ( .B1(n19017), .B2(BS16), .A(n19097), .ZN(n19096) );
  OAI21_X1 U19980 ( .B1(n19097), .B2(n19151), .A(n19096), .ZN(P3_U2636) );
  INV_X1 U19981 ( .A(n16810), .ZN(n16812) );
  NOR3_X1 U19982 ( .A1(n16813), .A2(n16812), .A3(n16811), .ZN(n18991) );
  NOR2_X1 U19983 ( .A1(n18991), .A2(n19149), .ZN(n19141) );
  OAI21_X1 U19984 ( .B1(n19141), .B2(n16815), .A(n16814), .ZN(P3_U2637) );
  NOR4_X1 U19985 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16819) );
  NOR4_X1 U19986 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16818) );
  NOR4_X1 U19987 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16817) );
  NOR4_X1 U19988 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16816) );
  NAND4_X1 U19989 ( .A1(n16819), .A2(n16818), .A3(n16817), .A4(n16816), .ZN(
        n16825) );
  NOR4_X1 U19990 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16823) );
  AOI211_X1 U19991 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_12__SCAN_IN), .B(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16822) );
  NOR4_X1 U19992 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16821) );
  NOR4_X1 U19993 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16820) );
  NAND4_X1 U19994 ( .A1(n16823), .A2(n16822), .A3(n16821), .A4(n16820), .ZN(
        n16824) );
  NOR2_X1 U19995 ( .A1(n16825), .A2(n16824), .ZN(n19134) );
  INV_X1 U19996 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16827) );
  NOR3_X1 U19997 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16828) );
  OAI21_X1 U19998 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16828), .A(n19134), .ZN(
        n16826) );
  OAI21_X1 U19999 ( .B1(n19134), .B2(n16827), .A(n16826), .ZN(P3_U2638) );
  INV_X1 U20000 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19130) );
  INV_X1 U20001 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19098) );
  AOI21_X1 U20002 ( .B1(n19130), .B2(n19098), .A(n16828), .ZN(n16830) );
  INV_X1 U20003 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16829) );
  INV_X1 U20004 ( .A(n19134), .ZN(n19137) );
  AOI22_X1 U20005 ( .A1(n19134), .A2(n16830), .B1(n16829), .B2(n19137), .ZN(
        P3_U2639) );
  NAND4_X1 U20006 ( .A1(n19005), .A2(n19099), .A3(n19151), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n19011) );
  NOR2_X1 U20007 ( .A1(n19102), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18844) );
  INV_X1 U20008 ( .A(n18844), .ZN(n19006) );
  NOR2_X1 U20009 ( .A1(n16831), .A2(n19006), .ZN(n19000) );
  NOR3_X1 U20010 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17174) );
  INV_X1 U20011 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n21367) );
  NAND2_X1 U20012 ( .A1(n17174), .A2(n21367), .ZN(n17164) );
  NOR2_X1 U20013 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17164), .ZN(n17140) );
  NAND2_X1 U20014 ( .A1(n17140), .A2(n17499), .ZN(n17136) );
  INV_X1 U20015 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17467) );
  NAND2_X1 U20016 ( .A1(n17116), .A2(n17467), .ZN(n17110) );
  NAND2_X1 U20017 ( .A1(n17093), .A2(n17085), .ZN(n17084) );
  NAND2_X1 U20018 ( .A1(n17069), .A2(n17429), .ZN(n17059) );
  NAND2_X1 U20019 ( .A1(n17044), .A2(n17396), .ZN(n17036) );
  INV_X1 U20020 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17013) );
  NAND2_X1 U20021 ( .A1(n17019), .A2(n17013), .ZN(n17011) );
  INV_X1 U20022 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17338) );
  NAND2_X1 U20023 ( .A1(n16998), .A2(n17338), .ZN(n16988) );
  INV_X1 U20024 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17324) );
  NAND2_X1 U20025 ( .A1(n16982), .A2(n17324), .ZN(n16970) );
  NAND2_X1 U20026 ( .A1(n16957), .A2(n17296), .ZN(n16953) );
  NAND2_X1 U20027 ( .A1(n16941), .A2(n17258), .ZN(n16931) );
  INV_X1 U20028 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17249) );
  NAND2_X1 U20029 ( .A1(n16921), .A2(n17249), .ZN(n16915) );
  NOR2_X1 U20030 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16915), .ZN(n16901) );
  NAND2_X1 U20031 ( .A1(n16901), .A2(n17242), .ZN(n16893) );
  NOR2_X1 U20032 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16893), .ZN(n16880) );
  INV_X1 U20033 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17237) );
  NAND2_X1 U20034 ( .A1(n16880), .A2(n17237), .ZN(n16874) );
  INV_X1 U20035 ( .A(n16874), .ZN(n16863) );
  NAND2_X1 U20036 ( .A1(n17683), .A2(n19168), .ZN(n19166) );
  NAND2_X1 U20037 ( .A1(n19151), .A2(n19153), .ZN(n16832) );
  NOR2_X1 U20038 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17194), .ZN(n16858) );
  INV_X1 U20039 ( .A(n19153), .ZN(n19146) );
  AOI211_X1 U20040 ( .C1(n19152), .C2(n19150), .A(n19146), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18995) );
  AOI211_X4 U20041 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18511), .A(n18995), .B(
        n19166), .ZN(n17154) );
  AOI22_X1 U20042 ( .A1(n16863), .A2(n16858), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17154), .ZN(n16856) );
  INV_X1 U20043 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19086) );
  NAND2_X1 U20044 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16886) );
  NOR2_X1 U20045 ( .A1(n19086), .A2(n16886), .ZN(n16839) );
  INV_X1 U20046 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19075) );
  INV_X1 U20047 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19068) );
  NAND3_X1 U20048 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16972) );
  NAND2_X1 U20049 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16960) );
  NOR3_X1 U20050 ( .A1(n19068), .A2(n16972), .A3(n16960), .ZN(n16834) );
  INV_X1 U20051 ( .A(n16834), .ZN(n16938) );
  INV_X1 U20052 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19054) );
  INV_X1 U20053 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19048) );
  INV_X1 U20054 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19041) );
  INV_X1 U20055 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19037) );
  NAND2_X1 U20056 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n17172) );
  NOR2_X1 U20057 ( .A1(n19037), .A2(n17172), .ZN(n17152) );
  NAND2_X1 U20058 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17152), .ZN(n17129) );
  NOR2_X1 U20059 ( .A1(n19041), .A2(n17129), .ZN(n17120) );
  NAND3_X1 U20060 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(n17120), .ZN(n17096) );
  NOR2_X1 U20061 ( .A1(n19048), .A2(n17096), .ZN(n17062) );
  NAND4_X1 U20062 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17062), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n17046) );
  NOR2_X1 U20063 ( .A1(n19054), .A2(n17046), .ZN(n17037) );
  NAND2_X1 U20064 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17037), .ZN(n16835) );
  NAND3_X1 U20065 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(n16952), .ZN(n16937) );
  NAND3_X1 U20066 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n16914), .ZN(n16898) );
  INV_X1 U20067 ( .A(n16898), .ZN(n16887) );
  AND2_X1 U20068 ( .A1(n16839), .A2(n16887), .ZN(n16854) );
  NOR2_X1 U20069 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n21437), .ZN(n16853) );
  NAND2_X1 U20070 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16838) );
  NAND4_X1 U20071 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n16834), .A4(P3_REIP_REG_22__SCAN_IN), .ZN(n16836) );
  INV_X1 U20072 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19059) );
  NOR3_X1 U20073 ( .A1(n17183), .A2(n19059), .A3(n16835), .ZN(n17021) );
  AOI21_X1 U20074 ( .B1(n16973), .B2(n16836), .A(n17024), .ZN(n16936) );
  INV_X1 U20075 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19076) );
  NAND2_X1 U20076 ( .A1(n16837), .A2(n19076), .ZN(n16927) );
  NAND2_X1 U20077 ( .A1(n16936), .A2(n16927), .ZN(n16913) );
  AOI21_X1 U20078 ( .B1(n16973), .B2(n16838), .A(n16913), .ZN(n16907) );
  OAI21_X1 U20079 ( .B1(n16839), .B2(n17187), .A(n16907), .ZN(n16862) );
  INV_X1 U20080 ( .A(n16862), .ZN(n16877) );
  NAND2_X1 U20081 ( .A1(n16854), .A2(n21437), .ZN(n16864) );
  AOI21_X1 U20082 ( .B1(n16877), .B2(n16864), .A(n19088), .ZN(n16852) );
  NAND2_X1 U20083 ( .A1(n16843), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16841) );
  AOI21_X1 U20084 ( .B1(n16882), .B2(n16841), .A(n16840), .ZN(n17790) );
  OAI21_X1 U20085 ( .B1(n16843), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16841), .ZN(n17809) );
  INV_X1 U20086 ( .A(n17809), .ZN(n16892) );
  INV_X1 U20087 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16902) );
  NAND2_X1 U20088 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17877) );
  NAND2_X1 U20089 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17874), .ZN(
        n16848) );
  NOR2_X1 U20090 ( .A1(n17877), .A2(n16848), .ZN(n17831) );
  NAND2_X1 U20091 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17834) );
  NOR2_X1 U20092 ( .A1(n16842), .A2(n17834), .ZN(n17820) );
  NAND2_X1 U20093 ( .A1(n17831), .A2(n17820), .ZN(n17789) );
  AOI21_X1 U20094 ( .B1(n16902), .B2(n17789), .A(n16843), .ZN(n17821) );
  INV_X1 U20095 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16923) );
  NAND2_X1 U20096 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17832), .ZN(
        n16845) );
  NOR2_X1 U20097 ( .A1(n16923), .A2(n16845), .ZN(n16844) );
  OAI21_X1 U20098 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16844), .A(
        n17789), .ZN(n17836) );
  INV_X1 U20099 ( .A(n17836), .ZN(n16911) );
  AOI21_X1 U20100 ( .B1(n16923), .B2(n16845), .A(n16844), .ZN(n17845) );
  OAI21_X1 U20101 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17831), .A(
        n16845), .ZN(n16846) );
  INV_X1 U20102 ( .A(n16846), .ZN(n17863) );
  INV_X1 U20103 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17875) );
  INV_X1 U20104 ( .A(n16848), .ZN(n16849) );
  NAND2_X1 U20105 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16849), .ZN(
        n16847) );
  AOI21_X1 U20106 ( .B1(n17875), .B2(n16847), .A(n17831), .ZN(n17873) );
  INV_X1 U20107 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17876) );
  OAI22_X1 U20108 ( .A1(n17876), .A2(n16849), .B1(n16848), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17889) );
  NOR2_X1 U20109 ( .A1(n21330), .A2(n17901), .ZN(n17871) );
  INV_X1 U20110 ( .A(n17871), .ZN(n16850) );
  AOI21_X1 U20111 ( .B1(n17900), .B2(n16850), .A(n16849), .ZN(n17903) );
  INV_X1 U20112 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17117) );
  NAND2_X1 U20113 ( .A1(n17117), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17168) );
  OAI21_X1 U20114 ( .B1(n17901), .B2(n17168), .A(n17157), .ZN(n16851) );
  INV_X1 U20115 ( .A(n16851), .ZN(n16962) );
  NOR2_X1 U20116 ( .A1(n17903), .A2(n16962), .ZN(n16961) );
  NOR2_X1 U20117 ( .A1(n16939), .A2(n17065), .ZN(n16930) );
  NOR2_X1 U20118 ( .A1(n17863), .A2(n16930), .ZN(n16929) );
  NOR2_X1 U20119 ( .A1(n16929), .A2(n17065), .ZN(n16920) );
  NOR2_X1 U20120 ( .A1(n17845), .A2(n16920), .ZN(n16919) );
  NOR2_X1 U20121 ( .A1(n16919), .A2(n17065), .ZN(n16910) );
  NOR2_X1 U20122 ( .A1(n16911), .A2(n16910), .ZN(n16909) );
  NOR2_X1 U20123 ( .A1(n16909), .A2(n17065), .ZN(n16900) );
  NOR2_X1 U20124 ( .A1(n17821), .A2(n16900), .ZN(n16899) );
  NOR2_X1 U20125 ( .A1(n16899), .A2(n17065), .ZN(n16891) );
  NOR2_X1 U20126 ( .A1(n16892), .A2(n16891), .ZN(n16890) );
  NOR2_X1 U20127 ( .A1(n16890), .A2(n17065), .ZN(n16879) );
  NOR2_X1 U20128 ( .A1(n17790), .A2(n16879), .ZN(n16878) );
  NOR2_X1 U20129 ( .A1(n16878), .A2(n17065), .ZN(n16869) );
  INV_X1 U20130 ( .A(n17147), .ZN(n17186) );
  OAI211_X1 U20131 ( .C1(n16857), .C2(n17184), .A(n16856), .B(n16855), .ZN(
        P3_U2640) );
  AOI22_X1 U20132 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n17115), .B1(
        n16858), .B2(n16874), .ZN(n16867) );
  XOR2_X1 U20133 ( .A(n16860), .B(n16859), .Z(n16861) );
  AOI22_X1 U20134 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16862), .B1(n17147), 
        .B2(n16861), .ZN(n16866) );
  OAI221_X1 U20135 ( .B1(n17154), .B2(n16863), .C1(n17154), .C2(n17176), .A(
        P3_EBX_REG_30__SCAN_IN), .ZN(n16865) );
  NAND4_X1 U20136 ( .A1(n16867), .A2(n16866), .A3(n16865), .A4(n16864), .ZN(
        P3_U2641) );
  AOI211_X1 U20137 ( .C1(n16870), .C2(n16869), .A(n16868), .B(n17186), .ZN(
        n16873) );
  NOR3_X1 U20138 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16886), .A3(n16898), 
        .ZN(n16872) );
  OAI22_X1 U20139 ( .A1(n10167), .A2(n17184), .B1(n17237), .B2(n17193), .ZN(
        n16871) );
  NOR3_X1 U20140 ( .A1(n16873), .A2(n16872), .A3(n16871), .ZN(n16876) );
  OAI211_X1 U20141 ( .C1(n16880), .C2(n17237), .A(n17176), .B(n16874), .ZN(
        n16875) );
  OAI211_X1 U20142 ( .C1(n16877), .C2(n19086), .A(n16876), .B(n16875), .ZN(
        P3_U2642) );
  INV_X1 U20143 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19084) );
  AOI211_X1 U20144 ( .C1(n17790), .C2(n16879), .A(n16878), .B(n17186), .ZN(
        n16885) );
  AOI211_X1 U20145 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16893), .A(n16880), .B(
        n17194), .ZN(n16884) );
  OAI22_X1 U20146 ( .A1(n16882), .A2(n17184), .B1(n16881), .B2(n17193), .ZN(
        n16883) );
  NOR3_X1 U20147 ( .A1(n16885), .A2(n16884), .A3(n16883), .ZN(n16889) );
  OAI211_X1 U20148 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16887), .B(n16886), .ZN(n16888) );
  OAI211_X1 U20149 ( .C1(n16907), .C2(n19084), .A(n16889), .B(n16888), .ZN(
        P3_U2643) );
  INV_X1 U20150 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19081) );
  AOI211_X1 U20151 ( .C1(n16892), .C2(n16891), .A(n16890), .B(n17186), .ZN(
        n16896) );
  OAI211_X1 U20152 ( .C1(n16901), .C2(n17242), .A(n17176), .B(n16893), .ZN(
        n16894) );
  OAI21_X1 U20153 ( .B1(n17193), .B2(n17242), .A(n16894), .ZN(n16895) );
  AOI211_X1 U20154 ( .C1(n17115), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16896), .B(n16895), .ZN(n16897) );
  OAI221_X1 U20155 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16898), .C1(n19081), 
        .C2(n16907), .A(n16897), .ZN(P3_U2644) );
  NAND2_X1 U20156 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16914), .ZN(n16908) );
  INV_X1 U20157 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21427) );
  AOI211_X1 U20158 ( .C1(n17821), .C2(n16900), .A(n16899), .B(n17186), .ZN(
        n16905) );
  AOI211_X1 U20159 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16915), .A(n16901), .B(
        n17194), .ZN(n16904) );
  INV_X1 U20160 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17253) );
  OAI22_X1 U20161 ( .A1(n16902), .A2(n17184), .B1(n17253), .B2(n17193), .ZN(
        n16903) );
  NOR3_X1 U20162 ( .A1(n16905), .A2(n16904), .A3(n16903), .ZN(n16906) );
  OAI221_X1 U20163 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n16908), .C1(n21427), 
        .C2(n16907), .A(n16906), .ZN(P3_U2645) );
  AOI22_X1 U20164 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17115), .B1(
        P3_EBX_REG_25__SCAN_IN), .B2(n17154), .ZN(n16918) );
  INV_X1 U20165 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19078) );
  AOI211_X1 U20166 ( .C1(n16911), .C2(n16910), .A(n16909), .B(n17186), .ZN(
        n16912) );
  AOI221_X1 U20167 ( .B1(n16914), .B2(n19078), .C1(n16913), .C2(
        P3_REIP_REG_25__SCAN_IN), .A(n16912), .ZN(n16917) );
  OAI211_X1 U20168 ( .C1(n16921), .C2(n17249), .A(n17176), .B(n16915), .ZN(
        n16916) );
  NAND3_X1 U20169 ( .A1(n16918), .A2(n16917), .A3(n16916), .ZN(P3_U2646) );
  AOI211_X1 U20170 ( .C1(n17845), .C2(n16920), .A(n16919), .B(n17186), .ZN(
        n16926) );
  AOI211_X1 U20171 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16931), .A(n16921), .B(
        n17194), .ZN(n16925) );
  OAI22_X1 U20172 ( .A1(n16923), .A2(n17184), .B1(n16922), .B2(n17193), .ZN(
        n16924) );
  NOR3_X1 U20173 ( .A1(n16926), .A2(n16925), .A3(n16924), .ZN(n16928) );
  OAI211_X1 U20174 ( .C1(n16936), .C2(n19076), .A(n16928), .B(n16927), .ZN(
        P3_U2647) );
  AOI211_X1 U20175 ( .C1(n17863), .C2(n16930), .A(n16929), .B(n17186), .ZN(
        n16934) );
  OAI211_X1 U20176 ( .C1(n16941), .C2(n17258), .A(n17176), .B(n16931), .ZN(
        n16932) );
  OAI21_X1 U20177 ( .B1(n17193), .B2(n17258), .A(n16932), .ZN(n16933) );
  AOI211_X1 U20178 ( .C1(n17115), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16934), .B(n16933), .ZN(n16935) );
  OAI221_X1 U20179 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n16937), .C1(n19075), 
        .C2(n16936), .A(n16935), .ZN(P3_U2648) );
  AOI21_X1 U20180 ( .B1(n16973), .B2(n16938), .A(n17024), .ZN(n16948) );
  INV_X1 U20181 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19072) );
  AOI211_X1 U20182 ( .C1(n17873), .C2(n16940), .A(n16939), .B(n17186), .ZN(
        n16944) );
  AOI211_X1 U20183 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16953), .A(n16941), .B(
        n17194), .ZN(n16943) );
  OAI22_X1 U20184 ( .A1(n17875), .A2(n17184), .B1(n17271), .B2(n17193), .ZN(
        n16942) );
  NOR3_X1 U20185 ( .A1(n16944), .A2(n16943), .A3(n16942), .ZN(n16947) );
  NAND2_X1 U20186 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n16945) );
  OAI211_X1 U20187 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(P3_REIP_REG_22__SCAN_IN), .A(n16952), .B(n16945), .ZN(n16946) );
  OAI211_X1 U20188 ( .C1(n16948), .C2(n19072), .A(n16947), .B(n16946), .ZN(
        P3_U2649) );
  AOI22_X1 U20189 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17115), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n17154), .ZN(n16956) );
  INV_X1 U20190 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19071) );
  INV_X1 U20191 ( .A(n16948), .ZN(n16964) );
  AOI211_X1 U20192 ( .C1(n17889), .C2(n16950), .A(n16949), .B(n17186), .ZN(
        n16951) );
  AOI221_X1 U20193 ( .B1(n16952), .B2(n19071), .C1(n16964), .C2(
        P3_REIP_REG_21__SCAN_IN), .A(n16951), .ZN(n16955) );
  OAI211_X1 U20194 ( .C1(n16957), .C2(n17296), .A(n17176), .B(n16953), .ZN(
        n16954) );
  NAND3_X1 U20195 ( .A1(n16956), .A2(n16955), .A3(n16954), .ZN(P3_U2650) );
  AOI211_X1 U20196 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16970), .A(n16957), .B(
        n17194), .ZN(n16958) );
  AOI21_X1 U20197 ( .B1(n17154), .B2(P3_EBX_REG_20__SCAN_IN), .A(n16958), .ZN(
        n16967) );
  INV_X1 U20198 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19062) );
  INV_X1 U20199 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19060) );
  NOR2_X1 U20200 ( .A1(n19062), .A2(n19060), .ZN(n17003) );
  INV_X1 U20201 ( .A(n17003), .ZN(n16959) );
  NOR2_X1 U20202 ( .A1(n16959), .A2(n17018), .ZN(n16993) );
  NAND2_X1 U20203 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16993), .ZN(n16987) );
  NOR2_X1 U20204 ( .A1(n16960), .A2(n16987), .ZN(n16965) );
  AOI211_X1 U20205 ( .C1(n17903), .C2(n16962), .A(n16961), .B(n17186), .ZN(
        n16963) );
  AOI221_X1 U20206 ( .B1(n16965), .B2(n19068), .C1(n16964), .C2(
        P3_REIP_REG_20__SCAN_IN), .A(n16963), .ZN(n16966) );
  OAI211_X1 U20207 ( .C1(n17900), .C2(n17184), .A(n16967), .B(n16966), .ZN(
        P3_U2651) );
  INV_X1 U20208 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17957) );
  NAND2_X1 U20209 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17990) );
  NOR2_X1 U20210 ( .A1(n21330), .A2(n18017), .ZN(n17053) );
  INV_X1 U20211 ( .A(n17053), .ZN(n17102) );
  NOR2_X1 U20212 ( .A1(n16968), .A2(n17102), .ZN(n17054) );
  INV_X1 U20213 ( .A(n17054), .ZN(n17987) );
  NOR2_X1 U20214 ( .A1(n17990), .A2(n17987), .ZN(n17029) );
  NAND2_X1 U20215 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17029), .ZN(
        n17942) );
  NOR2_X1 U20216 ( .A1(n17957), .A2(n17942), .ZN(n17008) );
  NAND2_X1 U20217 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17008), .ZN(
        n17000) );
  NOR2_X1 U20218 ( .A1(n21440), .A2(n17000), .ZN(n17909) );
  NAND2_X1 U20219 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17909), .ZN(
        n16979) );
  AOI21_X1 U20220 ( .B1(n17008), .B2(n17117), .A(n17065), .ZN(n17001) );
  AOI21_X1 U20221 ( .B1(n17157), .B2(n16979), .A(n17001), .ZN(n16969) );
  AOI21_X1 U20222 ( .B1(n10182), .B2(n16979), .A(n17871), .ZN(n17910) );
  XOR2_X1 U20223 ( .A(n16969), .B(n17910), .Z(n16978) );
  OAI211_X1 U20224 ( .C1(n16982), .C2(n17324), .A(n17176), .B(n16970), .ZN(
        n16971) );
  OAI211_X1 U20225 ( .C1(n17324), .C2(n17193), .A(n18484), .B(n16971), .ZN(
        n16976) );
  INV_X1 U20226 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19065) );
  XOR2_X1 U20227 ( .A(P3_REIP_REG_19__SCAN_IN), .B(n19065), .Z(n16974) );
  INV_X1 U20228 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n21473) );
  AOI21_X1 U20229 ( .B1(n16973), .B2(n16972), .A(n17024), .ZN(n16997) );
  OAI22_X1 U20230 ( .A1(n16987), .A2(n16974), .B1(n21473), .B2(n16997), .ZN(
        n16975) );
  AOI211_X1 U20231 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17115), .A(
        n16976), .B(n16975), .ZN(n16977) );
  OAI21_X1 U20232 ( .B1(n16978), .B2(n17186), .A(n16977), .ZN(P3_U2652) );
  OAI21_X1 U20233 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17909), .A(
        n16979), .ZN(n17919) );
  NAND3_X1 U20234 ( .A1(n17008), .A2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17117), .ZN(n16991) );
  OAI21_X1 U20235 ( .B1(n21440), .B2(n16991), .A(n17157), .ZN(n16981) );
  OAI21_X1 U20236 ( .B1(n17919), .B2(n16981), .A(n17147), .ZN(n16980) );
  AOI21_X1 U20237 ( .B1(n17919), .B2(n16981), .A(n16980), .ZN(n16985) );
  AOI211_X1 U20238 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16988), .A(n16982), .B(
        n17194), .ZN(n16984) );
  INV_X1 U20239 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17339) );
  OAI22_X1 U20240 ( .A1(n10181), .A2(n17184), .B1(n17339), .B2(n17193), .ZN(
        n16983) );
  NOR4_X1 U20241 ( .A1(n18479), .A2(n16985), .A3(n16984), .A4(n16983), .ZN(
        n16986) );
  OAI221_X1 U20242 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16987), .C1(n19065), 
        .C2(n16997), .A(n16986), .ZN(P3_U2653) );
  INV_X1 U20243 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19064) );
  OAI211_X1 U20244 ( .C1(n16998), .C2(n17338), .A(n17176), .B(n16988), .ZN(
        n16989) );
  OAI211_X1 U20245 ( .C1(n17338), .C2(n17193), .A(n18484), .B(n16989), .ZN(
        n16990) );
  AOI21_X1 U20246 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17115), .A(
        n16990), .ZN(n16996) );
  AOI21_X1 U20247 ( .B1(n21440), .B2(n17000), .A(n17909), .ZN(n17937) );
  NAND2_X1 U20248 ( .A1(n17157), .A2(n16991), .ZN(n16992) );
  XNOR2_X1 U20249 ( .A(n17937), .B(n16992), .ZN(n16994) );
  AOI22_X1 U20250 ( .A1(n17147), .A2(n16994), .B1(n16993), .B2(n19064), .ZN(
        n16995) );
  OAI211_X1 U20251 ( .C1(n16997), .C2(n19064), .A(n16996), .B(n16995), .ZN(
        P3_U2654) );
  INV_X1 U20252 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17945) );
  AOI211_X1 U20253 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17011), .A(n16998), .B(
        n17194), .ZN(n16999) );
  AOI211_X1 U20254 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17154), .A(n18479), .B(
        n16999), .ZN(n17007) );
  OAI21_X1 U20255 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17008), .A(
        n17000), .ZN(n17943) );
  INV_X1 U20256 ( .A(n17943), .ZN(n17002) );
  INV_X1 U20257 ( .A(n17001), .ZN(n17010) );
  AOI221_X1 U20258 ( .B1(n17002), .B2(n17001), .C1(n17943), .C2(n17010), .A(
        n17186), .ZN(n17005) );
  AOI211_X1 U20259 ( .C1(n19062), .C2(n19060), .A(n17003), .B(n17018), .ZN(
        n17004) );
  AOI211_X1 U20260 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n17024), .A(n17005), 
        .B(n17004), .ZN(n17006) );
  OAI211_X1 U20261 ( .C1(n17945), .C2(n17184), .A(n17007), .B(n17006), .ZN(
        P3_U2655) );
  AOI21_X1 U20262 ( .B1(n17957), .B2(n17942), .A(n17008), .ZN(n17960) );
  NAND2_X1 U20263 ( .A1(n17157), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17185) );
  NAND2_X1 U20264 ( .A1(n17147), .A2(n17185), .ZN(n17113) );
  AOI21_X1 U20265 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17157), .A(
        n17113), .ZN(n17009) );
  AOI22_X1 U20266 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17115), .B1(
        n17960), .B2(n17009), .ZN(n17017) );
  NOR3_X1 U20267 ( .A1(n17960), .A2(n17186), .A3(n17010), .ZN(n17015) );
  OAI211_X1 U20268 ( .C1(n17019), .C2(n17013), .A(n17176), .B(n17011), .ZN(
        n17012) );
  OAI211_X1 U20269 ( .C1(n17013), .C2(n17193), .A(n18484), .B(n17012), .ZN(
        n17014) );
  AOI211_X1 U20270 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n17024), .A(n17015), 
        .B(n17014), .ZN(n17016) );
  OAI211_X1 U20271 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n17018), .A(n17017), 
        .B(n17016), .ZN(P3_U2656) );
  AOI211_X1 U20272 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17036), .A(n17019), .B(
        n17194), .ZN(n17020) );
  AOI21_X1 U20273 ( .B1(n17115), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17020), .ZN(n17028) );
  INV_X1 U20274 ( .A(n17021), .ZN(n17022) );
  AOI22_X1 U20275 ( .A1(n17154), .A2(P3_EBX_REG_14__SCAN_IN), .B1(n17023), 
        .B2(n17022), .ZN(n17027) );
  OAI21_X1 U20276 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17029), .A(
        n17942), .ZN(n17975) );
  OAI21_X1 U20277 ( .B1(n17974), .B2(n17168), .A(n17157), .ZN(n17031) );
  XOR2_X1 U20278 ( .A(n17975), .B(n17031), .Z(n17025) );
  AOI22_X1 U20279 ( .A1(n17147), .A2(n17025), .B1(P3_REIP_REG_14__SCAN_IN), 
        .B2(n17024), .ZN(n17026) );
  NAND4_X1 U20280 ( .A1(n17028), .A2(n17027), .A3(n17026), .A4(n18484), .ZN(
        P3_U2657) );
  AOI22_X1 U20281 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17115), .B1(
        P3_EBX_REG_13__SCAN_IN), .B2(n17154), .ZN(n17041) );
  AOI21_X1 U20282 ( .B1(n17173), .B2(n17046), .A(n17183), .ZN(n17057) );
  NAND2_X1 U20283 ( .A1(n17173), .A2(n19054), .ZN(n17045) );
  INV_X1 U20284 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19056) );
  AOI21_X1 U20285 ( .B1(n17057), .B2(n17045), .A(n19056), .ZN(n17035) );
  INV_X1 U20286 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17992) );
  INV_X1 U20287 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18001) );
  NOR2_X1 U20288 ( .A1(n18001), .A2(n17987), .ZN(n17042) );
  INV_X1 U20289 ( .A(n17042), .ZN(n17030) );
  AOI21_X1 U20290 ( .B1(n17992), .B2(n17030), .A(n17029), .ZN(n17994) );
  NOR3_X1 U20291 ( .A1(n17994), .A2(n17186), .A3(n17031), .ZN(n17034) );
  INV_X1 U20292 ( .A(n17113), .ZN(n17190) );
  OAI211_X1 U20293 ( .C1(n17065), .C2(n17042), .A(n17994), .B(n17190), .ZN(
        n17032) );
  INV_X1 U20294 ( .A(n17032), .ZN(n17033) );
  NOR4_X1 U20295 ( .A1(n18479), .A2(n17035), .A3(n17034), .A4(n17033), .ZN(
        n17040) );
  OAI211_X1 U20296 ( .C1(n17044), .C2(n17396), .A(n17176), .B(n17036), .ZN(
        n17039) );
  NAND3_X1 U20297 ( .A1(n17173), .A2(n17037), .A3(n19056), .ZN(n17038) );
  NAND4_X1 U20298 ( .A1(n17041), .A2(n17040), .A3(n17039), .A4(n17038), .ZN(
        P3_U2658) );
  AOI22_X1 U20299 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17115), .B1(
        P3_EBX_REG_12__SCAN_IN), .B2(n17154), .ZN(n17051) );
  AOI21_X1 U20300 ( .B1(n18001), .B2(n17987), .A(n17042), .ZN(n18005) );
  NOR3_X1 U20301 ( .A1(n21330), .A2(n18097), .A3(n18098), .ZN(n17118) );
  AOI21_X1 U20302 ( .B1(n17118), .B2(n17117), .A(n17065), .ZN(n17104) );
  INV_X1 U20303 ( .A(n17104), .ZN(n17103) );
  OAI21_X1 U20304 ( .B1(n17065), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n17103), .ZN(n17091) );
  INV_X1 U20305 ( .A(n17091), .ZN(n17090) );
  OAI21_X1 U20306 ( .B1(n18019), .B2(n17065), .A(n17090), .ZN(n17043) );
  XOR2_X1 U20307 ( .A(n18005), .B(n17043), .Z(n17049) );
  AOI211_X1 U20308 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17059), .A(n17044), .B(
        n17194), .ZN(n17048) );
  OAI21_X1 U20309 ( .B1(n17046), .B2(n17045), .A(n18484), .ZN(n17047) );
  AOI211_X1 U20310 ( .C1(n17049), .C2(n17147), .A(n17048), .B(n17047), .ZN(
        n17050) );
  OAI211_X1 U20311 ( .C1(n17057), .C2(n19054), .A(n17051), .B(n17050), .ZN(
        P3_U2659) );
  INV_X1 U20312 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19050) );
  INV_X1 U20313 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19049) );
  NOR2_X1 U20314 ( .A1(n19050), .A2(n19049), .ZN(n17052) );
  NOR3_X1 U20315 ( .A1(n17187), .A2(n19048), .A3(n17096), .ZN(n17083) );
  AOI21_X1 U20316 ( .B1(n17052), .B2(n17083), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17056) );
  NOR2_X1 U20317 ( .A1(n18064), .A2(n18048), .ZN(n17066) );
  NAND2_X1 U20318 ( .A1(n17066), .A2(n17053), .ZN(n17077) );
  INV_X1 U20319 ( .A(n17077), .ZN(n17064) );
  NAND2_X1 U20320 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17064), .ZN(
        n17063) );
  AOI21_X1 U20321 ( .B1(n21455), .B2(n17063), .A(n17054), .ZN(n18022) );
  OAI21_X1 U20322 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17063), .A(
        n17157), .ZN(n17068) );
  XOR2_X1 U20323 ( .A(n18022), .B(n17068), .Z(n17055) );
  OAI22_X1 U20324 ( .A1(n17057), .A2(n17056), .B1(n17186), .B2(n17055), .ZN(
        n17058) );
  AOI211_X1 U20325 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n17154), .A(n18479), .B(
        n17058), .ZN(n17061) );
  OAI211_X1 U20326 ( .C1(n17069), .C2(n17429), .A(n17176), .B(n17059), .ZN(
        n17060) );
  OAI211_X1 U20327 ( .C1(n17184), .C2(n21455), .A(n17061), .B(n17060), .ZN(
        P3_U2660) );
  NAND2_X1 U20328 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17083), .ZN(n17076) );
  OAI21_X1 U20329 ( .B1(n17062), .B2(n17187), .A(n17197), .ZN(n17097) );
  AOI21_X1 U20330 ( .B1(n17083), .B2(n19049), .A(n17097), .ZN(n17075) );
  OAI21_X1 U20331 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17064), .A(
        n17063), .ZN(n18035) );
  OAI21_X1 U20332 ( .B1(n17066), .B2(n17065), .A(n17090), .ZN(n17079) );
  INV_X1 U20333 ( .A(n18035), .ZN(n17067) );
  AOI221_X1 U20334 ( .B1(n17068), .B2(n18035), .C1(n17079), .C2(n17067), .A(
        n17186), .ZN(n17073) );
  AOI211_X1 U20335 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17084), .A(n17069), .B(
        n17194), .ZN(n17072) );
  INV_X1 U20336 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17448) );
  OAI22_X1 U20337 ( .A1(n17070), .A2(n17184), .B1(n17448), .B2(n17193), .ZN(
        n17071) );
  NOR4_X1 U20338 ( .A1(n18479), .A2(n17073), .A3(n17072), .A4(n17071), .ZN(
        n17074) );
  OAI221_X1 U20339 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n17076), .C1(n19050), 
        .C2(n17075), .A(n17074), .ZN(P3_U2661) );
  AOI22_X1 U20340 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17115), .B1(
        P3_EBX_REG_9__SCAN_IN), .B2(n17154), .ZN(n17088) );
  NOR2_X1 U20341 ( .A1(n18064), .A2(n17102), .ZN(n17089) );
  OAI21_X1 U20342 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17089), .A(
        n17077), .ZN(n17078) );
  AOI21_X1 U20343 ( .B1(n17089), .B2(n17117), .A(n17078), .ZN(n17081) );
  INV_X1 U20344 ( .A(n17078), .ZN(n18052) );
  NOR2_X1 U20345 ( .A1(n18052), .A2(n17079), .ZN(n17080) );
  AOI211_X1 U20346 ( .C1(n17157), .C2(n17081), .A(n17080), .B(n17186), .ZN(
        n17082) );
  AOI221_X1 U20347 ( .B1(n17083), .B2(n19049), .C1(n17097), .C2(
        P3_REIP_REG_9__SCAN_IN), .A(n17082), .ZN(n17087) );
  OAI211_X1 U20348 ( .C1(n17093), .C2(n17085), .A(n17176), .B(n17084), .ZN(
        n17086) );
  NAND4_X1 U20349 ( .A1(n17088), .A2(n17087), .A3(n18484), .A4(n17086), .ZN(
        P3_U2662) );
  AOI21_X1 U20350 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17154), .A(n18479), .ZN(
        n17101) );
  AOI21_X1 U20351 ( .B1(n18064), .B2(n17102), .A(n17089), .ZN(n17092) );
  INV_X1 U20352 ( .A(n17092), .ZN(n18061) );
  AOI221_X1 U20353 ( .B1(n17092), .B2(n17091), .C1(n18061), .C2(n17090), .A(
        n17186), .ZN(n17095) );
  AOI211_X1 U20354 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17110), .A(n17093), .B(
        n17194), .ZN(n17094) );
  AOI211_X1 U20355 ( .C1(n17115), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17095), .B(n17094), .ZN(n17100) );
  NOR2_X1 U20356 ( .A1(n17187), .A2(n17096), .ZN(n17098) );
  OAI21_X1 U20357 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n17098), .A(n17097), .ZN(
        n17099) );
  NAND3_X1 U20358 ( .A1(n17101), .A2(n17100), .A3(n17099), .ZN(P3_U2663) );
  INV_X1 U20359 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18084) );
  OAI221_X1 U20360 ( .B1(n17187), .B2(P3_REIP_REG_6__SCAN_IN), .C1(n17187), 
        .C2(n17120), .A(n17197), .ZN(n17109) );
  OAI21_X1 U20361 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17118), .A(
        n17102), .ZN(n18080) );
  INV_X1 U20362 ( .A(n18080), .ZN(n17105) );
  AOI221_X1 U20363 ( .B1(n17105), .B2(n17104), .C1(n18080), .C2(n17103), .A(
        n17186), .ZN(n17108) );
  INV_X1 U20364 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19045) );
  NAND4_X1 U20365 ( .A1(n17173), .A2(P3_REIP_REG_6__SCAN_IN), .A3(n17120), 
        .A4(n19045), .ZN(n17106) );
  OAI211_X1 U20366 ( .C1(n17467), .C2(n17193), .A(n18484), .B(n17106), .ZN(
        n17107) );
  AOI211_X1 U20367 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n17109), .A(n17108), .B(
        n17107), .ZN(n17112) );
  OAI211_X1 U20368 ( .C1(n17116), .C2(n17467), .A(n17176), .B(n17110), .ZN(
        n17111) );
  OAI211_X1 U20369 ( .C1(n17184), .C2(n18084), .A(n17112), .B(n17111), .ZN(
        P3_U2664) );
  NOR2_X1 U20370 ( .A1(n17120), .A2(n17187), .ZN(n17130) );
  NOR2_X1 U20371 ( .A1(n17183), .A2(n17130), .ZN(n17133) );
  INV_X1 U20372 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19043) );
  OR2_X1 U20373 ( .A1(n21330), .A2(n18097), .ZN(n17127) );
  AOI21_X1 U20374 ( .B1(n18098), .B2(n17127), .A(n17118), .ZN(n18100) );
  AOI21_X1 U20375 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17157), .A(
        n17113), .ZN(n17114) );
  AOI22_X1 U20376 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17115), .B1(
        n18100), .B2(n17114), .ZN(n17126) );
  AOI211_X1 U20377 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17136), .A(n17116), .B(
        n17194), .ZN(n17124) );
  NAND2_X1 U20378 ( .A1(n17118), .A2(n17117), .ZN(n17119) );
  NAND3_X1 U20379 ( .A1(n17147), .A2(n17157), .A3(n17119), .ZN(n17122) );
  NAND3_X1 U20380 ( .A1(n17173), .A2(n17120), .A3(n19043), .ZN(n17121) );
  OAI211_X1 U20381 ( .C1(n18100), .C2(n17122), .A(n18484), .B(n17121), .ZN(
        n17123) );
  AOI211_X1 U20382 ( .C1(n17154), .C2(P3_EBX_REG_6__SCAN_IN), .A(n17124), .B(
        n17123), .ZN(n17125) );
  OAI211_X1 U20383 ( .C1(n17133), .C2(n19043), .A(n17126), .B(n17125), .ZN(
        P3_U2665) );
  NAND2_X1 U20384 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18106), .ZN(
        n17128) );
  INV_X1 U20385 ( .A(n17128), .ZN(n17139) );
  OAI21_X1 U20386 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17139), .A(
        n17127), .ZN(n18113) );
  OAI21_X1 U20387 ( .B1(n17128), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17157), .ZN(n17145) );
  XOR2_X1 U20388 ( .A(n18113), .B(n17145), .Z(n17135) );
  INV_X1 U20389 ( .A(n17129), .ZN(n17131) );
  AOI22_X1 U20390 ( .A1(n17131), .A2(n17130), .B1(P3_EBX_REG_5__SCAN_IN), .B2(
        n17154), .ZN(n17132) );
  OAI211_X1 U20391 ( .C1(n17133), .C2(n19041), .A(n17132), .B(n18484), .ZN(
        n17134) );
  AOI21_X1 U20392 ( .B1(n17135), .B2(n17147), .A(n17134), .ZN(n17138) );
  OAI211_X1 U20393 ( .C1(n17140), .C2(n17499), .A(n17176), .B(n17136), .ZN(
        n17137) );
  OAI211_X1 U20394 ( .C1(n17184), .C2(n10171), .A(n17138), .B(n17137), .ZN(
        P3_U2666) );
  AOI21_X1 U20395 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17154), .A(n18479), .ZN(
        n17151) );
  NOR2_X1 U20396 ( .A1(n17157), .A2(n17186), .ZN(n17171) );
  NAND2_X1 U20397 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17144), .ZN(
        n17155) );
  AOI21_X1 U20398 ( .B1(n18122), .B2(n17155), .A(n17139), .ZN(n18124) );
  AOI211_X1 U20399 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17164), .A(n17140), .B(
        n17194), .ZN(n17143) );
  INV_X1 U20400 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19039) );
  NAND3_X1 U20401 ( .A1(n17173), .A2(n17152), .A3(n19039), .ZN(n17141) );
  OAI21_X1 U20402 ( .B1(n17184), .B2(n18122), .A(n17141), .ZN(n17142) );
  AOI211_X1 U20403 ( .C1(n17171), .C2(n18124), .A(n17143), .B(n17142), .ZN(
        n17150) );
  NAND2_X1 U20404 ( .A1(n17144), .A2(n18122), .ZN(n18127) );
  OAI22_X1 U20405 ( .A1(n18124), .A2(n17145), .B1(n17168), .B2(n18127), .ZN(
        n17146) );
  OAI21_X1 U20406 ( .B1(n17152), .B2(n17187), .A(n17197), .ZN(n17163) );
  AOI22_X1 U20407 ( .A1(n17147), .A2(n17146), .B1(P3_REIP_REG_4__SCAN_IN), 
        .B2(n17163), .ZN(n17149) );
  INV_X1 U20408 ( .A(n19168), .ZN(n19164) );
  NOR2_X1 U20409 ( .A1(n17683), .A2(n19164), .ZN(n17195) );
  OAI21_X1 U20410 ( .B1(n17458), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n17195), .ZN(n17148) );
  NAND4_X1 U20411 ( .A1(n17151), .A2(n17150), .A3(n17149), .A4(n17148), .ZN(
        P3_U2667) );
  OR2_X1 U20412 ( .A1(n17187), .A2(n17152), .ZN(n17161) );
  NOR2_X1 U20413 ( .A1(n19128), .A2(n17153), .ZN(n18954) );
  OAI21_X1 U20414 ( .B1(n18954), .B2(n19108), .A(n17435), .ZN(n19105) );
  AOI22_X1 U20415 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17154), .B1(n17195), .B2(
        n19105), .ZN(n17160) );
  NOR2_X1 U20416 ( .A1(n21330), .A2(n18153), .ZN(n17156) );
  OAI21_X1 U20417 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17156), .A(
        n17155), .ZN(n18137) );
  OAI21_X1 U20418 ( .B1(n18153), .B2(n17168), .A(n17157), .ZN(n17167) );
  AOI21_X1 U20419 ( .B1(n18137), .B2(n17167), .A(n17186), .ZN(n17158) );
  OAI21_X1 U20420 ( .B1(n18137), .B2(n17167), .A(n17158), .ZN(n17159) );
  OAI211_X1 U20421 ( .C1(n17161), .C2(n17172), .A(n17160), .B(n17159), .ZN(
        n17162) );
  AOI21_X1 U20422 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n17163), .A(n17162), .ZN(
        n17166) );
  OAI211_X1 U20423 ( .C1(n17174), .C2(n21367), .A(n17176), .B(n17164), .ZN(
        n17165) );
  OAI211_X1 U20424 ( .C1(n17184), .C2(n18135), .A(n17166), .B(n17165), .ZN(
        P3_U2668) );
  AOI21_X1 U20425 ( .B1(n13017), .B2(n18976), .A(n18954), .ZN(n19111) );
  AOI22_X1 U20426 ( .A1(n17183), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n19111), 
        .B2(n17195), .ZN(n17181) );
  OAI22_X1 U20427 ( .A1(n21330), .A2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n18153), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18145) );
  AOI211_X1 U20428 ( .C1(n18145), .C2(n17168), .A(n17186), .B(n17167), .ZN(
        n17170) );
  OAI22_X1 U20429 ( .A1(n18153), .A2(n17184), .B1(n17512), .B2(n17193), .ZN(
        n17169) );
  AOI211_X1 U20430 ( .C1(n17171), .C2(n18145), .A(n17170), .B(n17169), .ZN(
        n17180) );
  OAI211_X1 U20431 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n17173), .B(n17172), .ZN(n17179) );
  NOR2_X1 U20432 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17177) );
  INV_X1 U20433 ( .A(n17174), .ZN(n17175) );
  OAI211_X1 U20434 ( .C1(n17177), .C2(n17512), .A(n17176), .B(n17175), .ZN(
        n17178) );
  NAND4_X1 U20435 ( .A1(n17181), .A2(n17180), .A3(n17179), .A4(n17178), .ZN(
        P3_U2669) );
  OAI21_X1 U20436 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17513), .ZN(n17521) );
  AND2_X1 U20437 ( .A1(n18976), .A2(n17182), .ZN(n19118) );
  AOI22_X1 U20438 ( .A1(n17183), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n19118), 
        .B2(n17195), .ZN(n17192) );
  OAI21_X1 U20439 ( .B1(n17186), .B2(n17185), .A(n17184), .ZN(n17189) );
  INV_X1 U20440 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17520) );
  OAI22_X1 U20441 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17187), .B1(n17520), 
        .B2(n17193), .ZN(n17188) );
  AOI221_X1 U20442 ( .B1(n17190), .B2(n21330), .C1(n17189), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17188), .ZN(n17191) );
  OAI211_X1 U20443 ( .C1(n17194), .C2(n17521), .A(n17192), .B(n17191), .ZN(
        P3_U2670) );
  INV_X1 U20444 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19136) );
  NAND2_X1 U20445 ( .A1(n17194), .A2(n17193), .ZN(n17196) );
  AOI22_X1 U20446 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17196), .B1(n17195), .B2(
        n19128), .ZN(n17200) );
  NAND3_X1 U20447 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17198), .A3(
        n17197), .ZN(n17199) );
  OAI211_X1 U20448 ( .C1(n17201), .C2(n19136), .A(n17200), .B(n17199), .ZN(
        P3_U2671) );
  INV_X1 U20449 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17207) );
  NOR4_X1 U20450 ( .A1(n17237), .A2(n17253), .A3(n17249), .A4(n17295), .ZN(
        n17202) );
  NAND3_X1 U20451 ( .A1(n17203), .A2(n17238), .A3(n17202), .ZN(n17206) );
  NOR2_X1 U20452 ( .A1(n17207), .A2(n17206), .ZN(n17232) );
  NAND2_X1 U20453 ( .A1(n17517), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17205) );
  NAND2_X1 U20454 ( .A1(n17232), .A2(n17612), .ZN(n17204) );
  OAI22_X1 U20455 ( .A1(n17232), .A2(n17205), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17204), .ZN(P3_U2672) );
  NAND2_X1 U20456 ( .A1(n17207), .A2(n17206), .ZN(n17208) );
  NAND2_X1 U20457 ( .A1(n17208), .A2(n17517), .ZN(n17231) );
  AOI22_X1 U20458 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20459 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17343), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17449), .ZN(n17211) );
  AOI22_X1 U20460 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n9822), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n13090), .ZN(n17210) );
  AOI22_X1 U20461 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17460), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17209) );
  NAND4_X1 U20462 ( .A1(n17212), .A2(n17211), .A3(n17210), .A4(n17209), .ZN(
        n17218) );
  AOI22_X1 U20463 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17417), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17450), .ZN(n17216) );
  AOI22_X1 U20464 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17456), .ZN(n17215) );
  AOI22_X1 U20465 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17457), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U20466 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17213) );
  NAND4_X1 U20467 ( .A1(n17216), .A2(n17215), .A3(n17214), .A4(n17213), .ZN(
        n17217) );
  NOR2_X1 U20468 ( .A1(n17218), .A2(n17217), .ZN(n17230) );
  AOI22_X1 U20469 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20470 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20471 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17219) );
  OAI21_X1 U20472 ( .B1(n17220), .B2(n21366), .A(n17219), .ZN(n17226) );
  AOI22_X1 U20473 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20474 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20475 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15918), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20476 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17221) );
  NAND4_X1 U20477 ( .A1(n17224), .A2(n17223), .A3(n17222), .A4(n17221), .ZN(
        n17225) );
  AOI211_X1 U20478 ( .C1(n17343), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17226), .B(n17225), .ZN(n17227) );
  NAND3_X1 U20479 ( .A1(n17229), .A2(n17228), .A3(n17227), .ZN(n17234) );
  NAND2_X1 U20480 ( .A1(n17235), .A2(n17234), .ZN(n17233) );
  XNOR2_X1 U20481 ( .A(n17230), .B(n17233), .ZN(n17534) );
  OAI22_X1 U20482 ( .A1(n17232), .A2(n17231), .B1(n17534), .B2(n17517), .ZN(
        P3_U2673) );
  OAI21_X1 U20483 ( .B1(n17235), .B2(n17234), .A(n17233), .ZN(n17542) );
  OAI222_X1 U20484 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17243), .B1(
        P3_EBX_REG_29__SCAN_IN), .B2(n17238), .C1(n17237), .C2(n17236), .ZN(
        n17239) );
  OAI21_X1 U20485 ( .B1(n17542), .B2(n17517), .A(n17239), .ZN(P3_U2674) );
  OAI21_X1 U20486 ( .B1(n17246), .B2(n17241), .A(n17240), .ZN(n17550) );
  AOI22_X1 U20487 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17244), .B1(n17243), 
        .B2(n17242), .ZN(n17245) );
  OAI21_X1 U20488 ( .B1(n17550), .B2(n17517), .A(n17245), .ZN(P3_U2676) );
  AOI21_X1 U20489 ( .B1(n17247), .B2(n17254), .A(n17246), .ZN(n17551) );
  NOR2_X1 U20490 ( .A1(n17249), .A2(n17248), .ZN(n17257) );
  AOI22_X1 U20491 ( .A1(n17551), .A2(n17523), .B1(n17257), .B2(n17250), .ZN(
        n17251) );
  OAI21_X1 U20492 ( .B1(n17253), .B2(n17252), .A(n17251), .ZN(P3_U2677) );
  AOI21_X1 U20493 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17517), .A(n17263), .ZN(
        n17256) );
  OAI21_X1 U20494 ( .B1(n17259), .B2(n17255), .A(n17254), .ZN(n17560) );
  OAI22_X1 U20495 ( .A1(n17257), .A2(n17256), .B1(n17560), .B2(n17517), .ZN(
        P3_U2678) );
  NAND2_X1 U20496 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17297), .ZN(n17270) );
  NOR3_X1 U20497 ( .A1(n17258), .A2(n17271), .A3(n17270), .ZN(n17268) );
  AOI21_X1 U20498 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17517), .A(n17268), .ZN(
        n17262) );
  AOI21_X1 U20499 ( .B1(n17260), .B2(n17264), .A(n17259), .ZN(n17561) );
  INV_X1 U20500 ( .A(n17561), .ZN(n17261) );
  OAI22_X1 U20501 ( .A1(n17263), .A2(n17262), .B1(n17261), .B2(n17517), .ZN(
        P3_U2679) );
  NOR2_X1 U20502 ( .A1(n17271), .A2(n17270), .ZN(n17269) );
  AOI21_X1 U20503 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17517), .A(n17269), .ZN(
        n17267) );
  OAI21_X1 U20504 ( .B1(n17266), .B2(n17265), .A(n17264), .ZN(n17573) );
  OAI22_X1 U20505 ( .A1(n17268), .A2(n17267), .B1(n17573), .B2(n17517), .ZN(
        P3_U2680) );
  INV_X1 U20506 ( .A(n17269), .ZN(n17283) );
  OAI21_X1 U20507 ( .B1(n17271), .B2(n17523), .A(n17270), .ZN(n17282) );
  AOI22_X1 U20508 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20509 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20510 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17272) );
  OAI21_X1 U20511 ( .B1(n10391), .B2(n21366), .A(n17272), .ZN(n17278) );
  AOI22_X1 U20512 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20513 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U20514 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U20515 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17273) );
  NAND4_X1 U20516 ( .A1(n17276), .A2(n17275), .A3(n17274), .A4(n17273), .ZN(
        n17277) );
  AOI211_X1 U20517 ( .C1(n17479), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n17278), .B(n17277), .ZN(n17279) );
  NAND3_X1 U20518 ( .A1(n17281), .A2(n17280), .A3(n17279), .ZN(n17575) );
  AOI22_X1 U20519 ( .A1(n17283), .A2(n17282), .B1(n17575), .B2(n17523), .ZN(
        n17284) );
  INV_X1 U20520 ( .A(n17284), .ZN(P3_U2681) );
  AOI22_X1 U20521 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U20522 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20523 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20524 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17285) );
  NAND4_X1 U20525 ( .A1(n17288), .A2(n17287), .A3(n17286), .A4(n17285), .ZN(
        n17294) );
  AOI22_X1 U20526 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U20527 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17458), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20528 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17290) );
  AOI22_X1 U20529 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17289) );
  NAND4_X1 U20530 ( .A1(n17292), .A2(n17291), .A3(n17290), .A4(n17289), .ZN(
        n17293) );
  NOR2_X1 U20531 ( .A1(n17294), .A2(n17293), .ZN(n17581) );
  AND2_X1 U20532 ( .A1(n17517), .A2(n17295), .ZN(n17310) );
  AOI22_X1 U20533 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17310), .B1(n17297), 
        .B2(n17296), .ZN(n17298) );
  OAI21_X1 U20534 ( .B1(n17581), .B2(n17517), .A(n17298), .ZN(P3_U2682) );
  AOI22_X1 U20535 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20536 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20537 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17299) );
  OAI21_X1 U20538 ( .B1(n10029), .B2(n17300), .A(n17299), .ZN(n17306) );
  AOI22_X1 U20539 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17458), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17304) );
  AOI22_X1 U20540 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17303) );
  AOI22_X1 U20541 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U20542 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17301) );
  NAND4_X1 U20543 ( .A1(n17304), .A2(n17303), .A3(n17302), .A4(n17301), .ZN(
        n17305) );
  AOI211_X1 U20544 ( .C1(n17479), .C2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n17306), .B(n17305), .ZN(n17307) );
  NAND3_X1 U20545 ( .A1(n17309), .A2(n17308), .A3(n17307), .ZN(n17585) );
  INV_X1 U20546 ( .A(n17585), .ZN(n17312) );
  AND2_X1 U20547 ( .A1(n17612), .A2(n17323), .ZN(n17325) );
  OAI221_X1 U20548 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(P3_EBX_REG_19__SCAN_IN), 
        .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17325), .A(n17310), .ZN(n17311) );
  OAI21_X1 U20549 ( .B1(n17312), .B2(n17517), .A(n17311), .ZN(P3_U2683) );
  AOI22_X1 U20550 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U20551 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U20552 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U20553 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17313) );
  NAND4_X1 U20554 ( .A1(n17316), .A2(n17315), .A3(n17314), .A4(n17313), .ZN(
        n17322) );
  AOI22_X1 U20555 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17320) );
  AOI22_X1 U20556 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17319) );
  AOI22_X1 U20557 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U20558 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17317) );
  NAND4_X1 U20559 ( .A1(n17320), .A2(n17319), .A3(n17318), .A4(n17317), .ZN(
        n17321) );
  NOR2_X1 U20560 ( .A1(n17322), .A2(n17321), .ZN(n17594) );
  NOR2_X1 U20561 ( .A1(n17523), .A2(n17323), .ZN(n17341) );
  AOI22_X1 U20562 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17341), .B1(n17325), 
        .B2(n17324), .ZN(n17326) );
  OAI21_X1 U20563 ( .B1(n17594), .B2(n17517), .A(n17326), .ZN(P3_U2684) );
  AOI22_X1 U20564 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U20565 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20566 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U20567 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17327) );
  NAND4_X1 U20568 ( .A1(n17330), .A2(n17329), .A3(n17328), .A4(n17327), .ZN(
        n17336) );
  AOI22_X1 U20569 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U20570 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17333) );
  AOI22_X1 U20571 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17332) );
  AOI22_X1 U20572 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17331) );
  NAND4_X1 U20573 ( .A1(n17334), .A2(n17333), .A3(n17332), .A4(n17331), .ZN(
        n17335) );
  NOR2_X1 U20574 ( .A1(n17336), .A2(n17335), .ZN(n17598) );
  NAND2_X1 U20575 ( .A1(n17612), .A2(n17411), .ZN(n17412) );
  NOR2_X1 U20576 ( .A1(n17337), .A2(n17412), .ZN(n17356) );
  NAND2_X1 U20577 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17356), .ZN(n17355) );
  NOR2_X1 U20578 ( .A1(n17338), .A2(n17355), .ZN(n17340) );
  AOI22_X1 U20579 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17341), .B1(n17340), 
        .B2(n17339), .ZN(n17342) );
  OAI21_X1 U20580 ( .B1(n17598), .B2(n17517), .A(n17342), .ZN(P3_U2685) );
  AOI22_X1 U20581 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17347) );
  AOI22_X1 U20582 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U20583 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17345) );
  AOI22_X1 U20584 ( .A1(n17343), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17344) );
  NAND4_X1 U20585 ( .A1(n17347), .A2(n17346), .A3(n17345), .A4(n17344), .ZN(
        n17353) );
  AOI22_X1 U20586 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17351) );
  AOI22_X1 U20587 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17350) );
  AOI22_X1 U20588 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17349) );
  AOI22_X1 U20589 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17348) );
  NAND4_X1 U20590 ( .A1(n17351), .A2(n17350), .A3(n17349), .A4(n17348), .ZN(
        n17352) );
  NOR2_X1 U20591 ( .A1(n17353), .A2(n17352), .ZN(n17605) );
  NAND3_X1 U20592 ( .A1(n17355), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17517), 
        .ZN(n17354) );
  OAI221_X1 U20593 ( .B1(n17355), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n17517), 
        .C2(n17605), .A(n17354), .ZN(P3_U2686) );
  INV_X1 U20594 ( .A(n17356), .ZN(n17381) );
  AOI22_X1 U20595 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17360) );
  AOI22_X1 U20596 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20597 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U20598 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17357) );
  NAND4_X1 U20599 ( .A1(n17360), .A2(n17359), .A3(n17358), .A4(n17357), .ZN(
        n17366) );
  AOI22_X1 U20600 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17364) );
  AOI22_X1 U20601 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U20602 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17362) );
  AOI22_X1 U20603 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17361) );
  NAND4_X1 U20604 ( .A1(n17364), .A2(n17363), .A3(n17362), .A4(n17361), .ZN(
        n17365) );
  NOR2_X1 U20605 ( .A1(n17366), .A2(n17365), .ZN(n17611) );
  NAND3_X1 U20606 ( .A1(n17381), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17517), 
        .ZN(n17367) );
  OAI221_X1 U20607 ( .B1(n17381), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17517), 
        .C2(n17611), .A(n17367), .ZN(P3_U2687) );
  AOI22_X1 U20608 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17368), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17460), .ZN(n17379) );
  AOI22_X1 U20609 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17450), .ZN(n17378) );
  AOI22_X1 U20610 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17449), .ZN(n17369) );
  OAI21_X1 U20611 ( .B1(n17370), .B2(n21409), .A(n17369), .ZN(n17376) );
  AOI22_X1 U20612 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17456), .ZN(n17374) );
  AOI22_X1 U20613 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17459), .ZN(n17373) );
  AOI22_X1 U20614 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17457), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17372) );
  AOI22_X1 U20615 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n9822), .ZN(n17371) );
  NAND4_X1 U20616 ( .A1(n17374), .A2(n17373), .A3(n17372), .A4(n17371), .ZN(
        n17375) );
  AOI211_X1 U20617 ( .C1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .C2(n17472), .A(
        n17376), .B(n17375), .ZN(n17377) );
  NAND3_X1 U20618 ( .A1(n17379), .A2(n17378), .A3(n17377), .ZN(n17615) );
  INV_X1 U20619 ( .A(n17615), .ZN(n17384) );
  INV_X1 U20620 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17400) );
  INV_X1 U20621 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17413) );
  NOR3_X1 U20622 ( .A1(n17400), .A2(n17396), .A3(n17413), .ZN(n17380) );
  AOI21_X1 U20623 ( .B1(n17411), .B2(n17380), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n17383) );
  NAND2_X1 U20624 ( .A1(n17517), .A2(n17381), .ZN(n17382) );
  OAI22_X1 U20625 ( .A1(n17384), .A2(n17517), .B1(n17383), .B2(n17382), .ZN(
        P3_U2688) );
  AOI22_X1 U20626 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20627 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U20628 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U20629 ( .B1(n9917), .B2(n21366), .A(n17385), .ZN(n17392) );
  AOI22_X1 U20630 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20631 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U20632 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U20633 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17387) );
  NAND4_X1 U20634 ( .A1(n17390), .A2(n17389), .A3(n17388), .A4(n17387), .ZN(
        n17391) );
  AOI211_X1 U20635 ( .C1(n17449), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n17392), .B(n17391), .ZN(n17393) );
  NAND3_X1 U20636 ( .A1(n17395), .A2(n17394), .A3(n17393), .ZN(n17619) );
  NOR4_X1 U20637 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17396), .A3(n17413), .A4(
        n17412), .ZN(n17397) );
  AOI21_X1 U20638 ( .B1(n17523), .B2(n17619), .A(n17397), .ZN(n17398) );
  OAI21_X1 U20639 ( .B1(n17400), .B2(n17399), .A(n17398), .ZN(P3_U2689) );
  AOI22_X1 U20640 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17404) );
  AOI22_X1 U20641 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17403) );
  AOI22_X1 U20642 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U20643 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17401) );
  NAND4_X1 U20644 ( .A1(n17404), .A2(n17403), .A3(n17402), .A4(n17401), .ZN(
        n17410) );
  AOI22_X1 U20645 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20646 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U20647 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U20648 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17405) );
  NAND4_X1 U20649 ( .A1(n17408), .A2(n17407), .A3(n17406), .A4(n17405), .ZN(
        n17409) );
  NOR2_X1 U20650 ( .A1(n17410), .A2(n17409), .ZN(n17628) );
  OR2_X1 U20651 ( .A1(n17523), .A2(n17411), .ZN(n17430) );
  OAI22_X1 U20652 ( .A1(n17413), .A2(n17430), .B1(n17412), .B2(
        P3_EBX_REG_12__SCAN_IN), .ZN(n17414) );
  INV_X1 U20653 ( .A(n17414), .ZN(n17415) );
  OAI21_X1 U20654 ( .B1(n17628), .B2(n17517), .A(n17415), .ZN(P3_U2691) );
  AOI22_X1 U20655 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U20656 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17425) );
  INV_X1 U20657 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n21397) );
  AOI22_X1 U20658 ( .A1(n13090), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17416) );
  OAI21_X1 U20659 ( .B1(n17435), .B2(n21397), .A(n17416), .ZN(n17423) );
  AOI22_X1 U20660 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17421) );
  AOI22_X1 U20661 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20662 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17419) );
  AOI22_X1 U20663 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17418) );
  NAND4_X1 U20664 ( .A1(n17421), .A2(n17420), .A3(n17419), .A4(n17418), .ZN(
        n17422) );
  AOI211_X1 U20665 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n17423), .B(n17422), .ZN(n17424) );
  NAND3_X1 U20666 ( .A1(n17426), .A2(n17425), .A3(n17424), .ZN(n17632) );
  NAND2_X1 U20667 ( .A1(n17523), .A2(n17632), .ZN(n17427) );
  OAI221_X1 U20668 ( .B1(n17430), .B2(n17429), .C1(n17430), .C2(n17428), .A(
        n17427), .ZN(P3_U2692) );
  INV_X1 U20669 ( .A(n17431), .ZN(n17445) );
  NAND2_X1 U20670 ( .A1(n17517), .A2(n17445), .ZN(n17468) );
  AOI22_X1 U20671 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20672 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20673 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17434) );
  OAI21_X1 U20674 ( .B1(n17435), .B2(n21467), .A(n17434), .ZN(n17441) );
  AOI22_X1 U20675 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17458), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U20676 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U20677 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U20678 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17436) );
  NAND4_X1 U20679 ( .A1(n17439), .A2(n17438), .A3(n17437), .A4(n17436), .ZN(
        n17440) );
  AOI211_X1 U20680 ( .C1(n17479), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n17441), .B(n17440), .ZN(n17442) );
  NAND3_X1 U20681 ( .A1(n17444), .A2(n17443), .A3(n17442), .ZN(n17635) );
  NOR3_X1 U20682 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18545), .A3(n17445), .ZN(
        n17446) );
  AOI21_X1 U20683 ( .B1(n17523), .B2(n17635), .A(n17446), .ZN(n17447) );
  OAI21_X1 U20684 ( .B1(n17448), .B2(n17468), .A(n17447), .ZN(P3_U2693) );
  AOI22_X1 U20685 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U20686 ( .A1(n17451), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20687 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U20688 ( .A1(n15908), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17452) );
  NAND4_X1 U20689 ( .A1(n17455), .A2(n17454), .A3(n17453), .A4(n17452), .ZN(
        n17466) );
  AOI22_X1 U20690 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17464) );
  AOI22_X1 U20691 ( .A1(n17458), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17432), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17463) );
  AOI22_X1 U20692 ( .A1(n17459), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U20693 ( .A1(n15918), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9849), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17461) );
  NAND4_X1 U20694 ( .A1(n17464), .A2(n17463), .A3(n17462), .A4(n17461), .ZN(
        n17465) );
  NOR2_X1 U20695 ( .A1(n17466), .A2(n17465), .ZN(n17639) );
  INV_X1 U20696 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17498) );
  NOR4_X1 U20697 ( .A1(n17467), .A2(n17498), .A3(n17499), .A4(n17502), .ZN(
        n17488) );
  AOI21_X1 U20698 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17488), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n17469) );
  OAI22_X1 U20699 ( .A1(n17639), .A2(n17517), .B1(n17469), .B2(n17468), .ZN(
        P3_U2694) );
  AOI22_X1 U20700 ( .A1(n9924), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U20701 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20702 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17475) );
  AOI22_X1 U20703 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17474) );
  NAND4_X1 U20704 ( .A1(n17477), .A2(n17476), .A3(n17475), .A4(n17474), .ZN(
        n17487) );
  AOI22_X1 U20705 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17478), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17485) );
  AOI22_X1 U20706 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U20707 ( .A1(n9849), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17483) );
  AOI22_X1 U20708 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17343), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17482) );
  NAND4_X1 U20709 ( .A1(n17485), .A2(n17484), .A3(n17483), .A4(n17482), .ZN(
        n17486) );
  NOR2_X1 U20710 ( .A1(n17487), .A2(n17486), .ZN(n17646) );
  NOR2_X1 U20711 ( .A1(n17523), .A2(n17488), .ZN(n17492) );
  INV_X1 U20712 ( .A(n17488), .ZN(n17489) );
  NOR3_X1 U20713 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18545), .A3(n17489), .ZN(
        n17490) );
  AOI21_X1 U20714 ( .B1(n17492), .B2(P3_EBX_REG_8__SCAN_IN), .A(n17490), .ZN(
        n17491) );
  OAI21_X1 U20715 ( .B1(n17646), .B2(n17517), .A(n17491), .ZN(P3_U2695) );
  NOR3_X1 U20716 ( .A1(n18545), .A2(n17499), .A3(n17502), .ZN(n17496) );
  AOI21_X1 U20717 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17496), .A(
        P3_EBX_REG_7__SCAN_IN), .ZN(n17495) );
  INV_X1 U20718 ( .A(n17492), .ZN(n17494) );
  INV_X1 U20719 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17493) );
  OAI22_X1 U20720 ( .A1(n17495), .A2(n17494), .B1(n17493), .B2(n17517), .ZN(
        P3_U2696) );
  OAI21_X1 U20721 ( .B1(n17499), .B2(n17502), .A(n17517), .ZN(n17500) );
  AOI22_X1 U20722 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17523), .B1(
        n17496), .B2(n17498), .ZN(n17497) );
  OAI21_X1 U20723 ( .B1(n17498), .B2(n17500), .A(n17497), .ZN(P3_U2697) );
  AND2_X1 U20724 ( .A1(n17499), .A2(n17502), .ZN(n17501) );
  INV_X1 U20725 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n21499) );
  OAI22_X1 U20726 ( .A1(n17501), .A2(n17500), .B1(n21499), .B2(n17517), .ZN(
        P3_U2698) );
  INV_X1 U20727 ( .A(n17502), .ZN(n17507) );
  INV_X1 U20728 ( .A(n17525), .ZN(n17503) );
  NAND2_X1 U20729 ( .A1(n17504), .A2(n17503), .ZN(n17514) );
  NOR2_X1 U20730 ( .A1(n21367), .A2(n17514), .ZN(n17511) );
  AOI21_X1 U20731 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17517), .A(n17511), .ZN(
        n17506) );
  INV_X1 U20732 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17505) );
  OAI22_X1 U20733 ( .A1(n17507), .A2(n17506), .B1(n17505), .B2(n17517), .ZN(
        P3_U2699) );
  INV_X1 U20734 ( .A(n17514), .ZN(n17508) );
  AOI21_X1 U20735 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17517), .A(n17508), .ZN(
        n17510) );
  INV_X1 U20736 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17509) );
  OAI22_X1 U20737 ( .A1(n17511), .A2(n17510), .B1(n17509), .B2(n17517), .ZN(
        P3_U2700) );
  OAI221_X1 U20738 ( .B1(n17513), .B2(n17522), .C1(n17612), .C2(n17522), .A(
        n17512), .ZN(n17515) );
  OAI211_X1 U20739 ( .C1(n17517), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17515), .B(n17514), .ZN(n17516) );
  INV_X1 U20740 ( .A(n17516), .ZN(P3_U2701) );
  OAI222_X1 U20741 ( .A1(n17521), .A2(n17525), .B1(n17520), .B2(n17519), .C1(
        n17518), .C2(n17517), .ZN(P3_U2702) );
  AOI22_X1 U20742 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17523), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17522), .ZN(n17524) );
  OAI21_X1 U20743 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17525), .A(n17524), .ZN(
        P3_U2703) );
  NOR2_X2 U20744 ( .A1(n17663), .A2(n17526), .ZN(n17606) );
  INV_X1 U20745 ( .A(n17606), .ZN(n17580) );
  INV_X1 U20746 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17745) );
  INV_X1 U20747 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17742) );
  INV_X1 U20748 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17740) );
  INV_X1 U20749 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17738) );
  NAND2_X1 U20750 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n17676) );
  NOR2_X1 U20751 ( .A1(n17674), .A2(n17676), .ZN(n17669) );
  INV_X1 U20752 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21531) );
  INV_X1 U20753 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17765) );
  INV_X1 U20754 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17758) );
  INV_X1 U20755 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17756) );
  NOR4_X1 U20756 ( .A1(n21531), .A2(n17765), .A3(n17758), .A4(n17756), .ZN(
        n17527) );
  NAND4_X1 U20757 ( .A1(n17669), .A2(P3_EAX_REG_6__SCAN_IN), .A3(
        P3_EAX_REG_5__SCAN_IN), .A4(n17527), .ZN(n17643) );
  INV_X1 U20758 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17772) );
  INV_X1 U20759 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17769) );
  INV_X1 U20760 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17767) );
  NOR2_X1 U20761 ( .A1(n17769), .A2(n17767), .ZN(n17618) );
  NAND4_X1 U20762 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_13__SCAN_IN), .A4(P3_EAX_REG_12__SCAN_IN), .ZN(n17528)
         );
  INV_X1 U20763 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17736) );
  INV_X1 U20764 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17730) );
  INV_X1 U20765 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17728) );
  INV_X1 U20766 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17726) );
  NOR4_X1 U20767 ( .A1(n17736), .A2(n17730), .A3(n17728), .A4(n17726), .ZN(
        n17529) );
  NAND4_X1 U20768 ( .A1(n17574), .A2(P3_EAX_REG_21__SCAN_IN), .A3(
        P3_EAX_REG_20__SCAN_IN), .A4(n17529), .ZN(n17569) );
  NAND2_X1 U20769 ( .A1(n17612), .A2(n17568), .ZN(n17562) );
  NAND2_X1 U20770 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17539), .ZN(n17538) );
  NOR2_X1 U20771 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17538), .ZN(n17531) );
  INV_X1 U20772 ( .A(n17677), .ZN(n17647) );
  NAND2_X1 U20773 ( .A1(n17663), .A2(n17538), .ZN(n17537) );
  OAI21_X1 U20774 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17647), .A(n17537), .ZN(
        n17530) );
  AOI22_X1 U20775 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17531), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17530), .ZN(n17532) );
  OAI21_X1 U20776 ( .B1(n18539), .B2(n17580), .A(n17532), .ZN(P3_U2704) );
  INV_X1 U20777 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17751) );
  NAND2_X1 U20778 ( .A1(n17533), .A2(n17614), .ZN(n17589) );
  OAI22_X1 U20779 ( .A1(n17534), .A2(n17680), .B1(n21395), .B2(n17580), .ZN(
        n17535) );
  AOI21_X1 U20780 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17607), .A(n17535), .ZN(
        n17536) );
  OAI221_X1 U20781 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17538), .C1(n17751), 
        .C2(n17537), .A(n17536), .ZN(P3_U2705) );
  AOI22_X1 U20782 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17607), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17606), .ZN(n17541) );
  OAI211_X1 U20783 ( .C1(n17539), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17663), .B(
        n17538), .ZN(n17540) );
  OAI211_X1 U20784 ( .C1(n17542), .C2(n17680), .A(n17541), .B(n17540), .ZN(
        P3_U2706) );
  INV_X1 U20785 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18526) );
  AOI22_X1 U20786 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17607), .B1(n17665), .B2(
        n17543), .ZN(n17546) );
  OAI211_X1 U20787 ( .C1(n9914), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17663), .B(
        n17544), .ZN(n17545) );
  OAI211_X1 U20788 ( .C1(n17580), .C2(n18526), .A(n17546), .B(n17545), .ZN(
        P3_U2707) );
  AOI22_X1 U20789 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17607), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17606), .ZN(n17549) );
  AOI211_X1 U20790 ( .C1(n17745), .C2(n17552), .A(n9914), .B(n17614), .ZN(
        n17547) );
  INV_X1 U20791 ( .A(n17547), .ZN(n17548) );
  OAI211_X1 U20792 ( .C1(n17550), .C2(n17680), .A(n17549), .B(n17548), .ZN(
        P3_U2708) );
  INV_X1 U20793 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17555) );
  AOI22_X1 U20794 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17606), .B1(n17665), .B2(
        n17551), .ZN(n17554) );
  OAI211_X1 U20795 ( .C1(n17556), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17663), .B(
        n17552), .ZN(n17553) );
  OAI211_X1 U20796 ( .C1(n17589), .C2(n17555), .A(n17554), .B(n17553), .ZN(
        P3_U2709) );
  AOI22_X1 U20797 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17607), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17606), .ZN(n17559) );
  AOI211_X1 U20798 ( .C1(n17742), .C2(n17563), .A(n17556), .B(n17614), .ZN(
        n17557) );
  INV_X1 U20799 ( .A(n17557), .ZN(n17558) );
  OAI211_X1 U20800 ( .C1(n17560), .C2(n17680), .A(n17559), .B(n17558), .ZN(
        P3_U2710) );
  INV_X1 U20801 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17567) );
  AOI22_X1 U20802 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17606), .B1(n17665), .B2(
        n17561), .ZN(n17566) );
  OAI21_X1 U20803 ( .B1(n17740), .B2(n17614), .A(n17562), .ZN(n17564) );
  NAND2_X1 U20804 ( .A1(n17564), .A2(n17563), .ZN(n17565) );
  OAI211_X1 U20805 ( .C1(n17589), .C2(n17567), .A(n17566), .B(n17565), .ZN(
        P3_U2711) );
  AOI211_X1 U20806 ( .C1(n17738), .C2(n17569), .A(n17614), .B(n17568), .ZN(
        n17570) );
  AOI21_X1 U20807 ( .B1(n17606), .B2(BUF2_REG_23__SCAN_IN), .A(n17570), .ZN(
        n17572) );
  NAND2_X1 U20808 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17607), .ZN(n17571) );
  OAI211_X1 U20809 ( .C1(n17573), .C2(n17680), .A(n17572), .B(n17571), .ZN(
        P3_U2712) );
  NAND2_X1 U20810 ( .A1(n17612), .A2(n17574), .ZN(n17599) );
  NAND2_X1 U20811 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17600), .ZN(n17595) );
  NAND3_X1 U20812 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(n17590), .ZN(n17579) );
  AOI22_X1 U20813 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17606), .B1(n17665), .B2(
        n17575), .ZN(n17578) );
  NAND2_X1 U20814 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17590), .ZN(n17586) );
  NAND2_X1 U20815 ( .A1(n17663), .A2(n17586), .ZN(n17584) );
  OAI21_X1 U20816 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17647), .A(n17584), .ZN(
        n17576) );
  AOI22_X1 U20817 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17607), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17576), .ZN(n17577) );
  OAI211_X1 U20818 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17579), .A(n17578), .B(
        n17577), .ZN(P3_U2713) );
  INV_X1 U20819 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17734) );
  OAI22_X1 U20820 ( .A1(n17581), .A2(n17680), .B1(n15357), .B2(n17580), .ZN(
        n17582) );
  AOI21_X1 U20821 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17607), .A(n17582), .ZN(
        n17583) );
  OAI221_X1 U20822 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17586), .C1(n17734), 
        .C2(n17584), .A(n17583), .ZN(P3_U2714) );
  INV_X1 U20823 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18527) );
  AOI22_X1 U20824 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17606), .B1(n17665), .B2(
        n17585), .ZN(n17588) );
  OAI211_X1 U20825 ( .C1(n17590), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17663), .B(
        n17586), .ZN(n17587) );
  OAI211_X1 U20826 ( .C1(n17589), .C2(n18527), .A(n17588), .B(n17587), .ZN(
        P3_U2715) );
  AOI22_X1 U20827 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17607), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17606), .ZN(n17593) );
  AOI211_X1 U20828 ( .C1(n17730), .C2(n17595), .A(n17590), .B(n17614), .ZN(
        n17591) );
  INV_X1 U20829 ( .A(n17591), .ZN(n17592) );
  OAI211_X1 U20830 ( .C1(n17594), .C2(n17680), .A(n17593), .B(n17592), .ZN(
        P3_U2716) );
  AOI22_X1 U20831 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17607), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17606), .ZN(n17597) );
  OAI211_X1 U20832 ( .C1(n17600), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17663), .B(
        n17595), .ZN(n17596) );
  OAI211_X1 U20833 ( .C1(n17598), .C2(n17680), .A(n17597), .B(n17596), .ZN(
        P3_U2717) );
  AOI22_X1 U20834 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17607), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17606), .ZN(n17604) );
  OAI21_X1 U20835 ( .B1(n17726), .B2(n17614), .A(n17599), .ZN(n17602) );
  INV_X1 U20836 ( .A(n17600), .ZN(n17601) );
  NAND2_X1 U20837 ( .A1(n17602), .A2(n17601), .ZN(n17603) );
  OAI211_X1 U20838 ( .C1(n17605), .C2(n17680), .A(n17604), .B(n17603), .ZN(
        P3_U2718) );
  AOI22_X1 U20839 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17607), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17606), .ZN(n17610) );
  OAI211_X1 U20840 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n9921), .A(n17663), .B(
        n17608), .ZN(n17609) );
  OAI211_X1 U20841 ( .C1(n17611), .C2(n17680), .A(n17610), .B(n17609), .ZN(
        P3_U2719) );
  NAND2_X1 U20842 ( .A1(n17612), .A2(n17613), .ZN(n17617) );
  INV_X1 U20843 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17785) );
  OR2_X1 U20844 ( .A1(n17614), .A2(n17613), .ZN(n17621) );
  AOI22_X1 U20845 ( .A1(n17665), .A2(n17615), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n17675), .ZN(n17616) );
  OAI221_X1 U20846 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17617), .C1(n17785), 
        .C2(n17621), .A(n17616), .ZN(P3_U2720) );
  NOR2_X1 U20847 ( .A1(n18545), .A2(n17643), .ZN(n17651) );
  NAND2_X1 U20848 ( .A1(n17618), .A2(n17651), .ZN(n17637) );
  INV_X1 U20849 ( .A(n17637), .ZN(n17641) );
  NAND2_X1 U20850 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17641), .ZN(n17634) );
  NOR2_X1 U20851 ( .A1(n17772), .A2(n17634), .ZN(n17627) );
  NAND2_X1 U20852 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17630), .ZN(n17622) );
  INV_X1 U20853 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17780) );
  AOI22_X1 U20854 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17675), .B1(n17665), .B2(
        n17619), .ZN(n17620) );
  OAI221_X1 U20855 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17622), .C1(n17780), 
        .C2(n17621), .A(n17620), .ZN(P3_U2721) );
  INV_X1 U20856 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17626) );
  INV_X1 U20857 ( .A(n17622), .ZN(n17625) );
  AOI21_X1 U20858 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17663), .A(n17630), .ZN(
        n17624) );
  OAI222_X1 U20859 ( .A1(n17673), .A2(n17626), .B1(n17625), .B2(n17624), .C1(
        n17680), .C2(n17623), .ZN(P3_U2722) );
  INV_X1 U20860 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17631) );
  AOI21_X1 U20861 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17663), .A(n17627), .ZN(
        n17629) );
  OAI222_X1 U20862 ( .A1(n17673), .A2(n17631), .B1(n17630), .B2(n17629), .C1(
        n17680), .C2(n17628), .ZN(P3_U2723) );
  NAND2_X1 U20863 ( .A1(n17663), .A2(n17634), .ZN(n17638) );
  AOI22_X1 U20864 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17675), .B1(n17665), .B2(
        n17632), .ZN(n17633) );
  OAI221_X1 U20865 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17634), .C1(n17772), 
        .C2(n17638), .A(n17633), .ZN(P3_U2724) );
  INV_X1 U20866 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n21523) );
  AOI22_X1 U20867 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17675), .B1(n17665), .B2(
        n17635), .ZN(n17636) );
  OAI221_X1 U20868 ( .B1(n17638), .B2(n21523), .C1(n17638), .C2(n17637), .A(
        n17636), .ZN(P3_U2725) );
  INV_X1 U20869 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17642) );
  AOI22_X1 U20870 ( .A1(n17651), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17663), .ZN(n17640) );
  OAI222_X1 U20871 ( .A1(n17673), .A2(n17642), .B1(n17641), .B2(n17640), .C1(
        n17680), .C2(n17639), .ZN(P3_U2726) );
  AOI22_X1 U20872 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17675), .B1(n17651), .B2(
        n17767), .ZN(n17645) );
  NAND3_X1 U20873 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17663), .A3(n17643), .ZN(
        n17644) );
  OAI211_X1 U20874 ( .C1(n17646), .C2(n17680), .A(n17645), .B(n17644), .ZN(
        P3_U2727) );
  INV_X1 U20875 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18542) );
  NAND2_X1 U20876 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n17648) );
  NOR3_X1 U20877 ( .A1(n17676), .A2(n17756), .A3(n17647), .ZN(n17658) );
  INV_X1 U20878 ( .A(n17658), .ZN(n17667) );
  NOR3_X1 U20879 ( .A1(n21531), .A2(n17758), .A3(n17667), .ZN(n17662) );
  INV_X1 U20880 ( .A(n17662), .ZN(n17654) );
  NOR2_X1 U20881 ( .A1(n17648), .A2(n17654), .ZN(n17653) );
  AOI21_X1 U20882 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17663), .A(n17653), .ZN(
        n17650) );
  OAI222_X1 U20883 ( .A1(n17673), .A2(n18542), .B1(n17651), .B2(n17650), .C1(
        n17680), .C2(n17649), .ZN(P3_U2728) );
  INV_X1 U20884 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18536) );
  AOI22_X1 U20885 ( .A1(n17662), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17663), .ZN(n17652) );
  INV_X1 U20886 ( .A(n18089), .ZN(n18090) );
  OAI222_X1 U20887 ( .A1(n18536), .A2(n17673), .B1(n17653), .B2(n17652), .C1(
        n17680), .C2(n18090), .ZN(P3_U2729) );
  INV_X1 U20888 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18532) );
  INV_X1 U20889 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17761) );
  NOR2_X1 U20890 ( .A1(n17761), .A2(n17654), .ZN(n17657) );
  AOI21_X1 U20891 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17663), .A(n17662), .ZN(
        n17656) );
  OAI222_X1 U20892 ( .A1(n18532), .A2(n17673), .B1(n17657), .B2(n17656), .C1(
        n17680), .C2(n17655), .ZN(P3_U2730) );
  AOI22_X1 U20893 ( .A1(n17658), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n17663), .ZN(n17661) );
  INV_X1 U20894 ( .A(n17659), .ZN(n17660) );
  OAI222_X1 U20895 ( .A1(n18527), .A2(n17673), .B1(n17662), .B2(n17661), .C1(
        n17680), .C2(n17660), .ZN(P3_U2731) );
  NAND2_X1 U20896 ( .A1(n17663), .A2(n17667), .ZN(n17671) );
  AOI22_X1 U20897 ( .A1(n17675), .A2(BUF2_REG_3__SCAN_IN), .B1(n17665), .B2(
        n17664), .ZN(n17666) );
  OAI221_X1 U20898 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17667), .C1(n17758), 
        .C2(n17671), .A(n17666), .ZN(P3_U2732) );
  INV_X1 U20899 ( .A(n17668), .ZN(n17672) );
  NOR2_X1 U20900 ( .A1(n17669), .A2(P3_EAX_REG_2__SCAN_IN), .ZN(n17670) );
  OAI222_X1 U20901 ( .A1(n17673), .A2(n18517), .B1(n17680), .B2(n17672), .C1(
        n17671), .C2(n17670), .ZN(P3_U2733) );
  AOI22_X1 U20902 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17675), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n17674), .ZN(n17679) );
  OAI211_X1 U20903 ( .C1(P3_EAX_REG_0__SCAN_IN), .C2(P3_EAX_REG_1__SCAN_IN), 
        .A(n17677), .B(n17676), .ZN(n17678) );
  OAI211_X1 U20904 ( .C1(n17681), .C2(n17680), .A(n17679), .B(n17678), .ZN(
        P3_U2734) );
  OR2_X1 U20905 ( .A1(n19109), .A2(n18165), .ZN(n19145) );
  INV_X2 U20906 ( .A(n19145), .ZN(n18997) );
  AND2_X1 U20907 ( .A1(n17698), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20908 ( .A1(n17701), .A2(n17683), .ZN(n17700) );
  AOI22_X1 U20909 ( .A1(n18997), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17717), .ZN(n17684) );
  OAI21_X1 U20910 ( .B1(n17751), .B2(n17700), .A(n17684), .ZN(P3_U2737) );
  INV_X1 U20911 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U20912 ( .A1(n18997), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17685) );
  OAI21_X1 U20913 ( .B1(n17749), .B2(n17700), .A(n17685), .ZN(P3_U2738) );
  INV_X1 U20914 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U20915 ( .A1(n18997), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17686) );
  OAI21_X1 U20916 ( .B1(n17747), .B2(n17700), .A(n17686), .ZN(P3_U2739) );
  AOI22_X1 U20917 ( .A1(n18997), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17687) );
  OAI21_X1 U20918 ( .B1(n17745), .B2(n17700), .A(n17687), .ZN(P3_U2740) );
  AOI22_X1 U20919 ( .A1(n18997), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17688) );
  OAI21_X1 U20920 ( .B1(n10034), .B2(n17700), .A(n17688), .ZN(P3_U2741) );
  AOI22_X1 U20921 ( .A1(n18997), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17689) );
  OAI21_X1 U20922 ( .B1(n17742), .B2(n17700), .A(n17689), .ZN(P3_U2742) );
  AOI22_X1 U20923 ( .A1(n18997), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17690) );
  OAI21_X1 U20924 ( .B1(n17740), .B2(n17700), .A(n17690), .ZN(P3_U2743) );
  AOI22_X1 U20925 ( .A1(n18997), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17691) );
  OAI21_X1 U20926 ( .B1(n17738), .B2(n17700), .A(n17691), .ZN(P3_U2744) );
  AOI22_X1 U20927 ( .A1(n18997), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17692) );
  OAI21_X1 U20928 ( .B1(n17736), .B2(n17700), .A(n17692), .ZN(P3_U2745) );
  AOI22_X1 U20929 ( .A1(n18997), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17693) );
  OAI21_X1 U20930 ( .B1(n17734), .B2(n17700), .A(n17693), .ZN(P3_U2746) );
  INV_X1 U20931 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17732) );
  AOI22_X1 U20932 ( .A1(n18997), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17694) );
  OAI21_X1 U20933 ( .B1(n17732), .B2(n17700), .A(n17694), .ZN(P3_U2747) );
  AOI22_X1 U20934 ( .A1(n18997), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17695) );
  OAI21_X1 U20935 ( .B1(n17730), .B2(n17700), .A(n17695), .ZN(P3_U2748) );
  AOI22_X1 U20936 ( .A1(n18997), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17696) );
  OAI21_X1 U20937 ( .B1(n17728), .B2(n17700), .A(n17696), .ZN(P3_U2749) );
  AOI22_X1 U20938 ( .A1(n18997), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17697) );
  OAI21_X1 U20939 ( .B1(n17726), .B2(n17700), .A(n17697), .ZN(P3_U2750) );
  INV_X1 U20940 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17724) );
  AOI22_X1 U20941 ( .A1(n18997), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17698), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17699) );
  OAI21_X1 U20942 ( .B1(n17724), .B2(n17700), .A(n17699), .ZN(P3_U2751) );
  AOI22_X1 U20943 ( .A1(n18997), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17702) );
  OAI21_X1 U20944 ( .B1(n17785), .B2(n17719), .A(n17702), .ZN(P3_U2752) );
  AOI22_X1 U20945 ( .A1(n18997), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17703) );
  OAI21_X1 U20946 ( .B1(n17780), .B2(n17719), .A(n17703), .ZN(P3_U2753) );
  INV_X1 U20947 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U20948 ( .A1(n18997), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17704) );
  OAI21_X1 U20949 ( .B1(n17778), .B2(n17719), .A(n17704), .ZN(P3_U2754) );
  INV_X1 U20950 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17775) );
  AOI22_X1 U20951 ( .A1(n18997), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17705) );
  OAI21_X1 U20952 ( .B1(n17775), .B2(n17719), .A(n17705), .ZN(P3_U2755) );
  AOI22_X1 U20953 ( .A1(n18997), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17706) );
  OAI21_X1 U20954 ( .B1(n17772), .B2(n17719), .A(n17706), .ZN(P3_U2756) );
  AOI22_X1 U20955 ( .A1(n18997), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17707) );
  OAI21_X1 U20956 ( .B1(n21523), .B2(n17719), .A(n17707), .ZN(P3_U2757) );
  AOI22_X1 U20957 ( .A1(n18997), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17708) );
  OAI21_X1 U20958 ( .B1(n17769), .B2(n17719), .A(n17708), .ZN(P3_U2758) );
  AOI22_X1 U20959 ( .A1(n18997), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17709) );
  OAI21_X1 U20960 ( .B1(n17767), .B2(n17719), .A(n17709), .ZN(P3_U2759) );
  AOI22_X1 U20961 ( .A1(n18997), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17710) );
  OAI21_X1 U20962 ( .B1(n17765), .B2(n17719), .A(n17710), .ZN(P3_U2760) );
  INV_X1 U20963 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17763) );
  AOI22_X1 U20964 ( .A1(n18997), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17711) );
  OAI21_X1 U20965 ( .B1(n17763), .B2(n17719), .A(n17711), .ZN(P3_U2761) );
  AOI22_X1 U20966 ( .A1(n18997), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17712) );
  OAI21_X1 U20967 ( .B1(n17761), .B2(n17719), .A(n17712), .ZN(P3_U2762) );
  AOI22_X1 U20968 ( .A1(n18997), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17713) );
  OAI21_X1 U20969 ( .B1(n21531), .B2(n17719), .A(n17713), .ZN(P3_U2763) );
  AOI22_X1 U20970 ( .A1(n18997), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17714) );
  OAI21_X1 U20971 ( .B1(n17758), .B2(n17719), .A(n17714), .ZN(P3_U2764) );
  AOI22_X1 U20972 ( .A1(n18997), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17715) );
  OAI21_X1 U20973 ( .B1(n17756), .B2(n17719), .A(n17715), .ZN(P3_U2765) );
  INV_X1 U20974 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17754) );
  AOI22_X1 U20975 ( .A1(n18997), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17716) );
  OAI21_X1 U20976 ( .B1(n17754), .B2(n17719), .A(n17716), .ZN(P3_U2766) );
  AOI22_X1 U20977 ( .A1(n18997), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17717), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17718) );
  OAI21_X1 U20978 ( .B1(n21494), .B2(n17719), .A(n17718), .ZN(P3_U2767) );
  NAND2_X2 U20979 ( .A1(n19152), .A2(n17722), .ZN(n17784) );
  AOI22_X1 U20980 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17782), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17781), .ZN(n17723) );
  OAI21_X1 U20981 ( .B1(n17724), .B2(n17784), .A(n17723), .ZN(P3_U2768) );
  AOI22_X1 U20982 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17782), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17781), .ZN(n17725) );
  OAI21_X1 U20983 ( .B1(n17726), .B2(n17784), .A(n17725), .ZN(P3_U2769) );
  AOI22_X1 U20984 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17782), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17781), .ZN(n17727) );
  OAI21_X1 U20985 ( .B1(n17728), .B2(n17784), .A(n17727), .ZN(P3_U2770) );
  AOI22_X1 U20986 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17773), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17781), .ZN(n17729) );
  OAI21_X1 U20987 ( .B1(n17730), .B2(n17784), .A(n17729), .ZN(P3_U2771) );
  AOI22_X1 U20988 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17773), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17781), .ZN(n17731) );
  OAI21_X1 U20989 ( .B1(n17732), .B2(n17784), .A(n17731), .ZN(P3_U2772) );
  AOI22_X1 U20990 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17773), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17781), .ZN(n17733) );
  OAI21_X1 U20991 ( .B1(n17734), .B2(n17784), .A(n17733), .ZN(P3_U2773) );
  AOI22_X1 U20992 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17773), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17781), .ZN(n17735) );
  OAI21_X1 U20993 ( .B1(n17736), .B2(n17784), .A(n17735), .ZN(P3_U2774) );
  AOI22_X1 U20994 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17773), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17781), .ZN(n17737) );
  OAI21_X1 U20995 ( .B1(n17738), .B2(n17784), .A(n17737), .ZN(P3_U2775) );
  AOI22_X1 U20996 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17773), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17781), .ZN(n17739) );
  OAI21_X1 U20997 ( .B1(n17740), .B2(n17784), .A(n17739), .ZN(P3_U2776) );
  AOI22_X1 U20998 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17773), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17781), .ZN(n17741) );
  OAI21_X1 U20999 ( .B1(n17742), .B2(n17784), .A(n17741), .ZN(P3_U2777) );
  AOI22_X1 U21000 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17773), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17781), .ZN(n17743) );
  OAI21_X1 U21001 ( .B1(n10034), .B2(n17784), .A(n17743), .ZN(P3_U2778) );
  AOI22_X1 U21002 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17773), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17781), .ZN(n17744) );
  OAI21_X1 U21003 ( .B1(n17745), .B2(n17784), .A(n17744), .ZN(P3_U2779) );
  AOI22_X1 U21004 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17782), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17781), .ZN(n17746) );
  OAI21_X1 U21005 ( .B1(n17747), .B2(n17784), .A(n17746), .ZN(P3_U2780) );
  AOI22_X1 U21006 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17782), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17781), .ZN(n17748) );
  OAI21_X1 U21007 ( .B1(n17749), .B2(n17784), .A(n17748), .ZN(P3_U2781) );
  AOI22_X1 U21008 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17782), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17781), .ZN(n17750) );
  OAI21_X1 U21009 ( .B1(n17751), .B2(n17784), .A(n17750), .ZN(P3_U2782) );
  AOI22_X1 U21010 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17781), .ZN(n17752) );
  OAI21_X1 U21011 ( .B1(n21494), .B2(n17784), .A(n17752), .ZN(P3_U2783) );
  AOI22_X1 U21012 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17781), .ZN(n17753) );
  OAI21_X1 U21013 ( .B1(n17754), .B2(n17784), .A(n17753), .ZN(P3_U2784) );
  AOI22_X1 U21014 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17781), .ZN(n17755) );
  OAI21_X1 U21015 ( .B1(n17756), .B2(n17784), .A(n17755), .ZN(P3_U2785) );
  AOI22_X1 U21016 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17781), .ZN(n17757) );
  OAI21_X1 U21017 ( .B1(n17758), .B2(n17784), .A(n17757), .ZN(P3_U2786) );
  AOI22_X1 U21018 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17776), .ZN(n17759) );
  OAI21_X1 U21019 ( .B1(n21531), .B2(n17784), .A(n17759), .ZN(P3_U2787) );
  AOI22_X1 U21020 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17776), .ZN(n17760) );
  OAI21_X1 U21021 ( .B1(n17761), .B2(n17784), .A(n17760), .ZN(P3_U2788) );
  AOI22_X1 U21022 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17776), .ZN(n17762) );
  OAI21_X1 U21023 ( .B1(n17763), .B2(n17784), .A(n17762), .ZN(P3_U2789) );
  AOI22_X1 U21024 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17776), .ZN(n17764) );
  OAI21_X1 U21025 ( .B1(n17765), .B2(n17784), .A(n17764), .ZN(P3_U2790) );
  AOI22_X1 U21026 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17776), .ZN(n17766) );
  OAI21_X1 U21027 ( .B1(n17767), .B2(n17784), .A(n17766), .ZN(P3_U2791) );
  AOI22_X1 U21028 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17776), .ZN(n17768) );
  OAI21_X1 U21029 ( .B1(n17769), .B2(n17784), .A(n17768), .ZN(P3_U2792) );
  AOI22_X1 U21030 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17773), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17776), .ZN(n17770) );
  OAI21_X1 U21031 ( .B1(n21523), .B2(n17784), .A(n17770), .ZN(P3_U2793) );
  AOI22_X1 U21032 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17776), .ZN(n17771) );
  OAI21_X1 U21033 ( .B1(n17772), .B2(n17784), .A(n17771), .ZN(P3_U2794) );
  AOI22_X1 U21034 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17773), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17776), .ZN(n17774) );
  OAI21_X1 U21035 ( .B1(n17775), .B2(n17784), .A(n17774), .ZN(P3_U2795) );
  AOI22_X1 U21036 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17776), .ZN(n17777) );
  OAI21_X1 U21037 ( .B1(n17778), .B2(n17784), .A(n17777), .ZN(P3_U2796) );
  AOI22_X1 U21038 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17781), .ZN(n17779) );
  OAI21_X1 U21039 ( .B1(n17780), .B2(n17784), .A(n17779), .ZN(P3_U2797) );
  AOI22_X1 U21040 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17782), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17781), .ZN(n17783) );
  OAI21_X1 U21041 ( .B1(n17785), .B2(n17784), .A(n17783), .ZN(P3_U2798) );
  AOI21_X1 U21042 ( .B1(n17786), .B2(n19013), .A(n18117), .ZN(n17787) );
  INV_X1 U21043 ( .A(n17787), .ZN(n17788) );
  AOI21_X1 U21044 ( .B1(n17986), .B2(n17789), .A(n17788), .ZN(n17825) );
  OAI21_X1 U21045 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17898), .A(
        n17825), .ZN(n17811) );
  AOI22_X1 U21046 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17811), .B1(
        n18006), .B2(n17790), .ZN(n17805) );
  NOR2_X1 U21047 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18170), .ZN(
        n17799) );
  NOR2_X1 U21048 ( .A1(n18070), .A2(n18157), .ZN(n17904) );
  OAI22_X1 U21049 ( .A1(n17791), .A2(n18025), .B1(n18177), .B2(n13159), .ZN(
        n17827) );
  NOR2_X1 U21050 ( .A1(n18170), .A2(n17827), .ZN(n17793) );
  NOR3_X1 U21051 ( .A1(n17904), .A2(n17793), .A3(n17792), .ZN(n17798) );
  AOI211_X1 U21052 ( .C1(n17796), .C2(n17795), .A(n17794), .B(n18057), .ZN(
        n17797) );
  AOI211_X1 U21053 ( .C1(n17799), .C2(n17814), .A(n17798), .B(n17797), .ZN(
        n17804) );
  NAND3_X1 U21054 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17800) );
  NAND2_X1 U21055 ( .A1(n17832), .A2(n17988), .ZN(n17847) );
  NOR2_X1 U21056 ( .A1(n17800), .A2(n17847), .ZN(n17813) );
  OAI211_X1 U21057 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17813), .B(n17801), .ZN(n17802) );
  NAND4_X1 U21058 ( .A1(n17805), .A2(n17804), .A3(n17803), .A4(n17802), .ZN(
        P3_U2802) );
  NAND2_X1 U21059 ( .A1(n17807), .A2(n17806), .ZN(n17808) );
  XOR2_X1 U21060 ( .A(n17808), .B(n18030), .Z(n18184) );
  OAI22_X1 U21061 ( .A1(n18484), .A2(n19081), .B1(n17944), .B2(n17809), .ZN(
        n17810) );
  AOI221_X1 U21062 ( .B1(n17813), .B2(n17812), .C1(n17811), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17810), .ZN(n17816) );
  AOI22_X1 U21063 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17827), .B1(
        n17814), .B2(n18170), .ZN(n17815) );
  OAI211_X1 U21064 ( .C1(n18184), .C2(n18057), .A(n17816), .B(n17815), .ZN(
        P3_U2803) );
  AOI21_X1 U21065 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17818), .A(
        n17817), .ZN(n18192) );
  NOR2_X1 U21066 ( .A1(n17931), .A2(n18187), .ZN(n17828) );
  NOR2_X1 U21067 ( .A1(n17819), .A2(n18540), .ZN(n17862) );
  AOI21_X1 U21068 ( .B1(n17820), .B2(n17862), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17824) );
  INV_X1 U21069 ( .A(n17898), .ZN(n17822) );
  OAI21_X1 U21070 ( .B1(n18006), .B2(n17822), .A(n17821), .ZN(n17823) );
  NAND2_X1 U21071 ( .A1(n18479), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18191) );
  OAI211_X1 U21072 ( .C1(n17825), .C2(n17824), .A(n17823), .B(n18191), .ZN(
        n17826) );
  AOI221_X1 U21073 ( .B1(n17828), .B2(n18186), .C1(n17827), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17826), .ZN(n17829) );
  OAI21_X1 U21074 ( .B1(n18192), .B2(n18057), .A(n17829), .ZN(P3_U2804) );
  OR2_X1 U21075 ( .A1(n18305), .A2(n17853), .ZN(n18210) );
  OAI21_X1 U21076 ( .B1(n17856), .B2(n18210), .A(n21488), .ZN(n17830) );
  OAI21_X1 U21077 ( .B1(n18187), .B2(n18305), .A(n17830), .ZN(n18205) );
  OAI22_X1 U21078 ( .A1(n17832), .A2(n18540), .B1(n17831), .B2(n18165), .ZN(
        n17833) );
  NOR2_X1 U21079 ( .A1(n18117), .A2(n17833), .ZN(n17866) );
  OAI21_X1 U21080 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17898), .A(
        n17866), .ZN(n17850) );
  NOR2_X1 U21081 ( .A1(n18484), .A2(n19078), .ZN(n18200) );
  OAI21_X1 U21082 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17834), .ZN(n17835) );
  OAI22_X1 U21083 ( .A1(n17944), .A2(n17836), .B1(n17847), .B2(n17835), .ZN(
        n17837) );
  AOI211_X1 U21084 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17850), .A(
        n18200), .B(n17837), .ZN(n17843) );
  NAND3_X1 U21085 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17964), .A3(
        n18196), .ZN(n17838) );
  XOR2_X1 U21086 ( .A(n17838), .B(n21488), .Z(n18202) );
  OAI21_X1 U21087 ( .B1(n18030), .B2(n17840), .A(n17839), .ZN(n17841) );
  XOR2_X1 U21088 ( .A(n17841), .B(n21488), .Z(n18201) );
  AOI22_X1 U21089 ( .A1(n18157), .A2(n18202), .B1(n18069), .B2(n18201), .ZN(
        n17842) );
  OAI211_X1 U21090 ( .C1(n18025), .C2(n18205), .A(n17843), .B(n17842), .ZN(
        P3_U2805) );
  NOR2_X1 U21091 ( .A1(n17853), .A2(n18306), .ZN(n18212) );
  INV_X1 U21092 ( .A(n18212), .ZN(n17844) );
  AOI22_X1 U21093 ( .A1(n18070), .A2(n18210), .B1(n18157), .B2(n17844), .ZN(
        n17870) );
  NAND2_X1 U21094 ( .A1(n18479), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18218) );
  INV_X1 U21095 ( .A(n18218), .ZN(n17849) );
  INV_X1 U21096 ( .A(n17845), .ZN(n17846) );
  OAI22_X1 U21097 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17847), .B1(
        n17846), .B2(n17944), .ZN(n17848) );
  AOI211_X1 U21098 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17850), .A(
        n17849), .B(n17848), .ZN(n17855) );
  OAI21_X1 U21099 ( .B1(n17852), .B2(n17856), .A(n17851), .ZN(n18208) );
  NOR2_X1 U21100 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17853), .ZN(
        n18206) );
  AOI22_X1 U21101 ( .A1(n18069), .A2(n18208), .B1(n18206), .B2(n17951), .ZN(
        n17854) );
  OAI211_X1 U21102 ( .C1(n17870), .C2(n17856), .A(n17855), .B(n17854), .ZN(
        P3_U2806) );
  AOI21_X1 U21103 ( .B1(n17858), .B2(n17928), .A(n17880), .ZN(n17859) );
  AOI211_X1 U21104 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18030), .A(
        n17859), .B(n17896), .ZN(n17860) );
  XOR2_X1 U21105 ( .A(n17860), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n18220) );
  NOR4_X1 U21106 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17931), .A3(
        n17861), .A4(n18245), .ZN(n17868) );
  NOR2_X1 U21107 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17862), .ZN(
        n17865) );
  OAI21_X1 U21108 ( .B1(n18006), .B2(n17822), .A(n17863), .ZN(n17864) );
  NAND2_X1 U21109 ( .A1(n18479), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18225) );
  OAI211_X1 U21110 ( .C1(n17866), .C2(n17865), .A(n17864), .B(n18225), .ZN(
        n17867) );
  AOI211_X1 U21111 ( .C1(n18069), .C2(n18220), .A(n17868), .B(n17867), .ZN(
        n17869) );
  OAI21_X1 U21112 ( .B1(n17870), .B2(n18213), .A(n17869), .ZN(P3_U2807) );
  OAI22_X1 U21113 ( .A1(n17874), .A2(n17984), .B1(n17871), .B2(n18165), .ZN(
        n17872) );
  NOR2_X1 U21114 ( .A1(n18117), .A2(n17872), .ZN(n17899) );
  OAI21_X1 U21115 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17898), .A(
        n17899), .ZN(n17892) );
  AOI22_X1 U21116 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17892), .B1(
        n18006), .B2(n17873), .ZN(n17885) );
  NAND2_X1 U21117 ( .A1(n17874), .A2(n17988), .ZN(n17890) );
  AOI21_X1 U21118 ( .B1(n17876), .B2(n17875), .A(n17890), .ZN(n17878) );
  AOI22_X1 U21119 ( .A1(n18479), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17878), 
        .B2(n17877), .ZN(n17884) );
  INV_X1 U21120 ( .A(n18171), .ZN(n18232) );
  NOR2_X1 U21121 ( .A1(n18232), .A2(n18245), .ZN(n18237) );
  AOI22_X1 U21122 ( .A1(n18070), .A2(n18305), .B1(n18157), .B2(n18306), .ZN(
        n17954) );
  OAI21_X1 U21123 ( .B1(n17904), .B2(n18237), .A(n17954), .ZN(n17893) );
  OAI221_X1 U21124 ( .B1(n17880), .B2(n17949), .C1(n17880), .C2(n18237), .A(
        n17879), .ZN(n17881) );
  XOR2_X1 U21125 ( .A(n18244), .B(n17881), .Z(n18240) );
  AOI22_X1 U21126 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17893), .B1(
        n18069), .B2(n18240), .ZN(n17883) );
  NAND3_X1 U21127 ( .A1(n18171), .A2(n17916), .A3(n18244), .ZN(n17882) );
  NAND4_X1 U21128 ( .A1(n17885), .A2(n17884), .A3(n17883), .A4(n17882), .ZN(
        P3_U2808) );
  OAI22_X1 U21129 ( .A1(n18250), .A2(n17907), .B1(n17887), .B2(n17928), .ZN(
        n17888) );
  XOR2_X1 U21130 ( .A(n21522), .B(n17888), .Z(n18256) );
  NOR2_X1 U21131 ( .A1(n18484), .A2(n19071), .ZN(n18252) );
  OAI22_X1 U21132 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17890), .B1(
        n10175), .B2(n17944), .ZN(n17891) );
  AOI211_X1 U21133 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17892), .A(
        n18252), .B(n17891), .ZN(n17895) );
  NOR2_X1 U21134 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18250), .ZN(
        n18254) );
  AOI22_X1 U21135 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17893), .B1(
        n18254), .B2(n17916), .ZN(n17894) );
  OAI211_X1 U21136 ( .C1(n18256), .C2(n18057), .A(n17895), .B(n17894), .ZN(
        P3_U2809) );
  INV_X1 U21137 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18266) );
  AOI221_X1 U21138 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17907), 
        .C1(n18266), .C2(n17925), .A(n17896), .ZN(n17897) );
  XOR2_X1 U21139 ( .A(n18228), .B(n17897), .Z(n18265) );
  NAND2_X1 U21140 ( .A1(n17944), .A2(n17898), .ZN(n18158) );
  AOI221_X1 U21141 ( .B1(n17901), .B2(n17900), .C1(n18540), .C2(n17900), .A(
        n17899), .ZN(n17902) );
  NOR2_X1 U21142 ( .A1(n18484), .A2(n19068), .ZN(n18257) );
  AOI211_X1 U21143 ( .C1(n17903), .C2(n18158), .A(n17902), .B(n18257), .ZN(
        n17906) );
  NOR2_X1 U21144 ( .A1(n18266), .A2(n18245), .ZN(n18233) );
  OAI21_X1 U21145 ( .B1(n17904), .B2(n18233), .A(n17954), .ZN(n17915) );
  NOR2_X1 U21146 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18266), .ZN(
        n18258) );
  AOI22_X1 U21147 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17915), .B1(
        n17916), .B2(n18258), .ZN(n17905) );
  OAI211_X1 U21148 ( .C1(n18057), .C2(n18265), .A(n17906), .B(n17905), .ZN(
        P3_U2810) );
  OAI21_X1 U21149 ( .B1(n17928), .B2(n17925), .A(n17907), .ZN(n17908) );
  XOR2_X1 U21150 ( .A(n17908), .B(n18266), .Z(n18271) );
  NOR2_X1 U21151 ( .A1(n10181), .A2(n10182), .ZN(n17913) );
  OAI211_X1 U21152 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17918), .B(n17988), .ZN(n17912) );
  AOI21_X1 U21153 ( .B1(n19013), .B2(n10183), .A(n18117), .ZN(n17934) );
  OAI21_X1 U21154 ( .B1(n17909), .B2(n18165), .A(n17934), .ZN(n17923) );
  AOI22_X1 U21155 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17923), .B1(
        n18006), .B2(n17910), .ZN(n17911) );
  NAND2_X1 U21156 ( .A1(n18479), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18269) );
  OAI211_X1 U21157 ( .C1(n17913), .C2(n17912), .A(n17911), .B(n18269), .ZN(
        n17914) );
  AOI221_X1 U21158 ( .B1(n17916), .B2(n18266), .C1(n17915), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17914), .ZN(n17917) );
  OAI21_X1 U21159 ( .B1(n18271), .B2(n18057), .A(n17917), .ZN(P3_U2811) );
  NAND2_X1 U21160 ( .A1(n17924), .A2(n17926), .ZN(n18285) );
  NAND2_X1 U21161 ( .A1(n18479), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18283) );
  INV_X1 U21162 ( .A(n18283), .ZN(n17922) );
  NAND2_X1 U21163 ( .A1(n17918), .A2(n17988), .ZN(n17920) );
  OAI22_X1 U21164 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17920), .B1(
        n17919), .B2(n17944), .ZN(n17921) );
  AOI211_X1 U21165 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17923), .A(
        n17922), .B(n17921), .ZN(n17930) );
  OAI21_X1 U21166 ( .B1(n17924), .B2(n17931), .A(n17954), .ZN(n17938) );
  OAI21_X1 U21167 ( .B1(n18030), .B2(n17926), .A(n17925), .ZN(n17927) );
  XOR2_X1 U21168 ( .A(n17928), .B(n17927), .Z(n18281) );
  AOI22_X1 U21169 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17938), .B1(
        n18069), .B2(n18281), .ZN(n17929) );
  OAI211_X1 U21170 ( .C1(n17931), .C2(n18285), .A(n17930), .B(n17929), .ZN(
        P3_U2812) );
  AOI21_X1 U21171 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17933), .A(
        n17932), .ZN(n18291) );
  AOI221_X1 U21172 ( .B1(n17935), .B2(n21440), .C1(n18540), .C2(n21440), .A(
        n17934), .ZN(n17936) );
  NOR2_X1 U21173 ( .A1(n18484), .A2(n19064), .ZN(n18288) );
  AOI211_X1 U21174 ( .C1(n17937), .C2(n18158), .A(n17936), .B(n18288), .ZN(
        n17940) );
  OAI221_X1 U21175 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17951), .A(n17938), .ZN(
        n17939) );
  OAI211_X1 U21176 ( .C1(n18291), .C2(n18057), .A(n17940), .B(n17939), .ZN(
        P3_U2813) );
  NAND2_X1 U21177 ( .A1(n17941), .A2(n17988), .ZN(n17958) );
  AOI221_X1 U21178 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n17957), .C2(n17945), .A(
        n17958), .ZN(n17947) );
  OAI21_X1 U21179 ( .B1(n17941), .B2(n17984), .A(n18164), .ZN(n17978) );
  AOI21_X1 U21180 ( .B1(n17986), .B2(n17942), .A(n17978), .ZN(n17956) );
  OAI22_X1 U21181 ( .A1(n17956), .A2(n17945), .B1(n17944), .B2(n17943), .ZN(
        n17946) );
  AOI211_X1 U21182 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n18479), .A(n17947), 
        .B(n17946), .ZN(n17953) );
  OAI21_X1 U21183 ( .B1(n18030), .B2(n17949), .A(n17948), .ZN(n17950) );
  XOR2_X1 U21184 ( .A(n17950), .B(n18303), .Z(n18300) );
  AOI22_X1 U21185 ( .A1(n18300), .A2(n18069), .B1(n18303), .B2(n17951), .ZN(
        n17952) );
  OAI211_X1 U21186 ( .C1(n17954), .C2(n18303), .A(n17953), .B(n17952), .ZN(
        P3_U2814) );
  NOR2_X1 U21187 ( .A1(n18327), .A2(n17955), .ZN(n18298) );
  AOI21_X1 U21188 ( .B1(n18024), .B2(n18298), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18310) );
  NAND2_X1 U21189 ( .A1(n18070), .A2(n18305), .ZN(n17969) );
  NAND2_X1 U21190 ( .A1(n18479), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18315) );
  OAI221_X1 U21191 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17958), .C1(
        n17957), .C2(n17956), .A(n18315), .ZN(n17959) );
  AOI21_X1 U21192 ( .B1(n18006), .B2(n17960), .A(n17959), .ZN(n17968) );
  NAND4_X1 U21193 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18068), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(n17961), .ZN(n18044) );
  NOR2_X1 U21194 ( .A1(n17962), .A2(n18044), .ZN(n17970) );
  NAND2_X1 U21195 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18343), .ZN(
        n18350) );
  OAI221_X1 U21196 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17971), 
        .C1(n18327), .C2(n17970), .A(n18350), .ZN(n17963) );
  XOR2_X1 U21197 ( .A(n18296), .B(n17963), .Z(n18314) );
  NOR2_X1 U21198 ( .A1(n17964), .A2(n13159), .ZN(n17966) );
  INV_X1 U21199 ( .A(n17995), .ZN(n18338) );
  NOR3_X1 U21200 ( .A1(n18343), .A2(n18327), .A3(n18338), .ZN(n17980) );
  NOR2_X1 U21201 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17980), .ZN(
        n18308) );
  INV_X1 U21202 ( .A(n18308), .ZN(n17965) );
  AOI22_X1 U21203 ( .A1(n18069), .A2(n18314), .B1(n17966), .B2(n17965), .ZN(
        n17967) );
  OAI211_X1 U21204 ( .C1(n18310), .C2(n17969), .A(n17968), .B(n17967), .ZN(
        P3_U2815) );
  OAI21_X1 U21205 ( .B1(n17971), .B2(n17970), .A(n18350), .ZN(n17972) );
  XOR2_X1 U21206 ( .A(n17972), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18334) );
  OAI21_X1 U21207 ( .B1(n17974), .B2(n18540), .A(n17973), .ZN(n17977) );
  OAI22_X1 U21208 ( .A1(n18150), .A2(n17975), .B1(n18484), .B2(n19059), .ZN(
        n17976) );
  AOI21_X1 U21209 ( .B1(n17978), .B2(n17977), .A(n17976), .ZN(n17983) );
  AOI22_X1 U21210 ( .A1(n18024), .A2(n18298), .B1(n17979), .B2(n18327), .ZN(
        n18331) );
  NAND2_X1 U21211 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17995), .ZN(
        n17981) );
  AOI21_X1 U21212 ( .B1(n18327), .B2(n17981), .A(n17980), .ZN(n18330) );
  AOI22_X1 U21213 ( .A1(n18070), .A2(n18331), .B1(n18157), .B2(n18330), .ZN(
        n17982) );
  OAI211_X1 U21214 ( .C1(n18057), .C2(n18334), .A(n17983), .B(n17982), .ZN(
        P3_U2816) );
  OAI22_X1 U21215 ( .A1(n18362), .A2(n13159), .B1(n18025), .B2(n18360), .ZN(
        n18053) );
  NAND2_X1 U21216 ( .A1(n18337), .A2(n18053), .ZN(n18013) );
  NOR2_X1 U21217 ( .A1(n18484), .A2(n19056), .ZN(n18347) );
  NOR2_X1 U21218 ( .A1(n17989), .A2(n17984), .ZN(n17985) );
  AOI211_X1 U21219 ( .C1(n17987), .C2(n17986), .A(n18117), .B(n17985), .ZN(
        n18003) );
  NAND2_X1 U21220 ( .A1(n17989), .A2(n17988), .ZN(n18002) );
  OAI21_X1 U21221 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17990), .ZN(n17991) );
  OAI22_X1 U21222 ( .A1(n17992), .A2(n18003), .B1(n18002), .B2(n17991), .ZN(
        n17993) );
  AOI211_X1 U21223 ( .C1(n18006), .C2(n17994), .A(n18347), .B(n17993), .ZN(
        n18000) );
  OAI22_X1 U21224 ( .A1(n18341), .A2(n18025), .B1(n17995), .B2(n13159), .ZN(
        n18010) );
  AOI21_X1 U21225 ( .B1(n21466), .B2(n18030), .A(n17996), .ZN(n17997) );
  AOI21_X1 U21226 ( .B1(n18030), .B2(n18007), .A(n17997), .ZN(n17998) );
  XOR2_X1 U21227 ( .A(n17998), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18348) );
  AOI22_X1 U21228 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18010), .B1(
        n18069), .B2(n18348), .ZN(n17999) );
  OAI211_X1 U21229 ( .C1(n18350), .C2(n18013), .A(n18000), .B(n17999), .ZN(
        P3_U2817) );
  NOR2_X1 U21230 ( .A1(n18484), .A2(n19054), .ZN(n18355) );
  AOI22_X1 U21231 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18003), .B1(
        n18002), .B2(n18001), .ZN(n18004) );
  AOI211_X1 U21232 ( .C1(n18006), .C2(n18005), .A(n18355), .B(n18004), .ZN(
        n18012) );
  OAI21_X1 U21233 ( .B1(n18008), .B2(n18044), .A(n18007), .ZN(n18009) );
  XOR2_X1 U21234 ( .A(n18009), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18357) );
  AOI22_X1 U21235 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18010), .B1(
        n18069), .B2(n18357), .ZN(n18011) );
  OAI211_X1 U21236 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18013), .A(
        n18012), .B(n18011), .ZN(P3_U2818) );
  NOR2_X1 U21237 ( .A1(n18366), .A2(n18044), .ZN(n18015) );
  NOR2_X1 U21238 ( .A1(n18015), .A2(n18014), .ZN(n18016) );
  XOR2_X1 U21239 ( .A(n18016), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18371) );
  NOR2_X1 U21240 ( .A1(n18017), .A2(n18540), .ZN(n18065) );
  NAND2_X1 U21241 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18065), .ZN(
        n18049) );
  NOR2_X1 U21242 ( .A1(n18048), .A2(n18049), .ZN(n18046) );
  NAND2_X1 U21243 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18046), .ZN(
        n18033) );
  NOR2_X1 U21244 ( .A1(n18117), .A2(n19013), .ZN(n18047) );
  INV_X1 U21245 ( .A(n18047), .ZN(n18159) );
  NAND2_X1 U21246 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18159), .ZN(
        n18018) );
  AOI22_X1 U21247 ( .A1(n18019), .A2(n18065), .B1(n18033), .B2(n18018), .ZN(
        n18021) );
  INV_X1 U21248 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19052) );
  NOR2_X1 U21249 ( .A1(n18484), .A2(n19052), .ZN(n18020) );
  AOI211_X1 U21250 ( .C1(n18022), .C2(n18158), .A(n18021), .B(n18020), .ZN(
        n18029) );
  NOR2_X1 U21251 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18366), .ZN(
        n18359) );
  OAI22_X1 U21252 ( .A1(n18025), .A2(n18024), .B1(n13159), .B2(n18023), .ZN(
        n18054) );
  INV_X1 U21253 ( .A(n18054), .ZN(n18037) );
  NAND2_X1 U21254 ( .A1(n18366), .A2(n18053), .ZN(n18038) );
  AOI21_X1 U21255 ( .B1(n18037), .B2(n18038), .A(n18026), .ZN(n18027) );
  AOI21_X1 U21256 ( .B1(n18359), .B2(n18053), .A(n18027), .ZN(n18028) );
  OAI211_X1 U21257 ( .C1(n18371), .C2(n18057), .A(n18029), .B(n18028), .ZN(
        P3_U2819) );
  INV_X1 U21258 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18381) );
  INV_X1 U21259 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18036) );
  OAI221_X1 U21260 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18043), .C1(
        n18381), .C2(n18044), .A(n18036), .ZN(n18032) );
  NAND4_X1 U21261 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n9976), .A3(
        n18030), .A4(n18381), .ZN(n18031) );
  OAI211_X1 U21262 ( .C1(n18044), .C2(n18366), .A(n18032), .B(n18031), .ZN(
        n18379) );
  OAI211_X1 U21263 ( .C1(n18046), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18159), .B(n18033), .ZN(n18034) );
  OAI21_X1 U21264 ( .B1(n18150), .B2(n18035), .A(n18034), .ZN(n18041) );
  OAI22_X1 U21265 ( .A1(n18039), .A2(n18038), .B1(n18037), .B2(n18036), .ZN(
        n18040) );
  AOI211_X1 U21266 ( .C1(n18479), .C2(P3_REIP_REG_10__SCAN_IN), .A(n18041), 
        .B(n18040), .ZN(n18042) );
  OAI21_X1 U21267 ( .B1(n18057), .B2(n18379), .A(n18042), .ZN(P3_U2820) );
  NAND2_X1 U21268 ( .A1(n18044), .A2(n18043), .ZN(n18045) );
  XOR2_X1 U21269 ( .A(n18045), .B(n18381), .Z(n18391) );
  AOI211_X1 U21270 ( .C1(n18049), .C2(n18048), .A(n18047), .B(n18046), .ZN(
        n18051) );
  NOR2_X1 U21271 ( .A1(n18484), .A2(n19049), .ZN(n18050) );
  AOI211_X1 U21272 ( .C1(n18052), .C2(n18158), .A(n18051), .B(n18050), .ZN(
        n18056) );
  AOI22_X1 U21273 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18054), .B1(
        n18053), .B2(n18381), .ZN(n18055) );
  OAI211_X1 U21274 ( .C1(n18391), .C2(n18057), .A(n18056), .B(n18055), .ZN(
        P3_U2821) );
  OAI21_X1 U21275 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18059), .A(
        n18058), .ZN(n18409) );
  INV_X1 U21276 ( .A(n18074), .ZN(n18060) );
  AOI21_X1 U21277 ( .B1(n19013), .B2(n18060), .A(n18117), .ZN(n18085) );
  OAI21_X1 U21278 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18540), .A(
        n18085), .ZN(n18063) );
  OAI22_X1 U21279 ( .A1(n18150), .A2(n18061), .B1(n18484), .B2(n19048), .ZN(
        n18062) );
  AOI221_X1 U21280 ( .B1(n18065), .B2(n18064), .C1(n18063), .C2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(n18062), .ZN(n18072) );
  INV_X1 U21281 ( .A(n18067), .ZN(n18406) );
  AOI21_X1 U21282 ( .B1(n18068), .B2(n18067), .A(n18066), .ZN(n18403) );
  AOI22_X1 U21283 ( .A1(n18070), .A2(n18406), .B1(n18069), .B2(n18403), .ZN(
        n18071) );
  OAI211_X1 U21284 ( .C1(n13159), .C2(n18409), .A(n18072), .B(n18071), .ZN(
        P3_U2822) );
  NOR2_X1 U21285 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18540), .ZN(
        n18073) );
  AOI22_X1 U21286 ( .A1(n18479), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n18074), 
        .B2(n18073), .ZN(n18083) );
  NOR2_X1 U21287 ( .A1(n18076), .A2(n18075), .ZN(n18077) );
  XOR2_X1 U21288 ( .A(n18077), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18414) );
  OAI21_X1 U21289 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18079), .A(
        n18078), .ZN(n18417) );
  OAI22_X1 U21290 ( .A1(n18150), .A2(n18080), .B1(n18168), .B2(n18417), .ZN(
        n18081) );
  AOI21_X1 U21291 ( .B1(n18157), .B2(n18414), .A(n18081), .ZN(n18082) );
  OAI211_X1 U21292 ( .C1(n18085), .C2(n18084), .A(n18083), .B(n18082), .ZN(
        P3_U2823) );
  AOI22_X1 U21293 ( .A1(n18088), .A2(n18103), .B1(n18087), .B2(n18086), .ZN(
        n18092) );
  AOI22_X1 U21294 ( .A1(n18090), .A2(n18418), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18089), .ZN(n18091) );
  XNOR2_X1 U21295 ( .A(n18092), .B(n18091), .ZN(n18423) );
  NOR2_X1 U21296 ( .A1(n18097), .A2(n18540), .ZN(n18093) );
  AOI22_X1 U21297 ( .A1(n18479), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18093), 
        .B2(n18098), .ZN(n18102) );
  OAI21_X1 U21298 ( .B1(n18096), .B2(n18095), .A(n18094), .ZN(n18421) );
  OAI21_X1 U21299 ( .B1(n18540), .B2(n18097), .A(n18159), .ZN(n18109) );
  OAI22_X1 U21300 ( .A1(n18168), .A2(n18421), .B1(n18098), .B2(n18109), .ZN(
        n18099) );
  AOI21_X1 U21301 ( .B1(n18100), .B2(n18158), .A(n18099), .ZN(n18101) );
  OAI211_X1 U21302 ( .C1(n18423), .C2(n13159), .A(n18102), .B(n18101), .ZN(
        P3_U2824) );
  AOI21_X1 U21303 ( .B1(n18105), .B2(n18104), .A(n18103), .ZN(n18430) );
  NOR2_X1 U21304 ( .A1(n18484), .A2(n19041), .ZN(n18429) );
  AOI21_X1 U21305 ( .B1(n18106), .B2(n18164), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18110) );
  OAI21_X1 U21306 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18108), .A(
        n18107), .ZN(n18434) );
  OAI22_X1 U21307 ( .A1(n18110), .A2(n18109), .B1(n18168), .B2(n18434), .ZN(
        n18111) );
  AOI211_X1 U21308 ( .C1(n18157), .C2(n18430), .A(n18429), .B(n18111), .ZN(
        n18112) );
  OAI21_X1 U21309 ( .B1(n18150), .B2(n18113), .A(n18112), .ZN(P3_U2825) );
  AOI21_X1 U21310 ( .B1(n18116), .B2(n18115), .A(n18114), .ZN(n18441) );
  AOI22_X1 U21311 ( .A1(n18157), .A2(n18441), .B1(n18479), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n18126) );
  AOI21_X1 U21312 ( .B1(n19013), .B2(n18139), .A(n18117), .ZN(n18136) );
  OAI21_X1 U21313 ( .B1(n18121), .B2(n18120), .A(n18119), .ZN(n18439) );
  OAI22_X1 U21314 ( .A1(n18136), .A2(n18122), .B1(n18168), .B2(n18439), .ZN(
        n18123) );
  AOI21_X1 U21315 ( .B1(n18124), .B2(n18158), .A(n18123), .ZN(n18125) );
  OAI211_X1 U21316 ( .C1(n18540), .C2(n18127), .A(n18126), .B(n18125), .ZN(
        P3_U2826) );
  OAI21_X1 U21317 ( .B1(n18130), .B2(n18129), .A(n18128), .ZN(n18131) );
  XOR2_X1 U21318 ( .A(n18131), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n18454) );
  AOI21_X1 U21319 ( .B1(n18134), .B2(n18133), .A(n18132), .ZN(n18449) );
  NOR2_X1 U21320 ( .A1(n18484), .A2(n19037), .ZN(n18448) );
  OAI22_X1 U21321 ( .A1(n18150), .A2(n18137), .B1(n18136), .B2(n18135), .ZN(
        n18138) );
  AOI211_X1 U21322 ( .C1(n18157), .C2(n18449), .A(n18448), .B(n18138), .ZN(
        n18141) );
  NAND4_X1 U21323 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19013), .A3(
        n18164), .A4(n18139), .ZN(n18140) );
  OAI211_X1 U21324 ( .C1(n18454), .C2(n18168), .A(n18141), .B(n18140), .ZN(
        P3_U2827) );
  AOI21_X1 U21325 ( .B1(n18144), .B2(n18143), .A(n18142), .ZN(n18467) );
  INV_X1 U21326 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n21516) );
  NOR2_X1 U21327 ( .A1(n18484), .A2(n21516), .ZN(n18455) );
  INV_X1 U21328 ( .A(n18145), .ZN(n18149) );
  OAI21_X1 U21329 ( .B1(n18148), .B2(n18147), .A(n18146), .ZN(n18471) );
  OAI22_X1 U21330 ( .A1(n18150), .A2(n18149), .B1(n18168), .B2(n18471), .ZN(
        n18151) );
  AOI211_X1 U21331 ( .C1(n18157), .C2(n18467), .A(n18455), .B(n18151), .ZN(
        n18152) );
  OAI221_X1 U21332 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18540), .C1(
        n18153), .C2(n18164), .A(n18152), .ZN(P3_U2828) );
  OAI21_X1 U21333 ( .B1(n18162), .B2(n18155), .A(n18154), .ZN(n18483) );
  NAND2_X1 U21334 ( .A1(n19125), .A2(n18163), .ZN(n18156) );
  XNOR2_X1 U21335 ( .A(n18156), .B(n18155), .ZN(n18478) );
  AOI22_X1 U21336 ( .A1(n18157), .A2(n18478), .B1(n18479), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U21337 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18159), .B1(
        n18158), .B2(n21330), .ZN(n18160) );
  OAI211_X1 U21338 ( .C1(n18168), .C2(n18483), .A(n18161), .B(n18160), .ZN(
        P3_U2829) );
  AOI21_X1 U21339 ( .B1(n18163), .B2(n19125), .A(n18162), .ZN(n18486) );
  INV_X1 U21340 ( .A(n18486), .ZN(n18488) );
  NAND3_X1 U21341 ( .A1(n19109), .A2(n18165), .A3(n18164), .ZN(n18166) );
  AOI22_X1 U21342 ( .A1(n18479), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18166), .ZN(n18167) );
  OAI221_X1 U21343 ( .B1(n18486), .B2(n13159), .C1(n18488), .C2(n18168), .A(
        n18167), .ZN(P3_U2830) );
  NAND2_X1 U21344 ( .A1(n18484), .A2(n18490), .ZN(n18474) );
  AOI221_X1 U21345 ( .B1(n18246), .B2(n18170), .C1(n18169), .C2(n18170), .A(
        n18490), .ZN(n18181) );
  NOR3_X1 U21346 ( .A1(n19125), .A2(n18245), .A3(n18295), .ZN(n18248) );
  OAI221_X1 U21347 ( .B1(n18956), .B2(n18171), .C1(n18956), .C2(n18248), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18231) );
  INV_X1 U21348 ( .A(n18237), .ZN(n18221) );
  NOR3_X1 U21349 ( .A1(n18231), .A2(n18295), .A3(n18221), .ZN(n18172) );
  NOR2_X1 U21350 ( .A1(n18172), .A2(n18459), .ZN(n18209) );
  AOI21_X1 U21351 ( .B1(n18965), .B2(n18174), .A(n18173), .ZN(n18176) );
  OAI21_X1 U21352 ( .B1(n18194), .B2(n21488), .A(n18396), .ZN(n18175) );
  OAI211_X1 U21353 ( .C1(n18177), .C2(n18227), .A(n18176), .B(n18175), .ZN(
        n18178) );
  AOI211_X1 U21354 ( .C1(n18361), .C2(n18179), .A(n18209), .B(n18178), .ZN(
        n18185) );
  OAI211_X1 U21355 ( .C1(n18975), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n18185), .ZN(n18180) );
  AOI22_X1 U21356 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18456), .B1(
        n18181), .B2(n18180), .ZN(n18183) );
  NAND2_X1 U21357 ( .A1(n18479), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18182) );
  OAI211_X1 U21358 ( .C1(n18184), .C2(n18390), .A(n18183), .B(n18182), .ZN(
        P3_U2835) );
  AOI21_X1 U21359 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18185), .A(
        n18490), .ZN(n18189) );
  OAI21_X1 U21360 ( .B1(n18246), .B2(n18187), .A(n18186), .ZN(n18188) );
  OAI221_X1 U21361 ( .B1(n18189), .B2(n18456), .C1(n18189), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n18188), .ZN(n18190) );
  OAI211_X1 U21362 ( .C1(n18192), .C2(n18390), .A(n18191), .B(n18190), .ZN(
        P3_U2836) );
  NOR2_X1 U21363 ( .A1(n18193), .A2(n18981), .ZN(n18214) );
  AOI211_X1 U21364 ( .C1(n18393), .C2(n18194), .A(n18214), .B(n18209), .ZN(
        n18198) );
  NAND3_X1 U21365 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18196), .A3(
        n18195), .ZN(n18197) );
  AOI221_X1 U21366 ( .B1(n18198), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n18197), .C2(n21488), .A(n18490), .ZN(n18199) );
  AOI211_X1 U21367 ( .C1(n18456), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18200), .B(n18199), .ZN(n18204) );
  AOI22_X1 U21368 ( .A1(n18489), .A2(n18202), .B1(n18404), .B2(n18201), .ZN(
        n18203) );
  OAI211_X1 U21369 ( .C1(n18335), .C2(n18205), .A(n18204), .B(n18203), .ZN(
        P3_U2837) );
  NOR2_X1 U21370 ( .A1(n18246), .A2(n18490), .ZN(n18207) );
  AOI22_X1 U21371 ( .A1(n18404), .A2(n18208), .B1(n18207), .B2(n18206), .ZN(
        n18219) );
  AOI211_X1 U21372 ( .C1(n18361), .C2(n18210), .A(n18209), .B(n18456), .ZN(
        n18211) );
  OAI21_X1 U21373 ( .B1(n18212), .B2(n18227), .A(n18211), .ZN(n18216) );
  NOR3_X1 U21374 ( .A1(n18214), .A2(n18213), .A3(n18216), .ZN(n18215) );
  NOR2_X1 U21375 ( .A1(n18479), .A2(n18215), .ZN(n18222) );
  OAI211_X1 U21376 ( .C1(n18393), .C2(n18216), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18222), .ZN(n18217) );
  NAND3_X1 U21377 ( .A1(n18219), .A2(n18218), .A3(n18217), .ZN(P3_U2838) );
  INV_X1 U21378 ( .A(n18220), .ZN(n18226) );
  NOR4_X1 U21379 ( .A1(n18456), .A2(n18246), .A3(n18244), .A4(n18221), .ZN(
        n18223) );
  OAI21_X1 U21380 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18223), .A(
        n18222), .ZN(n18224) );
  OAI211_X1 U21381 ( .C1(n18226), .C2(n18390), .A(n18225), .B(n18224), .ZN(
        P3_U2839) );
  NAND2_X1 U21382 ( .A1(n18227), .A2(n18340), .ZN(n18365) );
  INV_X1 U21383 ( .A(n18365), .ZN(n18230) );
  AOI22_X1 U21384 ( .A1(n9866), .A2(n18306), .B1(n18361), .B2(n18305), .ZN(
        n18292) );
  NAND2_X1 U21385 ( .A1(n18967), .A2(n18228), .ZN(n18229) );
  OAI211_X1 U21386 ( .C1(n18237), .C2(n18230), .A(n18292), .B(n18229), .ZN(
        n18249) );
  AOI211_X1 U21387 ( .C1(n18342), .C2(n18232), .A(n18231), .B(n18249), .ZN(
        n18239) );
  INV_X1 U21388 ( .A(n18233), .ZN(n18260) );
  NOR2_X1 U21389 ( .A1(n18280), .A2(n18234), .ZN(n18277) );
  AOI21_X1 U21390 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18277), .A(
        n18981), .ZN(n18235) );
  AOI221_X1 U21391 ( .B1(n18295), .B2(n18967), .C1(n18260), .C2(n18967), .A(
        n18235), .ZN(n18247) );
  NAND2_X1 U21392 ( .A1(n18237), .A2(n18236), .ZN(n18238) );
  AOI22_X1 U21393 ( .A1(n18239), .A2(n18247), .B1(n18244), .B2(n18238), .ZN(
        n18241) );
  AOI22_X1 U21394 ( .A1(n18473), .A2(n18241), .B1(n18404), .B2(n18240), .ZN(
        n18243) );
  NAND2_X1 U21395 ( .A1(n18479), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18242) );
  OAI211_X1 U21396 ( .C1(n18474), .C2(n18244), .A(n18243), .B(n18242), .ZN(
        P3_U2840) );
  NOR3_X1 U21397 ( .A1(n18246), .A2(n18245), .A3(n18490), .ZN(n18267) );
  NOR2_X1 U21398 ( .A1(n18965), .A2(n18958), .ZN(n18318) );
  INV_X1 U21399 ( .A(n18318), .ZN(n18472) );
  OAI211_X1 U21400 ( .C1(n18956), .C2(n18248), .A(n18473), .B(n18247), .ZN(
        n18259) );
  AOI211_X1 U21401 ( .C1(n18250), .C2(n18472), .A(n18259), .B(n18249), .ZN(
        n18251) );
  NOR3_X1 U21402 ( .A1(n18479), .A2(n18251), .A3(n21522), .ZN(n18253) );
  AOI211_X1 U21403 ( .C1(n18254), .C2(n18267), .A(n18253), .B(n18252), .ZN(
        n18255) );
  OAI21_X1 U21404 ( .B1(n18256), .B2(n18390), .A(n18255), .ZN(P3_U2841) );
  AOI21_X1 U21405 ( .B1(n18258), .B2(n18267), .A(n18257), .ZN(n18264) );
  AOI21_X1 U21406 ( .B1(n18260), .B2(n18365), .A(n18259), .ZN(n18261) );
  AOI21_X1 U21407 ( .B1(n18292), .B2(n18261), .A(n18479), .ZN(n18268) );
  NOR3_X1 U21408 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18318), .A3(
        n19005), .ZN(n18262) );
  OAI21_X1 U21409 ( .B1(n18268), .B2(n18262), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18263) );
  OAI211_X1 U21410 ( .C1(n18265), .C2(n18390), .A(n18264), .B(n18263), .ZN(
        P3_U2842) );
  AOI22_X1 U21411 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18268), .B1(
        n18267), .B2(n18266), .ZN(n18270) );
  OAI211_X1 U21412 ( .C1(n18271), .C2(n18390), .A(n18270), .B(n18269), .ZN(
        P3_U2843) );
  OAI22_X1 U21413 ( .A1(n18462), .A2(n18981), .B1(n18272), .B2(n18466), .ZN(
        n18451) );
  NAND3_X1 U21414 ( .A1(n18274), .A2(n18273), .A3(n18451), .ZN(n18326) );
  NOR2_X1 U21415 ( .A1(n18327), .A2(n18326), .ZN(n18312) );
  OAI211_X1 U21416 ( .C1(n18275), .C2(n18312), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18473), .ZN(n18304) );
  AOI21_X1 U21417 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18276), .A(
        n18459), .ZN(n18279) );
  OAI211_X1 U21418 ( .C1(n18277), .C2(n18981), .A(n18473), .B(n18292), .ZN(
        n18278) );
  AOI211_X1 U21419 ( .C1(n18280), .C2(n18365), .A(n18279), .B(n18278), .ZN(
        n18286) );
  AOI221_X1 U21420 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18286), 
        .C1(n18459), .C2(n18286), .A(n18479), .ZN(n18282) );
  AOI22_X1 U21421 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18282), .B1(
        n18404), .B2(n18281), .ZN(n18284) );
  OAI211_X1 U21422 ( .C1(n18285), .C2(n18304), .A(n18284), .B(n18283), .ZN(
        P3_U2844) );
  NOR2_X1 U21423 ( .A1(n18479), .A2(n18286), .ZN(n18289) );
  NOR3_X1 U21424 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18303), .A3(
        n18304), .ZN(n18287) );
  AOI211_X1 U21425 ( .C1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18289), .A(
        n18288), .B(n18287), .ZN(n18290) );
  OAI21_X1 U21426 ( .B1(n18291), .B2(n18390), .A(n18290), .ZN(P3_U2845) );
  NAND2_X1 U21427 ( .A1(n18473), .A2(n18292), .ZN(n18299) );
  INV_X1 U21428 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18400) );
  NAND2_X1 U21429 ( .A1(n18419), .A2(n18437), .ZN(n18395) );
  NOR3_X1 U21430 ( .A1(n18418), .A2(n18411), .A3(n18395), .ZN(n18294) );
  OAI22_X1 U21431 ( .A1(n18975), .A2(n18294), .B1(n18293), .B2(n18981), .ZN(
        n18387) );
  AOI21_X1 U21432 ( .B1(n18967), .B2(n18400), .A(n18387), .ZN(n18374) );
  OAI22_X1 U21433 ( .A1(n18965), .A2(n18296), .B1(n19125), .B2(n18295), .ZN(
        n18297) );
  OAI211_X1 U21434 ( .C1(n18375), .C2(n18298), .A(n18374), .B(n18297), .ZN(
        n18313) );
  OAI221_X1 U21435 ( .B1(n18299), .B2(n18393), .C1(n18299), .C2(n18313), .A(
        n18484), .ZN(n18302) );
  AOI22_X1 U21436 ( .A1(n18479), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18404), 
        .B2(n18300), .ZN(n18301) );
  OAI221_X1 U21437 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18304), 
        .C1(n18303), .C2(n18302), .A(n18301), .ZN(P3_U2846) );
  NAND2_X1 U21438 ( .A1(n18361), .A2(n18305), .ZN(n18309) );
  NAND2_X1 U21439 ( .A1(n9866), .A2(n18306), .ZN(n18307) );
  OAI22_X1 U21440 ( .A1(n18310), .A2(n18309), .B1(n18308), .B2(n18307), .ZN(
        n18311) );
  AOI221_X1 U21441 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18313), 
        .C1(n18312), .C2(n18313), .A(n18311), .ZN(n18317) );
  AOI22_X1 U21442 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18456), .B1(
        n18404), .B2(n18314), .ZN(n18316) );
  OAI211_X1 U21443 ( .C1(n18317), .C2(n18490), .A(n18316), .B(n18315), .ZN(
        P3_U2847) );
  NOR2_X1 U21444 ( .A1(n18484), .A2(n19059), .ZN(n18329) );
  OAI22_X1 U21445 ( .A1(n18975), .A2(n18319), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18318), .ZN(n18324) );
  NOR2_X1 U21446 ( .A1(n19125), .A2(n18320), .ZN(n18385) );
  NAND2_X1 U21447 ( .A1(n18321), .A2(n18385), .ZN(n18352) );
  NAND2_X1 U21448 ( .A1(n18965), .A2(n18352), .ZN(n18344) );
  OAI211_X1 U21449 ( .C1(n18322), .C2(n18981), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18344), .ZN(n18323) );
  OAI21_X1 U21450 ( .B1(n18324), .B2(n18323), .A(n18473), .ZN(n18325) );
  AOI21_X1 U21451 ( .B1(n18327), .B2(n18326), .A(n18325), .ZN(n18328) );
  AOI211_X1 U21452 ( .C1(n18456), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18329), .B(n18328), .ZN(n18333) );
  AOI22_X1 U21453 ( .A1(n18405), .A2(n18331), .B1(n18489), .B2(n18330), .ZN(
        n18332) );
  OAI211_X1 U21454 ( .C1(n18390), .C2(n18334), .A(n18333), .B(n18332), .ZN(
        P3_U2848) );
  NAND2_X1 U21455 ( .A1(n18473), .A2(n18451), .ZN(n18435) );
  OAI222_X1 U21456 ( .A1(n18435), .A2(n18336), .B1(n18422), .B2(n18362), .C1(
        n18360), .C2(n18335), .ZN(n18380) );
  NAND2_X1 U21457 ( .A1(n18337), .A2(n18380), .ZN(n18354) );
  AOI21_X1 U21458 ( .B1(n18337), .B2(n18374), .A(n18375), .ZN(n18368) );
  AOI21_X1 U21459 ( .B1(n9866), .B2(n18338), .A(n18368), .ZN(n18339) );
  OAI21_X1 U21460 ( .B1(n18341), .B2(n18340), .A(n18339), .ZN(n18351) );
  AOI211_X1 U21461 ( .C1(n18342), .C2(n21466), .A(n18490), .B(n18351), .ZN(
        n18345) );
  AOI211_X1 U21462 ( .C1(n18345), .C2(n18344), .A(n18479), .B(n18343), .ZN(
        n18346) );
  AOI211_X1 U21463 ( .C1(n18348), .C2(n18404), .A(n18347), .B(n18346), .ZN(
        n18349) );
  OAI21_X1 U21464 ( .B1(n18350), .B2(n18354), .A(n18349), .ZN(P3_U2849) );
  AOI211_X1 U21465 ( .C1(n18352), .C2(n18965), .A(n18351), .B(n21466), .ZN(
        n18353) );
  AOI211_X1 U21466 ( .C1(n18354), .C2(n21466), .A(n18490), .B(n18353), .ZN(
        n18356) );
  AOI211_X1 U21467 ( .C1(n18404), .C2(n18357), .A(n18356), .B(n18355), .ZN(
        n18358) );
  OAI21_X1 U21468 ( .B1(n21466), .B2(n18474), .A(n18358), .ZN(P3_U2850) );
  AOI22_X1 U21469 ( .A1(n18479), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18359), 
        .B2(n18380), .ZN(n18370) );
  AOI21_X1 U21470 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18385), .A(
        n18956), .ZN(n18364) );
  AOI22_X1 U21471 ( .A1(n9866), .A2(n18362), .B1(n18361), .B2(n18360), .ZN(
        n18363) );
  NAND2_X1 U21472 ( .A1(n18473), .A2(n18363), .ZN(n18382) );
  AOI211_X1 U21473 ( .C1(n18366), .C2(n18365), .A(n18364), .B(n18382), .ZN(
        n18373) );
  OAI21_X1 U21474 ( .B1(n18956), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18373), .ZN(n18367) );
  OAI211_X1 U21475 ( .C1(n18368), .C2(n18367), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18484), .ZN(n18369) );
  OAI211_X1 U21476 ( .C1(n18371), .C2(n18390), .A(n18370), .B(n18369), .ZN(
        P3_U2851) );
  NOR2_X1 U21477 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18381), .ZN(
        n18372) );
  AOI22_X1 U21478 ( .A1(n18479), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18372), 
        .B2(n18380), .ZN(n18378) );
  OAI211_X1 U21479 ( .C1(n18375), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18374), .B(n18373), .ZN(n18376) );
  NAND3_X1 U21480 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18484), .A3(
        n18376), .ZN(n18377) );
  OAI211_X1 U21481 ( .C1(n18390), .C2(n18379), .A(n18378), .B(n18377), .ZN(
        P3_U2852) );
  AOI22_X1 U21482 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18479), .B1(n18381), 
        .B2(n18380), .ZN(n18389) );
  NAND2_X1 U21483 ( .A1(n18967), .A2(n18400), .ZN(n18384) );
  INV_X1 U21484 ( .A(n18382), .ZN(n18383) );
  OAI211_X1 U21485 ( .C1(n18385), .C2(n18956), .A(n18384), .B(n18383), .ZN(
        n18386) );
  OAI211_X1 U21486 ( .C1(n18387), .C2(n18386), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18484), .ZN(n18388) );
  OAI211_X1 U21487 ( .C1(n18391), .C2(n18390), .A(n18389), .B(n18388), .ZN(
        P3_U2853) );
  NAND2_X1 U21488 ( .A1(n18392), .A2(n18451), .ZN(n18410) );
  OAI21_X1 U21489 ( .B1(n18411), .B2(n18410), .A(n18400), .ZN(n18402) );
  INV_X1 U21490 ( .A(n18393), .ZN(n18398) );
  NOR2_X1 U21491 ( .A1(n18418), .A2(n18411), .ZN(n18397) );
  AOI21_X1 U21492 ( .B1(n18462), .B2(n18958), .A(n18461), .ZN(n18436) );
  OAI21_X1 U21493 ( .B1(n18419), .B2(n18981), .A(n18436), .ZN(n18394) );
  AOI21_X1 U21494 ( .B1(n18396), .B2(n18395), .A(n18394), .ZN(n18420) );
  OAI21_X1 U21495 ( .B1(n18398), .B2(n18397), .A(n18420), .ZN(n18412) );
  AOI22_X1 U21496 ( .A1(n18438), .A2(n18412), .B1(n18473), .B2(n18400), .ZN(
        n18399) );
  OAI21_X1 U21497 ( .B1(n18400), .B2(n18474), .A(n18399), .ZN(n18401) );
  AOI22_X1 U21498 ( .A1(n18479), .A2(P3_REIP_REG_8__SCAN_IN), .B1(n18402), 
        .B2(n18401), .ZN(n18408) );
  AOI22_X1 U21499 ( .A1(n18406), .A2(n18405), .B1(n18404), .B2(n18403), .ZN(
        n18407) );
  OAI211_X1 U21500 ( .C1(n18422), .C2(n18409), .A(n18408), .B(n18407), .ZN(
        P3_U2854) );
  AOI22_X1 U21501 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18456), .B1(
        n18479), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n18416) );
  AOI21_X1 U21502 ( .B1(n18411), .B2(n18410), .A(n18490), .ZN(n18413) );
  AOI22_X1 U21503 ( .A1(n18489), .A2(n18414), .B1(n18413), .B2(n18412), .ZN(
        n18415) );
  OAI211_X1 U21504 ( .C1(n18482), .C2(n18417), .A(n18416), .B(n18415), .ZN(
        P3_U2855) );
  NAND2_X1 U21505 ( .A1(n18419), .A2(n18418), .ZN(n18427) );
  OAI21_X1 U21506 ( .B1(n18420), .B2(n18490), .A(n18474), .ZN(n18431) );
  OAI22_X1 U21507 ( .A1(n18423), .A2(n18422), .B1(n18482), .B2(n18421), .ZN(
        n18424) );
  AOI21_X1 U21508 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18431), .A(
        n18424), .ZN(n18426) );
  NAND2_X1 U21509 ( .A1(n18479), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18425) );
  OAI211_X1 U21510 ( .C1(n18435), .C2(n18427), .A(n18426), .B(n18425), .ZN(
        P3_U2856) );
  NOR4_X1 U21511 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18446), .A3(
        n18444), .A4(n18435), .ZN(n18428) );
  AOI211_X1 U21512 ( .C1(n18489), .C2(n18430), .A(n18429), .B(n18428), .ZN(
        n18433) );
  NAND2_X1 U21513 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18431), .ZN(
        n18432) );
  OAI211_X1 U21514 ( .C1(n18434), .C2(n18482), .A(n18433), .B(n18432), .ZN(
        P3_U2857) );
  OR2_X1 U21515 ( .A1(n18446), .A2(n18435), .ZN(n18445) );
  OAI211_X1 U21516 ( .C1(n18459), .C2(n18437), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18436), .ZN(n18450) );
  AOI21_X1 U21517 ( .B1(n18438), .B2(n18450), .A(n18456), .ZN(n18443) );
  OAI22_X1 U21518 ( .A1(n18484), .A2(n19039), .B1(n18482), .B2(n18439), .ZN(
        n18440) );
  AOI21_X1 U21519 ( .B1(n18489), .B2(n18441), .A(n18440), .ZN(n18442) );
  OAI221_X1 U21520 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18445), .C1(
        n18444), .C2(n18443), .A(n18442), .ZN(P3_U2858) );
  NOR2_X1 U21521 ( .A1(n18446), .A2(n18474), .ZN(n18447) );
  AOI211_X1 U21522 ( .C1(n18489), .C2(n18449), .A(n18448), .B(n18447), .ZN(
        n18453) );
  OAI211_X1 U21523 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18451), .A(
        n18473), .B(n18450), .ZN(n18452) );
  OAI211_X1 U21524 ( .C1(n18454), .C2(n18482), .A(n18453), .B(n18452), .ZN(
        P3_U2859) );
  AOI21_X1 U21525 ( .B1(n18456), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18455), .ZN(n18470) );
  NAND2_X1 U21526 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18457), .ZN(
        n18465) );
  NAND2_X1 U21527 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18458) );
  OAI22_X1 U21528 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18459), .B1(
        n18981), .B2(n18458), .ZN(n18460) );
  OAI21_X1 U21529 ( .B1(n18461), .B2(n18460), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18464) );
  NAND2_X1 U21530 ( .A1(n18958), .A2(n18462), .ZN(n18463) );
  OAI211_X1 U21531 ( .C1(n18466), .C2(n18465), .A(n18464), .B(n18463), .ZN(
        n18468) );
  AOI22_X1 U21532 ( .A1(n18473), .A2(n18468), .B1(n18489), .B2(n18467), .ZN(
        n18469) );
  OAI211_X1 U21533 ( .C1(n18482), .C2(n18471), .A(n18470), .B(n18469), .ZN(
        P3_U2860) );
  NAND3_X1 U21534 ( .A1(n18473), .A2(n19125), .A3(n18472), .ZN(n18492) );
  INV_X1 U21535 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19110) );
  AOI21_X1 U21536 ( .B1(n18474), .B2(n18492), .A(n19110), .ZN(n18477) );
  AOI211_X1 U21537 ( .C1(n18975), .C2(n19125), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18475), .ZN(n18476) );
  AOI211_X1 U21538 ( .C1(n18489), .C2(n18478), .A(n18477), .B(n18476), .ZN(
        n18481) );
  NAND2_X1 U21539 ( .A1(n18479), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18480) );
  OAI211_X1 U21540 ( .C1(n18483), .C2(n18482), .A(n18481), .B(n18480), .ZN(
        P3_U2861) );
  NOR2_X1 U21541 ( .A1(n18484), .A2(n19136), .ZN(n18485) );
  AOI221_X1 U21542 ( .B1(n18489), .B2(n18488), .C1(n18487), .C2(n18486), .A(
        n18485), .ZN(n18493) );
  OAI211_X1 U21543 ( .C1(n18967), .C2(n18490), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18484), .ZN(n18491) );
  NAND3_X1 U21544 ( .A1(n18493), .A2(n18492), .A3(n18491), .ZN(P3_U2862) );
  OAI211_X1 U21545 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18494), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n19004)
         );
  OAI21_X1 U21546 ( .B1(n18496), .B2(n19148), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18495) );
  OAI221_X1 U21547 ( .B1(n18496), .B2(n19004), .C1(n18496), .C2(n18549), .A(
        n18495), .ZN(P3_U2863) );
  INV_X1 U21548 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18987) );
  NAND2_X1 U21549 ( .A1(n18497), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18772) );
  INV_X1 U21550 ( .A(n18772), .ZN(n18794) );
  NOR2_X1 U21551 ( .A1(n18497), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18681) );
  NOR2_X1 U21552 ( .A1(n18794), .A2(n18681), .ZN(n18499) );
  OAI22_X1 U21553 ( .A1(n18500), .A2(n18987), .B1(n18499), .B2(n18498), .ZN(
        P3_U2866) );
  NOR2_X1 U21554 ( .A1(n18502), .A2(n18501), .ZN(P3_U2867) );
  NAND2_X1 U21555 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18883), .ZN(n18855) );
  NAND2_X1 U21556 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18504) );
  NOR2_X1 U21557 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18504), .ZN(
        n18882) );
  INV_X1 U21558 ( .A(n18882), .ZN(n18821) );
  NOR2_X2 U21559 ( .A1(n18968), .A2(n18821), .ZN(n18929) );
  INV_X1 U21560 ( .A(n18929), .ZN(n18887) );
  NAND2_X1 U21561 ( .A1(n18883), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18888) );
  INV_X1 U21562 ( .A(n18888), .ZN(n18845) );
  NAND2_X1 U21563 ( .A1(n18968), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18749) );
  NOR2_X2 U21564 ( .A1(n18749), .A2(n18504), .ZN(n18851) );
  NOR2_X2 U21565 ( .A1(n18541), .A2(n18503), .ZN(n18878) );
  NOR2_X1 U21566 ( .A1(n18987), .A2(n18679), .ZN(n18881) );
  NAND2_X1 U21567 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18881), .ZN(
        n18925) );
  NOR2_X1 U21568 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18972) );
  NOR2_X1 U21569 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18590) );
  NAND2_X1 U21570 ( .A1(n18972), .A2(n18590), .ZN(n18610) );
  NAND2_X1 U21571 ( .A1(n18925), .A2(n18610), .ZN(n18505) );
  INV_X1 U21572 ( .A(n18505), .ZN(n18569) );
  NOR2_X1 U21573 ( .A1(n18844), .A2(n18569), .ZN(n18543) );
  AOI22_X1 U21574 ( .A1(n18845), .A2(n18851), .B1(n18878), .B2(n18543), .ZN(
        n18510) );
  INV_X1 U21575 ( .A(n18749), .ZN(n18568) );
  NAND2_X1 U21576 ( .A1(n18969), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18635) );
  INV_X1 U21577 ( .A(n18635), .ZN(n18728) );
  NOR2_X1 U21578 ( .A1(n18568), .A2(n18728), .ZN(n18797) );
  NOR2_X1 U21579 ( .A1(n18797), .A2(n18504), .ZN(n18843) );
  AOI21_X1 U21580 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18541), .ZN(n18702) );
  AOI22_X1 U21581 ( .A1(n18883), .A2(n18843), .B1(n18702), .B2(n18505), .ZN(
        n18546) );
  NOR2_X1 U21582 ( .A1(n18507), .A2(n18506), .ZN(n18544) );
  INV_X1 U21583 ( .A(n18544), .ZN(n18522) );
  NOR2_X2 U21584 ( .A1(n18508), .A2(n18522), .ZN(n18884) );
  INV_X1 U21585 ( .A(n18610), .ZN(n18603) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18546), .B1(
        n18884), .B2(n18603), .ZN(n18509) );
  OAI211_X1 U21587 ( .C1(n18855), .C2(n18887), .A(n18510), .B(n18509), .ZN(
        P3_U2868) );
  NAND2_X1 U21588 ( .A1(n18544), .A2(n18511), .ZN(n18894) );
  NOR2_X2 U21589 ( .A1(n18541), .A2(n18512), .ZN(n18890) );
  NOR2_X2 U21590 ( .A1(n18513), .A2(n18540), .ZN(n18889) );
  AOI22_X1 U21591 ( .A1(n18890), .A2(n18543), .B1(n18889), .B2(n18929), .ZN(
        n18515) );
  AND2_X1 U21592 ( .A1(n18883), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18891) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18546), .B1(
        n18891), .B2(n18851), .ZN(n18514) );
  OAI211_X1 U21594 ( .C1(n18894), .C2(n18610), .A(n18515), .B(n18514), .ZN(
        P3_U2869) );
  NOR2_X1 U21595 ( .A1(n18516), .A2(n18522), .ZN(n18803) );
  INV_X1 U21596 ( .A(n18803), .ZN(n18900) );
  NOR2_X1 U21597 ( .A1(n21500), .A2(n18540), .ZN(n18896) );
  NOR2_X2 U21598 ( .A1(n18541), .A2(n18517), .ZN(n18895) );
  AOI22_X1 U21599 ( .A1(n18896), .A2(n18929), .B1(n18895), .B2(n18543), .ZN(
        n18520) );
  NOR2_X2 U21600 ( .A1(n18540), .A2(n18518), .ZN(n18897) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18546), .B1(
        n18897), .B2(n18851), .ZN(n18519) );
  OAI211_X1 U21602 ( .C1(n18900), .C2(n18610), .A(n18520), .B(n18519), .ZN(
        P3_U2870) );
  OR2_X1 U21603 ( .A1(n18522), .A2(n18521), .ZN(n18906) );
  AND2_X1 U21604 ( .A1(n18883), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18903) );
  AND2_X1 U21605 ( .A1(n18850), .A2(BUF2_REG_3__SCAN_IN), .ZN(n18902) );
  AOI22_X1 U21606 ( .A1(n18903), .A2(n18851), .B1(n18902), .B2(n18543), .ZN(
        n18525) );
  INV_X1 U21607 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18523) );
  NOR2_X2 U21608 ( .A1(n18523), .A2(n18540), .ZN(n18901) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18546), .B1(
        n18901), .B2(n18929), .ZN(n18524) );
  OAI211_X1 U21610 ( .C1(n18906), .C2(n18610), .A(n18525), .B(n18524), .ZN(
        P3_U2871) );
  NOR2_X1 U21611 ( .A1(n18526), .A2(n18540), .ZN(n18862) );
  AND2_X1 U21612 ( .A1(n18883), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18908) );
  NOR2_X2 U21613 ( .A1(n18541), .A2(n18527), .ZN(n18907) );
  AOI22_X1 U21614 ( .A1(n18908), .A2(n18851), .B1(n18907), .B2(n18543), .ZN(
        n18530) );
  NAND2_X1 U21615 ( .A1(n18528), .A2(n18544), .ZN(n18865) );
  INV_X1 U21616 ( .A(n18865), .ZN(n18909) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18546), .B1(
        n18909), .B2(n18603), .ZN(n18529) );
  OAI211_X1 U21618 ( .C1(n18912), .C2(n18887), .A(n18530), .B(n18529), .ZN(
        P3_U2872) );
  NAND2_X1 U21619 ( .A1(n18544), .A2(n18531), .ZN(n18918) );
  AND2_X1 U21620 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18883), .ZN(n18915) );
  NOR2_X2 U21621 ( .A1(n18541), .A2(n18532), .ZN(n18913) );
  AOI22_X1 U21622 ( .A1(n18915), .A2(n18929), .B1(n18913), .B2(n18543), .ZN(
        n18534) );
  NOR2_X2 U21623 ( .A1(n18540), .A2(n15357), .ZN(n18914) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18546), .B1(
        n18914), .B2(n18851), .ZN(n18533) );
  OAI211_X1 U21625 ( .C1(n18918), .C2(n18610), .A(n18534), .B(n18533), .ZN(
        P3_U2873) );
  NAND2_X1 U21626 ( .A1(n18544), .A2(n18535), .ZN(n18926) );
  NOR2_X2 U21627 ( .A1(n21395), .A2(n18540), .ZN(n18922) );
  NOR2_X2 U21628 ( .A1(n18541), .A2(n18536), .ZN(n18919) );
  AOI22_X1 U21629 ( .A1(n18922), .A2(n18929), .B1(n18919), .B2(n18543), .ZN(
        n18538) );
  INV_X1 U21630 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19560) );
  NOR2_X2 U21631 ( .A1(n18540), .A2(n19560), .ZN(n18920) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18546), .B1(
        n18920), .B2(n18851), .ZN(n18537) );
  OAI211_X1 U21633 ( .C1(n18926), .C2(n18610), .A(n18538), .B(n18537), .ZN(
        P3_U2874) );
  NOR2_X1 U21634 ( .A1(n18540), .A2(n18539), .ZN(n18872) );
  INV_X1 U21635 ( .A(n18872), .ZN(n18937) );
  AND2_X1 U21636 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18883), .ZN(n18930) );
  NOR2_X2 U21637 ( .A1(n18542), .A2(n18541), .ZN(n18928) );
  AOI22_X1 U21638 ( .A1(n18930), .A2(n18851), .B1(n18928), .B2(n18543), .ZN(
        n18548) );
  NAND2_X1 U21639 ( .A1(n18545), .A2(n18544), .ZN(n18877) );
  INV_X1 U21640 ( .A(n18877), .ZN(n18932) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18546), .B1(
        n18932), .B2(n18603), .ZN(n18547) );
  OAI211_X1 U21642 ( .C1(n18937), .C2(n18887), .A(n18548), .B(n18547), .ZN(
        P3_U2875) );
  INV_X1 U21643 ( .A(n18851), .ZN(n18876) );
  INV_X1 U21644 ( .A(n18925), .ZN(n18931) );
  INV_X1 U21645 ( .A(n18590), .ZN(n18589) );
  NAND2_X1 U21646 ( .A1(n18969), .A2(n19006), .ZN(n18725) );
  NOR2_X1 U21647 ( .A1(n18589), .A2(n18725), .ZN(n18564) );
  AOI22_X1 U21648 ( .A1(n18845), .A2(n18931), .B1(n18878), .B2(n18564), .ZN(
        n18551) );
  NAND2_X1 U21649 ( .A1(n18850), .A2(n18549), .ZN(n18726) );
  NOR2_X1 U21650 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18726), .ZN(
        n18633) );
  AOI22_X1 U21651 ( .A1(n18883), .A2(n18881), .B1(n18590), .B2(n18633), .ZN(
        n18565) );
  NAND2_X1 U21652 ( .A1(n18728), .A2(n18590), .ZN(n18632) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18565), .B1(
        n18884), .B2(n18625), .ZN(n18550) );
  OAI211_X1 U21654 ( .C1(n18855), .C2(n18876), .A(n18551), .B(n18550), .ZN(
        P3_U2876) );
  AOI22_X1 U21655 ( .A1(n18890), .A2(n18564), .B1(n18889), .B2(n18851), .ZN(
        n18553) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18565), .B1(
        n18891), .B2(n18931), .ZN(n18552) );
  OAI211_X1 U21657 ( .C1(n18894), .C2(n18632), .A(n18553), .B(n18552), .ZN(
        P3_U2877) );
  AOI22_X1 U21658 ( .A1(n18895), .A2(n18564), .B1(n18897), .B2(n18931), .ZN(
        n18555) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18565), .B1(
        n18803), .B2(n18625), .ZN(n18554) );
  OAI211_X1 U21660 ( .C1(n18806), .C2(n18876), .A(n18555), .B(n18554), .ZN(
        P3_U2878) );
  AOI22_X1 U21661 ( .A1(n18902), .A2(n18564), .B1(n18901), .B2(n18851), .ZN(
        n18557) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18565), .B1(
        n18903), .B2(n18931), .ZN(n18556) );
  OAI211_X1 U21663 ( .C1(n18906), .C2(n18632), .A(n18557), .B(n18556), .ZN(
        P3_U2879) );
  AOI22_X1 U21664 ( .A1(n18862), .A2(n18851), .B1(n18907), .B2(n18564), .ZN(
        n18559) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18565), .B1(
        n18908), .B2(n18931), .ZN(n18558) );
  OAI211_X1 U21666 ( .C1(n18865), .C2(n18632), .A(n18559), .B(n18558), .ZN(
        P3_U2880) );
  AOI22_X1 U21667 ( .A1(n18915), .A2(n18851), .B1(n18913), .B2(n18564), .ZN(
        n18561) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18565), .B1(
        n18914), .B2(n18931), .ZN(n18560) );
  OAI211_X1 U21669 ( .C1(n18918), .C2(n18632), .A(n18561), .B(n18560), .ZN(
        P3_U2881) );
  AOI22_X1 U21670 ( .A1(n18920), .A2(n18931), .B1(n18919), .B2(n18564), .ZN(
        n18563) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18565), .B1(
        n18922), .B2(n18851), .ZN(n18562) );
  OAI211_X1 U21672 ( .C1(n18926), .C2(n18632), .A(n18563), .B(n18562), .ZN(
        P3_U2882) );
  AOI22_X1 U21673 ( .A1(n18872), .A2(n18851), .B1(n18928), .B2(n18564), .ZN(
        n18567) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18565), .B1(
        n18930), .B2(n18931), .ZN(n18566) );
  OAI211_X1 U21675 ( .C1(n18877), .C2(n18632), .A(n18567), .B(n18566), .ZN(
        P3_U2883) );
  INV_X1 U21676 ( .A(n18855), .ZN(n18879) );
  NAND2_X1 U21677 ( .A1(n18568), .A2(n18590), .ZN(n18655) );
  NOR2_X1 U21678 ( .A1(n18625), .A2(n18648), .ZN(n18611) );
  NOR2_X1 U21679 ( .A1(n18844), .A2(n18611), .ZN(n18585) );
  AOI22_X1 U21680 ( .A1(n18879), .A2(n18931), .B1(n18878), .B2(n18585), .ZN(
        n18572) );
  OAI21_X1 U21681 ( .B1(n18569), .B2(n18847), .A(n18611), .ZN(n18570) );
  OAI211_X1 U21682 ( .C1(n18648), .C2(n19102), .A(n18850), .B(n18570), .ZN(
        n18586) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18586), .B1(
        n18884), .B2(n18648), .ZN(n18571) );
  OAI211_X1 U21684 ( .C1(n18888), .C2(n18610), .A(n18572), .B(n18571), .ZN(
        P3_U2884) );
  AOI22_X1 U21685 ( .A1(n18890), .A2(n18585), .B1(n18889), .B2(n18931), .ZN(
        n18574) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18586), .B1(
        n18891), .B2(n18603), .ZN(n18573) );
  OAI211_X1 U21687 ( .C1(n18894), .C2(n18655), .A(n18574), .B(n18573), .ZN(
        P3_U2885) );
  AOI22_X1 U21688 ( .A1(n18895), .A2(n18585), .B1(n18897), .B2(n18603), .ZN(
        n18576) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18586), .B1(
        n18896), .B2(n18931), .ZN(n18575) );
  OAI211_X1 U21690 ( .C1(n18900), .C2(n18655), .A(n18576), .B(n18575), .ZN(
        P3_U2886) );
  AOI22_X1 U21691 ( .A1(n18903), .A2(n18603), .B1(n18902), .B2(n18585), .ZN(
        n18578) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18586), .B1(
        n18901), .B2(n18931), .ZN(n18577) );
  OAI211_X1 U21693 ( .C1(n18906), .C2(n18655), .A(n18578), .B(n18577), .ZN(
        P3_U2887) );
  AOI22_X1 U21694 ( .A1(n18908), .A2(n18603), .B1(n18907), .B2(n18585), .ZN(
        n18580) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18586), .B1(
        n18862), .B2(n18931), .ZN(n18579) );
  OAI211_X1 U21696 ( .C1(n18865), .C2(n18655), .A(n18580), .B(n18579), .ZN(
        P3_U2888) );
  AOI22_X1 U21697 ( .A1(n18914), .A2(n18603), .B1(n18913), .B2(n18585), .ZN(
        n18582) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18586), .B1(
        n18915), .B2(n18931), .ZN(n18581) );
  OAI211_X1 U21699 ( .C1(n18918), .C2(n18655), .A(n18582), .B(n18581), .ZN(
        P3_U2889) );
  AOI22_X1 U21700 ( .A1(n18922), .A2(n18931), .B1(n18919), .B2(n18585), .ZN(
        n18584) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18586), .B1(
        n18920), .B2(n18603), .ZN(n18583) );
  OAI211_X1 U21702 ( .C1(n18926), .C2(n18655), .A(n18584), .B(n18583), .ZN(
        P3_U2890) );
  AOI22_X1 U21703 ( .A1(n18930), .A2(n18603), .B1(n18928), .B2(n18585), .ZN(
        n18588) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18586), .B1(
        n18872), .B2(n18931), .ZN(n18587) );
  OAI211_X1 U21705 ( .C1(n18877), .C2(n18655), .A(n18588), .B(n18587), .ZN(
        P3_U2891) );
  NOR2_X1 U21706 ( .A1(n18969), .A2(n18589), .ZN(n18634) );
  AND2_X1 U21707 ( .A1(n19006), .A2(n18634), .ZN(n18606) );
  AOI22_X1 U21708 ( .A1(n18845), .A2(n18625), .B1(n18878), .B2(n18606), .ZN(
        n18592) );
  AOI21_X1 U21709 ( .B1(n18969), .B2(n18847), .A(n18726), .ZN(n18680) );
  NAND2_X1 U21710 ( .A1(n18590), .A2(n18680), .ZN(n18607) );
  NAND2_X1 U21711 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18634), .ZN(
        n18678) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18607), .B1(
        n18671), .B2(n18884), .ZN(n18591) );
  OAI211_X1 U21713 ( .C1(n18855), .C2(n18610), .A(n18592), .B(n18591), .ZN(
        P3_U2892) );
  AOI22_X1 U21714 ( .A1(n18890), .A2(n18606), .B1(n18889), .B2(n18603), .ZN(
        n18594) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18607), .B1(
        n18891), .B2(n18625), .ZN(n18593) );
  OAI211_X1 U21716 ( .C1(n18678), .C2(n18894), .A(n18594), .B(n18593), .ZN(
        P3_U2893) );
  AOI22_X1 U21717 ( .A1(n18895), .A2(n18606), .B1(n18897), .B2(n18625), .ZN(
        n18596) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18607), .B1(
        n18671), .B2(n18803), .ZN(n18595) );
  OAI211_X1 U21719 ( .C1(n18806), .C2(n18610), .A(n18596), .B(n18595), .ZN(
        P3_U2894) );
  AOI22_X1 U21720 ( .A1(n18902), .A2(n18606), .B1(n18901), .B2(n18603), .ZN(
        n18598) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18607), .B1(
        n18903), .B2(n18625), .ZN(n18597) );
  OAI211_X1 U21722 ( .C1(n18678), .C2(n18906), .A(n18598), .B(n18597), .ZN(
        P3_U2895) );
  AOI22_X1 U21723 ( .A1(n18908), .A2(n18625), .B1(n18907), .B2(n18606), .ZN(
        n18600) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18607), .B1(
        n18671), .B2(n18909), .ZN(n18599) );
  OAI211_X1 U21725 ( .C1(n18912), .C2(n18610), .A(n18600), .B(n18599), .ZN(
        P3_U2896) );
  AOI22_X1 U21726 ( .A1(n18915), .A2(n18603), .B1(n18913), .B2(n18606), .ZN(
        n18602) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18607), .B1(
        n18914), .B2(n18625), .ZN(n18601) );
  OAI211_X1 U21728 ( .C1(n18678), .C2(n18918), .A(n18602), .B(n18601), .ZN(
        P3_U2897) );
  AOI22_X1 U21729 ( .A1(n18920), .A2(n18625), .B1(n18919), .B2(n18606), .ZN(
        n18605) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18607), .B1(
        n18922), .B2(n18603), .ZN(n18604) );
  OAI211_X1 U21731 ( .C1(n18678), .C2(n18926), .A(n18605), .B(n18604), .ZN(
        P3_U2898) );
  AOI22_X1 U21732 ( .A1(n18930), .A2(n18625), .B1(n18928), .B2(n18606), .ZN(
        n18609) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18607), .B1(
        n18671), .B2(n18932), .ZN(n18608) );
  OAI211_X1 U21734 ( .C1(n18937), .C2(n18610), .A(n18609), .B(n18608), .ZN(
        P3_U2899) );
  NAND2_X1 U21735 ( .A1(n18972), .A2(n18681), .ZN(n18701) );
  NOR2_X1 U21736 ( .A1(n18694), .A2(n18671), .ZN(n18657) );
  NOR2_X1 U21737 ( .A1(n18844), .A2(n18657), .ZN(n18628) );
  AOI22_X1 U21738 ( .A1(n18845), .A2(n18648), .B1(n18878), .B2(n18628), .ZN(
        n18614) );
  AOI221_X1 U21739 ( .B1(n18611), .B2(n18678), .C1(n18847), .C2(n18678), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18612) );
  OAI21_X1 U21740 ( .B1(n18694), .B2(n18612), .A(n18850), .ZN(n18629) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18629), .B1(
        n18694), .B2(n18884), .ZN(n18613) );
  OAI211_X1 U21742 ( .C1(n18855), .C2(n18632), .A(n18614), .B(n18613), .ZN(
        P3_U2900) );
  AOI22_X1 U21743 ( .A1(n18890), .A2(n18628), .B1(n18889), .B2(n18625), .ZN(
        n18616) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18629), .B1(
        n18891), .B2(n18648), .ZN(n18615) );
  OAI211_X1 U21745 ( .C1(n18701), .C2(n18894), .A(n18616), .B(n18615), .ZN(
        P3_U2901) );
  AOI22_X1 U21746 ( .A1(n18896), .A2(n18625), .B1(n18895), .B2(n18628), .ZN(
        n18618) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18629), .B1(
        n18897), .B2(n18648), .ZN(n18617) );
  OAI211_X1 U21748 ( .C1(n18701), .C2(n18900), .A(n18618), .B(n18617), .ZN(
        P3_U2902) );
  AOI22_X1 U21749 ( .A1(n18903), .A2(n18648), .B1(n18902), .B2(n18628), .ZN(
        n18620) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18629), .B1(
        n18901), .B2(n18625), .ZN(n18619) );
  OAI211_X1 U21751 ( .C1(n18701), .C2(n18906), .A(n18620), .B(n18619), .ZN(
        P3_U2903) );
  AOI22_X1 U21752 ( .A1(n18908), .A2(n18648), .B1(n18907), .B2(n18628), .ZN(
        n18622) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18629), .B1(
        n18694), .B2(n18909), .ZN(n18621) );
  OAI211_X1 U21754 ( .C1(n18912), .C2(n18632), .A(n18622), .B(n18621), .ZN(
        P3_U2904) );
  AOI22_X1 U21755 ( .A1(n18914), .A2(n18648), .B1(n18913), .B2(n18628), .ZN(
        n18624) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18629), .B1(
        n18915), .B2(n18625), .ZN(n18623) );
  OAI211_X1 U21757 ( .C1(n18701), .C2(n18918), .A(n18624), .B(n18623), .ZN(
        P3_U2905) );
  AOI22_X1 U21758 ( .A1(n18920), .A2(n18648), .B1(n18919), .B2(n18628), .ZN(
        n18627) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18629), .B1(
        n18922), .B2(n18625), .ZN(n18626) );
  OAI211_X1 U21760 ( .C1(n18701), .C2(n18926), .A(n18627), .B(n18626), .ZN(
        P3_U2906) );
  AOI22_X1 U21761 ( .A1(n18930), .A2(n18648), .B1(n18928), .B2(n18628), .ZN(
        n18631) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18629), .B1(
        n18694), .B2(n18932), .ZN(n18630) );
  OAI211_X1 U21763 ( .C1(n18937), .C2(n18632), .A(n18631), .B(n18630), .ZN(
        P3_U2907) );
  INV_X1 U21764 ( .A(n18681), .ZN(n18656) );
  NOR2_X1 U21765 ( .A1(n18656), .A2(n18725), .ZN(n18651) );
  AOI22_X1 U21766 ( .A1(n18671), .A2(n18845), .B1(n18878), .B2(n18651), .ZN(
        n18637) );
  AOI22_X1 U21767 ( .A1(n18883), .A2(n18634), .B1(n18681), .B2(n18633), .ZN(
        n18652) );
  NOR2_X2 U21768 ( .A1(n18656), .A2(n18635), .ZN(n18721) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18652), .B1(
        n18721), .B2(n18884), .ZN(n18636) );
  OAI211_X1 U21770 ( .C1(n18855), .C2(n18655), .A(n18637), .B(n18636), .ZN(
        P3_U2908) );
  AOI22_X1 U21771 ( .A1(n18890), .A2(n18651), .B1(n18889), .B2(n18648), .ZN(
        n18639) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18652), .B1(
        n18671), .B2(n18891), .ZN(n18638) );
  OAI211_X1 U21773 ( .C1(n18715), .C2(n18894), .A(n18639), .B(n18638), .ZN(
        P3_U2909) );
  AOI22_X1 U21774 ( .A1(n18671), .A2(n18897), .B1(n18895), .B2(n18651), .ZN(
        n18641) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18652), .B1(
        n18721), .B2(n18803), .ZN(n18640) );
  OAI211_X1 U21776 ( .C1(n18806), .C2(n18655), .A(n18641), .B(n18640), .ZN(
        P3_U2910) );
  AOI22_X1 U21777 ( .A1(n18902), .A2(n18651), .B1(n18901), .B2(n18648), .ZN(
        n18643) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18652), .B1(
        n18671), .B2(n18903), .ZN(n18642) );
  OAI211_X1 U21779 ( .C1(n18715), .C2(n18906), .A(n18643), .B(n18642), .ZN(
        P3_U2911) );
  AOI22_X1 U21780 ( .A1(n18671), .A2(n18908), .B1(n18907), .B2(n18651), .ZN(
        n18645) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18652), .B1(
        n18721), .B2(n18909), .ZN(n18644) );
  OAI211_X1 U21782 ( .C1(n18912), .C2(n18655), .A(n18645), .B(n18644), .ZN(
        P3_U2912) );
  AOI22_X1 U21783 ( .A1(n18915), .A2(n18648), .B1(n18913), .B2(n18651), .ZN(
        n18647) );
  AOI22_X1 U21784 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18652), .B1(
        n18671), .B2(n18914), .ZN(n18646) );
  OAI211_X1 U21785 ( .C1(n18715), .C2(n18918), .A(n18647), .B(n18646), .ZN(
        P3_U2913) );
  AOI22_X1 U21786 ( .A1(n18922), .A2(n18648), .B1(n18919), .B2(n18651), .ZN(
        n18650) );
  AOI22_X1 U21787 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18652), .B1(
        n18671), .B2(n18920), .ZN(n18649) );
  OAI211_X1 U21788 ( .C1(n18715), .C2(n18926), .A(n18650), .B(n18649), .ZN(
        P3_U2914) );
  AOI22_X1 U21789 ( .A1(n18671), .A2(n18930), .B1(n18928), .B2(n18651), .ZN(
        n18654) );
  AOI22_X1 U21790 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18652), .B1(
        n18721), .B2(n18932), .ZN(n18653) );
  OAI211_X1 U21791 ( .C1(n18937), .C2(n18655), .A(n18654), .B(n18653), .ZN(
        P3_U2915) );
  NOR2_X2 U21792 ( .A1(n18749), .A2(n18656), .ZN(n18741) );
  INV_X1 U21793 ( .A(n18741), .ZN(n18748) );
  AOI21_X1 U21794 ( .B1(n18748), .B2(n18715), .A(n18844), .ZN(n18674) );
  AOI22_X1 U21795 ( .A1(n18694), .A2(n18845), .B1(n18878), .B2(n18674), .ZN(
        n18660) );
  AOI221_X1 U21796 ( .B1(n18657), .B2(n18715), .C1(n18847), .C2(n18715), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18658) );
  OAI21_X1 U21797 ( .B1(n18741), .B2(n18658), .A(n18850), .ZN(n18675) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18675), .B1(
        n18741), .B2(n18884), .ZN(n18659) );
  OAI211_X1 U21799 ( .C1(n18678), .C2(n18855), .A(n18660), .B(n18659), .ZN(
        P3_U2916) );
  AOI22_X1 U21800 ( .A1(n18671), .A2(n18889), .B1(n18674), .B2(n18890), .ZN(
        n18662) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18675), .B1(
        n18694), .B2(n18891), .ZN(n18661) );
  OAI211_X1 U21802 ( .C1(n18748), .C2(n18894), .A(n18662), .B(n18661), .ZN(
        P3_U2917) );
  AOI22_X1 U21803 ( .A1(n18694), .A2(n18897), .B1(n18674), .B2(n18895), .ZN(
        n18664) );
  AOI22_X1 U21804 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18675), .B1(
        n18741), .B2(n18803), .ZN(n18663) );
  OAI211_X1 U21805 ( .C1(n18678), .C2(n18806), .A(n18664), .B(n18663), .ZN(
        P3_U2918) );
  AOI22_X1 U21806 ( .A1(n18671), .A2(n18901), .B1(n18674), .B2(n18902), .ZN(
        n18666) );
  AOI22_X1 U21807 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18675), .B1(
        n18694), .B2(n18903), .ZN(n18665) );
  OAI211_X1 U21808 ( .C1(n18748), .C2(n18906), .A(n18666), .B(n18665), .ZN(
        P3_U2919) );
  AOI22_X1 U21809 ( .A1(n18694), .A2(n18908), .B1(n18674), .B2(n18907), .ZN(
        n18668) );
  AOI22_X1 U21810 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18675), .B1(
        n18741), .B2(n18909), .ZN(n18667) );
  OAI211_X1 U21811 ( .C1(n18678), .C2(n18912), .A(n18668), .B(n18667), .ZN(
        P3_U2920) );
  AOI22_X1 U21812 ( .A1(n18671), .A2(n18915), .B1(n18674), .B2(n18913), .ZN(
        n18670) );
  AOI22_X1 U21813 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18675), .B1(
        n18694), .B2(n18914), .ZN(n18669) );
  OAI211_X1 U21814 ( .C1(n18748), .C2(n18918), .A(n18670), .B(n18669), .ZN(
        P3_U2921) );
  AOI22_X1 U21815 ( .A1(n18671), .A2(n18922), .B1(n18674), .B2(n18919), .ZN(
        n18673) );
  AOI22_X1 U21816 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18675), .B1(
        n18694), .B2(n18920), .ZN(n18672) );
  OAI211_X1 U21817 ( .C1(n18748), .C2(n18926), .A(n18673), .B(n18672), .ZN(
        P3_U2922) );
  AOI22_X1 U21818 ( .A1(n18694), .A2(n18930), .B1(n18674), .B2(n18928), .ZN(
        n18677) );
  AOI22_X1 U21819 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18675), .B1(
        n18741), .B2(n18932), .ZN(n18676) );
  OAI211_X1 U21820 ( .C1(n18678), .C2(n18937), .A(n18677), .B(n18676), .ZN(
        P3_U2923) );
  NOR2_X1 U21821 ( .A1(n18679), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18727) );
  AND2_X1 U21822 ( .A1(n19006), .A2(n18727), .ZN(n18697) );
  AOI22_X1 U21823 ( .A1(n18721), .A2(n18845), .B1(n18878), .B2(n18697), .ZN(
        n18683) );
  NAND2_X1 U21824 ( .A1(n18681), .A2(n18680), .ZN(n18698) );
  NAND2_X1 U21825 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18727), .ZN(
        n18771) );
  INV_X1 U21826 ( .A(n18771), .ZN(n18764) );
  AOI22_X1 U21827 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18698), .B1(
        n18884), .B2(n18764), .ZN(n18682) );
  OAI211_X1 U21828 ( .C1(n18701), .C2(n18855), .A(n18683), .B(n18682), .ZN(
        P3_U2924) );
  AOI22_X1 U21829 ( .A1(n18694), .A2(n18889), .B1(n18890), .B2(n18697), .ZN(
        n18685) );
  AOI22_X1 U21830 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18698), .B1(
        n18721), .B2(n18891), .ZN(n18684) );
  OAI211_X1 U21831 ( .C1(n18894), .C2(n18771), .A(n18685), .B(n18684), .ZN(
        P3_U2925) );
  AOI22_X1 U21832 ( .A1(n18721), .A2(n18897), .B1(n18895), .B2(n18697), .ZN(
        n18687) );
  AOI22_X1 U21833 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18698), .B1(
        n18803), .B2(n18764), .ZN(n18686) );
  OAI211_X1 U21834 ( .C1(n18701), .C2(n18806), .A(n18687), .B(n18686), .ZN(
        P3_U2926) );
  AOI22_X1 U21835 ( .A1(n18694), .A2(n18901), .B1(n18902), .B2(n18697), .ZN(
        n18689) );
  AOI22_X1 U21836 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18698), .B1(
        n18721), .B2(n18903), .ZN(n18688) );
  OAI211_X1 U21837 ( .C1(n18906), .C2(n18771), .A(n18689), .B(n18688), .ZN(
        P3_U2927) );
  AOI22_X1 U21838 ( .A1(n18721), .A2(n18908), .B1(n18907), .B2(n18697), .ZN(
        n18691) );
  AOI22_X1 U21839 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18698), .B1(
        n18909), .B2(n18764), .ZN(n18690) );
  OAI211_X1 U21840 ( .C1(n18701), .C2(n18912), .A(n18691), .B(n18690), .ZN(
        P3_U2928) );
  AOI22_X1 U21841 ( .A1(n18721), .A2(n18914), .B1(n18913), .B2(n18697), .ZN(
        n18693) );
  AOI22_X1 U21842 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18698), .B1(
        n18694), .B2(n18915), .ZN(n18692) );
  OAI211_X1 U21843 ( .C1(n18918), .C2(n18771), .A(n18693), .B(n18692), .ZN(
        P3_U2929) );
  AOI22_X1 U21844 ( .A1(n18694), .A2(n18922), .B1(n18919), .B2(n18697), .ZN(
        n18696) );
  AOI22_X1 U21845 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18698), .B1(
        n18721), .B2(n18920), .ZN(n18695) );
  OAI211_X1 U21846 ( .C1(n18926), .C2(n18771), .A(n18696), .B(n18695), .ZN(
        P3_U2930) );
  AOI22_X1 U21847 ( .A1(n18721), .A2(n18930), .B1(n18928), .B2(n18697), .ZN(
        n18700) );
  AOI22_X1 U21848 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18698), .B1(
        n18932), .B2(n18764), .ZN(n18699) );
  OAI211_X1 U21849 ( .C1(n18701), .C2(n18937), .A(n18700), .B(n18699), .ZN(
        P3_U2931) );
  NAND2_X1 U21850 ( .A1(n18972), .A2(n18794), .ZN(n18784) );
  NAND2_X1 U21851 ( .A1(n18771), .A2(n18784), .ZN(n18704) );
  INV_X1 U21852 ( .A(n18704), .ZN(n18750) );
  NOR2_X1 U21853 ( .A1(n18844), .A2(n18750), .ZN(n18720) );
  AOI22_X1 U21854 ( .A1(n18741), .A2(n18845), .B1(n18878), .B2(n18720), .ZN(
        n18706) );
  NAND2_X1 U21855 ( .A1(n18748), .A2(n18715), .ZN(n18703) );
  OAI221_X1 U21856 ( .B1(n18704), .B2(n18795), .C1(n18704), .C2(n18703), .A(
        n18702), .ZN(n18722) );
  INV_X1 U21857 ( .A(n18784), .ZN(n18790) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18722), .B1(
        n18884), .B2(n18790), .ZN(n18705) );
  OAI211_X1 U21859 ( .C1(n18715), .C2(n18855), .A(n18706), .B(n18705), .ZN(
        P3_U2932) );
  AOI22_X1 U21860 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18722), .B1(
        n18890), .B2(n18720), .ZN(n18708) );
  AOI22_X1 U21861 ( .A1(n18741), .A2(n18891), .B1(n18721), .B2(n18889), .ZN(
        n18707) );
  OAI211_X1 U21862 ( .C1(n18894), .C2(n18784), .A(n18708), .B(n18707), .ZN(
        P3_U2933) );
  AOI22_X1 U21863 ( .A1(n18741), .A2(n18897), .B1(n18895), .B2(n18720), .ZN(
        n18710) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18722), .B1(
        n18803), .B2(n18790), .ZN(n18709) );
  OAI211_X1 U21865 ( .C1(n18715), .C2(n18806), .A(n18710), .B(n18709), .ZN(
        P3_U2934) );
  AOI22_X1 U21866 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18722), .B1(
        n18902), .B2(n18720), .ZN(n18712) );
  AOI22_X1 U21867 ( .A1(n18741), .A2(n18903), .B1(n18721), .B2(n18901), .ZN(
        n18711) );
  OAI211_X1 U21868 ( .C1(n18906), .C2(n18784), .A(n18712), .B(n18711), .ZN(
        P3_U2935) );
  AOI22_X1 U21869 ( .A1(n18741), .A2(n18908), .B1(n18907), .B2(n18720), .ZN(
        n18714) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18722), .B1(
        n18909), .B2(n18790), .ZN(n18713) );
  OAI211_X1 U21871 ( .C1(n18715), .C2(n18912), .A(n18714), .B(n18713), .ZN(
        P3_U2936) );
  AOI22_X1 U21872 ( .A1(n18741), .A2(n18914), .B1(n18913), .B2(n18720), .ZN(
        n18717) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18722), .B1(
        n18721), .B2(n18915), .ZN(n18716) );
  OAI211_X1 U21874 ( .C1(n18918), .C2(n18784), .A(n18717), .B(n18716), .ZN(
        P3_U2937) );
  AOI22_X1 U21875 ( .A1(n18741), .A2(n18920), .B1(n18919), .B2(n18720), .ZN(
        n18719) );
  AOI22_X1 U21876 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18722), .B1(
        n18721), .B2(n18922), .ZN(n18718) );
  OAI211_X1 U21877 ( .C1(n18926), .C2(n18784), .A(n18719), .B(n18718), .ZN(
        P3_U2938) );
  AOI22_X1 U21878 ( .A1(n18721), .A2(n18872), .B1(n18928), .B2(n18720), .ZN(
        n18724) );
  AOI22_X1 U21879 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18722), .B1(
        n18741), .B2(n18930), .ZN(n18723) );
  OAI211_X1 U21880 ( .C1(n18877), .C2(n18784), .A(n18724), .B(n18723), .ZN(
        P3_U2939) );
  NOR2_X1 U21881 ( .A1(n18772), .A2(n18725), .ZN(n18744) );
  AOI22_X1 U21882 ( .A1(n18741), .A2(n18879), .B1(n18878), .B2(n18744), .ZN(
        n18730) );
  INV_X1 U21883 ( .A(n18726), .ZN(n18880) );
  NOR2_X1 U21884 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18772), .ZN(
        n18773) );
  AOI22_X1 U21885 ( .A1(n18883), .A2(n18727), .B1(n18880), .B2(n18773), .ZN(
        n18745) );
  NAND2_X1 U21886 ( .A1(n18728), .A2(n18794), .ZN(n18811) );
  INV_X1 U21887 ( .A(n18811), .ZN(n18817) );
  AOI22_X1 U21888 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18745), .B1(
        n18884), .B2(n18817), .ZN(n18729) );
  OAI211_X1 U21889 ( .C1(n18888), .C2(n18771), .A(n18730), .B(n18729), .ZN(
        P3_U2940) );
  AOI22_X1 U21890 ( .A1(n18741), .A2(n18889), .B1(n18890), .B2(n18744), .ZN(
        n18732) );
  AOI22_X1 U21891 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18745), .B1(
        n18891), .B2(n18764), .ZN(n18731) );
  OAI211_X1 U21892 ( .C1(n18894), .C2(n18811), .A(n18732), .B(n18731), .ZN(
        P3_U2941) );
  AOI22_X1 U21893 ( .A1(n18895), .A2(n18744), .B1(n18897), .B2(n18764), .ZN(
        n18734) );
  AOI22_X1 U21894 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18745), .B1(
        n18803), .B2(n18817), .ZN(n18733) );
  OAI211_X1 U21895 ( .C1(n18748), .C2(n18806), .A(n18734), .B(n18733), .ZN(
        P3_U2942) );
  AOI22_X1 U21896 ( .A1(n18741), .A2(n18901), .B1(n18902), .B2(n18744), .ZN(
        n18736) );
  AOI22_X1 U21897 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18745), .B1(
        n18903), .B2(n18764), .ZN(n18735) );
  OAI211_X1 U21898 ( .C1(n18906), .C2(n18811), .A(n18736), .B(n18735), .ZN(
        P3_U2943) );
  AOI22_X1 U21899 ( .A1(n18908), .A2(n18764), .B1(n18907), .B2(n18744), .ZN(
        n18738) );
  AOI22_X1 U21900 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18745), .B1(
        n18909), .B2(n18817), .ZN(n18737) );
  OAI211_X1 U21901 ( .C1(n18748), .C2(n18912), .A(n18738), .B(n18737), .ZN(
        P3_U2944) );
  AOI22_X1 U21902 ( .A1(n18914), .A2(n18764), .B1(n18913), .B2(n18744), .ZN(
        n18740) );
  AOI22_X1 U21903 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18745), .B1(
        n18741), .B2(n18915), .ZN(n18739) );
  OAI211_X1 U21904 ( .C1(n18918), .C2(n18811), .A(n18740), .B(n18739), .ZN(
        P3_U2945) );
  AOI22_X1 U21905 ( .A1(n18741), .A2(n18922), .B1(n18919), .B2(n18744), .ZN(
        n18743) );
  AOI22_X1 U21906 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18745), .B1(
        n18920), .B2(n18764), .ZN(n18742) );
  OAI211_X1 U21907 ( .C1(n18926), .C2(n18811), .A(n18743), .B(n18742), .ZN(
        P3_U2946) );
  AOI22_X1 U21908 ( .A1(n18930), .A2(n18764), .B1(n18928), .B2(n18744), .ZN(
        n18747) );
  AOI22_X1 U21909 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18745), .B1(
        n18932), .B2(n18817), .ZN(n18746) );
  OAI211_X1 U21910 ( .C1(n18748), .C2(n18937), .A(n18747), .B(n18746), .ZN(
        P3_U2947) );
  NOR2_X2 U21911 ( .A1(n18749), .A2(n18772), .ZN(n18835) );
  INV_X1 U21912 ( .A(n18835), .ZN(n18842) );
  AOI21_X1 U21913 ( .B1(n18811), .B2(n18842), .A(n18844), .ZN(n18767) );
  AOI22_X1 U21914 ( .A1(n18879), .A2(n18764), .B1(n18878), .B2(n18767), .ZN(
        n18753) );
  OAI211_X1 U21915 ( .C1(n18750), .C2(n18847), .A(n18811), .B(n18842), .ZN(
        n18751) );
  OAI211_X1 U21916 ( .C1(n18835), .C2(n19102), .A(n18850), .B(n18751), .ZN(
        n18768) );
  AOI22_X1 U21917 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18768), .B1(
        n18884), .B2(n18835), .ZN(n18752) );
  OAI211_X1 U21918 ( .C1(n18888), .C2(n18784), .A(n18753), .B(n18752), .ZN(
        P3_U2948) );
  AOI22_X1 U21919 ( .A1(n18890), .A2(n18767), .B1(n18889), .B2(n18764), .ZN(
        n18755) );
  AOI22_X1 U21920 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18768), .B1(
        n18891), .B2(n18790), .ZN(n18754) );
  OAI211_X1 U21921 ( .C1(n18894), .C2(n18842), .A(n18755), .B(n18754), .ZN(
        P3_U2949) );
  AOI22_X1 U21922 ( .A1(n18895), .A2(n18767), .B1(n18897), .B2(n18790), .ZN(
        n18757) );
  AOI22_X1 U21923 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18768), .B1(
        n18803), .B2(n18835), .ZN(n18756) );
  OAI211_X1 U21924 ( .C1(n18806), .C2(n18771), .A(n18757), .B(n18756), .ZN(
        P3_U2950) );
  AOI22_X1 U21925 ( .A1(n18902), .A2(n18767), .B1(n18901), .B2(n18764), .ZN(
        n18759) );
  AOI22_X1 U21926 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18768), .B1(
        n18903), .B2(n18790), .ZN(n18758) );
  OAI211_X1 U21927 ( .C1(n18906), .C2(n18842), .A(n18759), .B(n18758), .ZN(
        P3_U2951) );
  AOI22_X1 U21928 ( .A1(n18862), .A2(n18764), .B1(n18907), .B2(n18767), .ZN(
        n18761) );
  AOI22_X1 U21929 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18768), .B1(
        n18908), .B2(n18790), .ZN(n18760) );
  OAI211_X1 U21930 ( .C1(n18865), .C2(n18842), .A(n18761), .B(n18760), .ZN(
        P3_U2952) );
  AOI22_X1 U21931 ( .A1(n18914), .A2(n18790), .B1(n18913), .B2(n18767), .ZN(
        n18763) );
  AOI22_X1 U21932 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18768), .B1(
        n18915), .B2(n18764), .ZN(n18762) );
  OAI211_X1 U21933 ( .C1(n18918), .C2(n18842), .A(n18763), .B(n18762), .ZN(
        P3_U2953) );
  AOI22_X1 U21934 ( .A1(n18922), .A2(n18764), .B1(n18919), .B2(n18767), .ZN(
        n18766) );
  AOI22_X1 U21935 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18768), .B1(
        n18920), .B2(n18790), .ZN(n18765) );
  OAI211_X1 U21936 ( .C1(n18926), .C2(n18842), .A(n18766), .B(n18765), .ZN(
        P3_U2954) );
  AOI22_X1 U21937 ( .A1(n18930), .A2(n18790), .B1(n18928), .B2(n18767), .ZN(
        n18770) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18768), .B1(
        n18932), .B2(n18835), .ZN(n18769) );
  OAI211_X1 U21939 ( .C1(n18937), .C2(n18771), .A(n18770), .B(n18769), .ZN(
        P3_U2955) );
  NOR2_X1 U21940 ( .A1(n18969), .A2(n18772), .ZN(n18822) );
  AND2_X1 U21941 ( .A1(n19006), .A2(n18822), .ZN(n18789) );
  AOI22_X1 U21942 ( .A1(n18845), .A2(n18817), .B1(n18878), .B2(n18789), .ZN(
        n18775) );
  AOI22_X1 U21943 ( .A1(n18883), .A2(n18773), .B1(n18880), .B2(n18822), .ZN(
        n18791) );
  NAND2_X1 U21944 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18822), .ZN(
        n18854) );
  AOI22_X1 U21945 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18791), .B1(
        n18884), .B2(n18871), .ZN(n18774) );
  OAI211_X1 U21946 ( .C1(n18855), .C2(n18784), .A(n18775), .B(n18774), .ZN(
        P3_U2956) );
  AOI22_X1 U21947 ( .A1(n18891), .A2(n18817), .B1(n18890), .B2(n18789), .ZN(
        n18777) );
  AOI22_X1 U21948 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18791), .B1(
        n18889), .B2(n18790), .ZN(n18776) );
  OAI211_X1 U21949 ( .C1(n18894), .C2(n18854), .A(n18777), .B(n18776), .ZN(
        P3_U2957) );
  AOI22_X1 U21950 ( .A1(n18896), .A2(n18790), .B1(n18895), .B2(n18789), .ZN(
        n18779) );
  AOI22_X1 U21951 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18791), .B1(
        n18897), .B2(n18817), .ZN(n18778) );
  OAI211_X1 U21952 ( .C1(n18900), .C2(n18854), .A(n18779), .B(n18778), .ZN(
        P3_U2958) );
  AOI22_X1 U21953 ( .A1(n18903), .A2(n18817), .B1(n18902), .B2(n18789), .ZN(
        n18781) );
  AOI22_X1 U21954 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18791), .B1(
        n18901), .B2(n18790), .ZN(n18780) );
  OAI211_X1 U21955 ( .C1(n18906), .C2(n18854), .A(n18781), .B(n18780), .ZN(
        P3_U2959) );
  AOI22_X1 U21956 ( .A1(n18908), .A2(n18817), .B1(n18907), .B2(n18789), .ZN(
        n18783) );
  AOI22_X1 U21957 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18791), .B1(
        n18909), .B2(n18871), .ZN(n18782) );
  OAI211_X1 U21958 ( .C1(n18912), .C2(n18784), .A(n18783), .B(n18782), .ZN(
        P3_U2960) );
  AOI22_X1 U21959 ( .A1(n18914), .A2(n18817), .B1(n18913), .B2(n18789), .ZN(
        n18786) );
  AOI22_X1 U21960 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18791), .B1(
        n18915), .B2(n18790), .ZN(n18785) );
  OAI211_X1 U21961 ( .C1(n18918), .C2(n18854), .A(n18786), .B(n18785), .ZN(
        P3_U2961) );
  AOI22_X1 U21962 ( .A1(n18920), .A2(n18817), .B1(n18919), .B2(n18789), .ZN(
        n18788) );
  AOI22_X1 U21963 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18791), .B1(
        n18922), .B2(n18790), .ZN(n18787) );
  OAI211_X1 U21964 ( .C1(n18926), .C2(n18854), .A(n18788), .B(n18787), .ZN(
        P3_U2962) );
  AOI22_X1 U21965 ( .A1(n18872), .A2(n18790), .B1(n18928), .B2(n18789), .ZN(
        n18793) );
  AOI22_X1 U21966 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18791), .B1(
        n18930), .B2(n18817), .ZN(n18792) );
  OAI211_X1 U21967 ( .C1(n18877), .C2(n18854), .A(n18793), .B(n18792), .ZN(
        P3_U2963) );
  NAND2_X1 U21968 ( .A1(n18968), .A2(n18882), .ZN(n18936) );
  INV_X1 U21969 ( .A(n18936), .ZN(n18921) );
  NAND2_X1 U21970 ( .A1(n18795), .A2(n18794), .ZN(n18796) );
  NOR2_X1 U21971 ( .A1(n18871), .A2(n18921), .ZN(n18848) );
  OAI21_X1 U21972 ( .B1(n18797), .B2(n18796), .A(n18848), .ZN(n18798) );
  OAI211_X1 U21973 ( .C1(n18921), .C2(n19102), .A(n18850), .B(n18798), .ZN(
        n18818) );
  NOR2_X1 U21974 ( .A1(n18844), .A2(n18848), .ZN(n18816) );
  AOI22_X1 U21975 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18818), .B1(
        n18878), .B2(n18816), .ZN(n18800) );
  AOI22_X1 U21976 ( .A1(n18879), .A2(n18817), .B1(n18884), .B2(n18921), .ZN(
        n18799) );
  OAI211_X1 U21977 ( .C1(n18888), .C2(n18842), .A(n18800), .B(n18799), .ZN(
        P3_U2964) );
  AOI22_X1 U21978 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18818), .B1(
        n18890), .B2(n18816), .ZN(n18802) );
  AOI22_X1 U21979 ( .A1(n18891), .A2(n18835), .B1(n18889), .B2(n18817), .ZN(
        n18801) );
  OAI211_X1 U21980 ( .C1(n18894), .C2(n18936), .A(n18802), .B(n18801), .ZN(
        P3_U2965) );
  AOI22_X1 U21981 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18818), .B1(
        n18895), .B2(n18816), .ZN(n18805) );
  AOI22_X1 U21982 ( .A1(n18803), .A2(n18921), .B1(n18897), .B2(n18835), .ZN(
        n18804) );
  OAI211_X1 U21983 ( .C1(n18806), .C2(n18811), .A(n18805), .B(n18804), .ZN(
        P3_U2966) );
  AOI22_X1 U21984 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18818), .B1(
        n18902), .B2(n18816), .ZN(n18808) );
  AOI22_X1 U21985 ( .A1(n18903), .A2(n18835), .B1(n18901), .B2(n18817), .ZN(
        n18807) );
  OAI211_X1 U21986 ( .C1(n18906), .C2(n18936), .A(n18808), .B(n18807), .ZN(
        P3_U2967) );
  AOI22_X1 U21987 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18818), .B1(
        n18907), .B2(n18816), .ZN(n18810) );
  AOI22_X1 U21988 ( .A1(n18909), .A2(n18921), .B1(n18908), .B2(n18835), .ZN(
        n18809) );
  OAI211_X1 U21989 ( .C1(n18912), .C2(n18811), .A(n18810), .B(n18809), .ZN(
        P3_U2968) );
  AOI22_X1 U21990 ( .A1(n18914), .A2(n18835), .B1(n18913), .B2(n18816), .ZN(
        n18813) );
  AOI22_X1 U21991 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18818), .B1(
        n18915), .B2(n18817), .ZN(n18812) );
  OAI211_X1 U21992 ( .C1(n18918), .C2(n18936), .A(n18813), .B(n18812), .ZN(
        P3_U2969) );
  AOI22_X1 U21993 ( .A1(n18922), .A2(n18817), .B1(n18919), .B2(n18816), .ZN(
        n18815) );
  AOI22_X1 U21994 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18818), .B1(
        n18920), .B2(n18835), .ZN(n18814) );
  OAI211_X1 U21995 ( .C1(n18926), .C2(n18936), .A(n18815), .B(n18814), .ZN(
        P3_U2970) );
  AOI22_X1 U21996 ( .A1(n18872), .A2(n18817), .B1(n18928), .B2(n18816), .ZN(
        n18820) );
  AOI22_X1 U21997 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18818), .B1(
        n18930), .B2(n18835), .ZN(n18819) );
  OAI211_X1 U21998 ( .C1(n18877), .C2(n18936), .A(n18820), .B(n18819), .ZN(
        P3_U2971) );
  NOR2_X1 U21999 ( .A1(n18844), .A2(n18821), .ZN(n18838) );
  AOI22_X1 U22000 ( .A1(n18879), .A2(n18835), .B1(n18878), .B2(n18838), .ZN(
        n18824) );
  AOI22_X1 U22001 ( .A1(n18883), .A2(n18822), .B1(n18882), .B2(n18880), .ZN(
        n18839) );
  AOI22_X1 U22002 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18839), .B1(
        n18884), .B2(n18929), .ZN(n18823) );
  OAI211_X1 U22003 ( .C1(n18888), .C2(n18854), .A(n18824), .B(n18823), .ZN(
        P3_U2972) );
  AOI22_X1 U22004 ( .A1(n18890), .A2(n18838), .B1(n18889), .B2(n18835), .ZN(
        n18826) );
  AOI22_X1 U22005 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18839), .B1(
        n18891), .B2(n18871), .ZN(n18825) );
  OAI211_X1 U22006 ( .C1(n18894), .C2(n18887), .A(n18826), .B(n18825), .ZN(
        P3_U2973) );
  AOI22_X1 U22007 ( .A1(n18896), .A2(n18835), .B1(n18895), .B2(n18838), .ZN(
        n18828) );
  AOI22_X1 U22008 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18839), .B1(
        n18897), .B2(n18871), .ZN(n18827) );
  OAI211_X1 U22009 ( .C1(n18900), .C2(n18887), .A(n18828), .B(n18827), .ZN(
        P3_U2974) );
  AOI22_X1 U22010 ( .A1(n18903), .A2(n18871), .B1(n18902), .B2(n18838), .ZN(
        n18830) );
  AOI22_X1 U22011 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18839), .B1(
        n18901), .B2(n18835), .ZN(n18829) );
  OAI211_X1 U22012 ( .C1(n18906), .C2(n18887), .A(n18830), .B(n18829), .ZN(
        P3_U2975) );
  AOI22_X1 U22013 ( .A1(n18862), .A2(n18835), .B1(n18907), .B2(n18838), .ZN(
        n18832) );
  AOI22_X1 U22014 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18839), .B1(
        n18908), .B2(n18871), .ZN(n18831) );
  OAI211_X1 U22015 ( .C1(n18865), .C2(n18887), .A(n18832), .B(n18831), .ZN(
        P3_U2976) );
  AOI22_X1 U22016 ( .A1(n18914), .A2(n18871), .B1(n18913), .B2(n18838), .ZN(
        n18834) );
  AOI22_X1 U22017 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18839), .B1(
        n18915), .B2(n18835), .ZN(n18833) );
  OAI211_X1 U22018 ( .C1(n18918), .C2(n18887), .A(n18834), .B(n18833), .ZN(
        P3_U2977) );
  AOI22_X1 U22019 ( .A1(n18920), .A2(n18871), .B1(n18919), .B2(n18838), .ZN(
        n18837) );
  AOI22_X1 U22020 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18839), .B1(
        n18922), .B2(n18835), .ZN(n18836) );
  OAI211_X1 U22021 ( .C1(n18926), .C2(n18887), .A(n18837), .B(n18836), .ZN(
        P3_U2978) );
  AOI22_X1 U22022 ( .A1(n18930), .A2(n18871), .B1(n18928), .B2(n18838), .ZN(
        n18841) );
  AOI22_X1 U22023 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18839), .B1(
        n18932), .B2(n18929), .ZN(n18840) );
  OAI211_X1 U22024 ( .C1(n18937), .C2(n18842), .A(n18841), .B(n18840), .ZN(
        P3_U2979) );
  INV_X1 U22025 ( .A(n18843), .ZN(n18846) );
  NOR2_X1 U22026 ( .A1(n18844), .A2(n18846), .ZN(n18870) );
  AOI22_X1 U22027 ( .A1(n18845), .A2(n18921), .B1(n18878), .B2(n18870), .ZN(
        n18853) );
  OAI21_X1 U22028 ( .B1(n18848), .B2(n18847), .A(n18846), .ZN(n18849) );
  OAI211_X1 U22029 ( .C1(n18851), .C2(n19102), .A(n18850), .B(n18849), .ZN(
        n18873) );
  AOI22_X1 U22030 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18873), .B1(
        n18884), .B2(n18851), .ZN(n18852) );
  OAI211_X1 U22031 ( .C1(n18855), .C2(n18854), .A(n18853), .B(n18852), .ZN(
        P3_U2980) );
  AOI22_X1 U22032 ( .A1(n18890), .A2(n18870), .B1(n18889), .B2(n18871), .ZN(
        n18857) );
  AOI22_X1 U22033 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18873), .B1(
        n18891), .B2(n18921), .ZN(n18856) );
  OAI211_X1 U22034 ( .C1(n18894), .C2(n18876), .A(n18857), .B(n18856), .ZN(
        P3_U2981) );
  AOI22_X1 U22035 ( .A1(n18896), .A2(n18871), .B1(n18895), .B2(n18870), .ZN(
        n18859) );
  AOI22_X1 U22036 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18873), .B1(
        n18897), .B2(n18921), .ZN(n18858) );
  OAI211_X1 U22037 ( .C1(n18900), .C2(n18876), .A(n18859), .B(n18858), .ZN(
        P3_U2982) );
  AOI22_X1 U22038 ( .A1(n18902), .A2(n18870), .B1(n18901), .B2(n18871), .ZN(
        n18861) );
  AOI22_X1 U22039 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18873), .B1(
        n18903), .B2(n18921), .ZN(n18860) );
  OAI211_X1 U22040 ( .C1(n18906), .C2(n18876), .A(n18861), .B(n18860), .ZN(
        P3_U2983) );
  AOI22_X1 U22041 ( .A1(n18862), .A2(n18871), .B1(n18907), .B2(n18870), .ZN(
        n18864) );
  AOI22_X1 U22042 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18873), .B1(
        n18908), .B2(n18921), .ZN(n18863) );
  OAI211_X1 U22043 ( .C1(n18865), .C2(n18876), .A(n18864), .B(n18863), .ZN(
        P3_U2984) );
  AOI22_X1 U22044 ( .A1(n18914), .A2(n18921), .B1(n18913), .B2(n18870), .ZN(
        n18867) );
  AOI22_X1 U22045 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18873), .B1(
        n18915), .B2(n18871), .ZN(n18866) );
  OAI211_X1 U22046 ( .C1(n18918), .C2(n18876), .A(n18867), .B(n18866), .ZN(
        P3_U2985) );
  AOI22_X1 U22047 ( .A1(n18922), .A2(n18871), .B1(n18919), .B2(n18870), .ZN(
        n18869) );
  AOI22_X1 U22048 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18873), .B1(
        n18920), .B2(n18921), .ZN(n18868) );
  OAI211_X1 U22049 ( .C1(n18926), .C2(n18876), .A(n18869), .B(n18868), .ZN(
        P3_U2986) );
  AOI22_X1 U22050 ( .A1(n18872), .A2(n18871), .B1(n18928), .B2(n18870), .ZN(
        n18875) );
  AOI22_X1 U22051 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18873), .B1(
        n18930), .B2(n18921), .ZN(n18874) );
  OAI211_X1 U22052 ( .C1(n18877), .C2(n18876), .A(n18875), .B(n18874), .ZN(
        P3_U2987) );
  AND2_X1 U22053 ( .A1(n19006), .A2(n18881), .ZN(n18927) );
  AOI22_X1 U22054 ( .A1(n18879), .A2(n18921), .B1(n18878), .B2(n18927), .ZN(
        n18886) );
  AOI22_X1 U22055 ( .A1(n18883), .A2(n18882), .B1(n18881), .B2(n18880), .ZN(
        n18933) );
  AOI22_X1 U22056 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18933), .B1(
        n18884), .B2(n18931), .ZN(n18885) );
  OAI211_X1 U22057 ( .C1(n18888), .C2(n18887), .A(n18886), .B(n18885), .ZN(
        P3_U2988) );
  AOI22_X1 U22058 ( .A1(n18890), .A2(n18927), .B1(n18889), .B2(n18921), .ZN(
        n18893) );
  AOI22_X1 U22059 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18933), .B1(
        n18891), .B2(n18929), .ZN(n18892) );
  OAI211_X1 U22060 ( .C1(n18894), .C2(n18925), .A(n18893), .B(n18892), .ZN(
        P3_U2989) );
  AOI22_X1 U22061 ( .A1(n18896), .A2(n18921), .B1(n18895), .B2(n18927), .ZN(
        n18899) );
  AOI22_X1 U22062 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18933), .B1(
        n18897), .B2(n18929), .ZN(n18898) );
  OAI211_X1 U22063 ( .C1(n18900), .C2(n18925), .A(n18899), .B(n18898), .ZN(
        P3_U2990) );
  AOI22_X1 U22064 ( .A1(n18902), .A2(n18927), .B1(n18901), .B2(n18921), .ZN(
        n18905) );
  AOI22_X1 U22065 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18933), .B1(
        n18903), .B2(n18929), .ZN(n18904) );
  OAI211_X1 U22066 ( .C1(n18906), .C2(n18925), .A(n18905), .B(n18904), .ZN(
        P3_U2991) );
  AOI22_X1 U22067 ( .A1(n18908), .A2(n18929), .B1(n18907), .B2(n18927), .ZN(
        n18911) );
  AOI22_X1 U22068 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18933), .B1(
        n18909), .B2(n18931), .ZN(n18910) );
  OAI211_X1 U22069 ( .C1(n18912), .C2(n18936), .A(n18911), .B(n18910), .ZN(
        P3_U2992) );
  AOI22_X1 U22070 ( .A1(n18914), .A2(n18929), .B1(n18913), .B2(n18927), .ZN(
        n18917) );
  AOI22_X1 U22071 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18933), .B1(
        n18915), .B2(n18921), .ZN(n18916) );
  OAI211_X1 U22072 ( .C1(n18918), .C2(n18925), .A(n18917), .B(n18916), .ZN(
        P3_U2993) );
  AOI22_X1 U22073 ( .A1(n18920), .A2(n18929), .B1(n18919), .B2(n18927), .ZN(
        n18924) );
  AOI22_X1 U22074 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18933), .B1(
        n18922), .B2(n18921), .ZN(n18923) );
  OAI211_X1 U22075 ( .C1(n18926), .C2(n18925), .A(n18924), .B(n18923), .ZN(
        P3_U2994) );
  AOI22_X1 U22076 ( .A1(n18930), .A2(n18929), .B1(n18928), .B2(n18927), .ZN(
        n18935) );
  AOI22_X1 U22077 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18933), .B1(
        n18932), .B2(n18931), .ZN(n18934) );
  OAI211_X1 U22078 ( .C1(n18937), .C2(n18936), .A(n18935), .B(n18934), .ZN(
        P3_U2995) );
  AND2_X1 U22079 ( .A1(n18939), .A2(n18938), .ZN(n18940) );
  OAI22_X1 U22080 ( .A1(n18943), .A2(n18942), .B1(n18941), .B2(n18940), .ZN(
        n18944) );
  AOI221_X1 U22081 ( .B1(n18958), .B2(n18946), .C1(n9866), .C2(n18946), .A(
        n18944), .ZN(n19143) );
  AOI211_X1 U22082 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18983), .A(
        n18948), .B(n18947), .ZN(n18994) );
  AOI21_X1 U22083 ( .B1(n18950), .B2(n18949), .A(n18957), .ZN(n18963) );
  OAI21_X1 U22084 ( .B1(n18953), .B2(n18952), .A(n18951), .ZN(n18977) );
  INV_X1 U22085 ( .A(n18977), .ZN(n18955) );
  NAND2_X1 U22086 ( .A1(n13017), .A2(n18976), .ZN(n18959) );
  OAI211_X1 U22087 ( .C1(n18955), .C2(n18954), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n18959), .ZN(n18962) );
  OAI21_X1 U22088 ( .B1(n19128), .B2(n18956), .A(n18975), .ZN(n18974) );
  AOI22_X1 U22089 ( .A1(n18959), .A2(n18958), .B1(n18974), .B2(n18957), .ZN(
        n18960) );
  INV_X1 U22090 ( .A(n18960), .ZN(n18961) );
  OAI22_X1 U22091 ( .A1(n18963), .A2(n18962), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18961), .ZN(n19104) );
  INV_X1 U22092 ( .A(n18983), .ZN(n18982) );
  AOI22_X1 U22093 ( .A1(n18983), .A2(n19108), .B1(n19104), .B2(n18982), .ZN(
        n18990) );
  OR2_X1 U22094 ( .A1(n18965), .A2(n18964), .ZN(n18966) );
  AOI22_X1 U22095 ( .A1(n19118), .A2(n18966), .B1(n19121), .B2(n18974), .ZN(
        n19115) );
  AOI22_X1 U22096 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18967), .B1(
        n18966), .B2(n19128), .ZN(n18970) );
  INV_X1 U22097 ( .A(n18970), .ZN(n19123) );
  NOR3_X1 U22098 ( .A1(n18969), .A2(n18968), .A3(n19123), .ZN(n18971) );
  OAI22_X1 U22099 ( .A1(n19115), .A2(n18971), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18970), .ZN(n18973) );
  AOI21_X1 U22100 ( .B1(n18973), .B2(n18982), .A(n18972), .ZN(n18985) );
  NAND3_X1 U22101 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n13017), .A3(
        n18974), .ZN(n18980) );
  NOR2_X1 U22102 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18975), .ZN(
        n18978) );
  OAI211_X1 U22103 ( .C1(n18978), .C2(n18977), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18976), .ZN(n18979) );
  OAI211_X1 U22104 ( .C1(n19111), .C2(n18981), .A(n18980), .B(n18979), .ZN(
        n19113) );
  AOI22_X1 U22105 ( .A1(n18983), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19113), .B2(n18982), .ZN(n18986) );
  OR2_X1 U22106 ( .A1(n18986), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18984) );
  AOI221_X1 U22107 ( .B1(n18985), .B2(n18984), .C1(n18986), .C2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18989) );
  OAI21_X1 U22108 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18986), .ZN(n18988) );
  AOI222_X1 U22109 ( .A1(n18990), .A2(n18989), .B1(n18990), .B2(n18988), .C1(
        n18989), .C2(n18987), .ZN(n18993) );
  OAI21_X1 U22110 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18991), .ZN(n18992) );
  NAND4_X1 U22111 ( .A1(n19143), .A2(n18994), .A3(n18993), .A4(n18992), .ZN(
        n19001) );
  AOI211_X1 U22112 ( .C1(n18996), .C2(n18995), .A(n19149), .B(n19001), .ZN(
        n19100) );
  AOI21_X1 U22113 ( .B1(n19146), .B2(n19005), .A(n19100), .ZN(n19007) );
  NOR2_X1 U22114 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19156) );
  NAND2_X1 U22115 ( .A1(n19146), .A2(n18997), .ZN(n19010) );
  INV_X1 U22116 ( .A(n19010), .ZN(n18998) );
  AOI211_X1 U22117 ( .C1(n19122), .C2(n19156), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18998), .ZN(n18999) );
  AOI211_X1 U22118 ( .C1(n19002), .C2(n19001), .A(n19000), .B(n18999), .ZN(
        n19003) );
  OAI221_X1 U22119 ( .B1(n19099), .B2(n19007), .C1(n19099), .C2(n19004), .A(
        n19003), .ZN(P3_U2996) );
  NAND3_X1 U22120 ( .A1(n19146), .A2(n19012), .A3(n19005), .ZN(n19015) );
  NAND3_X1 U22121 ( .A1(n19008), .A2(n19007), .A3(n19006), .ZN(n19009) );
  NAND4_X1 U22122 ( .A1(n19011), .A2(n19010), .A3(n19015), .A4(n19009), .ZN(
        P3_U2997) );
  OR3_X1 U22123 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19013), .A3(n19012), 
        .ZN(n19014) );
  AND3_X1 U22124 ( .A1(n19015), .A2(n19101), .A3(n19014), .ZN(P3_U2998) );
  AND2_X1 U22125 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(
        P3_U2999) );
  AND2_X1 U22126 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(
        P3_U3000) );
  AND2_X1 U22127 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(
        P3_U3001) );
  AND2_X1 U22128 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_28__SCAN_IN), .ZN(
        P3_U3002) );
  AND2_X1 U22129 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(
        P3_U3003) );
  AND2_X1 U22130 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(
        P3_U3004) );
  AND2_X1 U22131 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(
        P3_U3005) );
  AND2_X1 U22132 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(
        P3_U3006) );
  AND2_X1 U22133 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(
        P3_U3007) );
  AND2_X1 U22134 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(
        P3_U3008) );
  AND2_X1 U22135 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(
        P3_U3009) );
  AND2_X1 U22136 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(
        P3_U3010) );
  AND2_X1 U22137 ( .A1(n19016), .A2(P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(
        P3_U3011) );
  AND2_X1 U22138 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(
        P3_U3012) );
  AND2_X1 U22139 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(
        P3_U3013) );
  AND2_X1 U22140 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(
        P3_U3014) );
  AND2_X1 U22141 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(
        P3_U3015) );
  AND2_X1 U22142 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(
        P3_U3016) );
  AND2_X1 U22143 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(
        P3_U3017) );
  AND2_X1 U22144 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(
        P3_U3019) );
  AND2_X1 U22145 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(
        P3_U3020) );
  AND2_X1 U22146 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(P3_U3021) );
  AND2_X1 U22147 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(P3_U3022) );
  AND2_X1 U22148 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(P3_U3023) );
  AND2_X1 U22149 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(P3_U3024) );
  INV_X1 U22150 ( .A(P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n21339) );
  NOR2_X1 U22151 ( .A1(n19097), .A2(n21339), .ZN(P3_U3025) );
  AND2_X1 U22152 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(P3_U3026) );
  AND2_X1 U22153 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(P3_U3027) );
  AND2_X1 U22154 ( .A1(n21240), .A2(P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(P3_U3028) );
  AOI221_X1 U22155 ( .B1(n19017), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20118), .C2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n19140), .ZN(n19020)
         );
  NAND2_X1 U22156 ( .A1(n19146), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19029) );
  INV_X1 U22157 ( .A(n19029), .ZN(n19025) );
  NOR2_X1 U22158 ( .A1(n19025), .A2(n21390), .ZN(n19019) );
  INV_X1 U22159 ( .A(NA), .ZN(n21130) );
  INV_X1 U22160 ( .A(n19018), .ZN(n19021) );
  OAI22_X1 U22161 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n19019), .B1(n21130), 
        .B2(n19021), .ZN(n19032) );
  OR2_X1 U22162 ( .A1(n19020), .A2(n19032), .ZN(P3_U3029) );
  NAND3_X1 U22163 ( .A1(n19034), .A2(P3_STATE_REG_1__SCAN_IN), .A3(HOLD), .ZN(
        n19024) );
  OAI211_X1 U22164 ( .C1(n19022), .C2(n20118), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .B(n19021), .ZN(n19023) );
  AND2_X1 U22165 ( .A1(n19024), .A2(n19023), .ZN(n19028) );
  NOR2_X1 U22166 ( .A1(n19026), .A2(n19025), .ZN(n19033) );
  AOI22_X1 U22167 ( .A1(n19028), .A2(n19033), .B1(n19027), .B2(n19153), .ZN(
        P3_U3030) );
  OAI222_X1 U22168 ( .A1(n20118), .A2(n19034), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n19029), .C2(NA), .ZN(n19030)
         );
  OAI211_X1 U22169 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n19030), .ZN(n19031) );
  OAI21_X1 U22170 ( .B1(n19033), .B2(n19032), .A(n19031), .ZN(P3_U3031) );
  OAI222_X1 U22171 ( .A1(n19083), .A2(n21516), .B1(n19035), .B2(n19140), .C1(
        n19130), .C2(n19090), .ZN(P3_U3032) );
  OAI222_X1 U22172 ( .A1(n19083), .A2(n19037), .B1(n19036), .B2(n19140), .C1(
        n21516), .C2(n19090), .ZN(P3_U3033) );
  OAI222_X1 U22173 ( .A1(n19083), .A2(n19039), .B1(n19038), .B2(n19140), .C1(
        n19037), .C2(n19090), .ZN(P3_U3034) );
  OAI222_X1 U22174 ( .A1(n19083), .A2(n19041), .B1(n19040), .B2(n19140), .C1(
        n19039), .C2(n19090), .ZN(P3_U3035) );
  OAI222_X1 U22175 ( .A1(n19083), .A2(n19043), .B1(n19042), .B2(n19140), .C1(
        n19041), .C2(n19090), .ZN(P3_U3036) );
  OAI222_X1 U22176 ( .A1(n19083), .A2(n19045), .B1(n19044), .B2(n19140), .C1(
        n19043), .C2(n19090), .ZN(P3_U3037) );
  OAI222_X1 U22177 ( .A1(n19083), .A2(n19048), .B1(n19046), .B2(n19140), .C1(
        n19045), .C2(n19090), .ZN(P3_U3038) );
  OAI222_X1 U22178 ( .A1(n19048), .A2(n19090), .B1(n19047), .B2(n19140), .C1(
        n19049), .C2(n19083), .ZN(P3_U3039) );
  OAI222_X1 U22179 ( .A1(n19083), .A2(n19050), .B1(n21503), .B2(n19140), .C1(
        n19049), .C2(n19090), .ZN(P3_U3040) );
  OAI222_X1 U22180 ( .A1(n19083), .A2(n19052), .B1(n19051), .B2(n19140), .C1(
        n19050), .C2(n19090), .ZN(P3_U3041) );
  OAI222_X1 U22181 ( .A1(n19083), .A2(n19054), .B1(n19053), .B2(n19140), .C1(
        n19052), .C2(n19090), .ZN(P3_U3042) );
  OAI222_X1 U22182 ( .A1(n19083), .A2(n19056), .B1(n19055), .B2(n19140), .C1(
        n19054), .C2(n19090), .ZN(P3_U3043) );
  OAI222_X1 U22183 ( .A1(n19083), .A2(n19059), .B1(n19057), .B2(n19140), .C1(
        n19056), .C2(n19090), .ZN(P3_U3044) );
  OAI222_X1 U22184 ( .A1(n19059), .A2(n19090), .B1(n19058), .B2(n19140), .C1(
        n19060), .C2(n19083), .ZN(P3_U3045) );
  OAI222_X1 U22185 ( .A1(n19083), .A2(n19062), .B1(n19061), .B2(n19140), .C1(
        n19060), .C2(n19090), .ZN(P3_U3046) );
  OAI222_X1 U22186 ( .A1(n19083), .A2(n19064), .B1(n21485), .B2(n19140), .C1(
        n19062), .C2(n19090), .ZN(P3_U3047) );
  OAI222_X1 U22187 ( .A1(n19064), .A2(n19090), .B1(n19063), .B2(n19140), .C1(
        n19065), .C2(n19083), .ZN(P3_U3048) );
  OAI222_X1 U22188 ( .A1(n19083), .A2(n21473), .B1(n19066), .B2(n19140), .C1(
        n19065), .C2(n19090), .ZN(P3_U3049) );
  OAI222_X1 U22189 ( .A1(n21473), .A2(n19090), .B1(n19067), .B2(n19140), .C1(
        n19068), .C2(n19083), .ZN(P3_U3050) );
  OAI222_X1 U22190 ( .A1(n19083), .A2(n19071), .B1(n19069), .B2(n19140), .C1(
        n19068), .C2(n19090), .ZN(P3_U3051) );
  OAI222_X1 U22191 ( .A1(n19071), .A2(n19090), .B1(n19070), .B2(n19140), .C1(
        n19072), .C2(n19083), .ZN(P3_U3052) );
  OAI222_X1 U22192 ( .A1(n19083), .A2(n19075), .B1(n19073), .B2(n19140), .C1(
        n19072), .C2(n19090), .ZN(P3_U3053) );
  OAI222_X1 U22193 ( .A1(n19075), .A2(n19090), .B1(n19074), .B2(n19140), .C1(
        n19076), .C2(n19083), .ZN(P3_U3054) );
  OAI222_X1 U22194 ( .A1(n19083), .A2(n19078), .B1(n19077), .B2(n19140), .C1(
        n19076), .C2(n19090), .ZN(P3_U3055) );
  OAI222_X1 U22195 ( .A1(n19083), .A2(n21427), .B1(n19079), .B2(n19140), .C1(
        n19078), .C2(n19090), .ZN(P3_U3056) );
  OAI222_X1 U22196 ( .A1(n19083), .A2(n19081), .B1(n19080), .B2(n19140), .C1(
        n21427), .C2(n19090), .ZN(P3_U3057) );
  OAI222_X1 U22197 ( .A1(n19083), .A2(n19084), .B1(n19082), .B2(n19140), .C1(
        n19081), .C2(n19090), .ZN(P3_U3058) );
  OAI222_X1 U22198 ( .A1(n19083), .A2(n19086), .B1(n19085), .B2(n19140), .C1(
        n19084), .C2(n19090), .ZN(P3_U3059) );
  OAI222_X1 U22199 ( .A1(n19083), .A2(n21437), .B1(n19087), .B2(n19140), .C1(
        n19086), .C2(n19090), .ZN(P3_U3060) );
  OAI222_X1 U22200 ( .A1(n19090), .A2(n21437), .B1(n19089), .B2(n19140), .C1(
        n19088), .C2(n19083), .ZN(P3_U3061) );
  OAI22_X1 U22201 ( .A1(n19161), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19140), .ZN(n19091) );
  INV_X1 U22202 ( .A(n19091), .ZN(P3_U3274) );
  OAI22_X1 U22203 ( .A1(n19161), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19140), .ZN(n19092) );
  INV_X1 U22204 ( .A(n19092), .ZN(P3_U3275) );
  OAI22_X1 U22205 ( .A1(n19161), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19140), .ZN(n19093) );
  INV_X1 U22206 ( .A(n19093), .ZN(P3_U3276) );
  OAI22_X1 U22207 ( .A1(n19161), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19140), .ZN(n19094) );
  INV_X1 U22208 ( .A(n19094), .ZN(P3_U3277) );
  OAI21_X1 U22209 ( .B1(n19097), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19096), 
        .ZN(n19095) );
  INV_X1 U22210 ( .A(n19095), .ZN(P3_U3280) );
  OAI21_X1 U22211 ( .B1(n19098), .B2(n19097), .A(n19096), .ZN(P3_U3281) );
  NOR2_X1 U22212 ( .A1(n19100), .A2(n19099), .ZN(n19103) );
  OAI21_X1 U22213 ( .B1(n19103), .B2(n19102), .A(n19101), .ZN(P3_U3282) );
  INV_X1 U22214 ( .A(n19104), .ZN(n19106) );
  AOI22_X1 U22215 ( .A1(n19124), .A2(n19106), .B1(n19122), .B2(n19105), .ZN(
        n19107) );
  AOI22_X1 U22216 ( .A1(n19129), .A2(n19108), .B1(n19107), .B2(n19126), .ZN(
        P3_U3285) );
  NOR2_X1 U22217 ( .A1(n19109), .A2(n19125), .ZN(n19116) );
  OAI22_X1 U22218 ( .A1(n13003), .A2(n19110), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19117) );
  INV_X1 U22219 ( .A(n19117), .ZN(n19112) );
  AOI222_X1 U22220 ( .A1(n19113), .A2(n19124), .B1(n19116), .B2(n19112), .C1(
        n19122), .C2(n19111), .ZN(n19114) );
  AOI22_X1 U22221 ( .A1(n19129), .A2(n13017), .B1(n19114), .B2(n19126), .ZN(
        P3_U3288) );
  INV_X1 U22222 ( .A(n19115), .ZN(n19119) );
  AOI222_X1 U22223 ( .A1(n19119), .A2(n19124), .B1(n19122), .B2(n19118), .C1(
        n19117), .C2(n19116), .ZN(n19120) );
  AOI22_X1 U22224 ( .A1(n19129), .A2(n19121), .B1(n19120), .B2(n19126), .ZN(
        P3_U3289) );
  AOI222_X1 U22225 ( .A1(n19125), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19124), 
        .B2(n19123), .C1(n19128), .C2(n19122), .ZN(n19127) );
  AOI22_X1 U22226 ( .A1(n19129), .A2(n19128), .B1(n19127), .B2(n19126), .ZN(
        P3_U3290) );
  AOI21_X1 U22227 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19131) );
  AOI22_X1 U22228 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19131), .B2(n19130), .ZN(n19133) );
  INV_X1 U22229 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19132) );
  AOI22_X1 U22230 ( .A1(n19134), .A2(n19133), .B1(n19132), .B2(n19137), .ZN(
        P3_U3292) );
  INV_X1 U22231 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19138) );
  NOR2_X1 U22232 ( .A1(n19137), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19135) );
  AOI22_X1 U22233 ( .A1(n19138), .A2(n19137), .B1(n19136), .B2(n19135), .ZN(
        P3_U3293) );
  INV_X1 U22234 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19139) );
  AOI22_X1 U22235 ( .A1(n19140), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19139), 
        .B2(n19161), .ZN(P3_U3294) );
  INV_X1 U22236 ( .A(n19141), .ZN(n19144) );
  NAND2_X1 U22237 ( .A1(n19144), .A2(P3_MORE_REG_SCAN_IN), .ZN(n19142) );
  OAI21_X1 U22238 ( .B1(n19144), .B2(n19143), .A(n19142), .ZN(P3_U3295) );
  OAI21_X1 U22239 ( .B1(n19146), .B2(n19145), .A(n19164), .ZN(n19147) );
  AOI21_X1 U22240 ( .B1(n19149), .B2(n19148), .A(n19147), .ZN(n19160) );
  AOI21_X1 U22241 ( .B1(n19152), .B2(n19151), .A(n19150), .ZN(n19154) );
  OAI211_X1 U22242 ( .C1(n19155), .C2(n19154), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19153), .ZN(n19157) );
  AOI21_X1 U22243 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19157), .A(n19156), 
        .ZN(n19159) );
  NAND2_X1 U22244 ( .A1(n19160), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19158) );
  OAI21_X1 U22245 ( .B1(n19160), .B2(n19159), .A(n19158), .ZN(P3_U3296) );
  MUX2_X1 U22246 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n19161), .Z(P3_U3297) );
  OAI21_X1 U22247 ( .B1(n19165), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19164), 
        .ZN(n19162) );
  OAI21_X1 U22248 ( .B1(n19164), .B2(n19163), .A(n19162), .ZN(P3_U3298) );
  NOR2_X1 U22249 ( .A1(n19165), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19167)
         );
  OAI21_X1 U22250 ( .B1(n19168), .B2(n19167), .A(n19166), .ZN(P3_U3299) );
  INV_X1 U22251 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20130) );
  NAND2_X1 U22252 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20130), .ZN(n20117) );
  INV_X1 U22253 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20109) );
  AOI22_X1 U22254 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20117), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n20109), .ZN(n20196) );
  AOI21_X1 U22255 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20196), .ZN(n19169) );
  INV_X1 U22256 ( .A(n19169), .ZN(P2_U2815) );
  INV_X1 U22257 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n21430) );
  OAI22_X1 U22258 ( .A1(n19170), .A2(n21430), .B1(n20200), .B2(n20100), .ZN(
        P2_U2816) );
  INV_X1 U22259 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20122) );
  INV_X2 U22260 ( .A(n20247), .ZN(n20246) );
  AOI21_X1 U22261 ( .B1(n20109), .B2(n20130), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19171) );
  AOI22_X1 U22262 ( .A1(n20246), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19171), 
        .B2(n20247), .ZN(P2_U2817) );
  OAI21_X1 U22263 ( .B1(n20121), .B2(BS16), .A(n20196), .ZN(n20194) );
  OAI21_X1 U22264 ( .B1(n20196), .B2(n20197), .A(n20194), .ZN(P2_U2818) );
  NOR2_X1 U22265 ( .A1(n19172), .A2(n20098), .ZN(n20235) );
  OAI21_X1 U22266 ( .B1(n20235), .B2(n19174), .A(n19173), .ZN(P2_U2819) );
  NOR4_X1 U22267 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19184) );
  NOR4_X1 U22268 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19183) );
  NOR4_X1 U22269 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19175) );
  INV_X1 U22270 ( .A(P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20106) );
  INV_X1 U22271 ( .A(P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21541) );
  NAND3_X1 U22272 ( .A1(n19175), .A2(n20106), .A3(n21541), .ZN(n19181) );
  NOR4_X1 U22273 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19179) );
  NOR4_X1 U22274 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19178) );
  NOR4_X1 U22275 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19177) );
  NOR4_X1 U22276 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19176) );
  NAND4_X1 U22277 ( .A1(n19179), .A2(n19178), .A3(n19177), .A4(n19176), .ZN(
        n19180) );
  AOI211_X1 U22278 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19181), .B(n19180), .ZN(n19182) );
  NAND3_X1 U22279 ( .A1(n19184), .A2(n19183), .A3(n19182), .ZN(n19193) );
  NOR2_X1 U22280 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19193), .ZN(n19187) );
  INV_X1 U22281 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19185) );
  AOI22_X1 U22282 ( .A1(n19187), .A2(n19188), .B1(n19193), .B2(n19185), .ZN(
        P2_U2820) );
  OR3_X1 U22283 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19192) );
  INV_X1 U22284 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19186) );
  AOI22_X1 U22285 ( .A1(n19187), .A2(n19192), .B1(n19193), .B2(n19186), .ZN(
        P2_U2821) );
  INV_X1 U22286 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20195) );
  NAND2_X1 U22287 ( .A1(n19187), .A2(n20195), .ZN(n19191) );
  INV_X1 U22288 ( .A(n19193), .ZN(n19195) );
  OAI21_X1 U22289 ( .B1(n19188), .B2(n20132), .A(n19195), .ZN(n19189) );
  OAI21_X1 U22290 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19195), .A(n19189), 
        .ZN(n19190) );
  OAI221_X1 U22291 ( .B1(n19191), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19191), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19190), .ZN(P2_U2822) );
  INV_X1 U22292 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19194) );
  OAI221_X1 U22293 ( .B1(n19195), .B2(n19194), .C1(n19193), .C2(n19192), .A(
        n19191), .ZN(P2_U2823) );
  OAI22_X1 U22294 ( .A1(n19353), .A2(n19197), .B1(n19196), .B2(n19378), .ZN(
        n19198) );
  AOI21_X1 U22295 ( .B1(P2_REIP_REG_21__SCAN_IN), .B2(n19369), .A(n19198), 
        .ZN(n19199) );
  OAI21_X1 U22296 ( .B1(n19200), .B2(n19343), .A(n19199), .ZN(n19201) );
  AOI21_X1 U22297 ( .B1(n19202), .B2(n19367), .A(n19201), .ZN(n19207) );
  OAI211_X1 U22298 ( .C1(n19205), .C2(n19204), .A(n20102), .B(n19203), .ZN(
        n19206) );
  OAI211_X1 U22299 ( .C1(n19371), .C2(n19208), .A(n19207), .B(n19206), .ZN(
        P2_U2834) );
  INV_X1 U22300 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20166) );
  AOI22_X1 U22301 ( .A1(n19209), .A2(n19367), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19356), .ZN(n19210) );
  OAI21_X1 U22302 ( .B1(n20166), .B2(n19349), .A(n19210), .ZN(n19211) );
  AOI211_X1 U22303 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19368), .A(n19247), .B(
        n19211), .ZN(n19220) );
  OAI22_X1 U22304 ( .A1(n19213), .A2(n19343), .B1(n19212), .B2(n19371), .ZN(
        n19214) );
  INV_X1 U22305 ( .A(n19214), .ZN(n19219) );
  OAI211_X1 U22306 ( .C1(n19217), .C2(n19216), .A(n20102), .B(n19215), .ZN(
        n19218) );
  NAND3_X1 U22307 ( .A1(n19220), .A2(n19219), .A3(n19218), .ZN(P2_U2836) );
  INV_X1 U22308 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n19221) );
  OAI222_X1 U22309 ( .A1(n19351), .A2(n19223), .B1(n19353), .B2(n19222), .C1(
        n19378), .C2(n19221), .ZN(n19224) );
  AOI211_X1 U22310 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19369), .A(n19247), 
        .B(n19224), .ZN(n19232) );
  AOI22_X1 U22311 ( .A1(n19226), .A2(n19364), .B1(n19225), .B2(n19275), .ZN(
        n19231) );
  OAI211_X1 U22312 ( .C1(n19229), .C2(n19228), .A(n20102), .B(n19227), .ZN(
        n19230) );
  NAND3_X1 U22313 ( .A1(n19232), .A2(n19231), .A3(n19230), .ZN(P2_U2837) );
  OAI21_X1 U22314 ( .B1(n20162), .B2(n19349), .A(n19233), .ZN(n19238) );
  INV_X1 U22315 ( .A(n19234), .ZN(n19236) );
  OAI22_X1 U22316 ( .A1(n19236), .A2(n19351), .B1(n19235), .B2(n19378), .ZN(
        n19237) );
  AOI211_X1 U22317 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19368), .A(n19238), .B(
        n19237), .ZN(n19246) );
  AOI22_X1 U22318 ( .A1(n19240), .A2(n19364), .B1(n19239), .B2(n19275), .ZN(
        n19245) );
  OAI211_X1 U22319 ( .C1(n19243), .C2(n19242), .A(n20102), .B(n19241), .ZN(
        n19244) );
  NAND3_X1 U22320 ( .A1(n19246), .A2(n19245), .A3(n19244), .ZN(P2_U2838) );
  AOI21_X1 U22321 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19356), .A(
        n19247), .ZN(n19249) );
  NAND2_X1 U22322 ( .A1(n19369), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n19248) );
  OAI211_X1 U22323 ( .C1(n19353), .C2(n19250), .A(n19249), .B(n19248), .ZN(
        n19253) );
  NOR2_X1 U22324 ( .A1(n19251), .A2(n19351), .ZN(n19252) );
  AOI211_X1 U22325 ( .C1(n19254), .C2(n19364), .A(n19253), .B(n19252), .ZN(
        n19259) );
  OAI211_X1 U22326 ( .C1(n19257), .C2(n19256), .A(n20102), .B(n19255), .ZN(
        n19258) );
  OAI211_X1 U22327 ( .C1(n19260), .C2(n19371), .A(n19259), .B(n19258), .ZN(
        P2_U2839) );
  XNOR2_X1 U22328 ( .A(n19262), .B(n19261), .ZN(n19269) );
  AOI22_X1 U22329 ( .A1(n19263), .A2(n19367), .B1(P2_REIP_REG_15__SCAN_IN), 
        .B2(n19369), .ZN(n19264) );
  OAI211_X1 U22330 ( .C1(n12412), .C2(n19353), .A(n19264), .B(n19348), .ZN(
        n19267) );
  OAI22_X1 U22331 ( .A1(n19265), .A2(n19343), .B1(n19371), .B2(n19391), .ZN(
        n19266) );
  AOI211_X1 U22332 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19356), .A(
        n19267), .B(n19266), .ZN(n19268) );
  OAI21_X1 U22333 ( .B1(n19334), .B2(n19269), .A(n19268), .ZN(P2_U2840) );
  NOR2_X1 U22334 ( .A1(n9824), .A2(n19270), .ZN(n19288) );
  XOR2_X1 U22335 ( .A(n19288), .B(n19271), .Z(n19279) );
  INV_X1 U22336 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20156) );
  AOI22_X1 U22337 ( .A1(n19272), .A2(n19367), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19356), .ZN(n19273) );
  OAI21_X1 U22338 ( .B1(n20156), .B2(n19349), .A(n19273), .ZN(n19274) );
  AOI211_X1 U22339 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n19368), .A(n19247), .B(
        n19274), .ZN(n19278) );
  AOI22_X1 U22340 ( .A1(n19276), .A2(n19364), .B1(n19275), .B2(n19392), .ZN(
        n19277) );
  OAI211_X1 U22341 ( .C1(n19334), .C2(n19279), .A(n19278), .B(n19277), .ZN(
        P2_U2841) );
  AOI22_X1 U22342 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19356), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19369), .ZN(n19280) );
  OAI211_X1 U22343 ( .C1(n19289), .C2(n19377), .A(n19348), .B(n19280), .ZN(
        n19282) );
  NOR2_X1 U22344 ( .A1(n19353), .A2(n12404), .ZN(n19281) );
  AOI211_X1 U22345 ( .C1(n19283), .C2(n19364), .A(n19282), .B(n19281), .ZN(
        n19284) );
  OAI21_X1 U22346 ( .B1(n19285), .B2(n19351), .A(n19284), .ZN(n19286) );
  INV_X1 U22347 ( .A(n19286), .ZN(n19292) );
  INV_X1 U22348 ( .A(n19287), .ZN(n19290) );
  OAI211_X1 U22349 ( .C1(n19290), .C2(n19289), .A(n20102), .B(n19288), .ZN(
        n19291) );
  OAI211_X1 U22350 ( .C1(n19397), .C2(n19371), .A(n19292), .B(n19291), .ZN(
        P2_U2842) );
  INV_X1 U22351 ( .A(n19300), .ZN(n19293) );
  OAI211_X1 U22352 ( .C1(n9824), .C2(n19294), .A(n20102), .B(n19293), .ZN(
        n19296) );
  AOI22_X1 U22353 ( .A1(n19368), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19356), .ZN(n19295) );
  OAI211_X1 U22354 ( .C1(n19297), .C2(n19351), .A(n19296), .B(n19295), .ZN(
        n19298) );
  AOI211_X1 U22355 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19369), .A(n19247), 
        .B(n19298), .ZN(n19303) );
  AOI22_X1 U22356 ( .A1(n19301), .A2(n19300), .B1(n19364), .B2(n19299), .ZN(
        n19302) );
  OAI211_X1 U22357 ( .C1(n19371), .C2(n19400), .A(n19303), .B(n19302), .ZN(
        P2_U2843) );
  OAI21_X1 U22358 ( .B1(n20148), .B2(n19349), .A(n19348), .ZN(n19306) );
  OAI22_X1 U22359 ( .A1(n19304), .A2(n19351), .B1(n10305), .B2(n19353), .ZN(
        n19305) );
  AOI211_X1 U22360 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19356), .A(
        n19306), .B(n19305), .ZN(n19313) );
  NOR2_X1 U22361 ( .A1(n9878), .A2(n19307), .ZN(n19309) );
  XNOR2_X1 U22362 ( .A(n19309), .B(n19308), .ZN(n19311) );
  AOI22_X1 U22363 ( .A1(n19311), .A2(n20102), .B1(n19364), .B2(n19310), .ZN(
        n19312) );
  OAI211_X1 U22364 ( .C1(n19371), .C2(n19405), .A(n19313), .B(n19312), .ZN(
        P2_U2845) );
  NAND2_X1 U22365 ( .A1(n9876), .A2(n19314), .ZN(n19316) );
  XOR2_X1 U22366 ( .A(n19316), .B(n19315), .Z(n19323) );
  AOI22_X1 U22367 ( .A1(n19317), .A2(n19367), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19356), .ZN(n19318) );
  OAI211_X1 U22368 ( .C1(n20146), .C2(n19349), .A(n19318), .B(n19348), .ZN(
        n19321) );
  OAI22_X1 U22369 ( .A1(n19319), .A2(n19343), .B1(n19371), .B2(n19407), .ZN(
        n19320) );
  AOI211_X1 U22370 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19368), .A(n19321), .B(
        n19320), .ZN(n19322) );
  OAI21_X1 U22371 ( .B1(n19323), .B2(n19334), .A(n19322), .ZN(P2_U2846) );
  NAND2_X1 U22372 ( .A1(n9875), .A2(n19324), .ZN(n19326) );
  XOR2_X1 U22373 ( .A(n19326), .B(n19325), .Z(n19335) );
  OAI22_X1 U22374 ( .A1(n19327), .A2(n19351), .B1(n12392), .B2(n19353), .ZN(
        n19328) );
  INV_X1 U22375 ( .A(n19328), .ZN(n19329) );
  OAI211_X1 U22376 ( .C1(n20143), .C2(n19349), .A(n19329), .B(n19348), .ZN(
        n19332) );
  OAI22_X1 U22377 ( .A1(n19413), .A2(n19371), .B1(n19343), .B2(n19330), .ZN(
        n19331) );
  AOI211_X1 U22378 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19356), .A(
        n19332), .B(n19331), .ZN(n19333) );
  OAI21_X1 U22379 ( .B1(n19335), .B2(n19334), .A(n19333), .ZN(P2_U2848) );
  OAI22_X1 U22380 ( .A1(n19337), .A2(n19351), .B1(n19336), .B2(n19378), .ZN(
        n19338) );
  AOI211_X1 U22381 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n19369), .A(n19247), .B(
        n19338), .ZN(n19347) );
  NOR2_X1 U22382 ( .A1(n9878), .A2(n19339), .ZN(n19340) );
  XNOR2_X1 U22383 ( .A(n19341), .B(n19340), .ZN(n19345) );
  OAI22_X1 U22384 ( .A1(n19414), .A2(n19371), .B1(n19343), .B2(n19342), .ZN(
        n19344) );
  AOI21_X1 U22385 ( .B1(n19345), .B2(n20102), .A(n19344), .ZN(n19346) );
  OAI211_X1 U22386 ( .C1(n12388), .C2(n19353), .A(n19347), .B(n19346), .ZN(
        P2_U2849) );
  OAI21_X1 U22387 ( .B1(n20139), .B2(n19349), .A(n19348), .ZN(n19355) );
  OAI22_X1 U22388 ( .A1(n19353), .A2(n19352), .B1(n19351), .B2(n19350), .ZN(
        n19354) );
  AOI211_X1 U22389 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19356), .A(
        n19355), .B(n19354), .ZN(n19363) );
  NAND2_X1 U22390 ( .A1(n9877), .A2(n19357), .ZN(n19358) );
  XNOR2_X1 U22391 ( .A(n19359), .B(n19358), .ZN(n19361) );
  AOI22_X1 U22392 ( .A1(n19361), .A2(n20102), .B1(n19364), .B2(n19360), .ZN(
        n19362) );
  OAI211_X1 U22393 ( .C1(n19371), .C2(n19422), .A(n19363), .B(n19362), .ZN(
        P2_U2850) );
  NAND2_X1 U22394 ( .A1(n19365), .A2(n19364), .ZN(n19375) );
  AOI22_X1 U22395 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(n19368), .B1(n19367), .B2(
        n19366), .ZN(n19374) );
  NAND2_X1 U22396 ( .A1(n19369), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19373) );
  OR2_X1 U22397 ( .A1(n19371), .A2(n19370), .ZN(n19372) );
  NAND4_X1 U22398 ( .A1(n19375), .A2(n19374), .A3(n19373), .A4(n19372), .ZN(
        n19380) );
  INV_X1 U22399 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19376) );
  AOI21_X1 U22400 ( .B1(n19378), .B2(n19377), .A(n19376), .ZN(n19379) );
  AOI211_X1 U22401 ( .C1(n19381), .C2(n19447), .A(n19380), .B(n19379), .ZN(
        n19382) );
  OAI21_X1 U22402 ( .B1(n19384), .B2(n19383), .A(n19382), .ZN(P2_U2855) );
  AOI22_X1 U22403 ( .A1(n19386), .A2(n19443), .B1(n19385), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19389) );
  AOI22_X1 U22404 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19442), .B1(n19387), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19388) );
  NAND2_X1 U22405 ( .A1(n19389), .A2(n19388), .ZN(P2_U2888) );
  INV_X1 U22406 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19454) );
  OAI222_X1 U22407 ( .A1(n19391), .A2(n19423), .B1(n19454), .B2(n19415), .C1(
        n19390), .C2(n19450), .ZN(P2_U2904) );
  INV_X1 U22408 ( .A(n19392), .ZN(n19395) );
  AOI22_X1 U22409 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19442), .B1(n19393), 
        .B2(n19409), .ZN(n19394) );
  OAI21_X1 U22410 ( .B1(n19423), .B2(n19395), .A(n19394), .ZN(P2_U2905) );
  INV_X1 U22411 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n21534) );
  OAI222_X1 U22412 ( .A1(n19397), .A2(n19423), .B1(n21534), .B2(n19415), .C1(
        n19450), .C2(n19396), .ZN(P2_U2906) );
  AOI22_X1 U22413 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19442), .B1(n19398), 
        .B2(n19409), .ZN(n19399) );
  OAI21_X1 U22414 ( .B1(n19423), .B2(n19400), .A(n19399), .ZN(P2_U2907) );
  INV_X1 U22415 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19461) );
  OAI222_X1 U22416 ( .A1(n19402), .A2(n19423), .B1(n19461), .B2(n19415), .C1(
        n19450), .C2(n19401), .ZN(P2_U2908) );
  AOI22_X1 U22417 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19442), .B1(n19403), 
        .B2(n19409), .ZN(n19404) );
  OAI21_X1 U22418 ( .B1(n19423), .B2(n19405), .A(n19404), .ZN(P2_U2909) );
  INV_X1 U22419 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19465) );
  OAI222_X1 U22420 ( .A1(n19407), .A2(n19423), .B1(n19465), .B2(n19415), .C1(
        n19450), .C2(n19406), .ZN(P2_U2910) );
  INV_X1 U22421 ( .A(n19408), .ZN(n19412) );
  AOI22_X1 U22422 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19442), .B1(n19410), .B2(
        n19409), .ZN(n19411) );
  OAI21_X1 U22423 ( .B1(n19423), .B2(n19412), .A(n19411), .ZN(P2_U2911) );
  OAI222_X1 U22424 ( .A1(n19413), .A2(n19423), .B1(n19470), .B2(n19415), .C1(
        n19450), .C2(n19572), .ZN(P2_U2912) );
  INV_X1 U22425 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19472) );
  OAI222_X1 U22426 ( .A1(n19414), .A2(n19423), .B1(n19472), .B2(n19415), .C1(
        n19450), .C2(n19558), .ZN(P2_U2913) );
  INV_X1 U22427 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19474) );
  OAI22_X1 U22428 ( .A1(n19474), .A2(n19415), .B1(n19553), .B2(n19450), .ZN(
        n19416) );
  INV_X1 U22429 ( .A(n19416), .ZN(n19421) );
  OAI21_X1 U22430 ( .B1(n19677), .B2(n20214), .A(n19417), .ZN(n19431) );
  XOR2_X1 U22431 ( .A(n19429), .B(n20202), .Z(n19432) );
  NAND2_X1 U22432 ( .A1(n19431), .A2(n19432), .ZN(n19430) );
  NAND2_X1 U22433 ( .A1(n20202), .A2(n19429), .ZN(n19418) );
  AOI21_X1 U22434 ( .B1(n19430), .B2(n19418), .A(n19504), .ZN(n19424) );
  OR3_X1 U22435 ( .A1(n19424), .A2(n19425), .A3(n19419), .ZN(n19420) );
  OAI211_X1 U22436 ( .C1(n19423), .C2(n19422), .A(n19421), .B(n19420), .ZN(
        P2_U2914) );
  AOI22_X1 U22437 ( .A1(n19443), .A2(n19504), .B1(n19442), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19428) );
  XOR2_X1 U22438 ( .A(n19425), .B(n19424), .Z(n19426) );
  NAND2_X1 U22439 ( .A1(n19426), .A2(n19444), .ZN(n19427) );
  OAI211_X1 U22440 ( .C1(n19548), .C2(n19450), .A(n19428), .B(n19427), .ZN(
        P2_U2915) );
  INV_X1 U22441 ( .A(n19429), .ZN(n20207) );
  AOI22_X1 U22442 ( .A1(n20207), .A2(n19443), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19442), .ZN(n19435) );
  OAI21_X1 U22443 ( .B1(n19432), .B2(n19431), .A(n19430), .ZN(n19433) );
  NAND2_X1 U22444 ( .A1(n19433), .A2(n19444), .ZN(n19434) );
  OAI211_X1 U22445 ( .C1(n19542), .C2(n19450), .A(n19435), .B(n19434), .ZN(
        P2_U2916) );
  AOI22_X1 U22446 ( .A1(n19443), .A2(n20223), .B1(n19442), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19440) );
  OAI21_X1 U22447 ( .B1(n19437), .B2(n19445), .A(n19436), .ZN(n19438) );
  NAND2_X1 U22448 ( .A1(n19438), .A2(n19444), .ZN(n19439) );
  OAI211_X1 U22449 ( .C1(n19441), .C2(n19450), .A(n19440), .B(n19439), .ZN(
        P2_U2918) );
  AOI22_X1 U22450 ( .A1(n19443), .A2(n19446), .B1(n19442), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19449) );
  OAI211_X1 U22451 ( .C1(n19447), .C2(n19446), .A(n19445), .B(n19444), .ZN(
        n19448) );
  OAI211_X1 U22452 ( .C1(n19451), .C2(n19450), .A(n19449), .B(n19448), .ZN(
        P2_U2919) );
  AND2_X1 U22453 ( .A1(n19475), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22454 ( .A1(n19485), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19453) );
  OAI21_X1 U22455 ( .B1(n19454), .B2(n19487), .A(n19453), .ZN(P2_U2936) );
  AOI22_X1 U22456 ( .A1(n19466), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19455) );
  OAI21_X1 U22457 ( .B1(n19456), .B2(n19487), .A(n19455), .ZN(P2_U2937) );
  AOI22_X1 U22458 ( .A1(n19466), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19457) );
  OAI21_X1 U22459 ( .B1(n21534), .B2(n19487), .A(n19457), .ZN(P2_U2938) );
  AOI22_X1 U22460 ( .A1(n19466), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19458) );
  OAI21_X1 U22461 ( .B1(n19459), .B2(n19487), .A(n19458), .ZN(P2_U2939) );
  AOI22_X1 U22462 ( .A1(n19466), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19460) );
  OAI21_X1 U22463 ( .B1(n19461), .B2(n19487), .A(n19460), .ZN(P2_U2940) );
  AOI22_X1 U22464 ( .A1(n19466), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19462) );
  OAI21_X1 U22465 ( .B1(n19463), .B2(n19487), .A(n19462), .ZN(P2_U2941) );
  AOI22_X1 U22466 ( .A1(n19466), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19464) );
  OAI21_X1 U22467 ( .B1(n19465), .B2(n19487), .A(n19464), .ZN(P2_U2942) );
  AOI22_X1 U22468 ( .A1(n19466), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19467) );
  OAI21_X1 U22469 ( .B1(n19468), .B2(n19487), .A(n19467), .ZN(P2_U2943) );
  AOI22_X1 U22470 ( .A1(n19485), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19469) );
  OAI21_X1 U22471 ( .B1(n19470), .B2(n19487), .A(n19469), .ZN(P2_U2944) );
  AOI22_X1 U22472 ( .A1(n19485), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19471) );
  OAI21_X1 U22473 ( .B1(n19472), .B2(n19487), .A(n19471), .ZN(P2_U2945) );
  AOI22_X1 U22474 ( .A1(n19485), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19473) );
  OAI21_X1 U22475 ( .B1(n19474), .B2(n19487), .A(n19473), .ZN(P2_U2946) );
  INV_X1 U22476 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19477) );
  AOI22_X1 U22477 ( .A1(n19485), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19475), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19476) );
  OAI21_X1 U22478 ( .B1(n19477), .B2(n19487), .A(n19476), .ZN(P2_U2947) );
  INV_X1 U22479 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19479) );
  AOI22_X1 U22480 ( .A1(n19485), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19478) );
  OAI21_X1 U22481 ( .B1(n19479), .B2(n19487), .A(n19478), .ZN(P2_U2948) );
  INV_X1 U22482 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19481) );
  AOI22_X1 U22483 ( .A1(n19485), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19480) );
  OAI21_X1 U22484 ( .B1(n19481), .B2(n19487), .A(n19480), .ZN(P2_U2949) );
  INV_X1 U22485 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19483) );
  AOI22_X1 U22486 ( .A1(n19485), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19482) );
  OAI21_X1 U22487 ( .B1(n19483), .B2(n19487), .A(n19482), .ZN(P2_U2950) );
  AOI22_X1 U22488 ( .A1(n19485), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19486) );
  OAI21_X1 U22489 ( .B1(n12475), .B2(n19487), .A(n19486), .ZN(P2_U2951) );
  AOI22_X1 U22490 ( .A1(n19488), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19247), .ZN(n19497) );
  XNOR2_X1 U22491 ( .A(n19490), .B(n19502), .ZN(n19506) );
  XOR2_X1 U22492 ( .A(n19492), .B(n19491), .Z(n19507) );
  AOI222_X1 U22493 ( .A1(n19506), .A2(n19495), .B1(n19494), .B2(n19501), .C1(
        n19493), .C2(n19507), .ZN(n19496) );
  OAI211_X1 U22494 ( .C1(n19499), .C2(n19498), .A(n19497), .B(n19496), .ZN(
        P2_U3010) );
  AOI22_X1 U22495 ( .A1(n19503), .A2(n19502), .B1(n19501), .B2(n19500), .ZN(
        n19511) );
  AOI22_X1 U22496 ( .A1(n19505), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19517), .B2(n19504), .ZN(n19510) );
  AOI22_X1 U22497 ( .A1(n19507), .A2(n19526), .B1(n12862), .B2(n19506), .ZN(
        n19509) );
  NAND2_X1 U22498 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19247), .ZN(n19508) );
  NAND4_X1 U22499 ( .A1(n19511), .A2(n19510), .A3(n19509), .A4(n19508), .ZN(
        P2_U3042) );
  OR2_X1 U22500 ( .A1(n19512), .A2(n19519), .ZN(n19514) );
  OAI211_X1 U22501 ( .C1(n19523), .C2(n19515), .A(n19514), .B(n19513), .ZN(
        n19516) );
  INV_X1 U22502 ( .A(n19516), .ZN(n19538) );
  NAND2_X1 U22503 ( .A1(n20214), .A2(n19517), .ZN(n19532) );
  INV_X1 U22504 ( .A(n19518), .ZN(n19520) );
  NAND2_X1 U22505 ( .A1(n19520), .A2(n19519), .ZN(n19530) );
  AOI22_X1 U22506 ( .A1(n12862), .A2(n19521), .B1(n19247), .B2(
        P2_REIP_REG_2__SCAN_IN), .ZN(n19529) );
  OR2_X1 U22507 ( .A1(n19523), .A2(n19522), .ZN(n19528) );
  NAND3_X1 U22508 ( .A1(n19526), .A2(n19525), .A3(n19524), .ZN(n19527) );
  AND4_X1 U22509 ( .A1(n19530), .A2(n19529), .A3(n19528), .A4(n19527), .ZN(
        n19531) );
  OAI211_X1 U22510 ( .C1(n19534), .C2(n19533), .A(n19532), .B(n19531), .ZN(
        n19535) );
  INV_X1 U22511 ( .A(n19535), .ZN(n19536) );
  OAI21_X1 U22512 ( .B1(n19538), .B2(n19537), .A(n19536), .ZN(P2_U3044) );
  AOI22_X1 U22513 ( .A1(n19883), .A2(n20092), .B1(n19571), .B2(n20013), .ZN(
        n19540) );
  AOI22_X1 U22514 ( .A1(n14206), .A2(n19573), .B1(n19605), .B2(n20014), .ZN(
        n19539) );
  OAI211_X1 U22515 ( .C1(n19566), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3048) );
  AOI22_X1 U22516 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19568), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19567), .ZN(n20069) );
  NOR2_X2 U22517 ( .A1(n11681), .A2(n19546), .ZN(n20064) );
  AOI22_X1 U22518 ( .A1(n20092), .A2(n19994), .B1(n19571), .B2(n20064), .ZN(
        n19544) );
  NOR2_X2 U22519 ( .A1(n19542), .A2(n19981), .ZN(n20065) );
  AOI22_X1 U22520 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19568), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19567), .ZN(n19997) );
  INV_X1 U22521 ( .A(n19997), .ZN(n20066) );
  AOI22_X1 U22522 ( .A1(n20065), .A2(n19573), .B1(n19605), .B2(n20066), .ZN(
        n19543) );
  OAI211_X1 U22523 ( .C1(n19566), .C2(n19545), .A(n19544), .B(n19543), .ZN(
        P2_U3051) );
  AOI22_X1 U22524 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19568), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19567), .ZN(n20002) );
  AOI22_X1 U22525 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19568), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19567), .ZN(n20074) );
  INV_X1 U22526 ( .A(n20074), .ZN(n19998) );
  NOR2_X2 U22527 ( .A1(n19547), .A2(n19546), .ZN(n20070) );
  AOI22_X1 U22528 ( .A1(n19998), .A2(n20092), .B1(n19571), .B2(n20070), .ZN(
        n19551) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19574), .B1(
        n19549), .B2(n19573), .ZN(n19550) );
  OAI211_X1 U22530 ( .C1(n20002), .C2(n19617), .A(n19551), .B(n19550), .ZN(
        P2_U3052) );
  AOI22_X1 U22531 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19568), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19567), .ZN(n20080) );
  INV_X1 U22532 ( .A(n20080), .ZN(n19964) );
  AOI22_X1 U22533 ( .A1(n19964), .A2(n20092), .B1(n19571), .B2(n20075), .ZN(
        n19555) );
  NOR2_X2 U22534 ( .A1(n19553), .A2(n19981), .ZN(n20076) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19574), .B1(
        n20076), .B2(n19573), .ZN(n19554) );
  OAI211_X1 U22536 ( .C1(n19968), .C2(n19617), .A(n19555), .B(n19554), .ZN(
        P2_U3053) );
  OAI22_X1 U22537 ( .A1(n19556), .A2(n19561), .B1(n21395), .B2(n19559), .ZN(
        n19660) );
  AND2_X1 U22538 ( .A1(n19557), .A2(n19569), .ZN(n20081) );
  AOI22_X1 U22539 ( .A1(n19660), .A2(n20092), .B1(n19571), .B2(n20081), .ZN(
        n19564) );
  NOR2_X2 U22540 ( .A1(n19558), .A2(n19981), .ZN(n20082) );
  OAI22_X2 U22541 ( .A1(n19562), .A2(n19561), .B1(n19560), .B2(n19559), .ZN(
        n20083) );
  AOI22_X1 U22542 ( .A1(n20082), .A2(n19573), .B1(n19605), .B2(n20083), .ZN(
        n19563) );
  OAI211_X1 U22543 ( .C1(n19566), .C2(n19565), .A(n19564), .B(n19563), .ZN(
        P2_U3054) );
  AOI22_X1 U22544 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19568), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19567), .ZN(n19943) );
  AOI22_X1 U22545 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19568), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19567), .ZN(n20097) );
  INV_X1 U22546 ( .A(n20097), .ZN(n19938) );
  AND2_X1 U22547 ( .A1(n19570), .A2(n19569), .ZN(n20087) );
  AOI22_X1 U22548 ( .A1(n19938), .A2(n20092), .B1(n19571), .B2(n20087), .ZN(
        n19576) );
  NOR2_X2 U22549 ( .A1(n19572), .A2(n19981), .ZN(n20089) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19574), .B1(
        n20089), .B2(n19573), .ZN(n19575) );
  OAI211_X1 U22551 ( .C1(n19943), .C2(n19617), .A(n19576), .B(n19575), .ZN(
        P2_U3055) );
  NOR2_X1 U22552 ( .A1(n19577), .A2(n19620), .ZN(n19588) );
  OR2_X1 U22553 ( .A1(n19588), .A2(n19913), .ZN(n19578) );
  NOR2_X1 U22554 ( .A1(n19579), .A2(n19578), .ZN(n19584) );
  INV_X1 U22555 ( .A(n19585), .ZN(n19580) );
  NOR2_X1 U22556 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19580), .ZN(n19581) );
  INV_X1 U22557 ( .A(n14206), .ZN(n19772) );
  INV_X1 U22558 ( .A(n19588), .ZN(n19611) );
  OAI22_X1 U22559 ( .A1(n19612), .A2(n19772), .B1(n19771), .B2(n19611), .ZN(
        n19582) );
  INV_X1 U22560 ( .A(n19582), .ZN(n19591) );
  NAND2_X1 U22561 ( .A1(n19704), .A2(n19583), .ZN(n19586) );
  AOI21_X1 U22562 ( .B1(n19586), .B2(n19585), .A(n19584), .ZN(n19587) );
  OAI211_X1 U22563 ( .C1(n19588), .C2(n19873), .A(n19587), .B(n20020), .ZN(
        n19614) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19614), .B1(
        n19646), .B2(n20014), .ZN(n19590) );
  OAI211_X1 U22565 ( .C1(n20028), .C2(n19617), .A(n19591), .B(n19590), .ZN(
        P2_U3056) );
  INV_X1 U22566 ( .A(n14210), .ZN(n19784) );
  INV_X1 U22567 ( .A(n20051), .ZN(n19783) );
  OAI22_X1 U22568 ( .A1(n19612), .A2(n19784), .B1(n19783), .B2(n19611), .ZN(
        n19592) );
  INV_X1 U22569 ( .A(n19592), .ZN(n19594) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19614), .B1(
        n19605), .B2(n20053), .ZN(n19593) );
  OAI211_X1 U22571 ( .C1(n20031), .C2(n19643), .A(n19594), .B(n19593), .ZN(
        P2_U3057) );
  INV_X1 U22572 ( .A(n14355), .ZN(n19789) );
  INV_X1 U22573 ( .A(n20059), .ZN(n19788) );
  OAI22_X1 U22574 ( .A1(n19612), .A2(n19789), .B1(n19788), .B2(n19611), .ZN(
        n19595) );
  INV_X1 U22575 ( .A(n19595), .ZN(n19597) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19614), .B1(
        n19605), .B2(n20033), .ZN(n19596) );
  OAI211_X1 U22577 ( .C1(n20036), .C2(n19643), .A(n19597), .B(n19596), .ZN(
        P2_U3058) );
  INV_X1 U22578 ( .A(n20065), .ZN(n19795) );
  INV_X1 U22579 ( .A(n20064), .ZN(n19794) );
  OAI22_X1 U22580 ( .A1(n19612), .A2(n19795), .B1(n19794), .B2(n19611), .ZN(
        n19598) );
  INV_X1 U22581 ( .A(n19598), .ZN(n19600) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19614), .B1(
        n19605), .B2(n19994), .ZN(n19599) );
  OAI211_X1 U22583 ( .C1(n19997), .C2(n19643), .A(n19600), .B(n19599), .ZN(
        P2_U3059) );
  INV_X1 U22584 ( .A(n19549), .ZN(n19800) );
  INV_X1 U22585 ( .A(n20070), .ZN(n19799) );
  OAI22_X1 U22586 ( .A1(n19612), .A2(n19800), .B1(n19799), .B2(n19611), .ZN(
        n19601) );
  INV_X1 U22587 ( .A(n19601), .ZN(n19603) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19614), .B1(
        n19605), .B2(n19998), .ZN(n19602) );
  OAI211_X1 U22589 ( .C1(n20002), .C2(n19643), .A(n19603), .B(n19602), .ZN(
        P2_U3060) );
  INV_X1 U22590 ( .A(n20076), .ZN(n19805) );
  INV_X1 U22591 ( .A(n20075), .ZN(n19804) );
  OAI22_X1 U22592 ( .A1(n19612), .A2(n19805), .B1(n19804), .B2(n19611), .ZN(
        n19604) );
  INV_X1 U22593 ( .A(n19604), .ZN(n19607) );
  AOI22_X1 U22594 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19614), .B1(
        n19605), .B2(n19964), .ZN(n19606) );
  OAI211_X1 U22595 ( .C1(n19968), .C2(n19643), .A(n19607), .B(n19606), .ZN(
        P2_U3061) );
  INV_X1 U22596 ( .A(n20082), .ZN(n19810) );
  INV_X1 U22597 ( .A(n20081), .ZN(n19809) );
  OAI22_X1 U22598 ( .A1(n19612), .A2(n19810), .B1(n19809), .B2(n19611), .ZN(
        n19608) );
  INV_X1 U22599 ( .A(n19608), .ZN(n19610) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19614), .B1(
        n19646), .B2(n20083), .ZN(n19609) );
  OAI211_X1 U22601 ( .C1(n20086), .C2(n19617), .A(n19610), .B(n19609), .ZN(
        P2_U3062) );
  INV_X1 U22602 ( .A(n20089), .ZN(n19815) );
  INV_X1 U22603 ( .A(n20087), .ZN(n19814) );
  OAI22_X1 U22604 ( .A1(n19612), .A2(n19815), .B1(n19814), .B2(n19611), .ZN(
        n19613) );
  INV_X1 U22605 ( .A(n19613), .ZN(n19616) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19614), .B1(
        n19646), .B2(n20091), .ZN(n19615) );
  OAI211_X1 U22607 ( .C1(n20097), .C2(n19617), .A(n19616), .B(n19615), .ZN(
        P2_U3063) );
  INV_X1 U22608 ( .A(n19623), .ZN(n19619) );
  NOR2_X1 U22609 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21540), .ZN(
        n19876) );
  AND2_X1 U22610 ( .A1(n19876), .A2(n19618), .ZN(n19644) );
  OAI21_X1 U22611 ( .B1(n19619), .B2(n19644), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19621) );
  OR2_X1 U22612 ( .A1(n19882), .A2(n19620), .ZN(n19624) );
  NAND2_X1 U22613 ( .A1(n19621), .A2(n19624), .ZN(n19645) );
  AOI22_X1 U22614 ( .A1(n19645), .A2(n14206), .B1(n20013), .B2(n19644), .ZN(
        n19630) );
  INV_X1 U22615 ( .A(n19644), .ZN(n19622) );
  OAI21_X1 U22616 ( .B1(n19623), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19622), 
        .ZN(n19627) );
  OAI21_X1 U22617 ( .B1(n19659), .B2(n19646), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19625) );
  NAND2_X1 U22618 ( .A1(n19625), .A2(n19624), .ZN(n19626) );
  MUX2_X1 U22619 ( .A(n19627), .B(n19626), .S(n20206), .Z(n19628) );
  NAND2_X1 U22620 ( .A1(n19628), .A2(n20020), .ZN(n19647) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19647), .B1(
        n19659), .B2(n20014), .ZN(n19629) );
  OAI211_X1 U22622 ( .C1(n20028), .C2(n19643), .A(n19630), .B(n19629), .ZN(
        P2_U3064) );
  AOI22_X1 U22623 ( .A1(n19645), .A2(n14210), .B1(n20051), .B2(n19644), .ZN(
        n19632) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19647), .B1(
        n19646), .B2(n20053), .ZN(n19631) );
  OAI211_X1 U22625 ( .C1(n20031), .C2(n19670), .A(n19632), .B(n19631), .ZN(
        P2_U3065) );
  AOI22_X1 U22626 ( .A1(n19645), .A2(n14355), .B1(n20059), .B2(n19644), .ZN(
        n19634) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19647), .B1(
        n19646), .B2(n20033), .ZN(n19633) );
  OAI211_X1 U22628 ( .C1(n20036), .C2(n19670), .A(n19634), .B(n19633), .ZN(
        P2_U3066) );
  AOI22_X1 U22629 ( .A1(n19645), .A2(n20065), .B1(n20064), .B2(n19644), .ZN(
        n19636) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19647), .B1(
        n19646), .B2(n19994), .ZN(n19635) );
  OAI211_X1 U22631 ( .C1(n19997), .C2(n19670), .A(n19636), .B(n19635), .ZN(
        P2_U3067) );
  AOI22_X1 U22632 ( .A1(n19645), .A2(n19549), .B1(n20070), .B2(n19644), .ZN(
        n19638) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19647), .B1(
        n19646), .B2(n19998), .ZN(n19637) );
  OAI211_X1 U22634 ( .C1(n20002), .C2(n19670), .A(n19638), .B(n19637), .ZN(
        P2_U3068) );
  AOI22_X1 U22635 ( .A1(n19645), .A2(n20076), .B1(n20075), .B2(n19644), .ZN(
        n19640) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19647), .B1(
        n19646), .B2(n19964), .ZN(n19639) );
  OAI211_X1 U22637 ( .C1(n19968), .C2(n19670), .A(n19640), .B(n19639), .ZN(
        P2_U3069) );
  AOI22_X1 U22638 ( .A1(n19645), .A2(n20082), .B1(n20081), .B2(n19644), .ZN(
        n19642) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19647), .B1(
        n19659), .B2(n20083), .ZN(n19641) );
  OAI211_X1 U22640 ( .C1(n20086), .C2(n19643), .A(n19642), .B(n19641), .ZN(
        P2_U3070) );
  AOI22_X1 U22641 ( .A1(n19645), .A2(n20089), .B1(n20087), .B2(n19644), .ZN(
        n19649) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19647), .B1(
        n19646), .B2(n19938), .ZN(n19648) );
  OAI211_X1 U22643 ( .C1(n19943), .C2(n19670), .A(n19649), .B(n19648), .ZN(
        P2_U3071) );
  AOI22_X1 U22644 ( .A1(n20060), .A2(n19700), .B1(n20059), .B2(n19665), .ZN(
        n19651) );
  AOI22_X1 U22645 ( .A1(n14355), .A2(n19666), .B1(n19659), .B2(n20033), .ZN(
        n19650) );
  OAI211_X1 U22646 ( .C1(n19664), .C2(n19652), .A(n19651), .B(n19650), .ZN(
        P2_U3074) );
  AOI22_X1 U22647 ( .A1(n20066), .A2(n19700), .B1(n19665), .B2(n20064), .ZN(
        n19654) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19667), .B1(
        n20065), .B2(n19666), .ZN(n19653) );
  OAI211_X1 U22649 ( .C1(n20069), .C2(n19670), .A(n19654), .B(n19653), .ZN(
        P2_U3075) );
  INV_X1 U22650 ( .A(n20002), .ZN(n20071) );
  AOI22_X1 U22651 ( .A1(n20071), .A2(n19700), .B1(n19665), .B2(n20070), .ZN(
        n19656) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19667), .B1(
        n19549), .B2(n19666), .ZN(n19655) );
  OAI211_X1 U22653 ( .C1(n20074), .C2(n19670), .A(n19656), .B(n19655), .ZN(
        P2_U3076) );
  AOI22_X1 U22654 ( .A1(n19964), .A2(n19659), .B1(n19665), .B2(n20075), .ZN(
        n19658) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19667), .B1(
        n20076), .B2(n19666), .ZN(n19657) );
  OAI211_X1 U22656 ( .C1(n19968), .C2(n19697), .A(n19658), .B(n19657), .ZN(
        P2_U3077) );
  AOI22_X1 U22657 ( .A1(n19660), .A2(n19659), .B1(n19665), .B2(n20081), .ZN(
        n19662) );
  AOI22_X1 U22658 ( .A1(n20082), .A2(n19666), .B1(n19700), .B2(n20083), .ZN(
        n19661) );
  OAI211_X1 U22659 ( .C1(n19664), .C2(n19663), .A(n19662), .B(n19661), .ZN(
        P2_U3078) );
  AOI22_X1 U22660 ( .A1(n20091), .A2(n19700), .B1(n19665), .B2(n20087), .ZN(
        n19669) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19667), .B1(
        n20089), .B2(n19666), .ZN(n19668) );
  OAI211_X1 U22662 ( .C1(n20097), .C2(n19670), .A(n19669), .B(n19668), .ZN(
        P2_U3079) );
  NOR3_X1 U22663 ( .A1(n21487), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19707) );
  NAND2_X1 U22664 ( .A1(n20233), .A2(n19707), .ZN(n19679) );
  INV_X1 U22665 ( .A(n19679), .ZN(n19698) );
  NOR3_X1 U22666 ( .A1(n19671), .A2(n19698), .A3(n19913), .ZN(n19678) );
  AND2_X1 U22667 ( .A1(n19673), .A2(n19672), .ZN(n19950) );
  INV_X1 U22668 ( .A(n19950), .ZN(n19945) );
  NOR2_X1 U22669 ( .A1(n19945), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19682) );
  AOI21_X1 U22670 ( .B1(n19873), .B2(n19682), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19674) );
  NOR2_X1 U22671 ( .A1(n19678), .A2(n19674), .ZN(n19699) );
  AOI22_X1 U22672 ( .A1(n19699), .A2(n14206), .B1(n20013), .B2(n19698), .ZN(
        n19684) );
  AOI21_X1 U22673 ( .B1(n19697), .B2(n19731), .A(n20197), .ZN(n19681) );
  AOI211_X1 U22674 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19679), .A(n19981), 
        .B(n19678), .ZN(n19680) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19701), .B1(
        n19718), .B2(n20014), .ZN(n19683) );
  OAI211_X1 U22676 ( .C1(n20028), .C2(n19697), .A(n19684), .B(n19683), .ZN(
        P2_U3080) );
  AOI22_X1 U22677 ( .A1(n19699), .A2(n14210), .B1(n20051), .B2(n19698), .ZN(
        n19686) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19701), .B1(
        n19700), .B2(n20053), .ZN(n19685) );
  OAI211_X1 U22679 ( .C1(n20031), .C2(n19731), .A(n19686), .B(n19685), .ZN(
        P2_U3081) );
  AOI22_X1 U22680 ( .A1(n19699), .A2(n14355), .B1(n20059), .B2(n19698), .ZN(
        n19688) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19701), .B1(
        n19718), .B2(n20060), .ZN(n19687) );
  OAI211_X1 U22682 ( .C1(n20063), .C2(n19697), .A(n19688), .B(n19687), .ZN(
        P2_U3082) );
  AOI22_X1 U22683 ( .A1(n19699), .A2(n20065), .B1(n20064), .B2(n19698), .ZN(
        n19690) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19701), .B1(
        n19700), .B2(n19994), .ZN(n19689) );
  OAI211_X1 U22685 ( .C1(n19997), .C2(n19731), .A(n19690), .B(n19689), .ZN(
        P2_U3083) );
  AOI22_X1 U22686 ( .A1(n19699), .A2(n19549), .B1(n20070), .B2(n19698), .ZN(
        n19692) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19701), .B1(
        n19718), .B2(n20071), .ZN(n19691) );
  OAI211_X1 U22688 ( .C1(n20074), .C2(n19697), .A(n19692), .B(n19691), .ZN(
        P2_U3084) );
  AOI22_X1 U22689 ( .A1(n19699), .A2(n20076), .B1(n20075), .B2(n19698), .ZN(
        n19694) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19701), .B1(
        n19718), .B2(n20077), .ZN(n19693) );
  OAI211_X1 U22691 ( .C1(n20080), .C2(n19697), .A(n19694), .B(n19693), .ZN(
        P2_U3085) );
  AOI22_X1 U22692 ( .A1(n19699), .A2(n20082), .B1(n20081), .B2(n19698), .ZN(
        n19696) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19701), .B1(
        n19718), .B2(n20083), .ZN(n19695) );
  OAI211_X1 U22694 ( .C1(n20086), .C2(n19697), .A(n19696), .B(n19695), .ZN(
        P2_U3086) );
  AOI22_X1 U22695 ( .A1(n19699), .A2(n20089), .B1(n20087), .B2(n19698), .ZN(
        n19703) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19701), .B1(
        n19700), .B2(n19938), .ZN(n19702) );
  OAI211_X1 U22697 ( .C1(n19943), .C2(n19731), .A(n19703), .B(n19702), .ZN(
        P2_U3087) );
  INV_X1 U22698 ( .A(n19707), .ZN(n19710) );
  NOR2_X1 U22699 ( .A1(n20233), .A2(n19710), .ZN(n19739) );
  AOI22_X1 U22700 ( .A1(n20014), .A2(n19755), .B1(n20013), .B2(n19739), .ZN(
        n19713) );
  INV_X1 U22701 ( .A(n19704), .ZN(n19774) );
  OAI21_X1 U22702 ( .B1(n19774), .B2(n19947), .A(n20206), .ZN(n19711) );
  INV_X1 U22703 ( .A(n19739), .ZN(n19705) );
  OAI211_X1 U22704 ( .C1(n12006), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19705), 
        .B(n20198), .ZN(n19706) );
  OAI211_X1 U22705 ( .C1(n19711), .C2(n19707), .A(n20020), .B(n19706), .ZN(
        n19728) );
  OAI21_X1 U22706 ( .B1(n19708), .B2(n19739), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19709) );
  OAI21_X1 U22707 ( .B1(n19711), .B2(n19710), .A(n19709), .ZN(n19727) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19728), .B1(
        n14206), .B2(n19727), .ZN(n19712) );
  OAI211_X1 U22709 ( .C1(n20028), .C2(n19731), .A(n19713), .B(n19712), .ZN(
        P2_U3088) );
  AOI22_X1 U22710 ( .A1(n20053), .A2(n19718), .B1(n20051), .B2(n19739), .ZN(
        n19715) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19728), .B1(
        n14210), .B2(n19727), .ZN(n19714) );
  OAI211_X1 U22712 ( .C1(n20031), .C2(n19765), .A(n19715), .B(n19714), .ZN(
        P2_U3089) );
  AOI22_X1 U22713 ( .A1(n20033), .A2(n19718), .B1(n20059), .B2(n19739), .ZN(
        n19717) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19728), .B1(
        n14355), .B2(n19727), .ZN(n19716) );
  OAI211_X1 U22715 ( .C1(n20036), .C2(n19765), .A(n19717), .B(n19716), .ZN(
        P2_U3090) );
  AOI22_X1 U22716 ( .A1(n19718), .A2(n19994), .B1(n19739), .B2(n20064), .ZN(
        n19720) );
  AOI22_X1 U22717 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19728), .B1(
        n20065), .B2(n19727), .ZN(n19719) );
  OAI211_X1 U22718 ( .C1(n19997), .C2(n19765), .A(n19720), .B(n19719), .ZN(
        P2_U3091) );
  AOI22_X1 U22719 ( .A1(n20071), .A2(n19755), .B1(n19739), .B2(n20070), .ZN(
        n19722) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19728), .B1(
        n19549), .B2(n19727), .ZN(n19721) );
  OAI211_X1 U22721 ( .C1(n20074), .C2(n19731), .A(n19722), .B(n19721), .ZN(
        P2_U3092) );
  AOI22_X1 U22722 ( .A1(n20077), .A2(n19755), .B1(n19739), .B2(n20075), .ZN(
        n19724) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19728), .B1(
        n20076), .B2(n19727), .ZN(n19723) );
  OAI211_X1 U22724 ( .C1(n20080), .C2(n19731), .A(n19724), .B(n19723), .ZN(
        P2_U3093) );
  AOI22_X1 U22725 ( .A1(n20083), .A2(n19755), .B1(n19739), .B2(n20081), .ZN(
        n19726) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19728), .B1(
        n20082), .B2(n19727), .ZN(n19725) );
  OAI211_X1 U22727 ( .C1(n20086), .C2(n19731), .A(n19726), .B(n19725), .ZN(
        P2_U3094) );
  AOI22_X1 U22728 ( .A1(n20091), .A2(n19755), .B1(n19739), .B2(n20087), .ZN(
        n19730) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19728), .B1(
        n20089), .B2(n19727), .ZN(n19729) );
  OAI211_X1 U22730 ( .C1(n20097), .C2(n19731), .A(n19730), .B(n19729), .ZN(
        P2_U3095) );
  AOI21_X1 U22731 ( .B1(n19765), .B2(n19821), .A(n20197), .ZN(n19733) );
  NOR2_X1 U22732 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20012), .ZN(
        n19778) );
  INV_X1 U22733 ( .A(n19778), .ZN(n19766) );
  NOR2_X1 U22734 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19766), .ZN(
        n19760) );
  AOI221_X1 U22735 ( .B1(n19739), .B2(n19873), .C1(n19733), .C2(n19873), .A(
        n19760), .ZN(n19738) );
  INV_X1 U22736 ( .A(n19760), .ZN(n19734) );
  NAND2_X1 U22737 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19734), .ZN(n19735) );
  OR2_X1 U22738 ( .A1(n19736), .A2(n19735), .ZN(n19742) );
  NAND2_X1 U22739 ( .A1(n19742), .A2(n20020), .ZN(n19737) );
  INV_X1 U22740 ( .A(n19762), .ZN(n19746) );
  INV_X1 U22741 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19745) );
  NOR2_X1 U22742 ( .A1(n19739), .A2(n19760), .ZN(n19740) );
  OAI21_X1 U22743 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19740), .A(n19913), 
        .ZN(n19741) );
  AND2_X1 U22744 ( .A1(n19742), .A2(n19741), .ZN(n19761) );
  AOI22_X1 U22745 ( .A1(n19761), .A2(n14206), .B1(n20013), .B2(n19760), .ZN(
        n19744) );
  AOI22_X1 U22746 ( .A1(n19791), .A2(n20014), .B1(n19755), .B2(n19883), .ZN(
        n19743) );
  OAI211_X1 U22747 ( .C1(n19746), .C2(n19745), .A(n19744), .B(n19743), .ZN(
        P2_U3096) );
  AOI22_X1 U22748 ( .A1(n19761), .A2(n14210), .B1(n20051), .B2(n19760), .ZN(
        n19748) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19762), .B1(
        n19755), .B2(n20053), .ZN(n19747) );
  OAI211_X1 U22750 ( .C1(n20031), .C2(n19821), .A(n19748), .B(n19747), .ZN(
        P2_U3097) );
  AOI22_X1 U22751 ( .A1(n19761), .A2(n14355), .B1(n20059), .B2(n19760), .ZN(
        n19750) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19762), .B1(
        n19791), .B2(n20060), .ZN(n19749) );
  OAI211_X1 U22753 ( .C1(n20063), .C2(n19765), .A(n19750), .B(n19749), .ZN(
        P2_U3098) );
  AOI22_X1 U22754 ( .A1(n19761), .A2(n20065), .B1(n20064), .B2(n19760), .ZN(
        n19752) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19762), .B1(
        n19755), .B2(n19994), .ZN(n19751) );
  OAI211_X1 U22756 ( .C1(n19997), .C2(n19821), .A(n19752), .B(n19751), .ZN(
        P2_U3099) );
  AOI22_X1 U22757 ( .A1(n19761), .A2(n19549), .B1(n20070), .B2(n19760), .ZN(
        n19754) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19762), .B1(
        n19791), .B2(n20071), .ZN(n19753) );
  OAI211_X1 U22759 ( .C1(n20074), .C2(n19765), .A(n19754), .B(n19753), .ZN(
        P2_U3100) );
  AOI22_X1 U22760 ( .A1(n19761), .A2(n20076), .B1(n20075), .B2(n19760), .ZN(
        n19757) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19762), .B1(
        n19755), .B2(n19964), .ZN(n19756) );
  OAI211_X1 U22762 ( .C1(n19968), .C2(n19821), .A(n19757), .B(n19756), .ZN(
        P2_U3101) );
  AOI22_X1 U22763 ( .A1(n19761), .A2(n20082), .B1(n20081), .B2(n19760), .ZN(
        n19759) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19762), .B1(
        n19791), .B2(n20083), .ZN(n19758) );
  OAI211_X1 U22765 ( .C1(n20086), .C2(n19765), .A(n19759), .B(n19758), .ZN(
        P2_U3102) );
  AOI22_X1 U22766 ( .A1(n19761), .A2(n20089), .B1(n20087), .B2(n19760), .ZN(
        n19764) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19762), .B1(
        n19791), .B2(n20091), .ZN(n19763) );
  OAI211_X1 U22768 ( .C1(n20097), .C2(n19765), .A(n19764), .B(n19763), .ZN(
        P2_U3103) );
  NOR2_X1 U22769 ( .A1(n20233), .A2(n19766), .ZN(n19829) );
  INV_X1 U22770 ( .A(n19829), .ZN(n19826) );
  NAND2_X1 U22771 ( .A1(n12007), .A2(n19826), .ZN(n19767) );
  MUX2_X1 U22772 ( .A(n19767), .B(n19778), .S(n19913), .Z(n19770) );
  INV_X1 U22773 ( .A(n19768), .ZN(n19769) );
  NAND2_X1 U22774 ( .A1(n19770), .A2(n19769), .ZN(n19816) );
  OAI22_X1 U22775 ( .A1(n19816), .A2(n19772), .B1(n19771), .B2(n19826), .ZN(
        n19773) );
  INV_X1 U22776 ( .A(n19773), .ZN(n19782) );
  NOR2_X1 U22777 ( .A1(n19774), .A2(n19779), .ZN(n20205) );
  OAI21_X1 U22778 ( .B1(n19775), .B2(n19913), .A(n19873), .ZN(n19776) );
  AOI21_X1 U22779 ( .B1(n19776), .B2(n19826), .A(n19981), .ZN(n19777) );
  OAI21_X1 U22780 ( .B1(n20205), .B2(n19778), .A(n19777), .ZN(n19818) );
  AOI22_X1 U22781 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19818), .B1(
        n19848), .B2(n20014), .ZN(n19781) );
  OAI211_X1 U22782 ( .C1(n20028), .C2(n19821), .A(n19782), .B(n19781), .ZN(
        P2_U3104) );
  OAI22_X1 U22783 ( .A1(n19816), .A2(n19784), .B1(n19783), .B2(n19826), .ZN(
        n19785) );
  INV_X1 U22784 ( .A(n19785), .ZN(n19787) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19818), .B1(
        n19791), .B2(n20053), .ZN(n19786) );
  OAI211_X1 U22786 ( .C1(n20031), .C2(n19846), .A(n19787), .B(n19786), .ZN(
        P2_U3105) );
  OAI22_X1 U22787 ( .A1(n19816), .A2(n19789), .B1(n19788), .B2(n19826), .ZN(
        n19790) );
  INV_X1 U22788 ( .A(n19790), .ZN(n19793) );
  AOI22_X1 U22789 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19818), .B1(
        n19791), .B2(n20033), .ZN(n19792) );
  OAI211_X1 U22790 ( .C1(n20036), .C2(n19846), .A(n19793), .B(n19792), .ZN(
        P2_U3106) );
  OAI22_X1 U22791 ( .A1(n19816), .A2(n19795), .B1(n19794), .B2(n19826), .ZN(
        n19796) );
  INV_X1 U22792 ( .A(n19796), .ZN(n19798) );
  AOI22_X1 U22793 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19818), .B1(
        n19848), .B2(n20066), .ZN(n19797) );
  OAI211_X1 U22794 ( .C1(n20069), .C2(n19821), .A(n19798), .B(n19797), .ZN(
        P2_U3107) );
  OAI22_X1 U22795 ( .A1(n19816), .A2(n19800), .B1(n19799), .B2(n19826), .ZN(
        n19801) );
  INV_X1 U22796 ( .A(n19801), .ZN(n19803) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19818), .B1(
        n19848), .B2(n20071), .ZN(n19802) );
  OAI211_X1 U22798 ( .C1(n20074), .C2(n19821), .A(n19803), .B(n19802), .ZN(
        P2_U3108) );
  OAI22_X1 U22799 ( .A1(n19816), .A2(n19805), .B1(n19804), .B2(n19826), .ZN(
        n19806) );
  INV_X1 U22800 ( .A(n19806), .ZN(n19808) );
  AOI22_X1 U22801 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19818), .B1(
        n19848), .B2(n20077), .ZN(n19807) );
  OAI211_X1 U22802 ( .C1(n20080), .C2(n19821), .A(n19808), .B(n19807), .ZN(
        P2_U3109) );
  OAI22_X1 U22803 ( .A1(n19816), .A2(n19810), .B1(n19809), .B2(n19826), .ZN(
        n19811) );
  INV_X1 U22804 ( .A(n19811), .ZN(n19813) );
  AOI22_X1 U22805 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19818), .B1(
        n19848), .B2(n20083), .ZN(n19812) );
  OAI211_X1 U22806 ( .C1(n20086), .C2(n19821), .A(n19813), .B(n19812), .ZN(
        P2_U3110) );
  OAI22_X1 U22807 ( .A1(n19816), .A2(n19815), .B1(n19814), .B2(n19826), .ZN(
        n19817) );
  INV_X1 U22808 ( .A(n19817), .ZN(n19820) );
  AOI22_X1 U22809 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19818), .B1(
        n19848), .B2(n20091), .ZN(n19819) );
  OAI211_X1 U22810 ( .C1(n20097), .C2(n19821), .A(n19820), .B(n19819), .ZN(
        P2_U3111) );
  NOR2_X1 U22811 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19822), .ZN(
        n19847) );
  AOI22_X1 U22812 ( .A1(n20014), .A2(n19857), .B1(n20013), .B2(n19847), .ZN(
        n19833) );
  AOI21_X1 U22813 ( .B1(n19870), .B2(n19846), .A(n20197), .ZN(n19823) );
  NOR2_X1 U22814 ( .A1(n19823), .A2(n20198), .ZN(n19828) );
  OAI21_X1 U22815 ( .B1(n11885), .B2(n19913), .A(n19873), .ZN(n19825) );
  AOI21_X1 U22816 ( .B1(n19828), .B2(n19826), .A(n19825), .ZN(n19827) );
  OAI21_X1 U22817 ( .B1(n19847), .B2(n19827), .A(n20020), .ZN(n19850) );
  OAI21_X1 U22818 ( .B1(n19847), .B2(n19829), .A(n19828), .ZN(n19831) );
  OAI21_X1 U22819 ( .B1(n11885), .B2(n19847), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19830) );
  NAND2_X1 U22820 ( .A1(n19831), .A2(n19830), .ZN(n19849) );
  AOI22_X1 U22821 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19850), .B1(
        n14206), .B2(n19849), .ZN(n19832) );
  OAI211_X1 U22822 ( .C1(n20028), .C2(n19846), .A(n19833), .B(n19832), .ZN(
        P2_U3112) );
  AOI22_X1 U22823 ( .A1(n20053), .A2(n19848), .B1(n20051), .B2(n19847), .ZN(
        n19835) );
  AOI22_X1 U22824 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n14210), .ZN(n19834) );
  OAI211_X1 U22825 ( .C1(n20031), .C2(n19870), .A(n19835), .B(n19834), .ZN(
        P2_U3113) );
  AOI22_X1 U22826 ( .A1(n19857), .A2(n20060), .B1(n20059), .B2(n19847), .ZN(
        n19837) );
  AOI22_X1 U22827 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n14355), .ZN(n19836) );
  OAI211_X1 U22828 ( .C1(n20063), .C2(n19846), .A(n19837), .B(n19836), .ZN(
        P2_U3114) );
  AOI22_X1 U22829 ( .A1(n19994), .A2(n19848), .B1(n20064), .B2(n19847), .ZN(
        n19839) );
  AOI22_X1 U22830 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20065), .ZN(n19838) );
  OAI211_X1 U22831 ( .C1(n19997), .C2(n19870), .A(n19839), .B(n19838), .ZN(
        P2_U3115) );
  AOI22_X1 U22832 ( .A1(n19998), .A2(n19848), .B1(n20070), .B2(n19847), .ZN(
        n19841) );
  AOI22_X1 U22833 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n19549), .ZN(n19840) );
  OAI211_X1 U22834 ( .C1(n20002), .C2(n19870), .A(n19841), .B(n19840), .ZN(
        P2_U3116) );
  AOI22_X1 U22835 ( .A1(n19964), .A2(n19848), .B1(n20075), .B2(n19847), .ZN(
        n19843) );
  AOI22_X1 U22836 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20076), .ZN(n19842) );
  OAI211_X1 U22837 ( .C1(n19968), .C2(n19870), .A(n19843), .B(n19842), .ZN(
        P2_U3117) );
  AOI22_X1 U22838 ( .A1(n20083), .A2(n19857), .B1(n20081), .B2(n19847), .ZN(
        n19845) );
  AOI22_X1 U22839 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20082), .ZN(n19844) );
  OAI211_X1 U22840 ( .C1(n20086), .C2(n19846), .A(n19845), .B(n19844), .ZN(
        P2_U3118) );
  AOI22_X1 U22841 ( .A1(n19938), .A2(n19848), .B1(n20087), .B2(n19847), .ZN(
        n19852) );
  AOI22_X1 U22842 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20089), .ZN(n19851) );
  OAI211_X1 U22843 ( .C1(n19943), .C2(n19870), .A(n19852), .B(n19851), .ZN(
        P2_U3119) );
  AOI22_X1 U22844 ( .A1(n20053), .A2(n19857), .B1(n20051), .B2(n19872), .ZN(
        n19854) );
  AOI22_X1 U22845 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19867), .B1(
        n14210), .B2(n19866), .ZN(n19853) );
  OAI211_X1 U22846 ( .C1(n20031), .C2(n19900), .A(n19854), .B(n19853), .ZN(
        P2_U3121) );
  AOI22_X1 U22847 ( .A1(n20033), .A2(n19857), .B1(n20059), .B2(n19872), .ZN(
        n19856) );
  AOI22_X1 U22848 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19867), .B1(
        n14355), .B2(n19866), .ZN(n19855) );
  OAI211_X1 U22849 ( .C1(n20036), .C2(n19900), .A(n19856), .B(n19855), .ZN(
        P2_U3122) );
  AOI22_X1 U22850 ( .A1(n19857), .A2(n19994), .B1(n19872), .B2(n20064), .ZN(
        n19859) );
  AOI22_X1 U22851 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19867), .B1(
        n20065), .B2(n19866), .ZN(n19858) );
  OAI211_X1 U22852 ( .C1(n19997), .C2(n19900), .A(n19859), .B(n19858), .ZN(
        P2_U3123) );
  AOI22_X1 U22853 ( .A1(n20071), .A2(n19903), .B1(n19872), .B2(n20070), .ZN(
        n19861) );
  AOI22_X1 U22854 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19867), .B1(
        n19549), .B2(n19866), .ZN(n19860) );
  OAI211_X1 U22855 ( .C1(n20074), .C2(n19870), .A(n19861), .B(n19860), .ZN(
        P2_U3124) );
  AOI22_X1 U22856 ( .A1(n20077), .A2(n19903), .B1(n19872), .B2(n20075), .ZN(
        n19863) );
  AOI22_X1 U22857 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19867), .B1(
        n20076), .B2(n19866), .ZN(n19862) );
  OAI211_X1 U22858 ( .C1(n20080), .C2(n19870), .A(n19863), .B(n19862), .ZN(
        P2_U3125) );
  AOI22_X1 U22859 ( .A1(n20083), .A2(n19903), .B1(n19872), .B2(n20081), .ZN(
        n19865) );
  AOI22_X1 U22860 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19867), .B1(
        n20082), .B2(n19866), .ZN(n19864) );
  OAI211_X1 U22861 ( .C1(n20086), .C2(n19870), .A(n19865), .B(n19864), .ZN(
        P2_U3126) );
  AOI22_X1 U22862 ( .A1(n19903), .A2(n20091), .B1(n19872), .B2(n20087), .ZN(
        n19869) );
  AOI22_X1 U22863 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19867), .B1(
        n20089), .B2(n19866), .ZN(n19868) );
  OAI211_X1 U22864 ( .C1(n20097), .C2(n19870), .A(n19869), .B(n19868), .ZN(
        P2_U3127) );
  INV_X1 U22865 ( .A(n20199), .ZN(n19871) );
  AOI221_X1 U22866 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19939), .C1(
        P2_STATEBS16_REG_SCAN_IN), .C2(n19903), .A(n19872), .ZN(n19875) );
  INV_X1 U22867 ( .A(n12016), .ZN(n19880) );
  AOI21_X1 U22868 ( .B1(n19880), .B2(n19873), .A(n20206), .ZN(n19874) );
  OR2_X1 U22869 ( .A1(n19875), .A2(n19874), .ZN(n19877) );
  NAND2_X1 U22870 ( .A1(n19876), .A2(n19908), .ZN(n19879) );
  NAND2_X1 U22871 ( .A1(n19877), .A2(n19879), .ZN(n19878) );
  AND2_X1 U22872 ( .A1(n19878), .A2(n20020), .ZN(n19889) );
  INV_X1 U22873 ( .A(n19879), .ZN(n19901) );
  OAI21_X1 U22874 ( .B1(n19880), .B2(n19901), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19881) );
  OAI21_X1 U22875 ( .B1(n19912), .B2(n19882), .A(n19881), .ZN(n19902) );
  AOI22_X1 U22876 ( .A1(n19902), .A2(n14206), .B1(n20013), .B2(n19901), .ZN(
        n19885) );
  AOI22_X1 U22877 ( .A1(n19939), .A2(n20014), .B1(n19903), .B2(n19883), .ZN(
        n19884) );
  OAI211_X1 U22878 ( .C1(n19889), .C2(n19886), .A(n19885), .B(n19884), .ZN(
        P2_U3128) );
  AOI22_X1 U22879 ( .A1(n19902), .A2(n14210), .B1(n20051), .B2(n19901), .ZN(
        n19888) );
  AOI22_X1 U22880 ( .A1(n19903), .A2(n20053), .B1(n19939), .B2(n20052), .ZN(
        n19887) );
  OAI211_X1 U22881 ( .C1(n19889), .C2(n13466), .A(n19888), .B(n19887), .ZN(
        P2_U3129) );
  AOI22_X1 U22882 ( .A1(n19902), .A2(n14355), .B1(n20059), .B2(n19901), .ZN(
        n19891) );
  AOI22_X1 U22883 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19904), .B1(
        n19939), .B2(n20060), .ZN(n19890) );
  OAI211_X1 U22884 ( .C1(n20063), .C2(n19900), .A(n19891), .B(n19890), .ZN(
        P2_U3130) );
  AOI22_X1 U22885 ( .A1(n19902), .A2(n20065), .B1(n20064), .B2(n19901), .ZN(
        n19893) );
  AOI22_X1 U22886 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19904), .B1(
        n19903), .B2(n19994), .ZN(n19892) );
  OAI211_X1 U22887 ( .C1(n19997), .C2(n19935), .A(n19893), .B(n19892), .ZN(
        P2_U3131) );
  AOI22_X1 U22888 ( .A1(n19902), .A2(n19549), .B1(n20070), .B2(n19901), .ZN(
        n19895) );
  AOI22_X1 U22889 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19904), .B1(
        n19903), .B2(n19998), .ZN(n19894) );
  OAI211_X1 U22890 ( .C1(n20002), .C2(n19935), .A(n19895), .B(n19894), .ZN(
        P2_U3132) );
  AOI22_X1 U22891 ( .A1(n19902), .A2(n20076), .B1(n20075), .B2(n19901), .ZN(
        n19897) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19904), .B1(
        n19903), .B2(n19964), .ZN(n19896) );
  OAI211_X1 U22893 ( .C1(n19968), .C2(n19935), .A(n19897), .B(n19896), .ZN(
        P2_U3133) );
  AOI22_X1 U22894 ( .A1(n19902), .A2(n20082), .B1(n20081), .B2(n19901), .ZN(
        n19899) );
  AOI22_X1 U22895 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19904), .B1(
        n19939), .B2(n20083), .ZN(n19898) );
  OAI211_X1 U22896 ( .C1(n20086), .C2(n19900), .A(n19899), .B(n19898), .ZN(
        P2_U3134) );
  AOI22_X1 U22897 ( .A1(n19902), .A2(n20089), .B1(n20087), .B2(n19901), .ZN(
        n19906) );
  AOI22_X1 U22898 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19904), .B1(
        n19903), .B2(n19938), .ZN(n19905) );
  OAI211_X1 U22899 ( .C1(n19943), .C2(n19935), .A(n19906), .B(n19905), .ZN(
        P2_U3135) );
  INV_X1 U22900 ( .A(n19907), .ZN(n19909) );
  NAND2_X1 U22901 ( .A1(n19909), .A2(n19908), .ZN(n19916) );
  AND2_X1 U22902 ( .A1(n19916), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19910) );
  NAND2_X1 U22903 ( .A1(n19911), .A2(n19910), .ZN(n19917) );
  NOR2_X1 U22904 ( .A1(n21540), .A2(n19912), .ZN(n19920) );
  INV_X1 U22905 ( .A(n19920), .ZN(n19914) );
  OAI21_X1 U22906 ( .B1(n19914), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19913), 
        .ZN(n19915) );
  AND2_X1 U22907 ( .A1(n19917), .A2(n19915), .ZN(n19937) );
  INV_X1 U22908 ( .A(n19916), .ZN(n19936) );
  AOI22_X1 U22909 ( .A1(n19937), .A2(n14206), .B1(n20013), .B2(n19936), .ZN(
        n19922) );
  OAI211_X1 U22910 ( .C1(n19936), .C2(n19873), .A(n19917), .B(n20020), .ZN(
        n19918) );
  INV_X1 U22911 ( .A(n19918), .ZN(n19919) );
  OAI221_X1 U22912 ( .B1(n19920), .B2(n20199), .C1(n19920), .C2(n19984), .A(
        n19919), .ZN(n19940) );
  NAND2_X1 U22913 ( .A1(n19987), .A2(n20199), .ZN(n19976) );
  AOI22_X1 U22914 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19940), .B1(
        n19965), .B2(n20014), .ZN(n19921) );
  OAI211_X1 U22915 ( .C1(n20028), .C2(n19935), .A(n19922), .B(n19921), .ZN(
        P2_U3136) );
  AOI22_X1 U22916 ( .A1(n19937), .A2(n14210), .B1(n20051), .B2(n19936), .ZN(
        n19924) );
  AOI22_X1 U22917 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n20053), .ZN(n19923) );
  OAI211_X1 U22918 ( .C1(n20031), .C2(n19976), .A(n19924), .B(n19923), .ZN(
        P2_U3137) );
  AOI22_X1 U22919 ( .A1(n19937), .A2(n14355), .B1(n20059), .B2(n19936), .ZN(
        n19926) );
  AOI22_X1 U22920 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n20033), .ZN(n19925) );
  OAI211_X1 U22921 ( .C1(n20036), .C2(n19976), .A(n19926), .B(n19925), .ZN(
        P2_U3138) );
  AOI22_X1 U22922 ( .A1(n19937), .A2(n20065), .B1(n20064), .B2(n19936), .ZN(
        n19928) );
  AOI22_X1 U22923 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19940), .B1(
        n19965), .B2(n20066), .ZN(n19927) );
  OAI211_X1 U22924 ( .C1(n20069), .C2(n19935), .A(n19928), .B(n19927), .ZN(
        P2_U3139) );
  AOI22_X1 U22925 ( .A1(n19937), .A2(n19549), .B1(n20070), .B2(n19936), .ZN(
        n19930) );
  AOI22_X1 U22926 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n19998), .ZN(n19929) );
  OAI211_X1 U22927 ( .C1(n20002), .C2(n19976), .A(n19930), .B(n19929), .ZN(
        P2_U3140) );
  AOI22_X1 U22928 ( .A1(n19937), .A2(n20076), .B1(n20075), .B2(n19936), .ZN(
        n19932) );
  AOI22_X1 U22929 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19940), .B1(
        n19965), .B2(n20077), .ZN(n19931) );
  OAI211_X1 U22930 ( .C1(n20080), .C2(n19935), .A(n19932), .B(n19931), .ZN(
        P2_U3141) );
  AOI22_X1 U22931 ( .A1(n19937), .A2(n20082), .B1(n20081), .B2(n19936), .ZN(
        n19934) );
  AOI22_X1 U22932 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19940), .B1(
        n19965), .B2(n20083), .ZN(n19933) );
  OAI211_X1 U22933 ( .C1(n20086), .C2(n19935), .A(n19934), .B(n19933), .ZN(
        P2_U3142) );
  AOI22_X1 U22934 ( .A1(n19937), .A2(n20089), .B1(n20087), .B2(n19936), .ZN(
        n19942) );
  AOI22_X1 U22935 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n19938), .ZN(n19941) );
  OAI211_X1 U22936 ( .C1(n19943), .C2(n19976), .A(n19942), .B(n19941), .ZN(
        P2_U3143) );
  NAND3_X1 U22937 ( .A1(n21540), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19978) );
  NOR2_X1 U22938 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19978), .ZN(
        n19971) );
  NOR2_X1 U22939 ( .A1(n12015), .A2(n19971), .ZN(n19952) );
  INV_X1 U22940 ( .A(n19944), .ZN(n19946) );
  OAI22_X1 U22941 ( .A1(n19952), .A2(n19913), .B1(n19946), .B2(n19945), .ZN(
        n19972) );
  AOI22_X1 U22942 ( .A1(n19972), .A2(n14206), .B1(n20013), .B2(n19971), .ZN(
        n19955) );
  AOI21_X1 U22943 ( .B1(n20011), .B2(n19976), .A(n20197), .ZN(n19949) );
  AOI21_X1 U22944 ( .B1(n19950), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19949), .ZN(n19951) );
  AOI211_X1 U22945 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19952), .A(n19981), 
        .B(n19951), .ZN(n19953) );
  AOI22_X1 U22946 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19973), .B1(
        n19999), .B2(n20014), .ZN(n19954) );
  OAI211_X1 U22947 ( .C1(n20028), .C2(n19976), .A(n19955), .B(n19954), .ZN(
        P2_U3144) );
  AOI22_X1 U22948 ( .A1(n19972), .A2(n14210), .B1(n20051), .B2(n19971), .ZN(
        n19957) );
  AOI22_X1 U22949 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19973), .B1(
        n19965), .B2(n20053), .ZN(n19956) );
  OAI211_X1 U22950 ( .C1(n20031), .C2(n20011), .A(n19957), .B(n19956), .ZN(
        P2_U3145) );
  AOI22_X1 U22951 ( .A1(n19972), .A2(n14355), .B1(n20059), .B2(n19971), .ZN(
        n19959) );
  AOI22_X1 U22952 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19973), .B1(
        n19965), .B2(n20033), .ZN(n19958) );
  OAI211_X1 U22953 ( .C1(n20036), .C2(n20011), .A(n19959), .B(n19958), .ZN(
        P2_U3146) );
  AOI22_X1 U22954 ( .A1(n19972), .A2(n20065), .B1(n20064), .B2(n19971), .ZN(
        n19961) );
  AOI22_X1 U22955 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19973), .B1(
        n19965), .B2(n19994), .ZN(n19960) );
  OAI211_X1 U22956 ( .C1(n19997), .C2(n20011), .A(n19961), .B(n19960), .ZN(
        P2_U3147) );
  AOI22_X1 U22957 ( .A1(n19972), .A2(n19549), .B1(n20070), .B2(n19971), .ZN(
        n19963) );
  AOI22_X1 U22958 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19973), .B1(
        n19965), .B2(n19998), .ZN(n19962) );
  OAI211_X1 U22959 ( .C1(n20002), .C2(n20011), .A(n19963), .B(n19962), .ZN(
        P2_U3148) );
  AOI22_X1 U22960 ( .A1(n19972), .A2(n20076), .B1(n20075), .B2(n19971), .ZN(
        n19967) );
  AOI22_X1 U22961 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19973), .B1(
        n19965), .B2(n19964), .ZN(n19966) );
  OAI211_X1 U22962 ( .C1(n19968), .C2(n20011), .A(n19967), .B(n19966), .ZN(
        P2_U3149) );
  AOI22_X1 U22963 ( .A1(n19972), .A2(n20082), .B1(n20081), .B2(n19971), .ZN(
        n19970) );
  AOI22_X1 U22964 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19973), .B1(
        n19999), .B2(n20083), .ZN(n19969) );
  OAI211_X1 U22965 ( .C1(n20086), .C2(n19976), .A(n19970), .B(n19969), .ZN(
        P2_U3150) );
  AOI22_X1 U22966 ( .A1(n19972), .A2(n20089), .B1(n20087), .B2(n19971), .ZN(
        n19975) );
  AOI22_X1 U22967 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19973), .B1(
        n19999), .B2(n20091), .ZN(n19974) );
  OAI211_X1 U22968 ( .C1(n20097), .C2(n19976), .A(n19975), .B(n19974), .ZN(
        P2_U3151) );
  NOR2_X1 U22969 ( .A1(n20233), .A2(n19978), .ZN(n20016) );
  NOR3_X1 U22970 ( .A1(n19977), .A2(n20016), .A3(n19913), .ZN(n19980) );
  INV_X1 U22971 ( .A(n19978), .ZN(n19985) );
  AOI21_X1 U22972 ( .B1(n19873), .B2(n19985), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19979) );
  NOR2_X1 U22973 ( .A1(n19980), .A2(n19979), .ZN(n20007) );
  AOI22_X1 U22974 ( .A1(n20007), .A2(n14206), .B1(n20013), .B2(n20016), .ZN(
        n19989) );
  INV_X1 U22975 ( .A(n20016), .ZN(n19982) );
  AOI211_X1 U22976 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19982), .A(n19981), 
        .B(n19980), .ZN(n19983) );
  OAI221_X1 U22977 ( .B1(n19985), .B2(n19986), .C1(n19985), .C2(n19984), .A(
        n19983), .ZN(n20008) );
  AOI22_X1 U22978 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20008), .B1(
        n20032), .B2(n20014), .ZN(n19988) );
  OAI211_X1 U22979 ( .C1(n20028), .C2(n20011), .A(n19989), .B(n19988), .ZN(
        P2_U3152) );
  AOI22_X1 U22980 ( .A1(n20007), .A2(n14210), .B1(n20051), .B2(n20016), .ZN(
        n19991) );
  AOI22_X1 U22981 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20008), .B1(
        n19999), .B2(n20053), .ZN(n19990) );
  OAI211_X1 U22982 ( .C1(n20031), .C2(n20050), .A(n19991), .B(n19990), .ZN(
        P2_U3153) );
  AOI22_X1 U22983 ( .A1(n20007), .A2(n14355), .B1(n20059), .B2(n20016), .ZN(
        n19993) );
  AOI22_X1 U22984 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20008), .B1(
        n20032), .B2(n20060), .ZN(n19992) );
  OAI211_X1 U22985 ( .C1(n20063), .C2(n20011), .A(n19993), .B(n19992), .ZN(
        P2_U3154) );
  AOI22_X1 U22986 ( .A1(n20007), .A2(n20065), .B1(n20064), .B2(n20016), .ZN(
        n19996) );
  AOI22_X1 U22987 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20008), .B1(
        n19999), .B2(n19994), .ZN(n19995) );
  OAI211_X1 U22988 ( .C1(n19997), .C2(n20050), .A(n19996), .B(n19995), .ZN(
        P2_U3155) );
  AOI22_X1 U22989 ( .A1(n20007), .A2(n19549), .B1(n20070), .B2(n20016), .ZN(
        n20001) );
  AOI22_X1 U22990 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20008), .B1(
        n19999), .B2(n19998), .ZN(n20000) );
  OAI211_X1 U22991 ( .C1(n20002), .C2(n20050), .A(n20001), .B(n20000), .ZN(
        P2_U3156) );
  AOI22_X1 U22992 ( .A1(n20007), .A2(n20076), .B1(n20075), .B2(n20016), .ZN(
        n20004) );
  AOI22_X1 U22993 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20008), .B1(
        n20032), .B2(n20077), .ZN(n20003) );
  OAI211_X1 U22994 ( .C1(n20080), .C2(n20011), .A(n20004), .B(n20003), .ZN(
        P2_U3157) );
  AOI22_X1 U22995 ( .A1(n20007), .A2(n20082), .B1(n20081), .B2(n20016), .ZN(
        n20006) );
  AOI22_X1 U22996 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20008), .B1(
        n20032), .B2(n20083), .ZN(n20005) );
  OAI211_X1 U22997 ( .C1(n20086), .C2(n20011), .A(n20006), .B(n20005), .ZN(
        P2_U3158) );
  AOI22_X1 U22998 ( .A1(n20007), .A2(n20089), .B1(n20087), .B2(n20016), .ZN(
        n20010) );
  AOI22_X1 U22999 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20008), .B1(
        n20032), .B2(n20091), .ZN(n20009) );
  OAI211_X1 U23000 ( .C1(n20097), .C2(n20011), .A(n20010), .B(n20009), .ZN(
        P2_U3159) );
  NOR3_X2 U23001 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20209), .A3(
        n20012), .ZN(n20045) );
  AOI22_X1 U23002 ( .A1(n20014), .A2(n20054), .B1(n20013), .B2(n20045), .ZN(
        n20027) );
  OAI21_X1 U23003 ( .B1(n20032), .B2(n20054), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20015) );
  NAND2_X1 U23004 ( .A1(n20015), .A2(n20206), .ZN(n20025) );
  NOR2_X1 U23005 ( .A1(n20045), .A2(n20016), .ZN(n20024) );
  INV_X1 U23006 ( .A(n20024), .ZN(n20021) );
  INV_X1 U23007 ( .A(n20022), .ZN(n20018) );
  INV_X1 U23008 ( .A(n20045), .ZN(n20017) );
  OAI211_X1 U23009 ( .C1(n20018), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20017), 
        .B(n20198), .ZN(n20019) );
  OAI211_X1 U23010 ( .C1(n20025), .C2(n20021), .A(n20020), .B(n20019), .ZN(
        n20047) );
  OAI21_X1 U23011 ( .B1(n20022), .B2(n20045), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20023) );
  AOI22_X1 U23012 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20047), .B1(
        n14206), .B2(n20046), .ZN(n20026) );
  OAI211_X1 U23013 ( .C1(n20028), .C2(n20050), .A(n20027), .B(n20026), .ZN(
        P2_U3160) );
  AOI22_X1 U23014 ( .A1(n20053), .A2(n20032), .B1(n20051), .B2(n20045), .ZN(
        n20030) );
  AOI22_X1 U23015 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20047), .B1(
        n14210), .B2(n20046), .ZN(n20029) );
  OAI211_X1 U23016 ( .C1(n20031), .C2(n20096), .A(n20030), .B(n20029), .ZN(
        P2_U3161) );
  AOI22_X1 U23017 ( .A1(n20033), .A2(n20032), .B1(n20059), .B2(n20045), .ZN(
        n20035) );
  AOI22_X1 U23018 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20047), .B1(
        n14355), .B2(n20046), .ZN(n20034) );
  OAI211_X1 U23019 ( .C1(n20036), .C2(n20096), .A(n20035), .B(n20034), .ZN(
        P2_U3162) );
  AOI22_X1 U23020 ( .A1(n20066), .A2(n20054), .B1(n20064), .B2(n20045), .ZN(
        n20038) );
  AOI22_X1 U23021 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20047), .B1(
        n20065), .B2(n20046), .ZN(n20037) );
  OAI211_X1 U23022 ( .C1(n20069), .C2(n20050), .A(n20038), .B(n20037), .ZN(
        P2_U3163) );
  AOI22_X1 U23023 ( .A1(n20054), .A2(n20071), .B1(n20070), .B2(n20045), .ZN(
        n20040) );
  AOI22_X1 U23024 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20047), .B1(
        n19549), .B2(n20046), .ZN(n20039) );
  OAI211_X1 U23025 ( .C1(n20074), .C2(n20050), .A(n20040), .B(n20039), .ZN(
        P2_U3164) );
  AOI22_X1 U23026 ( .A1(n20077), .A2(n20054), .B1(n20075), .B2(n20045), .ZN(
        n20042) );
  AOI22_X1 U23027 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20047), .B1(
        n20076), .B2(n20046), .ZN(n20041) );
  OAI211_X1 U23028 ( .C1(n20080), .C2(n20050), .A(n20042), .B(n20041), .ZN(
        P2_U3165) );
  AOI22_X1 U23029 ( .A1(n20083), .A2(n20054), .B1(n20081), .B2(n20045), .ZN(
        n20044) );
  AOI22_X1 U23030 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20047), .B1(
        n20082), .B2(n20046), .ZN(n20043) );
  OAI211_X1 U23031 ( .C1(n20086), .C2(n20050), .A(n20044), .B(n20043), .ZN(
        P2_U3166) );
  AOI22_X1 U23032 ( .A1(n20054), .A2(n20091), .B1(n20087), .B2(n20045), .ZN(
        n20049) );
  AOI22_X1 U23033 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20047), .B1(
        n20089), .B2(n20046), .ZN(n20048) );
  OAI211_X1 U23034 ( .C1(n20097), .C2(n20050), .A(n20049), .B(n20048), .ZN(
        P2_U3167) );
  AOI22_X1 U23035 ( .A1(n20090), .A2(n14210), .B1(n20088), .B2(n20051), .ZN(
        n20056) );
  AOI22_X1 U23036 ( .A1(n20054), .A2(n20053), .B1(n20092), .B2(n20052), .ZN(
        n20055) );
  OAI211_X1 U23037 ( .C1(n20058), .C2(n20057), .A(n20056), .B(n20055), .ZN(
        P2_U3169) );
  AOI22_X1 U23038 ( .A1(n20090), .A2(n14355), .B1(n20088), .B2(n20059), .ZN(
        n20062) );
  AOI22_X1 U23039 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20093), .B1(
        n20092), .B2(n20060), .ZN(n20061) );
  OAI211_X1 U23040 ( .C1(n20063), .C2(n20096), .A(n20062), .B(n20061), .ZN(
        P2_U3170) );
  AOI22_X1 U23041 ( .A1(n20090), .A2(n20065), .B1(n20088), .B2(n20064), .ZN(
        n20068) );
  AOI22_X1 U23042 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20093), .B1(
        n20092), .B2(n20066), .ZN(n20067) );
  OAI211_X1 U23043 ( .C1(n20069), .C2(n20096), .A(n20068), .B(n20067), .ZN(
        P2_U3171) );
  AOI22_X1 U23044 ( .A1(n20090), .A2(n19549), .B1(n20088), .B2(n20070), .ZN(
        n20073) );
  AOI22_X1 U23045 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20093), .B1(
        n20092), .B2(n20071), .ZN(n20072) );
  OAI211_X1 U23046 ( .C1(n20074), .C2(n20096), .A(n20073), .B(n20072), .ZN(
        P2_U3172) );
  AOI22_X1 U23047 ( .A1(n20090), .A2(n20076), .B1(n20088), .B2(n20075), .ZN(
        n20079) );
  AOI22_X1 U23048 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20093), .B1(
        n20092), .B2(n20077), .ZN(n20078) );
  OAI211_X1 U23049 ( .C1(n20080), .C2(n20096), .A(n20079), .B(n20078), .ZN(
        P2_U3173) );
  AOI22_X1 U23050 ( .A1(n20090), .A2(n20082), .B1(n20088), .B2(n20081), .ZN(
        n20085) );
  AOI22_X1 U23051 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20093), .B1(
        n20092), .B2(n20083), .ZN(n20084) );
  OAI211_X1 U23052 ( .C1(n20086), .C2(n20096), .A(n20085), .B(n20084), .ZN(
        P2_U3174) );
  AOI22_X1 U23053 ( .A1(n20090), .A2(n20089), .B1(n20088), .B2(n20087), .ZN(
        n20095) );
  AOI22_X1 U23054 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20093), .B1(
        n20092), .B2(n20091), .ZN(n20094) );
  OAI211_X1 U23055 ( .C1(n20097), .C2(n20096), .A(n20095), .B(n20094), .ZN(
        P2_U3175) );
  OAI21_X1 U23056 ( .B1(n20200), .B2(n20099), .A(n20098), .ZN(n20103) );
  AOI211_X1 U23057 ( .C1(n20104), .C2(n20100), .A(n20108), .B(n15818), .ZN(
        n20101) );
  AOI211_X1 U23058 ( .C1(n20104), .C2(n20103), .A(n20102), .B(n20101), .ZN(
        n20105) );
  INV_X1 U23059 ( .A(n20105), .ZN(P2_U3177) );
  AND2_X1 U23060 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20107), .ZN(
        P2_U3179) );
  AND2_X1 U23061 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20107), .ZN(
        P2_U3180) );
  AND2_X1 U23062 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20107), .ZN(
        P2_U3181) );
  AND2_X1 U23063 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20107), .ZN(
        P2_U3182) );
  AND2_X1 U23064 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20107), .ZN(
        P2_U3183) );
  AND2_X1 U23065 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20107), .ZN(
        P2_U3184) );
  AND2_X1 U23066 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20107), .ZN(
        P2_U3185) );
  AND2_X1 U23067 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20107), .ZN(
        P2_U3186) );
  AND2_X1 U23068 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20107), .ZN(
        P2_U3187) );
  AND2_X1 U23069 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20107), .ZN(
        P2_U3188) );
  AND2_X1 U23070 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20107), .ZN(
        P2_U3189) );
  AND2_X1 U23071 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20107), .ZN(
        P2_U3190) );
  AND2_X1 U23072 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20107), .ZN(
        P2_U3191) );
  AND2_X1 U23073 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20107), .ZN(
        P2_U3192) );
  AND2_X1 U23074 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20107), .ZN(
        P2_U3193) );
  AND2_X1 U23075 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20107), .ZN(
        P2_U3194) );
  AND2_X1 U23076 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20107), .ZN(
        P2_U3195) );
  AND2_X1 U23077 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20107), .ZN(
        P2_U3196) );
  AND2_X1 U23078 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20107), .ZN(
        P2_U3197) );
  NOR2_X1 U23079 ( .A1(n21541), .A2(n20196), .ZN(P2_U3198) );
  AND2_X1 U23080 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20107), .ZN(
        P2_U3199) );
  NOR2_X1 U23081 ( .A1(n20106), .A2(n20196), .ZN(P2_U3200) );
  AND2_X1 U23082 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20107), .ZN(P2_U3201) );
  AND2_X1 U23083 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20107), .ZN(P2_U3202) );
  AND2_X1 U23084 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20107), .ZN(P2_U3203) );
  AND2_X1 U23085 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20107), .ZN(P2_U3204) );
  AND2_X1 U23086 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20107), .ZN(P2_U3205) );
  AND2_X1 U23087 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20107), .ZN(P2_U3206) );
  AND2_X1 U23088 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20107), .ZN(P2_U3207) );
  AND2_X1 U23089 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20107), .ZN(P2_U3208) );
  NOR2_X1 U23090 ( .A1(n20108), .A2(n20122), .ZN(n20119) );
  OR3_X1 U23091 ( .A1(n20119), .A2(n20120), .A3(n20109), .ZN(n20111) );
  AOI211_X1 U23092 ( .C1(n20118), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n20121), .B(n20246), .ZN(n20110) );
  NOR3_X1 U23093 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21130), .ZN(n20127) );
  AOI211_X1 U23094 ( .C1(n20130), .C2(n20111), .A(n20110), .B(n20127), .ZN(
        n20112) );
  INV_X1 U23095 ( .A(n20112), .ZN(P2_U3209) );
  AOI21_X1 U23096 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20118), .A(n20130), 
        .ZN(n20123) );
  NOR3_X1 U23097 ( .A1(n20123), .A2(n20120), .A3(n20109), .ZN(n20113) );
  NOR2_X1 U23098 ( .A1(n20113), .A2(n20119), .ZN(n20116) );
  INV_X1 U23099 ( .A(n20114), .ZN(n20115) );
  OAI211_X1 U23100 ( .C1(n20118), .C2(n20117), .A(n20116), .B(n20115), .ZN(
        P2_U3210) );
  AOI22_X1 U23101 ( .A1(n20121), .A2(n20120), .B1(n20119), .B2(n21130), .ZN(
        n20129) );
  OAI21_X1 U23102 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20128) );
  NOR2_X1 U23103 ( .A1(n20122), .A2(n20130), .ZN(n20125) );
  AOI21_X1 U23104 ( .B1(n20125), .B2(n20124), .A(n20123), .ZN(n20126) );
  OAI22_X1 U23105 ( .A1(n20129), .A2(n20128), .B1(n20127), .B2(n20126), .ZN(
        P2_U3211) );
  OAI222_X1 U23106 ( .A1(n20186), .A2(n20132), .B1(n20131), .B2(n20246), .C1(
        n20133), .C2(n20185), .ZN(P2_U3212) );
  OAI222_X1 U23107 ( .A1(n20185), .A2(n20135), .B1(n20134), .B2(n20246), .C1(
        n20133), .C2(n20186), .ZN(P2_U3213) );
  INV_X1 U23108 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20137) );
  OAI222_X1 U23109 ( .A1(n20185), .A2(n20137), .B1(n20136), .B2(n20246), .C1(
        n20135), .C2(n20186), .ZN(P2_U3214) );
  OAI222_X1 U23110 ( .A1(n20185), .A2(n20139), .B1(n20138), .B2(n20246), .C1(
        n20137), .C2(n20186), .ZN(P2_U3215) );
  OAI222_X1 U23111 ( .A1(n20185), .A2(n20141), .B1(n20140), .B2(n20246), .C1(
        n20139), .C2(n20186), .ZN(P2_U3216) );
  OAI222_X1 U23112 ( .A1(n20185), .A2(n20143), .B1(n20142), .B2(n20246), .C1(
        n20141), .C2(n20186), .ZN(P2_U3217) );
  INV_X1 U23113 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20144) );
  OAI222_X1 U23114 ( .A1(n20185), .A2(n20144), .B1(n21517), .B2(n20246), .C1(
        n20143), .C2(n20186), .ZN(P2_U3218) );
  OAI222_X1 U23115 ( .A1(n20185), .A2(n20146), .B1(n20145), .B2(n20246), .C1(
        n20144), .C2(n20186), .ZN(P2_U3219) );
  OAI222_X1 U23116 ( .A1(n20185), .A2(n20148), .B1(n20147), .B2(n20246), .C1(
        n20146), .C2(n20186), .ZN(P2_U3220) );
  OAI222_X1 U23117 ( .A1(n20185), .A2(n20150), .B1(n20149), .B2(n20246), .C1(
        n20148), .C2(n20186), .ZN(P2_U3221) );
  OAI222_X1 U23118 ( .A1(n20185), .A2(n20152), .B1(n20151), .B2(n20246), .C1(
        n20150), .C2(n20186), .ZN(P2_U3222) );
  OAI222_X1 U23119 ( .A1(n20185), .A2(n20154), .B1(n20153), .B2(n20246), .C1(
        n20152), .C2(n20186), .ZN(P2_U3223) );
  OAI222_X1 U23120 ( .A1(n20185), .A2(n20156), .B1(n20155), .B2(n20246), .C1(
        n20154), .C2(n20186), .ZN(P2_U3224) );
  OAI222_X1 U23121 ( .A1(n20185), .A2(n20158), .B1(n20157), .B2(n20246), .C1(
        n20156), .C2(n20186), .ZN(P2_U3225) );
  INV_X1 U23122 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20160) );
  OAI222_X1 U23123 ( .A1(n20185), .A2(n20160), .B1(n20159), .B2(n20246), .C1(
        n20158), .C2(n20186), .ZN(P2_U3226) );
  OAI222_X1 U23124 ( .A1(n20185), .A2(n20162), .B1(n20161), .B2(n20246), .C1(
        n20160), .C2(n20186), .ZN(P2_U3227) );
  OAI222_X1 U23125 ( .A1(n20185), .A2(n20164), .B1(n20163), .B2(n20246), .C1(
        n20162), .C2(n20186), .ZN(P2_U3228) );
  OAI222_X1 U23126 ( .A1(n20185), .A2(n20166), .B1(n20165), .B2(n20246), .C1(
        n20164), .C2(n20186), .ZN(P2_U3229) );
  INV_X1 U23127 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20167) );
  OAI222_X1 U23128 ( .A1(n20185), .A2(n20167), .B1(n21378), .B2(n20246), .C1(
        n20166), .C2(n20186), .ZN(P2_U3230) );
  INV_X1 U23129 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20169) );
  OAI222_X1 U23130 ( .A1(n20185), .A2(n20169), .B1(n20168), .B2(n20246), .C1(
        n20167), .C2(n20186), .ZN(P2_U3231) );
  OAI222_X1 U23131 ( .A1(n20185), .A2(n20171), .B1(n20170), .B2(n20246), .C1(
        n20169), .C2(n20186), .ZN(P2_U3232) );
  OAI222_X1 U23132 ( .A1(n20185), .A2(n20173), .B1(n20172), .B2(n20246), .C1(
        n20171), .C2(n20186), .ZN(P2_U3233) );
  OAI222_X1 U23133 ( .A1(n20185), .A2(n20175), .B1(n20174), .B2(n20246), .C1(
        n20173), .C2(n20186), .ZN(P2_U3234) );
  OAI222_X1 U23134 ( .A1(n20185), .A2(n20177), .B1(n20176), .B2(n20246), .C1(
        n20175), .C2(n20186), .ZN(P2_U3235) );
  INV_X1 U23135 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20178) );
  OAI222_X1 U23136 ( .A1(n20185), .A2(n20178), .B1(n21436), .B2(n20246), .C1(
        n20177), .C2(n20186), .ZN(P2_U3236) );
  INV_X1 U23137 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20181) );
  OAI222_X1 U23138 ( .A1(n20185), .A2(n20181), .B1(n20179), .B2(n20246), .C1(
        n20178), .C2(n20186), .ZN(P2_U3237) );
  OAI222_X1 U23139 ( .A1(n20186), .A2(n20181), .B1(n20180), .B2(n20246), .C1(
        n20182), .C2(n20185), .ZN(P2_U3238) );
  OAI222_X1 U23140 ( .A1(n20185), .A2(n21456), .B1(n20183), .B2(n20246), .C1(
        n20182), .C2(n20186), .ZN(P2_U3239) );
  INV_X1 U23141 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20187) );
  OAI222_X1 U23142 ( .A1(n20185), .A2(n20187), .B1(n20184), .B2(n20246), .C1(
        n21456), .C2(n20186), .ZN(P2_U3240) );
  INV_X1 U23143 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20189) );
  OAI222_X1 U23144 ( .A1(n20185), .A2(n20189), .B1(n20188), .B2(n20246), .C1(
        n20187), .C2(n20186), .ZN(P2_U3241) );
  OAI22_X1 U23145 ( .A1(n20247), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20246), .ZN(n20190) );
  INV_X1 U23146 ( .A(n20190), .ZN(P2_U3585) );
  MUX2_X1 U23147 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20247), .Z(P2_U3586) );
  OAI22_X1 U23148 ( .A1(n20247), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20246), .ZN(n20191) );
  INV_X1 U23149 ( .A(n20191), .ZN(P2_U3587) );
  OAI22_X1 U23150 ( .A1(n20247), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20246), .ZN(n20192) );
  INV_X1 U23151 ( .A(n20192), .ZN(P2_U3588) );
  OAI21_X1 U23152 ( .B1(n20196), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20194), 
        .ZN(n20193) );
  INV_X1 U23153 ( .A(n20193), .ZN(P2_U3591) );
  OAI21_X1 U23154 ( .B1(n20196), .B2(n20195), .A(n20194), .ZN(P2_U3592) );
  INV_X1 U23155 ( .A(n20232), .ZN(n20231) );
  NOR2_X1 U23156 ( .A1(n20198), .A2(n20197), .ZN(n20216) );
  NAND2_X1 U23157 ( .A1(n20199), .A2(n20216), .ZN(n20210) );
  NAND3_X1 U23158 ( .A1(n20221), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20200), 
        .ZN(n20201) );
  NAND2_X1 U23159 ( .A1(n20201), .A2(n20225), .ZN(n20211) );
  NAND2_X1 U23160 ( .A1(n20210), .A2(n20211), .ZN(n20204) );
  INV_X1 U23161 ( .A(n20202), .ZN(n20203) );
  AOI222_X1 U23162 ( .A1(n20207), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n20206), 
        .B2(n20205), .C1(n20204), .C2(n20203), .ZN(n20208) );
  AOI22_X1 U23163 ( .A1(n20231), .A2(n20209), .B1(n20208), .B2(n20232), .ZN(
        P2_U3602) );
  OAI21_X1 U23164 ( .B1(n20212), .B2(n20211), .A(n20210), .ZN(n20213) );
  AOI21_X1 U23165 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20214), .A(n20213), 
        .ZN(n20215) );
  AOI22_X1 U23166 ( .A1(n20231), .A2(n21487), .B1(n20215), .B2(n20232), .ZN(
        P2_U3603) );
  INV_X1 U23167 ( .A(n20216), .ZN(n20220) );
  INV_X1 U23168 ( .A(n20217), .ZN(n20218) );
  NAND3_X1 U23169 ( .A1(n20221), .A2(n20225), .A3(n20218), .ZN(n20219) );
  OAI21_X1 U23170 ( .B1(n20221), .B2(n20220), .A(n20219), .ZN(n20222) );
  AOI21_X1 U23171 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20223), .A(n20222), 
        .ZN(n20224) );
  AOI22_X1 U23172 ( .A1(n20231), .A2(n21540), .B1(n20224), .B2(n20232), .ZN(
        P2_U3604) );
  INV_X1 U23173 ( .A(n20225), .ZN(n20227) );
  OAI21_X1 U23174 ( .B1(n20228), .B2(n20227), .A(n20226), .ZN(n20229) );
  AOI21_X1 U23175 ( .B1(n20233), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20229), 
        .ZN(n20230) );
  OAI22_X1 U23176 ( .A1(n20233), .A2(n20232), .B1(n20231), .B2(n20230), .ZN(
        P2_U3605) );
  AOI22_X1 U23177 ( .A1(n20246), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20234), 
        .B2(n20247), .ZN(P2_U3608) );
  INV_X1 U23178 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n20245) );
  INV_X1 U23179 ( .A(n20235), .ZN(n20244) );
  INV_X1 U23180 ( .A(n20236), .ZN(n20238) );
  AOI22_X1 U23181 ( .A1(n20240), .A2(n20239), .B1(n20238), .B2(n20237), .ZN(
        n20243) );
  NOR2_X1 U23182 ( .A1(n20244), .A2(n20241), .ZN(n20242) );
  AOI22_X1 U23183 ( .A1(n20245), .A2(n20244), .B1(n20243), .B2(n20242), .ZN(
        P2_U3609) );
  OAI22_X1 U23184 ( .A1(n20247), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20246), .ZN(n20248) );
  INV_X1 U23185 ( .A(n20248), .ZN(P2_U3611) );
  AOI21_X1 U23186 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21137), .A(n21136), 
        .ZN(n20256) );
  INV_X1 U23187 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20249) );
  INV_X1 U23188 ( .A(n21222), .ZN(n21223) );
  AOI21_X1 U23189 ( .B1(n20256), .B2(n20249), .A(n21223), .ZN(P1_U2802) );
  INV_X1 U23190 ( .A(n20250), .ZN(n20252) );
  OAI21_X1 U23191 ( .B1(n20252), .B2(n20251), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20253) );
  OAI21_X1 U23192 ( .B1(n20254), .B2(n20500), .A(n20253), .ZN(P1_U2803) );
  NOR2_X1 U23193 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20257) );
  INV_X1 U23194 ( .A(n21223), .ZN(n21239) );
  OAI21_X1 U23195 ( .B1(n20257), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21239), .ZN(
        n20255) );
  OAI21_X1 U23196 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21222), .A(n20255), 
        .ZN(P1_U2804) );
  NOR2_X1 U23197 ( .A1(n21223), .A2(n20256), .ZN(n21186) );
  OAI21_X1 U23198 ( .B1(BS16), .B2(n20257), .A(n21186), .ZN(n21184) );
  OAI21_X1 U23199 ( .B1(n21186), .B2(n20927), .A(n21184), .ZN(P1_U2805) );
  OAI21_X1 U23200 ( .B1(n20259), .B2(n16029), .A(n20258), .ZN(P1_U2806) );
  NOR4_X1 U23201 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20263) );
  NOR4_X1 U23202 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20262) );
  NOR4_X1 U23203 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20261) );
  NOR4_X1 U23204 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20260) );
  NAND4_X1 U23205 ( .A1(n20263), .A2(n20262), .A3(n20261), .A4(n20260), .ZN(
        n20269) );
  NOR4_X1 U23206 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20267) );
  AOI211_X1 U23207 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20266) );
  NOR4_X1 U23208 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20265) );
  NOR4_X1 U23209 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20264) );
  NAND4_X1 U23210 ( .A1(n20267), .A2(n20266), .A3(n20265), .A4(n20264), .ZN(
        n20268) );
  NOR2_X1 U23211 ( .A1(n20269), .A2(n20268), .ZN(n21221) );
  INV_X1 U23212 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20271) );
  NOR3_X1 U23213 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20272) );
  OAI21_X1 U23214 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20272), .A(n21221), .ZN(
        n20270) );
  OAI21_X1 U23215 ( .B1(n21221), .B2(n20271), .A(n20270), .ZN(P1_U2807) );
  INV_X1 U23216 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21185) );
  AOI21_X1 U23217 ( .B1(n20273), .B2(n21185), .A(n20272), .ZN(n20275) );
  INV_X1 U23218 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20274) );
  INV_X1 U23219 ( .A(n21221), .ZN(n21219) );
  AOI22_X1 U23220 ( .A1(n21221), .A2(n20275), .B1(n20274), .B2(n21219), .ZN(
        P1_U2808) );
  NAND2_X1 U23221 ( .A1(n20276), .A2(n20324), .ZN(n20293) );
  OAI21_X1 U23222 ( .B1(n20342), .B2(n20277), .A(n20447), .ZN(n20281) );
  INV_X1 U23223 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20278) );
  OAI22_X1 U23224 ( .A1(n20279), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n20278), 
        .B2(n20330), .ZN(n20280) );
  AOI211_X1 U23225 ( .C1(n20345), .C2(n20282), .A(n20281), .B(n20280), .ZN(
        n20287) );
  INV_X1 U23226 ( .A(n20283), .ZN(n20285) );
  AOI22_X1 U23227 ( .A1(n20285), .A2(n20307), .B1(n20350), .B2(n20284), .ZN(
        n20286) );
  OAI211_X1 U23228 ( .C1(n20288), .C2(n20293), .A(n20287), .B(n20286), .ZN(
        P1_U2831) );
  OAI21_X1 U23229 ( .B1(n20342), .B2(n20289), .A(n20447), .ZN(n20292) );
  NOR3_X1 U23230 ( .A1(n20318), .A2(P1_REIP_REG_8__SCAN_IN), .A3(n20290), .ZN(
        n20291) );
  AOI211_X1 U23231 ( .C1(n20344), .C2(P1_EBX_REG_8__SCAN_IN), .A(n20292), .B(
        n20291), .ZN(n20299) );
  OAI22_X1 U23232 ( .A1(n20295), .A2(n20294), .B1(n14444), .B2(n20293), .ZN(
        n20296) );
  AOI21_X1 U23233 ( .B1(n20297), .B2(n20350), .A(n20296), .ZN(n20298) );
  OAI211_X1 U23234 ( .C1(n20301), .C2(n20300), .A(n20299), .B(n20298), .ZN(
        P1_U2832) );
  INV_X1 U23235 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20315) );
  NOR3_X1 U23236 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20302), .A3(n20318), .ZN(
        n20303) );
  AOI211_X1 U23237 ( .C1(n20351), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20487), .B(n20303), .ZN(n20312) );
  INV_X1 U23238 ( .A(n20304), .ZN(n20305) );
  AOI22_X1 U23239 ( .A1(n20344), .A2(P1_EBX_REG_6__SCAN_IN), .B1(n20305), .B2(
        n20350), .ZN(n20311) );
  NAND2_X1 U23240 ( .A1(n20306), .A2(n20345), .ZN(n20310) );
  NAND2_X1 U23241 ( .A1(n20308), .A2(n20307), .ZN(n20309) );
  AND4_X1 U23242 ( .A1(n20312), .A2(n20311), .A3(n20310), .A4(n20309), .ZN(
        n20313) );
  OAI21_X1 U23243 ( .B1(n20315), .B2(n20314), .A(n20313), .ZN(P1_U2834) );
  OAI21_X1 U23244 ( .B1(n20342), .B2(n20316), .A(n20447), .ZN(n20320) );
  INV_X1 U23245 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20317) );
  OAI22_X1 U23246 ( .A1(n20318), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20317), 
        .B2(n20330), .ZN(n20319) );
  AOI211_X1 U23247 ( .C1(n20345), .C2(n20321), .A(n20320), .B(n20319), .ZN(
        n20327) );
  INV_X1 U23248 ( .A(n20322), .ZN(n20325) );
  AND2_X1 U23249 ( .A1(n20324), .A2(n20323), .ZN(n20339) );
  AOI22_X1 U23250 ( .A1(n20325), .A2(n20357), .B1(n20339), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20326) );
  OAI211_X1 U23251 ( .C1(n20328), .C2(n20333), .A(n20327), .B(n20326), .ZN(
        P1_U2835) );
  INV_X1 U23252 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20343) );
  NOR3_X1 U23253 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20346), .A3(n20354), .ZN(
        n20329) );
  AOI211_X1 U23254 ( .C1(n20345), .C2(n20444), .A(n20487), .B(n20329), .ZN(
        n20341) );
  OAI22_X1 U23255 ( .A1(n20332), .A2(n20331), .B1(n11463), .B2(n20330), .ZN(
        n20338) );
  OAI22_X1 U23256 ( .A1(n20336), .A2(n20335), .B1(n20334), .B2(n20333), .ZN(
        n20337) );
  AOI211_X1 U23257 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n20339), .A(n20338), .B(
        n20337), .ZN(n20340) );
  OAI211_X1 U23258 ( .C1(n20343), .C2(n20342), .A(n20341), .B(n20340), .ZN(
        P1_U2836) );
  INV_X1 U23259 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21142) );
  AOI22_X1 U23260 ( .A1(n20345), .A2(n20453), .B1(n20344), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n20360) );
  OAI21_X1 U23261 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20346), .ZN(n20355) );
  NAND2_X1 U23262 ( .A1(n14039), .A2(n20347), .ZN(n20353) );
  INV_X1 U23263 ( .A(n20348), .ZN(n20349) );
  AOI22_X1 U23264 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20351), .B1(
        n20350), .B2(n20349), .ZN(n20352) );
  OAI211_X1 U23265 ( .C1(n20355), .C2(n20354), .A(n20353), .B(n20352), .ZN(
        n20356) );
  AOI21_X1 U23266 ( .B1(n20358), .B2(n20357), .A(n20356), .ZN(n20359) );
  OAI211_X1 U23267 ( .C1(n20361), .C2(n21142), .A(n20360), .B(n20359), .ZN(
        P1_U2837) );
  INV_X1 U23268 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n21426) );
  OAI22_X1 U23269 ( .A1(n20379), .A2(n16802), .B1(n20362), .B2(n20365), .ZN(
        n20363) );
  INV_X1 U23270 ( .A(n20363), .ZN(n20364) );
  OAI21_X1 U23271 ( .B1(n21426), .B2(n20380), .A(n20364), .ZN(P1_U2906) );
  INV_X1 U23272 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n21318) );
  INV_X1 U23273 ( .A(n20365), .ZN(n20366) );
  AOI22_X1 U23274 ( .A1(n20366), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20387), .ZN(n20367) );
  OAI21_X1 U23275 ( .B1(n20379), .B2(n21318), .A(n20367), .ZN(P1_U2907) );
  AOI22_X1 U23276 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20368) );
  OAI21_X1 U23277 ( .B1(n13979), .B2(n20389), .A(n20368), .ZN(P1_U2921) );
  AOI22_X1 U23278 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20369) );
  OAI21_X1 U23279 ( .B1(n14506), .B2(n20389), .A(n20369), .ZN(P1_U2922) );
  AOI22_X1 U23280 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20370) );
  OAI21_X1 U23281 ( .B1(n14532), .B2(n20389), .A(n20370), .ZN(P1_U2923) );
  AOI22_X1 U23282 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20371) );
  OAI21_X1 U23283 ( .B1(n14495), .B2(n20389), .A(n20371), .ZN(P1_U2924) );
  INV_X1 U23284 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20373) );
  AOI22_X1 U23285 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20372) );
  OAI21_X1 U23286 ( .B1(n20373), .B2(n20389), .A(n20372), .ZN(P1_U2925) );
  AOI22_X1 U23287 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20374) );
  OAI21_X1 U23288 ( .B1(n14476), .B2(n20389), .A(n20374), .ZN(P1_U2926) );
  AOI22_X1 U23289 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20375) );
  OAI21_X1 U23290 ( .B1(n14450), .B2(n20389), .A(n20375), .ZN(P1_U2927) );
  AOI22_X1 U23291 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20376) );
  OAI21_X1 U23292 ( .B1(n14363), .B2(n20389), .A(n20376), .ZN(P1_U2928) );
  AOI22_X1 U23293 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20377) );
  OAI21_X1 U23294 ( .B1(n10783), .B2(n20389), .A(n20377), .ZN(P1_U2929) );
  AOI22_X1 U23295 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20378) );
  OAI21_X1 U23296 ( .B1(n10773), .B2(n20389), .A(n20378), .ZN(P1_U2930) );
  INV_X1 U23297 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n21444) );
  OAI222_X1 U23298 ( .A1(n20380), .A2(n21444), .B1(n20389), .B2(n14187), .C1(
        n20379), .C2(n21439), .ZN(P1_U2931) );
  AOI22_X1 U23299 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20381) );
  OAI21_X1 U23300 ( .B1(n20382), .B2(n20389), .A(n20381), .ZN(P1_U2932) );
  AOI22_X1 U23301 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20383) );
  OAI21_X1 U23302 ( .B1(n10709), .B2(n20389), .A(n20383), .ZN(P1_U2933) );
  AOI22_X1 U23303 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20384) );
  OAI21_X1 U23304 ( .B1(n10658), .B2(n20389), .A(n20384), .ZN(P1_U2934) );
  AOI22_X1 U23305 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20385) );
  OAI21_X1 U23306 ( .B1(n10664), .B2(n20389), .A(n20385), .ZN(P1_U2935) );
  AOI22_X1 U23307 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20387), .B1(n20386), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20388) );
  OAI21_X1 U23308 ( .B1(n10672), .B2(n20389), .A(n20388), .ZN(P1_U2936) );
  AOI22_X1 U23309 ( .A1(n20426), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20397), .ZN(n20392) );
  INV_X1 U23310 ( .A(n20390), .ZN(n20391) );
  NAND2_X1 U23311 ( .A1(n20411), .A2(n20391), .ZN(n20413) );
  NAND2_X1 U23312 ( .A1(n20392), .A2(n20413), .ZN(P1_U2945) );
  AOI22_X1 U23313 ( .A1(n20393), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20397), .ZN(n20396) );
  INV_X1 U23314 ( .A(n20394), .ZN(n20395) );
  NAND2_X1 U23315 ( .A1(n20411), .A2(n20395), .ZN(n20415) );
  NAND2_X1 U23316 ( .A1(n20396), .A2(n20415), .ZN(P1_U2946) );
  AOI22_X1 U23317 ( .A1(n20426), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20397), .ZN(n20400) );
  INV_X1 U23318 ( .A(n20398), .ZN(n20399) );
  NAND2_X1 U23319 ( .A1(n20411), .A2(n20399), .ZN(n20417) );
  NAND2_X1 U23320 ( .A1(n20400), .A2(n20417), .ZN(P1_U2947) );
  AOI22_X1 U23321 ( .A1(n20426), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20425), .ZN(n20402) );
  NAND2_X1 U23322 ( .A1(n20411), .A2(n20401), .ZN(n20419) );
  NAND2_X1 U23323 ( .A1(n20402), .A2(n20419), .ZN(P1_U2948) );
  AOI22_X1 U23324 ( .A1(n20426), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20425), .ZN(n20405) );
  INV_X1 U23325 ( .A(n20403), .ZN(n20404) );
  NAND2_X1 U23326 ( .A1(n20411), .A2(n20404), .ZN(n20421) );
  NAND2_X1 U23327 ( .A1(n20405), .A2(n20421), .ZN(P1_U2949) );
  AOI22_X1 U23328 ( .A1(n20426), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20425), .ZN(n20408) );
  INV_X1 U23329 ( .A(n20406), .ZN(n20407) );
  NAND2_X1 U23330 ( .A1(n20411), .A2(n20407), .ZN(n20423) );
  NAND2_X1 U23331 ( .A1(n20408), .A2(n20423), .ZN(P1_U2950) );
  AOI22_X1 U23332 ( .A1(n20426), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20397), .ZN(n20412) );
  INV_X1 U23333 ( .A(n20409), .ZN(n20410) );
  NAND2_X1 U23334 ( .A1(n20411), .A2(n20410), .ZN(n20427) );
  NAND2_X1 U23335 ( .A1(n20412), .A2(n20427), .ZN(P1_U2951) );
  AOI22_X1 U23336 ( .A1(n20426), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20425), .ZN(n20414) );
  NAND2_X1 U23337 ( .A1(n20414), .A2(n20413), .ZN(P1_U2960) );
  AOI22_X1 U23338 ( .A1(n20426), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20397), .ZN(n20416) );
  NAND2_X1 U23339 ( .A1(n20416), .A2(n20415), .ZN(P1_U2961) );
  AOI22_X1 U23340 ( .A1(n20426), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20425), .ZN(n20418) );
  NAND2_X1 U23341 ( .A1(n20418), .A2(n20417), .ZN(P1_U2962) );
  AOI22_X1 U23342 ( .A1(n20426), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20397), .ZN(n20420) );
  NAND2_X1 U23343 ( .A1(n20420), .A2(n20419), .ZN(P1_U2963) );
  AOI22_X1 U23344 ( .A1(n20426), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20425), .ZN(n20422) );
  NAND2_X1 U23345 ( .A1(n20422), .A2(n20421), .ZN(P1_U2964) );
  AOI22_X1 U23346 ( .A1(n20426), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20425), .ZN(n20424) );
  NAND2_X1 U23347 ( .A1(n20424), .A2(n20423), .ZN(P1_U2965) );
  AOI22_X1 U23348 ( .A1(n20426), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20425), .ZN(n20428) );
  NAND2_X1 U23349 ( .A1(n20428), .A2(n20427), .ZN(P1_U2966) );
  INV_X1 U23350 ( .A(n20429), .ZN(n20431) );
  AOI21_X1 U23351 ( .B1(n20431), .B2(n20473), .A(n20430), .ZN(n20488) );
  NAND2_X1 U23352 ( .A1(n20433), .A2(n20432), .ZN(n20434) );
  AOI22_X1 U23353 ( .A1(n20435), .A2(n20488), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20434), .ZN(n20437) );
  NAND2_X1 U23354 ( .A1(n20487), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20436) );
  OAI211_X1 U23355 ( .C1(n20438), .C2(n20496), .A(n20437), .B(n20436), .ZN(
        P1_U2999) );
  OAI21_X1 U23356 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20439), .ZN(n20446) );
  OAI22_X1 U23357 ( .A1(n20456), .A2(n20441), .B1(n20440), .B2(n20449), .ZN(
        n20442) );
  AOI211_X1 U23358 ( .C1(n20486), .C2(n20444), .A(n20443), .B(n20442), .ZN(
        n20445) );
  OAI21_X1 U23359 ( .B1(n20448), .B2(n20446), .A(n20445), .ZN(P1_U3027) );
  NOR2_X1 U23360 ( .A1(n20447), .A2(n21142), .ZN(n20452) );
  OAI22_X1 U23361 ( .A1(n20450), .A2(n20449), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20448), .ZN(n20451) );
  AOI211_X1 U23362 ( .C1(n20486), .C2(n20453), .A(n20452), .B(n20451), .ZN(
        n20454) );
  OAI21_X1 U23363 ( .B1(n20456), .B2(n20455), .A(n20454), .ZN(P1_U3028) );
  AOI21_X1 U23364 ( .B1(n14133), .B2(n20458), .A(n20457), .ZN(n20469) );
  INV_X1 U23365 ( .A(n20459), .ZN(n20467) );
  NAND2_X1 U23366 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20461) );
  OAI21_X1 U23367 ( .B1(n20470), .B2(n20461), .A(n20460), .ZN(n20462) );
  AOI22_X1 U23368 ( .A1(n20463), .A2(n20462), .B1(n20487), .B2(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20464) );
  OAI21_X1 U23369 ( .B1(n20479), .B2(n20465), .A(n20464), .ZN(n20466) );
  AOI21_X1 U23370 ( .B1(n20467), .B2(n20489), .A(n20466), .ZN(n20468) );
  OAI221_X1 U23371 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20471), .C1(
        n20470), .C2(n20469), .A(n20468), .ZN(P1_U3029) );
  NAND2_X1 U23372 ( .A1(n20473), .A2(n20472), .ZN(n20491) );
  INV_X1 U23373 ( .A(n20474), .ZN(n20476) );
  NOR3_X1 U23374 ( .A1(n20476), .A2(n20475), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20481) );
  OAI21_X1 U23375 ( .B1(n20479), .B2(n20478), .A(n20477), .ZN(n20480) );
  AOI211_X1 U23376 ( .C1(n20482), .C2(n20489), .A(n20481), .B(n20480), .ZN(
        n20483) );
  OAI221_X1 U23377 ( .B1(n14133), .B2(n20484), .C1(n14133), .C2(n20491), .A(
        n20483), .ZN(P1_U3030) );
  AOI22_X1 U23378 ( .A1(n20487), .A2(P1_REIP_REG_0__SCAN_IN), .B1(n20486), 
        .B2(n20485), .ZN(n20493) );
  AOI22_X1 U23379 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20490), .B1(
        n20489), .B2(n20488), .ZN(n20492) );
  NAND3_X1 U23380 ( .A1(n20493), .A2(n20492), .A3(n20491), .ZN(P1_U3031) );
  NOR2_X1 U23381 ( .A1(n20494), .A2(n21212), .ZN(P1_U3032) );
  NAND2_X1 U23382 ( .A1(n20551), .A2(n20501), .ZN(n20925) );
  NAND3_X1 U23383 ( .A1(n21205), .A2(n20922), .A3(n20850), .ZN(n20564) );
  NOR2_X1 U23384 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20564), .ZN(
        n20509) );
  INV_X1 U23385 ( .A(n20509), .ZN(n20554) );
  AOI22_X1 U23386 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20552), .B1(DATAI_24_), 
        .B2(n20498), .ZN(n21077) );
  OR2_X1 U23387 ( .A1(n21073), .A2(n21077), .ZN(n20503) );
  OAI21_X1 U23388 ( .B1(n20925), .B2(n20554), .A(n20503), .ZN(n20504) );
  INV_X1 U23389 ( .A(n20504), .ZN(n20516) );
  NAND2_X1 U23390 ( .A1(n20512), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21012) );
  NAND3_X1 U23391 ( .A1(n20587), .A2(n21206), .A3(n21073), .ZN(n20506) );
  NAND2_X1 U23392 ( .A1(n20506), .A2(n21199), .ZN(n20511) );
  OR2_X1 U23393 ( .A1(n14039), .A2(n20507), .ZN(n20627) );
  OR2_X1 U23394 ( .A1(n20627), .A2(n21016), .ZN(n20513) );
  NAND2_X1 U23395 ( .A1(n20853), .A2(n20798), .ZN(n20667) );
  AOI22_X1 U23396 ( .A1(n20511), .A2(n20513), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20667), .ZN(n20508) );
  OAI211_X1 U23397 ( .C1(n20509), .C2(n20931), .A(n20856), .B(n20508), .ZN(
        n20558) );
  NOR2_X2 U23398 ( .A1(n20510), .A2(n20670), .ZN(n21064) );
  INV_X1 U23399 ( .A(n20511), .ZN(n20514) );
  NOR2_X1 U23400 ( .A1(n20512), .A2(n20980), .ZN(n20671) );
  INV_X1 U23401 ( .A(n20671), .ZN(n20859) );
  OAI22_X1 U23402 ( .A1(n20514), .A2(n20513), .B1(n20667), .B2(n20859), .ZN(
        n20557) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20558), .B1(
        n21064), .B2(n20557), .ZN(n20515) );
  OAI211_X1 U23404 ( .C1(n21026), .C2(n20587), .A(n20516), .B(n20515), .ZN(
        P1_U3033) );
  AOI22_X1 U23405 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20552), .B1(DATAI_17_), 
        .B2(n20498), .ZN(n21030) );
  NAND2_X1 U23406 ( .A1(n20551), .A2(n20517), .ZN(n20940) );
  AOI22_X1 U23407 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20552), .B1(DATAI_25_), 
        .B2(n20498), .ZN(n21082) );
  OR2_X1 U23408 ( .A1(n21073), .A2(n21082), .ZN(n20518) );
  OAI21_X1 U23409 ( .B1(n20940), .B2(n20554), .A(n20518), .ZN(n20519) );
  INV_X1 U23410 ( .A(n20519), .ZN(n20522) );
  NOR2_X2 U23411 ( .A1(n20520), .A2(n20670), .ZN(n21078) );
  AOI22_X1 U23412 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20558), .B1(
        n21078), .B2(n20557), .ZN(n20521) );
  OAI211_X1 U23413 ( .C1(n10000), .C2(n20587), .A(n20522), .B(n20521), .ZN(
        P1_U3034) );
  AOI22_X1 U23414 ( .A1(DATAI_18_), .A2(n20498), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20552), .ZN(n21034) );
  NAND2_X1 U23415 ( .A1(n20551), .A2(n20523), .ZN(n20945) );
  AOI22_X1 U23416 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20552), .B1(DATAI_26_), 
        .B2(n20498), .ZN(n21087) );
  OR2_X1 U23417 ( .A1(n21073), .A2(n21087), .ZN(n20524) );
  OAI21_X1 U23418 ( .B1(n20945), .B2(n20554), .A(n20524), .ZN(n20525) );
  INV_X1 U23419 ( .A(n20525), .ZN(n20528) );
  NOR2_X2 U23420 ( .A1(n20526), .A2(n20670), .ZN(n21083) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20558), .B1(
        n21083), .B2(n20557), .ZN(n20527) );
  OAI211_X1 U23422 ( .C1(n10002), .C2(n20587), .A(n20528), .B(n20527), .ZN(
        P1_U3035) );
  AOI22_X1 U23423 ( .A1(DATAI_19_), .A2(n20498), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20552), .ZN(n21038) );
  NAND2_X1 U23424 ( .A1(n20551), .A2(n10546), .ZN(n20950) );
  AOI22_X1 U23425 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20552), .B1(DATAI_27_), 
        .B2(n20498), .ZN(n21092) );
  OR2_X1 U23426 ( .A1(n21073), .A2(n21092), .ZN(n20529) );
  OAI21_X1 U23427 ( .B1(n20950), .B2(n20554), .A(n20529), .ZN(n20530) );
  INV_X1 U23428 ( .A(n20530), .ZN(n20533) );
  NOR2_X2 U23429 ( .A1(n20531), .A2(n20670), .ZN(n21088) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20558), .B1(
        n21088), .B2(n20557), .ZN(n20532) );
  OAI211_X1 U23431 ( .C1(n10004), .C2(n20587), .A(n20533), .B(n20532), .ZN(
        P1_U3036) );
  NAND2_X1 U23432 ( .A1(n20551), .A2(n20534), .ZN(n20955) );
  AOI22_X1 U23433 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20552), .B1(DATAI_28_), 
        .B2(n20498), .ZN(n21097) );
  OR2_X1 U23434 ( .A1(n21073), .A2(n9994), .ZN(n20535) );
  OAI21_X1 U23435 ( .B1(n20955), .B2(n20554), .A(n20535), .ZN(n20536) );
  INV_X1 U23436 ( .A(n20536), .ZN(n20539) );
  NOR2_X2 U23437 ( .A1(n20537), .A2(n20670), .ZN(n21093) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20558), .B1(
        n21093), .B2(n20557), .ZN(n20538) );
  OAI211_X1 U23439 ( .C1(n21041), .C2(n20587), .A(n20539), .B(n20538), .ZN(
        P1_U3037) );
  AOI22_X1 U23440 ( .A1(DATAI_21_), .A2(n20498), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20552), .ZN(n21045) );
  NAND2_X1 U23441 ( .A1(n20551), .A2(n11248), .ZN(n20960) );
  AOI22_X1 U23442 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20552), .B1(DATAI_29_), 
        .B2(n20498), .ZN(n21102) );
  OR2_X1 U23443 ( .A1(n21073), .A2(n21102), .ZN(n20540) );
  OAI21_X1 U23444 ( .B1(n20960), .B2(n20554), .A(n20540), .ZN(n20541) );
  INV_X1 U23445 ( .A(n20541), .ZN(n20544) );
  NOR2_X2 U23446 ( .A1(n20542), .A2(n20670), .ZN(n21098) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20558), .B1(
        n21098), .B2(n20557), .ZN(n20543) );
  OAI211_X1 U23448 ( .C1(n10006), .C2(n20587), .A(n20544), .B(n20543), .ZN(
        P1_U3038) );
  AOI22_X1 U23449 ( .A1(DATAI_22_), .A2(n20498), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20552), .ZN(n21049) );
  NAND2_X1 U23450 ( .A1(n20551), .A2(n10553), .ZN(n20965) );
  AOI22_X1 U23451 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20552), .B1(DATAI_30_), 
        .B2(n20498), .ZN(n21107) );
  OR2_X1 U23452 ( .A1(n21073), .A2(n21107), .ZN(n20545) );
  OAI21_X1 U23453 ( .B1(n20965), .B2(n20554), .A(n20545), .ZN(n20546) );
  INV_X1 U23454 ( .A(n20546), .ZN(n20549) );
  NOR2_X2 U23455 ( .A1(n20547), .A2(n20670), .ZN(n21103) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20558), .B1(
        n21103), .B2(n20557), .ZN(n20548) );
  OAI211_X1 U23457 ( .C1(n9998), .C2(n20587), .A(n20549), .B(n20548), .ZN(
        P1_U3039) );
  NAND2_X1 U23458 ( .A1(n20551), .A2(n20550), .ZN(n20971) );
  AOI22_X1 U23459 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20552), .B1(DATAI_31_), 
        .B2(n20498), .ZN(n21118) );
  OR2_X1 U23460 ( .A1(n21073), .A2(n9996), .ZN(n20553) );
  OAI21_X1 U23461 ( .B1(n20971), .B2(n20554), .A(n20553), .ZN(n20555) );
  INV_X1 U23462 ( .A(n20555), .ZN(n20560) );
  NOR2_X2 U23463 ( .A1(n20670), .A2(n20556), .ZN(n21109) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20558), .B1(
        n21109), .B2(n20557), .ZN(n20559) );
  OAI211_X1 U23465 ( .C1(n21056), .C2(n20587), .A(n20560), .B(n20559), .ZN(
        P1_U3040) );
  NOR2_X1 U23466 ( .A1(n21214), .A2(n20564), .ZN(n20582) );
  OR2_X1 U23467 ( .A1(n20561), .A2(n21194), .ZN(n20978) );
  INV_X1 U23468 ( .A(n20582), .ZN(n20562) );
  OAI222_X1 U23469 ( .A1(n20978), .A2(n20627), .B1(n20980), .B2(n20564), .C1(
        n21194), .C2(n20562), .ZN(n20581) );
  AOI22_X1 U23470 ( .A1(n21065), .A2(n20582), .B1(n21064), .B2(n20581), .ZN(
        n20567) );
  INV_X1 U23471 ( .A(n20563), .ZN(n20985) );
  OAI21_X1 U23472 ( .B1(n20631), .B2(n20985), .A(n20564), .ZN(n20565) );
  NAND2_X1 U23473 ( .A1(n20565), .A2(n21070), .ZN(n20584) );
  INV_X1 U23474 ( .A(n21077), .ZN(n21023) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20584), .B1(
        n20578), .B2(n21023), .ZN(n20566) );
  OAI211_X1 U23476 ( .C1(n21026), .C2(n20625), .A(n20567), .B(n20566), .ZN(
        P1_U3041) );
  AOI22_X1 U23477 ( .A1(n21079), .A2(n20582), .B1(n21078), .B2(n20581), .ZN(
        n20569) );
  INV_X1 U23478 ( .A(n21082), .ZN(n21027) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20584), .B1(
        n20578), .B2(n21027), .ZN(n20568) );
  OAI211_X1 U23480 ( .C1(n10000), .C2(n20625), .A(n20569), .B(n20568), .ZN(
        P1_U3042) );
  AOI22_X1 U23481 ( .A1(n21084), .A2(n20582), .B1(n21083), .B2(n20581), .ZN(
        n20571) );
  INV_X1 U23482 ( .A(n21087), .ZN(n21031) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20584), .B1(
        n20578), .B2(n21031), .ZN(n20570) );
  OAI211_X1 U23484 ( .C1(n10002), .C2(n20625), .A(n20571), .B(n20570), .ZN(
        P1_U3043) );
  AOI22_X1 U23485 ( .A1(n21089), .A2(n20582), .B1(n21088), .B2(n20581), .ZN(
        n20573) );
  INV_X1 U23486 ( .A(n21092), .ZN(n21035) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20584), .B1(
        n20578), .B2(n21035), .ZN(n20572) );
  OAI211_X1 U23488 ( .C1(n10004), .C2(n20625), .A(n20573), .B(n20572), .ZN(
        P1_U3044) );
  AOI22_X1 U23489 ( .A1(n21094), .A2(n20582), .B1(n21093), .B2(n20581), .ZN(
        n20575) );
  INV_X1 U23490 ( .A(n20625), .ZN(n20583) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n9990), .ZN(n20574) );
  OAI211_X1 U23492 ( .C1(n9994), .C2(n20587), .A(n20575), .B(n20574), .ZN(
        P1_U3045) );
  AOI22_X1 U23493 ( .A1(n21099), .A2(n20582), .B1(n21098), .B2(n20581), .ZN(
        n20577) );
  INV_X1 U23494 ( .A(n21102), .ZN(n21042) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20584), .B1(
        n20578), .B2(n21042), .ZN(n20576) );
  OAI211_X1 U23496 ( .C1(n10006), .C2(n20625), .A(n20577), .B(n20576), .ZN(
        P1_U3046) );
  AOI22_X1 U23497 ( .A1(n21104), .A2(n20582), .B1(n21103), .B2(n20581), .ZN(
        n20580) );
  INV_X1 U23498 ( .A(n21107), .ZN(n21046) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20584), .B1(
        n20578), .B2(n21046), .ZN(n20579) );
  OAI211_X1 U23500 ( .C1(n9998), .C2(n20625), .A(n20580), .B(n20579), .ZN(
        P1_U3047) );
  AOI22_X1 U23501 ( .A1(n21111), .A2(n20582), .B1(n21109), .B2(n20581), .ZN(
        n20586) );
  INV_X1 U23502 ( .A(n21056), .ZN(n21112) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n21112), .ZN(n20585) );
  OAI211_X1 U23504 ( .C1(n9996), .C2(n20587), .A(n20586), .B(n20585), .ZN(
        P1_U3048) );
  NAND3_X1 U23505 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21205), .A3(
        n20922), .ZN(n20635) );
  NOR2_X1 U23506 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20635), .ZN(
        n20592) );
  INV_X1 U23507 ( .A(n20592), .ZN(n20619) );
  OAI22_X1 U23508 ( .A1(n20625), .A2(n21077), .B1(n20925), .B2(n20619), .ZN(
        n20589) );
  INV_X1 U23509 ( .A(n20589), .ZN(n20600) );
  NAND2_X1 U23510 ( .A1(n20987), .A2(n21008), .ZN(n20590) );
  NAND2_X1 U23511 ( .A1(n20590), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21014) );
  OR2_X1 U23512 ( .A1(n20631), .A2(n21014), .ZN(n20591) );
  AND2_X1 U23513 ( .A1(n20591), .A2(n21206), .ZN(n20595) );
  OR2_X1 U23514 ( .A1(n20627), .A2(n14077), .ZN(n20597) );
  NOR2_X1 U23515 ( .A1(n20592), .A2(n20931), .ZN(n20593) );
  AOI21_X1 U23516 ( .B1(n20595), .B2(n20597), .A(n20593), .ZN(n20594) );
  OAI21_X1 U23517 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20853), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20723) );
  NAND3_X1 U23518 ( .A1(n20856), .A2(n20594), .A3(n20723), .ZN(n20622) );
  INV_X1 U23519 ( .A(n20595), .ZN(n20598) );
  INV_X1 U23520 ( .A(n20853), .ZN(n20596) );
  NAND2_X1 U23521 ( .A1(n20596), .A2(n21205), .ZN(n20726) );
  OAI22_X1 U23522 ( .A1(n20598), .A2(n20597), .B1(n20859), .B2(n20726), .ZN(
        n20621) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20622), .B1(
        n21064), .B2(n20621), .ZN(n20599) );
  OAI211_X1 U23524 ( .C1(n21026), .C2(n20664), .A(n20600), .B(n20599), .ZN(
        P1_U3049) );
  OAI22_X1 U23525 ( .A1(n20664), .A2(n10000), .B1(n20940), .B2(n20619), .ZN(
        n20601) );
  INV_X1 U23526 ( .A(n20601), .ZN(n20603) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20622), .B1(
        n21078), .B2(n20621), .ZN(n20602) );
  OAI211_X1 U23528 ( .C1(n21082), .C2(n20625), .A(n20603), .B(n20602), .ZN(
        P1_U3050) );
  OAI22_X1 U23529 ( .A1(n20664), .A2(n10002), .B1(n20945), .B2(n20619), .ZN(
        n20604) );
  INV_X1 U23530 ( .A(n20604), .ZN(n20606) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20622), .B1(
        n21083), .B2(n20621), .ZN(n20605) );
  OAI211_X1 U23532 ( .C1(n21087), .C2(n20625), .A(n20606), .B(n20605), .ZN(
        P1_U3051) );
  OAI22_X1 U23533 ( .A1(n20625), .A2(n21092), .B1(n20950), .B2(n20619), .ZN(
        n20607) );
  INV_X1 U23534 ( .A(n20607), .ZN(n20609) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20622), .B1(
        n21088), .B2(n20621), .ZN(n20608) );
  OAI211_X1 U23536 ( .C1(n10004), .C2(n20664), .A(n20609), .B(n20608), .ZN(
        P1_U3052) );
  OAI22_X1 U23537 ( .A1(n20625), .A2(n9994), .B1(n20955), .B2(n20619), .ZN(
        n20610) );
  INV_X1 U23538 ( .A(n20610), .ZN(n20612) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20622), .B1(
        n21093), .B2(n20621), .ZN(n20611) );
  OAI211_X1 U23540 ( .C1(n21041), .C2(n20664), .A(n20612), .B(n20611), .ZN(
        P1_U3053) );
  OAI22_X1 U23541 ( .A1(n20625), .A2(n21102), .B1(n20960), .B2(n20619), .ZN(
        n20613) );
  INV_X1 U23542 ( .A(n20613), .ZN(n20615) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20622), .B1(
        n21098), .B2(n20621), .ZN(n20614) );
  OAI211_X1 U23544 ( .C1(n10006), .C2(n20664), .A(n20615), .B(n20614), .ZN(
        P1_U3054) );
  OAI22_X1 U23545 ( .A1(n20664), .A2(n9998), .B1(n20965), .B2(n20619), .ZN(
        n20616) );
  INV_X1 U23546 ( .A(n20616), .ZN(n20618) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20622), .B1(
        n21103), .B2(n20621), .ZN(n20617) );
  OAI211_X1 U23548 ( .C1(n21107), .C2(n20625), .A(n20618), .B(n20617), .ZN(
        P1_U3055) );
  OAI22_X1 U23549 ( .A1(n20664), .A2(n21056), .B1(n20971), .B2(n20619), .ZN(
        n20620) );
  INV_X1 U23550 ( .A(n20620), .ZN(n20624) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20622), .B1(
        n21109), .B2(n20621), .ZN(n20623) );
  OAI211_X1 U23552 ( .C1(n9996), .C2(n20625), .A(n20624), .B(n20623), .ZN(
        P1_U3056) );
  OR2_X1 U23553 ( .A1(n20891), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20658) );
  OAI22_X1 U23554 ( .A1(n20693), .A2(n21026), .B1(n20925), .B2(n20658), .ZN(
        n20626) );
  INV_X1 U23555 ( .A(n20626), .ZN(n20639) );
  INV_X1 U23556 ( .A(n20627), .ZN(n20630) );
  AND2_X1 U23557 ( .A1(n20628), .A2(n21209), .ZN(n21057) );
  INV_X1 U23558 ( .A(n20658), .ZN(n20629) );
  AOI21_X1 U23559 ( .B1(n20630), .B2(n21057), .A(n20629), .ZN(n20637) );
  OR2_X1 U23560 ( .A1(n20631), .A2(n21068), .ZN(n20632) );
  AOI22_X1 U23561 ( .A1(n20637), .A2(n20634), .B1(n21194), .B2(n20635), .ZN(
        n20633) );
  NAND2_X1 U23562 ( .A1(n21070), .A2(n20633), .ZN(n20661) );
  INV_X1 U23563 ( .A(n20634), .ZN(n20636) );
  OAI22_X1 U23564 ( .A1(n20637), .A2(n20636), .B1(n20980), .B2(n20635), .ZN(
        n20660) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20661), .B1(
        n21064), .B2(n20660), .ZN(n20638) );
  OAI211_X1 U23566 ( .C1(n21077), .C2(n20664), .A(n20639), .B(n20638), .ZN(
        P1_U3057) );
  OAI22_X1 U23567 ( .A1(n20693), .A2(n10000), .B1(n20940), .B2(n20658), .ZN(
        n20640) );
  INV_X1 U23568 ( .A(n20640), .ZN(n20642) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20661), .B1(
        n21078), .B2(n20660), .ZN(n20641) );
  OAI211_X1 U23570 ( .C1(n21082), .C2(n20664), .A(n20642), .B(n20641), .ZN(
        P1_U3058) );
  OAI22_X1 U23571 ( .A1(n20693), .A2(n10002), .B1(n20945), .B2(n20658), .ZN(
        n20643) );
  INV_X1 U23572 ( .A(n20643), .ZN(n20645) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20661), .B1(
        n21083), .B2(n20660), .ZN(n20644) );
  OAI211_X1 U23574 ( .C1(n21087), .C2(n20664), .A(n20645), .B(n20644), .ZN(
        P1_U3059) );
  OAI22_X1 U23575 ( .A1(n20693), .A2(n10004), .B1(n20950), .B2(n20658), .ZN(
        n20646) );
  INV_X1 U23576 ( .A(n20646), .ZN(n20648) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20661), .B1(
        n21088), .B2(n20660), .ZN(n20647) );
  OAI211_X1 U23578 ( .C1(n21092), .C2(n20664), .A(n20648), .B(n20647), .ZN(
        P1_U3060) );
  OAI22_X1 U23579 ( .A1(n20693), .A2(n21041), .B1(n20955), .B2(n20658), .ZN(
        n20649) );
  INV_X1 U23580 ( .A(n20649), .ZN(n20651) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20661), .B1(
        n21093), .B2(n20660), .ZN(n20650) );
  OAI211_X1 U23582 ( .C1(n9994), .C2(n20664), .A(n20651), .B(n20650), .ZN(
        P1_U3061) );
  OAI22_X1 U23583 ( .A1(n20693), .A2(n10006), .B1(n20960), .B2(n20658), .ZN(
        n20652) );
  INV_X1 U23584 ( .A(n20652), .ZN(n20654) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20661), .B1(
        n21098), .B2(n20660), .ZN(n20653) );
  OAI211_X1 U23586 ( .C1(n21102), .C2(n20664), .A(n20654), .B(n20653), .ZN(
        P1_U3062) );
  OAI22_X1 U23587 ( .A1(n20693), .A2(n9998), .B1(n20965), .B2(n20658), .ZN(
        n20655) );
  INV_X1 U23588 ( .A(n20655), .ZN(n20657) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20661), .B1(
        n21103), .B2(n20660), .ZN(n20656) );
  OAI211_X1 U23590 ( .C1(n21107), .C2(n20664), .A(n20657), .B(n20656), .ZN(
        P1_U3063) );
  OAI22_X1 U23591 ( .A1(n20693), .A2(n21056), .B1(n20971), .B2(n20658), .ZN(
        n20659) );
  INV_X1 U23592 ( .A(n20659), .ZN(n20663) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20661), .B1(
        n21109), .B2(n20660), .ZN(n20662) );
  OAI211_X1 U23594 ( .C1(n9996), .C2(n20664), .A(n20663), .B(n20662), .ZN(
        P1_U3064) );
  NOR3_X1 U23595 ( .A1(n20922), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20699) );
  INV_X1 U23596 ( .A(n20699), .ZN(n20695) );
  NOR2_X1 U23597 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20695), .ZN(
        n20689) );
  NOR2_X1 U23598 ( .A1(n13832), .A2(n20665), .ZN(n20765) );
  NAND3_X1 U23599 ( .A1(n20765), .A2(n21206), .A3(n14077), .ZN(n20666) );
  OAI21_X1 U23600 ( .B1(n20667), .B2(n21012), .A(n20666), .ZN(n20688) );
  AOI22_X1 U23601 ( .A1(n21065), .A2(n20689), .B1(n21064), .B2(n20688), .ZN(
        n20675) );
  AOI21_X1 U23602 ( .B1(n20693), .B2(n20673), .A(n20927), .ZN(n20668) );
  AOI21_X1 U23603 ( .B1(n20765), .B2(n14077), .A(n20668), .ZN(n20669) );
  NOR2_X1 U23604 ( .A1(n20669), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20672) );
  INV_X1 U23605 ( .A(n21026), .ZN(n21074) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20690), .B1(
        n20716), .B2(n21074), .ZN(n20674) );
  OAI211_X1 U23607 ( .C1(n21077), .C2(n20693), .A(n20675), .B(n20674), .ZN(
        P1_U3065) );
  AOI22_X1 U23608 ( .A1(n21079), .A2(n20689), .B1(n21078), .B2(n20688), .ZN(
        n20677) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20690), .B1(
        n20716), .B2(n9999), .ZN(n20676) );
  OAI211_X1 U23610 ( .C1(n21082), .C2(n20693), .A(n20677), .B(n20676), .ZN(
        P1_U3066) );
  AOI22_X1 U23611 ( .A1(n21084), .A2(n20689), .B1(n21083), .B2(n20688), .ZN(
        n20679) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20690), .B1(
        n20716), .B2(n10001), .ZN(n20678) );
  OAI211_X1 U23613 ( .C1(n21087), .C2(n20693), .A(n20679), .B(n20678), .ZN(
        P1_U3067) );
  AOI22_X1 U23614 ( .A1(n21089), .A2(n20689), .B1(n21088), .B2(n20688), .ZN(
        n20681) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20690), .B1(
        n20716), .B2(n10003), .ZN(n20680) );
  OAI211_X1 U23616 ( .C1(n21092), .C2(n20693), .A(n20681), .B(n20680), .ZN(
        P1_U3068) );
  AOI22_X1 U23617 ( .A1(n21094), .A2(n20689), .B1(n21093), .B2(n20688), .ZN(
        n20683) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20690), .B1(
        n20716), .B2(n9990), .ZN(n20682) );
  OAI211_X1 U23619 ( .C1(n9994), .C2(n20693), .A(n20683), .B(n20682), .ZN(
        P1_U3069) );
  AOI22_X1 U23620 ( .A1(n21099), .A2(n20689), .B1(n21098), .B2(n20688), .ZN(
        n20685) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20690), .B1(
        n20716), .B2(n10005), .ZN(n20684) );
  OAI211_X1 U23622 ( .C1(n21102), .C2(n20693), .A(n20685), .B(n20684), .ZN(
        P1_U3070) );
  AOI22_X1 U23623 ( .A1(n21104), .A2(n20689), .B1(n21103), .B2(n20688), .ZN(
        n20687) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20690), .B1(
        n20716), .B2(n9997), .ZN(n20686) );
  OAI211_X1 U23625 ( .C1(n21107), .C2(n20693), .A(n20687), .B(n20686), .ZN(
        P1_U3071) );
  AOI22_X1 U23626 ( .A1(n21111), .A2(n20689), .B1(n21109), .B2(n20688), .ZN(
        n20692) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20690), .B1(
        n20716), .B2(n21112), .ZN(n20691) );
  OAI211_X1 U23628 ( .C1(n9996), .C2(n20693), .A(n20692), .B(n20691), .ZN(
        P1_U3072) );
  NOR2_X1 U23629 ( .A1(n21214), .A2(n20695), .ZN(n20715) );
  INV_X1 U23630 ( .A(n20561), .ZN(n20694) );
  AOI21_X1 U23631 ( .B1(n20765), .B2(n20694), .A(n20715), .ZN(n20696) );
  OAI22_X1 U23632 ( .A1(n20696), .A2(n21194), .B1(n20695), .B2(n20980), .ZN(
        n20714) );
  AOI22_X1 U23633 ( .A1(n21065), .A2(n20715), .B1(n21064), .B2(n20714), .ZN(
        n20701) );
  INV_X1 U23634 ( .A(n20764), .ZN(n20771) );
  NAND2_X1 U23635 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20771), .ZN(n20697) );
  NAND2_X1 U23636 ( .A1(n20697), .A2(n20696), .ZN(n20698) );
  OAI221_X1 U23637 ( .B1(n21206), .B2(n20699), .C1(n21194), .C2(n20698), .A(
        n21070), .ZN(n20717) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n21023), .ZN(n20700) );
  OAI211_X1 U23639 ( .C1(n21026), .C2(n20762), .A(n20701), .B(n20700), .ZN(
        P1_U3073) );
  AOI22_X1 U23640 ( .A1(n21079), .A2(n20715), .B1(n21078), .B2(n20714), .ZN(
        n20703) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n21027), .ZN(n20702) );
  OAI211_X1 U23642 ( .C1(n10000), .C2(n20762), .A(n20703), .B(n20702), .ZN(
        P1_U3074) );
  AOI22_X1 U23643 ( .A1(n21084), .A2(n20715), .B1(n21083), .B2(n20714), .ZN(
        n20705) );
  AOI22_X1 U23644 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n21031), .ZN(n20704) );
  OAI211_X1 U23645 ( .C1(n10002), .C2(n20762), .A(n20705), .B(n20704), .ZN(
        P1_U3075) );
  AOI22_X1 U23646 ( .A1(n21089), .A2(n20715), .B1(n21088), .B2(n20714), .ZN(
        n20707) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n21035), .ZN(n20706) );
  OAI211_X1 U23648 ( .C1(n10004), .C2(n20762), .A(n20707), .B(n20706), .ZN(
        P1_U3076) );
  AOI22_X1 U23649 ( .A1(n21094), .A2(n20715), .B1(n21093), .B2(n20714), .ZN(
        n20709) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n9993), .ZN(n20708) );
  OAI211_X1 U23651 ( .C1(n21041), .C2(n20762), .A(n20709), .B(n20708), .ZN(
        P1_U3077) );
  AOI22_X1 U23652 ( .A1(n21099), .A2(n20715), .B1(n21098), .B2(n20714), .ZN(
        n20711) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n21042), .ZN(n20710) );
  OAI211_X1 U23654 ( .C1(n10006), .C2(n20762), .A(n20711), .B(n20710), .ZN(
        P1_U3078) );
  AOI22_X1 U23655 ( .A1(n21104), .A2(n20715), .B1(n21103), .B2(n20714), .ZN(
        n20713) );
  AOI22_X1 U23656 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n21046), .ZN(n20712) );
  OAI211_X1 U23657 ( .C1(n9998), .C2(n20762), .A(n20713), .B(n20712), .ZN(
        P1_U3079) );
  AOI22_X1 U23658 ( .A1(n21111), .A2(n20715), .B1(n21109), .B2(n20714), .ZN(
        n20719) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20717), .B1(
        n20716), .B2(n9995), .ZN(n20718) );
  OAI211_X1 U23660 ( .C1(n21056), .C2(n20762), .A(n20719), .B(n20718), .ZN(
        P1_U3080) );
  NAND2_X1 U23661 ( .A1(n21214), .A2(n10375), .ZN(n20756) );
  OR2_X1 U23662 ( .A1(n20762), .A2(n21077), .ZN(n20720) );
  OAI21_X1 U23663 ( .B1(n20925), .B2(n20756), .A(n20720), .ZN(n20721) );
  INV_X1 U23664 ( .A(n20721), .ZN(n20730) );
  OR2_X1 U23665 ( .A1(n20764), .A2(n21014), .ZN(n20722) );
  AND2_X1 U23666 ( .A1(n20722), .A2(n21206), .ZN(n20725) );
  NAND2_X1 U23667 ( .A1(n20765), .A2(n21016), .ZN(n20727) );
  AOI22_X1 U23668 ( .A1(n20725), .A2(n20727), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20756), .ZN(n20724) );
  NAND3_X1 U23669 ( .A1(n21021), .A2(n20724), .A3(n20723), .ZN(n20759) );
  INV_X1 U23670 ( .A(n20725), .ZN(n20728) );
  OAI22_X1 U23671 ( .A1(n20728), .A2(n20727), .B1(n21012), .B2(n20726), .ZN(
        n20758) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20759), .B1(
        n21064), .B2(n20758), .ZN(n20729) );
  OAI211_X1 U23673 ( .C1(n21026), .C2(n20775), .A(n20730), .B(n20729), .ZN(
        P1_U3081) );
  OR2_X1 U23674 ( .A1(n20775), .A2(n10000), .ZN(n20731) );
  OAI21_X1 U23675 ( .B1(n20940), .B2(n20756), .A(n20731), .ZN(n20732) );
  INV_X1 U23676 ( .A(n20732), .ZN(n20734) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20759), .B1(
        n21078), .B2(n20758), .ZN(n20733) );
  OAI211_X1 U23678 ( .C1(n21082), .C2(n20762), .A(n20734), .B(n20733), .ZN(
        P1_U3082) );
  OR2_X1 U23679 ( .A1(n20775), .A2(n10002), .ZN(n20735) );
  OAI21_X1 U23680 ( .B1(n20945), .B2(n20756), .A(n20735), .ZN(n20736) );
  INV_X1 U23681 ( .A(n20736), .ZN(n20738) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20759), .B1(
        n21083), .B2(n20758), .ZN(n20737) );
  OAI211_X1 U23683 ( .C1(n21087), .C2(n20762), .A(n20738), .B(n20737), .ZN(
        P1_U3083) );
  OR2_X1 U23684 ( .A1(n20762), .A2(n21092), .ZN(n20739) );
  OAI21_X1 U23685 ( .B1(n20950), .B2(n20756), .A(n20739), .ZN(n20740) );
  INV_X1 U23686 ( .A(n20740), .ZN(n20742) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20759), .B1(
        n21088), .B2(n20758), .ZN(n20741) );
  OAI211_X1 U23688 ( .C1(n10004), .C2(n20775), .A(n20742), .B(n20741), .ZN(
        P1_U3084) );
  OR2_X1 U23689 ( .A1(n20775), .A2(n21041), .ZN(n20743) );
  OAI21_X1 U23690 ( .B1(n20955), .B2(n20756), .A(n20743), .ZN(n20744) );
  INV_X1 U23691 ( .A(n20744), .ZN(n20746) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20759), .B1(
        n21093), .B2(n20758), .ZN(n20745) );
  OAI211_X1 U23693 ( .C1(n9994), .C2(n20762), .A(n20746), .B(n20745), .ZN(
        P1_U3085) );
  OR2_X1 U23694 ( .A1(n20762), .A2(n21102), .ZN(n20747) );
  OAI21_X1 U23695 ( .B1(n20960), .B2(n20756), .A(n20747), .ZN(n20748) );
  INV_X1 U23696 ( .A(n20748), .ZN(n20750) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20759), .B1(
        n21098), .B2(n20758), .ZN(n20749) );
  OAI211_X1 U23698 ( .C1(n10006), .C2(n20775), .A(n20750), .B(n20749), .ZN(
        P1_U3086) );
  OR2_X1 U23699 ( .A1(n20775), .A2(n9998), .ZN(n20751) );
  OAI21_X1 U23700 ( .B1(n20965), .B2(n20756), .A(n20751), .ZN(n20752) );
  INV_X1 U23701 ( .A(n20752), .ZN(n20754) );
  AOI22_X1 U23702 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20759), .B1(
        n21103), .B2(n20758), .ZN(n20753) );
  OAI211_X1 U23703 ( .C1(n21107), .C2(n20762), .A(n20754), .B(n20753), .ZN(
        P1_U3087) );
  OR2_X1 U23704 ( .A1(n20775), .A2(n21056), .ZN(n20755) );
  OAI21_X1 U23705 ( .B1(n20971), .B2(n20756), .A(n20755), .ZN(n20757) );
  INV_X1 U23706 ( .A(n20757), .ZN(n20761) );
  AOI22_X1 U23707 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20759), .B1(
        n21109), .B2(n20758), .ZN(n20760) );
  OAI211_X1 U23708 ( .C1(n9996), .C2(n20762), .A(n20761), .B(n20760), .ZN(
        P1_U3088) );
  INV_X1 U23709 ( .A(n20766), .ZN(n20791) );
  NAND2_X1 U23710 ( .A1(n20765), .A2(n21057), .ZN(n20767) );
  NAND2_X1 U23711 ( .A1(n20767), .A2(n20766), .ZN(n20772) );
  NAND2_X1 U23712 ( .A1(n20772), .A2(n21206), .ZN(n20769) );
  NAND2_X1 U23713 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n10375), .ZN(n20768) );
  NAND2_X1 U23714 ( .A1(n20769), .A2(n20768), .ZN(n20790) );
  AOI22_X1 U23715 ( .A1(n21065), .A2(n20791), .B1(n21064), .B2(n20790), .ZN(
        n20777) );
  INV_X1 U23716 ( .A(n21068), .ZN(n20770) );
  NAND2_X1 U23717 ( .A1(n20771), .A2(n20770), .ZN(n21196) );
  INV_X1 U23718 ( .A(n20772), .ZN(n20773) );
  NAND2_X1 U23719 ( .A1(n21196), .A2(n20773), .ZN(n20774) );
  OAI221_X1 U23720 ( .B1(n21206), .B2(n10375), .C1(n21194), .C2(n20774), .A(
        n21070), .ZN(n20793) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21023), .ZN(n20776) );
  OAI211_X1 U23722 ( .C1(n21026), .C2(n20800), .A(n20777), .B(n20776), .ZN(
        P1_U3089) );
  AOI22_X1 U23723 ( .A1(n21079), .A2(n20791), .B1(n21078), .B2(n20790), .ZN(
        n20779) );
  AOI22_X1 U23724 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21027), .ZN(n20778) );
  OAI211_X1 U23725 ( .C1(n10000), .C2(n20800), .A(n20779), .B(n20778), .ZN(
        P1_U3090) );
  AOI22_X1 U23726 ( .A1(n21084), .A2(n20791), .B1(n21083), .B2(n20790), .ZN(
        n20781) );
  AOI22_X1 U23727 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21031), .ZN(n20780) );
  OAI211_X1 U23728 ( .C1(n10002), .C2(n20800), .A(n20781), .B(n20780), .ZN(
        P1_U3091) );
  AOI22_X1 U23729 ( .A1(n21089), .A2(n20791), .B1(n21088), .B2(n20790), .ZN(
        n20783) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21035), .ZN(n20782) );
  OAI211_X1 U23731 ( .C1(n10004), .C2(n20800), .A(n20783), .B(n20782), .ZN(
        P1_U3092) );
  AOI22_X1 U23732 ( .A1(n21094), .A2(n20791), .B1(n21093), .B2(n20790), .ZN(
        n20785) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n9993), .ZN(n20784) );
  OAI211_X1 U23734 ( .C1(n21041), .C2(n20800), .A(n20785), .B(n20784), .ZN(
        P1_U3093) );
  AOI22_X1 U23735 ( .A1(n21099), .A2(n20791), .B1(n21098), .B2(n20790), .ZN(
        n20787) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21042), .ZN(n20786) );
  OAI211_X1 U23737 ( .C1(n10006), .C2(n20800), .A(n20787), .B(n20786), .ZN(
        P1_U3094) );
  AOI22_X1 U23738 ( .A1(n21104), .A2(n20791), .B1(n21103), .B2(n20790), .ZN(
        n20789) );
  AOI22_X1 U23739 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21046), .ZN(n20788) );
  OAI211_X1 U23740 ( .C1(n9998), .C2(n20800), .A(n20789), .B(n20788), .ZN(
        P1_U3095) );
  AOI22_X1 U23741 ( .A1(n21111), .A2(n20791), .B1(n21109), .B2(n20790), .ZN(
        n20795) );
  AOI22_X1 U23742 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n9995), .ZN(n20794) );
  OAI211_X1 U23743 ( .C1(n21056), .C2(n20800), .A(n20795), .B(n20794), .ZN(
        P1_U3096) );
  INV_X1 U23744 ( .A(n15120), .ZN(n20796) );
  INV_X1 U23745 ( .A(n20923), .ZN(n20797) );
  NAND3_X1 U23746 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20922), .A3(
        n20850), .ZN(n20827) );
  NOR2_X1 U23747 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20827), .ZN(
        n20820) );
  AND2_X1 U23748 ( .A1(n14039), .A2(n13832), .ZN(n20892) );
  AOI21_X1 U23749 ( .B1(n20892), .B2(n14077), .A(n20820), .ZN(n20802) );
  INV_X1 U23750 ( .A(n20798), .ZN(n20799) );
  NAND2_X1 U23751 ( .A1(n20799), .A2(n20853), .ZN(n20934) );
  OAI22_X1 U23752 ( .A1(n20802), .A2(n21194), .B1(n20934), .B2(n20859), .ZN(
        n20819) );
  AOI22_X1 U23753 ( .A1(n21065), .A2(n20820), .B1(n21064), .B2(n20819), .ZN(
        n20806) );
  INV_X1 U23754 ( .A(n20849), .ZN(n20801) );
  OAI21_X1 U23755 ( .B1(n20801), .B2(n20821), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20803) );
  NAND2_X1 U23756 ( .A1(n20803), .A2(n20802), .ZN(n20804) );
  AOI22_X1 U23757 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20822), .B1(
        n20821), .B2(n21023), .ZN(n20805) );
  OAI211_X1 U23758 ( .C1(n21026), .C2(n20849), .A(n20806), .B(n20805), .ZN(
        P1_U3097) );
  AOI22_X1 U23759 ( .A1(n21079), .A2(n20820), .B1(n21078), .B2(n20819), .ZN(
        n20808) );
  AOI22_X1 U23760 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20822), .B1(
        n20821), .B2(n21027), .ZN(n20807) );
  OAI211_X1 U23761 ( .C1(n10000), .C2(n20849), .A(n20808), .B(n20807), .ZN(
        P1_U3098) );
  AOI22_X1 U23762 ( .A1(n21084), .A2(n20820), .B1(n21083), .B2(n20819), .ZN(
        n20810) );
  AOI22_X1 U23763 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20822), .B1(
        n20821), .B2(n21031), .ZN(n20809) );
  OAI211_X1 U23764 ( .C1(n10002), .C2(n20849), .A(n20810), .B(n20809), .ZN(
        P1_U3099) );
  AOI22_X1 U23765 ( .A1(n21089), .A2(n20820), .B1(n21088), .B2(n20819), .ZN(
        n20812) );
  AOI22_X1 U23766 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20822), .B1(
        n20821), .B2(n21035), .ZN(n20811) );
  OAI211_X1 U23767 ( .C1(n10004), .C2(n20849), .A(n20812), .B(n20811), .ZN(
        P1_U3100) );
  AOI22_X1 U23768 ( .A1(n21094), .A2(n20820), .B1(n21093), .B2(n20819), .ZN(
        n20814) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20822), .B1(
        n20821), .B2(n9993), .ZN(n20813) );
  OAI211_X1 U23770 ( .C1(n21041), .C2(n20849), .A(n20814), .B(n20813), .ZN(
        P1_U3101) );
  AOI22_X1 U23771 ( .A1(n21099), .A2(n20820), .B1(n21098), .B2(n20819), .ZN(
        n20816) );
  AOI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20822), .B1(
        n20821), .B2(n21042), .ZN(n20815) );
  OAI211_X1 U23773 ( .C1(n10006), .C2(n20849), .A(n20816), .B(n20815), .ZN(
        P1_U3102) );
  AOI22_X1 U23774 ( .A1(n21104), .A2(n20820), .B1(n21103), .B2(n20819), .ZN(
        n20818) );
  AOI22_X1 U23775 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20822), .B1(
        n20821), .B2(n21046), .ZN(n20817) );
  OAI211_X1 U23776 ( .C1(n9998), .C2(n20849), .A(n20818), .B(n20817), .ZN(
        P1_U3103) );
  AOI22_X1 U23777 ( .A1(n21111), .A2(n20820), .B1(n21109), .B2(n20819), .ZN(
        n20824) );
  AOI22_X1 U23778 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20822), .B1(
        n20821), .B2(n9995), .ZN(n20823) );
  OAI211_X1 U23779 ( .C1(n21056), .C2(n20849), .A(n20824), .B(n20823), .ZN(
        P1_U3104) );
  NOR2_X1 U23780 ( .A1(n21214), .A2(n20827), .ZN(n20844) );
  INV_X1 U23781 ( .A(n20892), .ZN(n20826) );
  INV_X1 U23782 ( .A(n20844), .ZN(n20825) );
  OAI222_X1 U23783 ( .A1(n20978), .A2(n20826), .B1(n20980), .B2(n20827), .C1(
        n21194), .C2(n20825), .ZN(n20843) );
  AOI22_X1 U23784 ( .A1(n21065), .A2(n20844), .B1(n21064), .B2(n20843), .ZN(
        n20830) );
  OAI21_X1 U23785 ( .B1(n21195), .B2(n20985), .A(n20827), .ZN(n20828) );
  NAND2_X1 U23786 ( .A1(n20828), .A2(n21070), .ZN(n20846) );
  AOI22_X1 U23787 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20846), .B1(
        n20845), .B2(n21074), .ZN(n20829) );
  OAI211_X1 U23788 ( .C1(n21077), .C2(n20849), .A(n20830), .B(n20829), .ZN(
        P1_U3105) );
  AOI22_X1 U23789 ( .A1(n21079), .A2(n20844), .B1(n21078), .B2(n20843), .ZN(
        n20832) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20846), .B1(
        n20845), .B2(n9999), .ZN(n20831) );
  OAI211_X1 U23791 ( .C1(n21082), .C2(n20849), .A(n20832), .B(n20831), .ZN(
        P1_U3106) );
  AOI22_X1 U23792 ( .A1(n21084), .A2(n20844), .B1(n21083), .B2(n20843), .ZN(
        n20834) );
  AOI22_X1 U23793 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20846), .B1(
        n20845), .B2(n10001), .ZN(n20833) );
  OAI211_X1 U23794 ( .C1(n21087), .C2(n20849), .A(n20834), .B(n20833), .ZN(
        P1_U3107) );
  AOI22_X1 U23795 ( .A1(n21089), .A2(n20844), .B1(n21088), .B2(n20843), .ZN(
        n20836) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20846), .B1(
        n20845), .B2(n10003), .ZN(n20835) );
  OAI211_X1 U23797 ( .C1(n21092), .C2(n20849), .A(n20836), .B(n20835), .ZN(
        P1_U3108) );
  AOI22_X1 U23798 ( .A1(n21094), .A2(n20844), .B1(n21093), .B2(n20843), .ZN(
        n20838) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20846), .B1(
        n20845), .B2(n9990), .ZN(n20837) );
  OAI211_X1 U23800 ( .C1(n9994), .C2(n20849), .A(n20838), .B(n20837), .ZN(
        P1_U3109) );
  AOI22_X1 U23801 ( .A1(n21099), .A2(n20844), .B1(n21098), .B2(n20843), .ZN(
        n20840) );
  AOI22_X1 U23802 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20846), .B1(
        n20845), .B2(n10005), .ZN(n20839) );
  OAI211_X1 U23803 ( .C1(n21102), .C2(n20849), .A(n20840), .B(n20839), .ZN(
        P1_U3110) );
  AOI22_X1 U23804 ( .A1(n21104), .A2(n20844), .B1(n21103), .B2(n20843), .ZN(
        n20842) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20846), .B1(
        n20845), .B2(n9997), .ZN(n20841) );
  OAI211_X1 U23806 ( .C1(n21107), .C2(n20849), .A(n20842), .B(n20841), .ZN(
        P1_U3111) );
  AOI22_X1 U23807 ( .A1(n21111), .A2(n20844), .B1(n21109), .B2(n20843), .ZN(
        n20848) );
  AOI22_X1 U23808 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20846), .B1(
        n20845), .B2(n21112), .ZN(n20847) );
  OAI211_X1 U23809 ( .C1(n9996), .C2(n20849), .A(n20848), .B(n20847), .ZN(
        P1_U3112) );
  NOR3_X1 U23810 ( .A1(n21205), .A2(n20850), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20900) );
  INV_X1 U23811 ( .A(n20900), .ZN(n20851) );
  NOR2_X1 U23812 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20851), .ZN(
        n20854) );
  INV_X1 U23813 ( .A(n20854), .ZN(n20882) );
  OAI22_X1 U23814 ( .A1(n20901), .A2(n21026), .B1(n20925), .B2(n20882), .ZN(
        n20852) );
  INV_X1 U23815 ( .A(n20852), .ZN(n20863) );
  OAI21_X1 U23816 ( .B1(n21195), .B2(n21014), .A(n21206), .ZN(n20861) );
  AND2_X1 U23817 ( .A1(n20892), .A2(n21016), .ZN(n20858) );
  OR2_X1 U23818 ( .A1(n20853), .A2(n21205), .ZN(n21011) );
  NAND2_X1 U23819 ( .A1(n21011), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21020) );
  OAI21_X1 U23820 ( .B1(n20931), .B2(n20854), .A(n21020), .ZN(n20855) );
  INV_X1 U23821 ( .A(n20855), .ZN(n20857) );
  OAI211_X1 U23822 ( .C1(n20861), .C2(n20858), .A(n20857), .B(n20856), .ZN(
        n20886) );
  INV_X1 U23823 ( .A(n20858), .ZN(n20860) );
  OAI22_X1 U23824 ( .A1(n20861), .A2(n20860), .B1(n20859), .B2(n21011), .ZN(
        n20885) );
  AOI22_X1 U23825 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20886), .B1(
        n21064), .B2(n20885), .ZN(n20862) );
  OAI211_X1 U23826 ( .C1(n21077), .C2(n20883), .A(n20863), .B(n20862), .ZN(
        P1_U3113) );
  OAI22_X1 U23827 ( .A1(n20901), .A2(n10000), .B1(n20882), .B2(n20940), .ZN(
        n20864) );
  INV_X1 U23828 ( .A(n20864), .ZN(n20866) );
  AOI22_X1 U23829 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20886), .B1(
        n21078), .B2(n20885), .ZN(n20865) );
  OAI211_X1 U23830 ( .C1(n21082), .C2(n20883), .A(n20866), .B(n20865), .ZN(
        P1_U3114) );
  OAI22_X1 U23831 ( .A1(n20901), .A2(n10002), .B1(n20882), .B2(n20945), .ZN(
        n20867) );
  INV_X1 U23832 ( .A(n20867), .ZN(n20869) );
  AOI22_X1 U23833 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20886), .B1(
        n21083), .B2(n20885), .ZN(n20868) );
  OAI211_X1 U23834 ( .C1(n21087), .C2(n20883), .A(n20869), .B(n20868), .ZN(
        P1_U3115) );
  OAI22_X1 U23835 ( .A1(n20883), .A2(n21092), .B1(n20882), .B2(n20950), .ZN(
        n20870) );
  INV_X1 U23836 ( .A(n20870), .ZN(n20872) );
  AOI22_X1 U23837 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20886), .B1(
        n21088), .B2(n20885), .ZN(n20871) );
  OAI211_X1 U23838 ( .C1(n10004), .C2(n20901), .A(n20872), .B(n20871), .ZN(
        P1_U3116) );
  OAI22_X1 U23839 ( .A1(n20883), .A2(n9994), .B1(n20882), .B2(n20955), .ZN(
        n20873) );
  INV_X1 U23840 ( .A(n20873), .ZN(n20875) );
  AOI22_X1 U23841 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20886), .B1(
        n21093), .B2(n20885), .ZN(n20874) );
  OAI211_X1 U23842 ( .C1(n21041), .C2(n20901), .A(n20875), .B(n20874), .ZN(
        P1_U3117) );
  OAI22_X1 U23843 ( .A1(n20901), .A2(n10006), .B1(n20960), .B2(n20882), .ZN(
        n20876) );
  INV_X1 U23844 ( .A(n20876), .ZN(n20878) );
  AOI22_X1 U23845 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20886), .B1(
        n21098), .B2(n20885), .ZN(n20877) );
  OAI211_X1 U23846 ( .C1(n21102), .C2(n20883), .A(n20878), .B(n20877), .ZN(
        P1_U3118) );
  OAI22_X1 U23847 ( .A1(n20883), .A2(n21107), .B1(n20965), .B2(n20882), .ZN(
        n20879) );
  INV_X1 U23848 ( .A(n20879), .ZN(n20881) );
  AOI22_X1 U23849 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20886), .B1(
        n21103), .B2(n20885), .ZN(n20880) );
  OAI211_X1 U23850 ( .C1(n9998), .C2(n20901), .A(n20881), .B(n20880), .ZN(
        P1_U3119) );
  OAI22_X1 U23851 ( .A1(n20883), .A2(n9996), .B1(n20971), .B2(n20882), .ZN(
        n20884) );
  INV_X1 U23852 ( .A(n20884), .ZN(n20888) );
  AOI22_X1 U23853 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20886), .B1(
        n21109), .B2(n20885), .ZN(n20887) );
  OAI211_X1 U23854 ( .C1(n21056), .C2(n20901), .A(n20888), .B(n20887), .ZN(
        P1_U3120) );
  OR2_X1 U23855 ( .A1(n20891), .A2(n21205), .ZN(n20893) );
  INV_X1 U23856 ( .A(n20893), .ZN(n20917) );
  NAND2_X1 U23857 ( .A1(n20892), .A2(n21057), .ZN(n20894) );
  NAND2_X1 U23858 ( .A1(n20894), .A2(n20893), .ZN(n20897) );
  NAND2_X1 U23859 ( .A1(n20897), .A2(n21206), .ZN(n20896) );
  NAND2_X1 U23860 ( .A1(n20900), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20895) );
  NAND2_X1 U23861 ( .A1(n20896), .A2(n20895), .ZN(n20916) );
  AOI22_X1 U23862 ( .A1(n21065), .A2(n20917), .B1(n21064), .B2(n20916), .ZN(
        n20903) );
  INV_X1 U23863 ( .A(n20897), .ZN(n20898) );
  OAI21_X1 U23864 ( .B1(n21195), .B2(n21068), .A(n20898), .ZN(n20899) );
  OAI221_X1 U23865 ( .B1(n21206), .B2(n20900), .C1(n21194), .C2(n20899), .A(
        n21070), .ZN(n20919) );
  AOI22_X1 U23866 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20919), .B1(
        n20918), .B2(n21023), .ZN(n20902) );
  OAI211_X1 U23867 ( .C1(n21026), .C2(n20977), .A(n20903), .B(n20902), .ZN(
        P1_U3121) );
  AOI22_X1 U23868 ( .A1(n21079), .A2(n20917), .B1(n21078), .B2(n20916), .ZN(
        n20905) );
  AOI22_X1 U23869 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20919), .B1(
        n20918), .B2(n21027), .ZN(n20904) );
  OAI211_X1 U23870 ( .C1(n10000), .C2(n20977), .A(n20905), .B(n20904), .ZN(
        P1_U3122) );
  AOI22_X1 U23871 ( .A1(n21084), .A2(n20917), .B1(n21083), .B2(n20916), .ZN(
        n20907) );
  AOI22_X1 U23872 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20919), .B1(
        n20918), .B2(n21031), .ZN(n20906) );
  OAI211_X1 U23873 ( .C1(n10002), .C2(n20977), .A(n20907), .B(n20906), .ZN(
        P1_U3123) );
  AOI22_X1 U23874 ( .A1(n21089), .A2(n20917), .B1(n21088), .B2(n20916), .ZN(
        n20909) );
  AOI22_X1 U23875 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20919), .B1(
        n20918), .B2(n21035), .ZN(n20908) );
  OAI211_X1 U23876 ( .C1(n10004), .C2(n20977), .A(n20909), .B(n20908), .ZN(
        P1_U3124) );
  AOI22_X1 U23877 ( .A1(n21094), .A2(n20917), .B1(n21093), .B2(n20916), .ZN(
        n20911) );
  AOI22_X1 U23878 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20919), .B1(
        n20918), .B2(n9993), .ZN(n20910) );
  OAI211_X1 U23879 ( .C1(n21041), .C2(n20977), .A(n20911), .B(n20910), .ZN(
        P1_U3125) );
  AOI22_X1 U23880 ( .A1(n21099), .A2(n20917), .B1(n21098), .B2(n20916), .ZN(
        n20913) );
  AOI22_X1 U23881 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20919), .B1(
        n20918), .B2(n21042), .ZN(n20912) );
  OAI211_X1 U23882 ( .C1(n10006), .C2(n20977), .A(n20913), .B(n20912), .ZN(
        P1_U3126) );
  AOI22_X1 U23883 ( .A1(n21104), .A2(n20917), .B1(n21103), .B2(n20916), .ZN(
        n20915) );
  AOI22_X1 U23884 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20919), .B1(
        n20918), .B2(n21046), .ZN(n20914) );
  OAI211_X1 U23885 ( .C1(n9998), .C2(n20977), .A(n20915), .B(n20914), .ZN(
        P1_U3127) );
  AOI22_X1 U23886 ( .A1(n21111), .A2(n20917), .B1(n21109), .B2(n20916), .ZN(
        n20921) );
  AOI22_X1 U23887 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20919), .B1(
        n20918), .B2(n9995), .ZN(n20920) );
  OAI211_X1 U23888 ( .C1(n21056), .C2(n20977), .A(n20921), .B(n20920), .ZN(
        P1_U3128) );
  NOR3_X1 U23889 ( .A1(n20922), .A2(n21205), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20986) );
  INV_X1 U23890 ( .A(n20986), .ZN(n20981) );
  NOR2_X1 U23891 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20981), .ZN(
        n20932) );
  INV_X1 U23892 ( .A(n20932), .ZN(n20970) );
  OR2_X1 U23893 ( .A1(n21007), .A2(n21026), .ZN(n20924) );
  OAI21_X1 U23894 ( .B1(n20925), .B2(n20970), .A(n20924), .ZN(n20926) );
  INV_X1 U23895 ( .A(n20926), .ZN(n20938) );
  AOI21_X1 U23896 ( .B1(n20977), .B2(n21007), .A(n20927), .ZN(n20928) );
  NOR2_X1 U23897 ( .A1(n20928), .A2(n21194), .ZN(n20933) );
  OR2_X1 U23898 ( .A1(n13832), .A2(n20929), .ZN(n21059) );
  OR2_X1 U23899 ( .A1(n21059), .A2(n21016), .ZN(n20935) );
  AOI22_X1 U23900 ( .A1(n20933), .A2(n20935), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20934), .ZN(n20930) );
  OAI211_X1 U23901 ( .C1(n20932), .C2(n20931), .A(n21021), .B(n20930), .ZN(
        n20974) );
  INV_X1 U23902 ( .A(n20933), .ZN(n20936) );
  AOI22_X1 U23903 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20974), .B1(
        n21064), .B2(n20973), .ZN(n20937) );
  OAI211_X1 U23904 ( .C1(n21077), .C2(n20977), .A(n20938), .B(n20937), .ZN(
        P1_U3129) );
  OR2_X1 U23905 ( .A1(n21007), .A2(n10000), .ZN(n20939) );
  OAI21_X1 U23906 ( .B1(n20940), .B2(n20970), .A(n20939), .ZN(n20941) );
  INV_X1 U23907 ( .A(n20941), .ZN(n20943) );
  AOI22_X1 U23908 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20974), .B1(
        n21078), .B2(n20973), .ZN(n20942) );
  OAI211_X1 U23909 ( .C1(n21082), .C2(n20977), .A(n20943), .B(n20942), .ZN(
        P1_U3130) );
  OR2_X1 U23910 ( .A1(n21007), .A2(n10002), .ZN(n20944) );
  OAI21_X1 U23911 ( .B1(n20945), .B2(n20970), .A(n20944), .ZN(n20946) );
  INV_X1 U23912 ( .A(n20946), .ZN(n20948) );
  AOI22_X1 U23913 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20974), .B1(
        n21083), .B2(n20973), .ZN(n20947) );
  OAI211_X1 U23914 ( .C1(n21087), .C2(n20977), .A(n20948), .B(n20947), .ZN(
        P1_U3131) );
  OR2_X1 U23915 ( .A1(n21007), .A2(n10004), .ZN(n20949) );
  OAI21_X1 U23916 ( .B1(n20950), .B2(n20970), .A(n20949), .ZN(n20951) );
  INV_X1 U23917 ( .A(n20951), .ZN(n20953) );
  AOI22_X1 U23918 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20974), .B1(
        n21088), .B2(n20973), .ZN(n20952) );
  OAI211_X1 U23919 ( .C1(n21092), .C2(n20977), .A(n20953), .B(n20952), .ZN(
        P1_U3132) );
  OR2_X1 U23920 ( .A1(n21007), .A2(n21041), .ZN(n20954) );
  OAI21_X1 U23921 ( .B1(n20955), .B2(n20970), .A(n20954), .ZN(n20956) );
  INV_X1 U23922 ( .A(n20956), .ZN(n20958) );
  AOI22_X1 U23923 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20974), .B1(
        n21093), .B2(n20973), .ZN(n20957) );
  OAI211_X1 U23924 ( .C1(n9994), .C2(n20977), .A(n20958), .B(n20957), .ZN(
        P1_U3133) );
  OR2_X1 U23925 ( .A1(n21007), .A2(n10006), .ZN(n20959) );
  OAI21_X1 U23926 ( .B1(n20960), .B2(n20970), .A(n20959), .ZN(n20961) );
  INV_X1 U23927 ( .A(n20961), .ZN(n20963) );
  AOI22_X1 U23928 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20974), .B1(
        n21098), .B2(n20973), .ZN(n20962) );
  OAI211_X1 U23929 ( .C1(n21102), .C2(n20977), .A(n20963), .B(n20962), .ZN(
        P1_U3134) );
  OR2_X1 U23930 ( .A1(n21007), .A2(n9998), .ZN(n20964) );
  OAI21_X1 U23931 ( .B1(n20965), .B2(n20970), .A(n20964), .ZN(n20966) );
  INV_X1 U23932 ( .A(n20966), .ZN(n20968) );
  AOI22_X1 U23933 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20974), .B1(
        n21103), .B2(n20973), .ZN(n20967) );
  OAI211_X1 U23934 ( .C1(n21107), .C2(n20977), .A(n20968), .B(n20967), .ZN(
        P1_U3135) );
  OR2_X1 U23935 ( .A1(n21007), .A2(n21056), .ZN(n20969) );
  OAI21_X1 U23936 ( .B1(n20971), .B2(n20970), .A(n20969), .ZN(n20972) );
  INV_X1 U23937 ( .A(n20972), .ZN(n20976) );
  AOI22_X1 U23938 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20974), .B1(
        n21109), .B2(n20973), .ZN(n20975) );
  OAI211_X1 U23939 ( .C1(n9996), .C2(n20977), .A(n20976), .B(n20975), .ZN(
        P1_U3136) );
  NOR2_X1 U23940 ( .A1(n21214), .A2(n20981), .ZN(n21003) );
  OR2_X1 U23941 ( .A1(n21059), .A2(n20978), .ZN(n20984) );
  INV_X1 U23942 ( .A(n21003), .ZN(n20979) );
  OAI22_X1 U23943 ( .A1(n20981), .A2(n20980), .B1(n21194), .B2(n20979), .ZN(
        n20982) );
  INV_X1 U23944 ( .A(n20982), .ZN(n20983) );
  NAND2_X1 U23945 ( .A1(n20984), .A2(n20983), .ZN(n21002) );
  AOI22_X1 U23946 ( .A1(n21065), .A2(n21003), .B1(n21064), .B2(n21002), .ZN(
        n20989) );
  NOR2_X1 U23947 ( .A1(n21069), .A2(n20985), .ZN(n21202) );
  OAI21_X1 U23948 ( .B1(n20986), .B2(n21202), .A(n21070), .ZN(n21004) );
  NOR2_X2 U23949 ( .A1(n21069), .A2(n20987), .ZN(n21052) );
  AOI22_X1 U23950 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21004), .B1(
        n21052), .B2(n21074), .ZN(n20988) );
  OAI211_X1 U23951 ( .C1(n21077), .C2(n21007), .A(n20989), .B(n20988), .ZN(
        P1_U3137) );
  AOI22_X1 U23952 ( .A1(n21079), .A2(n21003), .B1(n21078), .B2(n21002), .ZN(
        n20991) );
  AOI22_X1 U23953 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21004), .B1(
        n21052), .B2(n9999), .ZN(n20990) );
  OAI211_X1 U23954 ( .C1(n21082), .C2(n21007), .A(n20991), .B(n20990), .ZN(
        P1_U3138) );
  AOI22_X1 U23955 ( .A1(n21084), .A2(n21003), .B1(n21083), .B2(n21002), .ZN(
        n20993) );
  AOI22_X1 U23956 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21004), .B1(
        n21052), .B2(n10001), .ZN(n20992) );
  OAI211_X1 U23957 ( .C1(n21087), .C2(n21007), .A(n20993), .B(n20992), .ZN(
        P1_U3139) );
  AOI22_X1 U23958 ( .A1(n21089), .A2(n21003), .B1(n21088), .B2(n21002), .ZN(
        n20995) );
  AOI22_X1 U23959 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21004), .B1(
        n21052), .B2(n10003), .ZN(n20994) );
  OAI211_X1 U23960 ( .C1(n21092), .C2(n21007), .A(n20995), .B(n20994), .ZN(
        P1_U3140) );
  AOI22_X1 U23961 ( .A1(n21094), .A2(n21003), .B1(n21093), .B2(n21002), .ZN(
        n20997) );
  AOI22_X1 U23962 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21004), .B1(
        n21052), .B2(n9990), .ZN(n20996) );
  OAI211_X1 U23963 ( .C1(n9994), .C2(n21007), .A(n20997), .B(n20996), .ZN(
        P1_U3141) );
  AOI22_X1 U23964 ( .A1(n21099), .A2(n21003), .B1(n21098), .B2(n21002), .ZN(
        n20999) );
  AOI22_X1 U23965 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21004), .B1(
        n21052), .B2(n10005), .ZN(n20998) );
  OAI211_X1 U23966 ( .C1(n21102), .C2(n21007), .A(n20999), .B(n20998), .ZN(
        P1_U3142) );
  AOI22_X1 U23967 ( .A1(n21104), .A2(n21003), .B1(n21103), .B2(n21002), .ZN(
        n21001) );
  AOI22_X1 U23968 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21004), .B1(
        n21052), .B2(n9997), .ZN(n21000) );
  OAI211_X1 U23969 ( .C1(n21107), .C2(n21007), .A(n21001), .B(n21000), .ZN(
        P1_U3143) );
  AOI22_X1 U23970 ( .A1(n21111), .A2(n21003), .B1(n21109), .B2(n21002), .ZN(
        n21006) );
  AOI22_X1 U23971 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21004), .B1(
        n21052), .B2(n21112), .ZN(n21005) );
  OAI211_X1 U23972 ( .C1(n9996), .C2(n21007), .A(n21006), .B(n21005), .ZN(
        P1_U3144) );
  INV_X1 U23973 ( .A(n21069), .ZN(n21018) );
  INV_X1 U23974 ( .A(n21008), .ZN(n21009) );
  INV_X1 U23975 ( .A(n21072), .ZN(n21010) );
  NOR2_X1 U23976 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21010), .ZN(
        n21051) );
  NAND2_X1 U23977 ( .A1(n21016), .A2(n21206), .ZN(n21013) );
  OAI22_X1 U23978 ( .A1(n21059), .A2(n21013), .B1(n21012), .B2(n21011), .ZN(
        n21050) );
  AOI22_X1 U23979 ( .A1(n21065), .A2(n21051), .B1(n21064), .B2(n21050), .ZN(
        n21025) );
  INV_X1 U23980 ( .A(n21014), .ZN(n21017) );
  INV_X1 U23981 ( .A(n21059), .ZN(n21015) );
  AOI22_X1 U23982 ( .A1(n21018), .A2(n21017), .B1(n21016), .B2(n21015), .ZN(
        n21019) );
  NOR2_X1 U23983 ( .A1(n21019), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21022) );
  AOI22_X1 U23984 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21053), .B1(
        n21052), .B2(n21023), .ZN(n21024) );
  OAI211_X1 U23985 ( .C1(n21026), .C2(n21117), .A(n21025), .B(n21024), .ZN(
        P1_U3145) );
  AOI22_X1 U23986 ( .A1(n21079), .A2(n21051), .B1(n21078), .B2(n21050), .ZN(
        n21029) );
  AOI22_X1 U23987 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21053), .B1(
        n21052), .B2(n21027), .ZN(n21028) );
  OAI211_X1 U23988 ( .C1(n10000), .C2(n21117), .A(n21029), .B(n21028), .ZN(
        P1_U3146) );
  AOI22_X1 U23989 ( .A1(n21084), .A2(n21051), .B1(n21083), .B2(n21050), .ZN(
        n21033) );
  AOI22_X1 U23990 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21053), .B1(
        n21052), .B2(n21031), .ZN(n21032) );
  OAI211_X1 U23991 ( .C1(n10002), .C2(n21117), .A(n21033), .B(n21032), .ZN(
        P1_U3147) );
  AOI22_X1 U23992 ( .A1(n21089), .A2(n21051), .B1(n21088), .B2(n21050), .ZN(
        n21037) );
  AOI22_X1 U23993 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21053), .B1(
        n21052), .B2(n21035), .ZN(n21036) );
  OAI211_X1 U23994 ( .C1(n10004), .C2(n21117), .A(n21037), .B(n21036), .ZN(
        P1_U3148) );
  AOI22_X1 U23995 ( .A1(n21094), .A2(n21051), .B1(n21093), .B2(n21050), .ZN(
        n21040) );
  AOI22_X1 U23996 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21053), .B1(
        n21052), .B2(n9993), .ZN(n21039) );
  OAI211_X1 U23997 ( .C1(n21041), .C2(n21117), .A(n21040), .B(n21039), .ZN(
        P1_U3149) );
  AOI22_X1 U23998 ( .A1(n21099), .A2(n21051), .B1(n21098), .B2(n21050), .ZN(
        n21044) );
  AOI22_X1 U23999 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21053), .B1(
        n21052), .B2(n21042), .ZN(n21043) );
  OAI211_X1 U24000 ( .C1(n10006), .C2(n21117), .A(n21044), .B(n21043), .ZN(
        P1_U3150) );
  AOI22_X1 U24001 ( .A1(n21104), .A2(n21051), .B1(n21103), .B2(n21050), .ZN(
        n21048) );
  AOI22_X1 U24002 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21053), .B1(
        n21052), .B2(n21046), .ZN(n21047) );
  OAI211_X1 U24003 ( .C1(n9998), .C2(n21117), .A(n21048), .B(n21047), .ZN(
        P1_U3151) );
  AOI22_X1 U24004 ( .A1(n21111), .A2(n21051), .B1(n21109), .B2(n21050), .ZN(
        n21055) );
  AOI22_X1 U24005 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21053), .B1(
        n21052), .B2(n9995), .ZN(n21054) );
  OAI211_X1 U24006 ( .C1(n21056), .C2(n21117), .A(n21055), .B(n21054), .ZN(
        P1_U3152) );
  INV_X1 U24007 ( .A(n21060), .ZN(n21110) );
  INV_X1 U24008 ( .A(n21057), .ZN(n21058) );
  OR2_X1 U24009 ( .A1(n21059), .A2(n21058), .ZN(n21061) );
  NAND2_X1 U24010 ( .A1(n21061), .A2(n21060), .ZN(n21066) );
  NAND2_X1 U24011 ( .A1(n21066), .A2(n21206), .ZN(n21063) );
  NAND2_X1 U24012 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21072), .ZN(n21062) );
  NAND2_X1 U24013 ( .A1(n21063), .A2(n21062), .ZN(n21108) );
  AOI22_X1 U24014 ( .A1(n21065), .A2(n21110), .B1(n21064), .B2(n21108), .ZN(
        n21076) );
  INV_X1 U24015 ( .A(n21066), .ZN(n21067) );
  OAI21_X1 U24016 ( .B1(n21069), .B2(n21068), .A(n21067), .ZN(n21071) );
  OAI221_X1 U24017 ( .B1(n21206), .B2(n21072), .C1(n21194), .C2(n21071), .A(
        n21070), .ZN(n21114) );
  AOI22_X1 U24018 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n21074), .ZN(n21075) );
  OAI211_X1 U24019 ( .C1(n21077), .C2(n21117), .A(n21076), .B(n21075), .ZN(
        P1_U3153) );
  AOI22_X1 U24020 ( .A1(n21079), .A2(n21110), .B1(n21078), .B2(n21108), .ZN(
        n21081) );
  AOI22_X1 U24021 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n9999), .ZN(n21080) );
  OAI211_X1 U24022 ( .C1(n21082), .C2(n21117), .A(n21081), .B(n21080), .ZN(
        P1_U3154) );
  AOI22_X1 U24023 ( .A1(n21084), .A2(n21110), .B1(n21083), .B2(n21108), .ZN(
        n21086) );
  AOI22_X1 U24024 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n10001), .ZN(n21085) );
  OAI211_X1 U24025 ( .C1(n21087), .C2(n21117), .A(n21086), .B(n21085), .ZN(
        P1_U3155) );
  AOI22_X1 U24026 ( .A1(n21089), .A2(n21110), .B1(n21088), .B2(n21108), .ZN(
        n21091) );
  AOI22_X1 U24027 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n10003), .ZN(n21090) );
  OAI211_X1 U24028 ( .C1(n21092), .C2(n21117), .A(n21091), .B(n21090), .ZN(
        P1_U3156) );
  AOI22_X1 U24029 ( .A1(n21094), .A2(n21110), .B1(n21093), .B2(n21108), .ZN(
        n21096) );
  AOI22_X1 U24030 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n9990), .ZN(n21095) );
  OAI211_X1 U24031 ( .C1(n9994), .C2(n21117), .A(n21096), .B(n21095), .ZN(
        P1_U3157) );
  AOI22_X1 U24032 ( .A1(n21099), .A2(n21110), .B1(n21098), .B2(n21108), .ZN(
        n21101) );
  AOI22_X1 U24033 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n10005), .ZN(n21100) );
  OAI211_X1 U24034 ( .C1(n21102), .C2(n21117), .A(n21101), .B(n21100), .ZN(
        P1_U3158) );
  AOI22_X1 U24035 ( .A1(n21104), .A2(n21110), .B1(n21103), .B2(n21108), .ZN(
        n21106) );
  AOI22_X1 U24036 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n9997), .ZN(n21105) );
  OAI211_X1 U24037 ( .C1(n21107), .C2(n21117), .A(n21106), .B(n21105), .ZN(
        P1_U3159) );
  AOI22_X1 U24038 ( .A1(n21111), .A2(n21110), .B1(n21109), .B2(n21108), .ZN(
        n21116) );
  AOI22_X1 U24039 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n21112), .ZN(n21115) );
  OAI211_X1 U24040 ( .C1(n9996), .C2(n21117), .A(n21116), .B(n21115), .ZN(
        P1_U3160) );
  NAND3_X1 U24041 ( .A1(n21121), .A2(n21120), .A3(n21119), .ZN(P1_U3163) );
  AND2_X1 U24042 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21122), .ZN(
        P1_U3164) );
  AND2_X1 U24043 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21122), .ZN(
        P1_U3165) );
  AND2_X1 U24044 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21122), .ZN(
        P1_U3166) );
  INV_X1 U24045 ( .A(P1_DATAWIDTH_REG_28__SCAN_IN), .ZN(n21393) );
  NOR2_X1 U24046 ( .A1(n21186), .A2(n21393), .ZN(P1_U3167) );
  AND2_X1 U24047 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21122), .ZN(
        P1_U3168) );
  AND2_X1 U24048 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21122), .ZN(
        P1_U3169) );
  AND2_X1 U24049 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21122), .ZN(
        P1_U3170) );
  AND2_X1 U24050 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21122), .ZN(
        P1_U3171) );
  AND2_X1 U24051 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21122), .ZN(
        P1_U3172) );
  AND2_X1 U24052 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21122), .ZN(
        P1_U3173) );
  AND2_X1 U24053 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21122), .ZN(
        P1_U3174) );
  AND2_X1 U24054 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21122), .ZN(
        P1_U3175) );
  AND2_X1 U24055 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21122), .ZN(
        P1_U3176) );
  AND2_X1 U24056 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21122), .ZN(
        P1_U3177) );
  AND2_X1 U24057 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21122), .ZN(
        P1_U3178) );
  AND2_X1 U24058 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21122), .ZN(
        P1_U3179) );
  AND2_X1 U24059 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21122), .ZN(
        P1_U3180) );
  AND2_X1 U24060 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21122), .ZN(
        P1_U3181) );
  AND2_X1 U24061 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21122), .ZN(
        P1_U3182) );
  AND2_X1 U24062 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21122), .ZN(
        P1_U3183) );
  INV_X1 U24063 ( .A(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n21532) );
  NOR2_X1 U24064 ( .A1(n21186), .A2(n21532), .ZN(P1_U3184) );
  AND2_X1 U24065 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21122), .ZN(
        P1_U3185) );
  AND2_X1 U24066 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21122), .ZN(P1_U3186) );
  AND2_X1 U24067 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21122), .ZN(P1_U3187) );
  AND2_X1 U24068 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21122), .ZN(P1_U3188) );
  AND2_X1 U24069 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21122), .ZN(P1_U3189) );
  AND2_X1 U24070 ( .A1(n21122), .A2(P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(P1_U3190) );
  AND2_X1 U24071 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21122), .ZN(P1_U3191) );
  AND2_X1 U24072 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21122), .ZN(P1_U3192) );
  AND2_X1 U24073 ( .A1(n21122), .A2(P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(P1_U3193) );
  AOI21_X1 U24074 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21132), .A(n21136), 
        .ZN(n21127) );
  OAI21_X1 U24075 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21130), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21123) );
  AOI211_X1 U24076 ( .C1(HOLD), .C2(P1_STATE_REG_2__SCAN_IN), .A(n21124), .B(
        n21123), .ZN(n21125) );
  OAI22_X1 U24077 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21127), .B1(n21223), 
        .B2(n21125), .ZN(P1_U3194) );
  OAI211_X1 U24078 ( .C1(NA), .C2(n21224), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n21137), .ZN(n21126) );
  OAI211_X1 U24079 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21452), .A(HOLD), .B(
        n21126), .ZN(n21135) );
  AOI211_X1 U24080 ( .C1(n21128), .C2(NA), .A(n21137), .B(n21127), .ZN(n21129)
         );
  INV_X1 U24081 ( .A(n21129), .ZN(n21134) );
  NAND4_X1 U24082 ( .A1(n21132), .A2(P1_STATE_REG_1__SCAN_IN), .A3(n21131), 
        .A4(n21130), .ZN(n21133) );
  OAI211_X1 U24083 ( .C1(n21136), .C2(n21135), .A(n21134), .B(n21133), .ZN(
        P1_U3196) );
  NOR2_X1 U24084 ( .A1(n21239), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21175) );
  OR2_X1 U24085 ( .A1(n21137), .A2(n21239), .ZN(n21166) );
  AOI222_X1 U24086 ( .A1(n21175), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n9827), .ZN(n21138) );
  INV_X1 U24087 ( .A(n21138), .ZN(P1_U3197) );
  INV_X1 U24088 ( .A(n21175), .ZN(n21168) );
  INV_X1 U24089 ( .A(n21168), .ZN(n21177) );
  AOI222_X1 U24090 ( .A1(n9827), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21239), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21177), .ZN(n21139) );
  INV_X1 U24091 ( .A(n21139), .ZN(P1_U3198) );
  OAI222_X1 U24092 ( .A1(n21166), .A2(n21142), .B1(n21141), .B2(n21223), .C1(
        n21140), .C2(n21168), .ZN(P1_U3199) );
  AOI222_X1 U24093 ( .A1(n21175), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n21239), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n9827), .ZN(n21143) );
  INV_X1 U24094 ( .A(n21143), .ZN(P1_U3200) );
  AOI222_X1 U24095 ( .A1(n9827), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n21239), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n21177), .ZN(n21144) );
  INV_X1 U24096 ( .A(n21144), .ZN(P1_U3201) );
  AOI222_X1 U24097 ( .A1(n9827), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n21177), .ZN(n21145) );
  INV_X1 U24098 ( .A(n21145), .ZN(P1_U3202) );
  AOI222_X1 U24099 ( .A1(n9827), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21177), .ZN(n21146) );
  INV_X1 U24100 ( .A(n21146), .ZN(P1_U3203) );
  AOI222_X1 U24101 ( .A1(n21175), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n9827), .ZN(n21147) );
  INV_X1 U24102 ( .A(n21147), .ZN(P1_U3204) );
  AOI222_X1 U24103 ( .A1(n9827), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21177), .ZN(n21148) );
  INV_X1 U24104 ( .A(n21148), .ZN(P1_U3205) );
  AOI22_X1 U24105 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n21239), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n21177), .ZN(n21149) );
  OAI21_X1 U24106 ( .B1(n21150), .B2(n21166), .A(n21149), .ZN(P1_U3206) );
  AOI22_X1 U24107 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21239), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n9827), .ZN(n21151) );
  OAI21_X1 U24108 ( .B1(n21152), .B2(n21168), .A(n21151), .ZN(P1_U3207) );
  AOI222_X1 U24109 ( .A1(n21175), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n9827), .ZN(n21153) );
  INV_X1 U24110 ( .A(n21153), .ZN(P1_U3208) );
  AOI222_X1 U24111 ( .A1(n9827), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21177), .ZN(n21154) );
  INV_X1 U24112 ( .A(n21154), .ZN(P1_U3209) );
  AOI222_X1 U24113 ( .A1(n21175), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n9827), .ZN(n21155) );
  INV_X1 U24114 ( .A(n21155), .ZN(P1_U3210) );
  AOI222_X1 U24115 ( .A1(n9827), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n21177), .ZN(n21156) );
  INV_X1 U24116 ( .A(n21156), .ZN(P1_U3211) );
  AOI22_X1 U24117 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21239), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21175), .ZN(n21157) );
  OAI21_X1 U24118 ( .B1(n21158), .B2(n21166), .A(n21157), .ZN(P1_U3212) );
  AOI22_X1 U24119 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21239), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n9827), .ZN(n21159) );
  OAI21_X1 U24120 ( .B1(n21160), .B2(n21168), .A(n21159), .ZN(P1_U3213) );
  AOI222_X1 U24121 ( .A1(n9827), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n21177), .ZN(n21161) );
  INV_X1 U24122 ( .A(n21161), .ZN(P1_U3214) );
  AOI222_X1 U24123 ( .A1(n9827), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n21177), .ZN(n21162) );
  INV_X1 U24124 ( .A(n21162), .ZN(P1_U3215) );
  AOI222_X1 U24125 ( .A1(n9827), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21177), .ZN(n21163) );
  INV_X1 U24126 ( .A(n21163), .ZN(P1_U3216) );
  AOI222_X1 U24127 ( .A1(n21175), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n9827), .ZN(n21164) );
  INV_X1 U24128 ( .A(n21164), .ZN(P1_U3217) );
  AOI22_X1 U24129 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21239), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21177), .ZN(n21165) );
  OAI21_X1 U24130 ( .B1(n14934), .B2(n21166), .A(n21165), .ZN(P1_U3218) );
  AOI22_X1 U24131 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21239), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n9827), .ZN(n21167) );
  OAI21_X1 U24132 ( .B1(n21169), .B2(n21168), .A(n21167), .ZN(P1_U3219) );
  AOI222_X1 U24133 ( .A1(n9827), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21177), .ZN(n21170) );
  INV_X1 U24134 ( .A(n21170), .ZN(P1_U3220) );
  AOI222_X1 U24135 ( .A1(n21175), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n9827), .ZN(n21171) );
  INV_X1 U24136 ( .A(n21171), .ZN(P1_U3221) );
  AOI222_X1 U24137 ( .A1(n9827), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21177), .ZN(n21172) );
  INV_X1 U24138 ( .A(n21172), .ZN(P1_U3222) );
  AOI222_X1 U24139 ( .A1(n9827), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n21177), .ZN(n21173) );
  INV_X1 U24140 ( .A(n21173), .ZN(P1_U3223) );
  AOI222_X1 U24141 ( .A1(n9827), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21175), .ZN(n21174) );
  INV_X1 U24142 ( .A(n21174), .ZN(P1_U3224) );
  AOI222_X1 U24143 ( .A1(n21175), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n9827), .ZN(n21176) );
  INV_X1 U24144 ( .A(n21176), .ZN(P1_U3225) );
  AOI222_X1 U24145 ( .A1(n9827), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21222), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21177), .ZN(n21178) );
  INV_X1 U24146 ( .A(n21178), .ZN(P1_U3226) );
  OAI22_X1 U24147 ( .A1(n21239), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21223), .ZN(n21179) );
  INV_X1 U24148 ( .A(n21179), .ZN(P1_U3458) );
  OAI22_X1 U24149 ( .A1(n21239), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21223), .ZN(n21180) );
  INV_X1 U24150 ( .A(n21180), .ZN(P1_U3459) );
  OAI22_X1 U24151 ( .A1(n21239), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21223), .ZN(n21181) );
  INV_X1 U24152 ( .A(n21181), .ZN(P1_U3460) );
  OAI22_X1 U24153 ( .A1(n21239), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21223), .ZN(n21182) );
  INV_X1 U24154 ( .A(n21182), .ZN(P1_U3461) );
  OAI21_X1 U24155 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21186), .A(n21184), 
        .ZN(n21183) );
  INV_X1 U24156 ( .A(n21183), .ZN(P1_U3464) );
  OAI21_X1 U24157 ( .B1(n21186), .B2(n21185), .A(n21184), .ZN(P1_U3465) );
  AOI22_X1 U24158 ( .A1(n21190), .A2(n21189), .B1(n21188), .B2(n21187), .ZN(
        n21191) );
  INV_X1 U24159 ( .A(n21191), .ZN(n21193) );
  MUX2_X1 U24160 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21193), .S(
        n21192), .Z(P1_U3469) );
  INV_X1 U24161 ( .A(n21212), .ZN(n21215) );
  AOI21_X1 U24162 ( .B1(n21196), .B2(n21195), .A(n21194), .ZN(n21203) );
  INV_X1 U24163 ( .A(n14039), .ZN(n21198) );
  OAI22_X1 U24164 ( .A1(n21200), .A2(n21199), .B1(n21198), .B2(n21197), .ZN(
        n21201) );
  NOR3_X1 U24165 ( .A1(n21203), .A2(n21202), .A3(n21201), .ZN(n21204) );
  AOI22_X1 U24166 ( .A1(n21215), .A2(n21205), .B1(n21204), .B2(n21212), .ZN(
        P1_U3475) );
  AOI22_X1 U24167 ( .A1(n21209), .A2(n21208), .B1(n21207), .B2(n21206), .ZN(
        n21210) );
  AND2_X1 U24168 ( .A1(n21211), .A2(n21210), .ZN(n21213) );
  AOI22_X1 U24169 ( .A1(n21215), .A2(n21214), .B1(n21213), .B2(n21212), .ZN(
        P1_U3478) );
  AOI211_X1 U24170 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21216) );
  AOI21_X1 U24171 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21216), .ZN(n21218) );
  INV_X1 U24172 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21217) );
  AOI22_X1 U24173 ( .A1(n21221), .A2(n21218), .B1(n21217), .B2(n21219), .ZN(
        P1_U3481) );
  NOR2_X1 U24174 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21220) );
  INV_X1 U24175 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21349) );
  AOI22_X1 U24176 ( .A1(n21221), .A2(n21220), .B1(n21349), .B2(n21219), .ZN(
        P1_U3482) );
  AOI22_X1 U24177 ( .A1(n21223), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21525), 
        .B2(n21222), .ZN(P1_U3483) );
  NAND2_X1 U24178 ( .A1(n21224), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21233) );
  INV_X1 U24179 ( .A(n21233), .ZN(n21227) );
  AOI211_X1 U24180 ( .C1(n21228), .C2(n21227), .A(n21226), .B(n21225), .ZN(
        n21238) );
  INV_X1 U24181 ( .A(n21229), .ZN(n21232) );
  AOI22_X1 U24182 ( .A1(n21232), .A2(n21231), .B1(P1_STATEBS16_REG_SCAN_IN), 
        .B2(n21230), .ZN(n21234) );
  OAI21_X1 U24183 ( .B1(n21234), .B2(n21233), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n21237) );
  NOR2_X1 U24184 ( .A1(n21238), .A2(n21235), .ZN(n21236) );
  AOI22_X1 U24185 ( .A1(n21452), .A2(n21238), .B1(n21237), .B2(n21236), .ZN(
        P1_U3485) );
  MUX2_X1 U24186 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21239), .Z(P1_U3486) );
  NAND2_X1 U24187 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n21240), .ZN(n21629) );
  AOI22_X1 U24188 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(keyinput182), 
        .B1(P2_EBX_REG_11__SCAN_IN), .B2(keyinput214), .ZN(n21241) );
  OAI221_X1 U24189 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput182), 
        .C1(P2_EBX_REG_11__SCAN_IN), .C2(keyinput214), .A(n21241), .ZN(n21248)
         );
  AOI22_X1 U24190 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput211), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput235), .ZN(n21242) );
  OAI221_X1 U24191 ( .B1(P2_DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput211), .C1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(keyinput235), .A(n21242), .ZN(
        n21247) );
  AOI22_X1 U24192 ( .A1(P1_EAX_REG_19__SCAN_IN), .A2(keyinput190), .B1(
        P2_INSTQUEUE_REG_3__0__SCAN_IN), .B2(keyinput192), .ZN(n21243) );
  OAI221_X1 U24193 ( .B1(P1_EAX_REG_19__SCAN_IN), .B2(keyinput190), .C1(
        P2_INSTQUEUE_REG_3__0__SCAN_IN), .C2(keyinput192), .A(n21243), .ZN(
        n21246) );
  AOI22_X1 U24194 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(keyinput231), .B1(
        P3_EAX_REG_25__SCAN_IN), .B2(keyinput147), .ZN(n21244) );
  OAI221_X1 U24195 ( .B1(P1_DATAWIDTH_REG_2__SCAN_IN), .B2(keyinput231), .C1(
        P3_EAX_REG_25__SCAN_IN), .C2(keyinput147), .A(n21244), .ZN(n21245) );
  NOR4_X1 U24196 ( .A1(n21248), .A2(n21247), .A3(n21246), .A4(n21245), .ZN(
        n21276) );
  AOI22_X1 U24197 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(keyinput241), 
        .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput152), .ZN(n21249) );
  OAI221_X1 U24198 ( .B1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput241), 
        .C1(P1_REIP_REG_19__SCAN_IN), .C2(keyinput152), .A(n21249), .ZN(n21256) );
  AOI22_X1 U24199 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(keyinput198), .B1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .B2(keyinput178), .ZN(n21250) );
  OAI221_X1 U24200 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(keyinput198), .C1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .C2(keyinput178), .A(n21250), .ZN(
        n21255) );
  AOI22_X1 U24201 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(keyinput141), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(keyinput228), .ZN(n21251) );
  OAI221_X1 U24202 ( .B1(P1_DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput141), .C1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .C2(keyinput228), .A(n21251), .ZN(
        n21254) );
  AOI22_X1 U24203 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(keyinput157), 
        .B1(P2_ADDRESS_REG_7__SCAN_IN), .B2(keyinput253), .ZN(n21252) );
  OAI221_X1 U24204 ( .B1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B2(keyinput157), 
        .C1(P2_ADDRESS_REG_7__SCAN_IN), .C2(keyinput253), .A(n21252), .ZN(
        n21253) );
  NOR4_X1 U24205 ( .A1(n21256), .A2(n21255), .A3(n21254), .A4(n21253), .ZN(
        n21275) );
  AOI22_X1 U24206 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(keyinput246), .B1(
        P2_ADDRESS_REG_24__SCAN_IN), .B2(keyinput140), .ZN(n21257) );
  OAI221_X1 U24207 ( .B1(P3_REIP_REG_2__SCAN_IN), .B2(keyinput246), .C1(
        P2_ADDRESS_REG_24__SCAN_IN), .C2(keyinput140), .A(n21257), .ZN(n21264)
         );
  AOI22_X1 U24208 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput195), 
        .B1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput191), .ZN(n21258) );
  OAI221_X1 U24209 ( .B1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput195), 
        .C1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .C2(keyinput191), .A(n21258), 
        .ZN(n21263) );
  AOI22_X1 U24210 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(keyinput167), .B1(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput200), .ZN(n21259) );
  OAI221_X1 U24211 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(keyinput167), .C1(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput200), .A(n21259), 
        .ZN(n21262) );
  AOI22_X1 U24212 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(keyinput217), .B1(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput221), .ZN(n21260) );
  OAI221_X1 U24213 ( .B1(P3_EAX_REG_27__SCAN_IN), .B2(keyinput217), .C1(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput221), .A(n21260), .ZN(
        n21261) );
  NOR4_X1 U24214 ( .A1(n21264), .A2(n21263), .A3(n21262), .A4(n21261), .ZN(
        n21274) );
  AOI22_X1 U24215 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(keyinput139), .B1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(keyinput164), .ZN(n21265) );
  OAI221_X1 U24216 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(keyinput139), .C1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .C2(keyinput164), .A(n21265), .ZN(
        n21272) );
  AOI22_X1 U24217 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(keyinput232), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(keyinput222), .ZN(n21266) );
  OAI221_X1 U24218 ( .B1(P2_UWORD_REG_3__SCAN_IN), .B2(keyinput232), .C1(
        P1_REIP_REG_6__SCAN_IN), .C2(keyinput222), .A(n21266), .ZN(n21271) );
  AOI22_X1 U24219 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(keyinput150), .B1(
        BUF1_REG_9__SCAN_IN), .B2(keyinput128), .ZN(n21267) );
  OAI221_X1 U24220 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(keyinput150), .C1(
        BUF1_REG_9__SCAN_IN), .C2(keyinput128), .A(n21267), .ZN(n21270) );
  AOI22_X1 U24221 ( .A1(BUF2_REG_26__SCAN_IN), .A2(keyinput158), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(keyinput181), .ZN(n21268) );
  OAI221_X1 U24222 ( .B1(BUF2_REG_26__SCAN_IN), .B2(keyinput158), .C1(
        P2_ADDRESS_REG_5__SCAN_IN), .C2(keyinput181), .A(n21268), .ZN(n21269)
         );
  NOR4_X1 U24223 ( .A1(n21272), .A2(n21271), .A3(n21270), .A4(n21269), .ZN(
        n21273) );
  NAND4_X1 U24224 ( .A1(n21276), .A2(n21275), .A3(n21274), .A4(n21273), .ZN(
        n21422) );
  AOI22_X1 U24225 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput215), .B1(
        P3_REIP_REG_26__SCAN_IN), .B2(keyinput148), .ZN(n21277) );
  OAI221_X1 U24226 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput215), 
        .C1(P3_REIP_REG_26__SCAN_IN), .C2(keyinput148), .A(n21277), .ZN(n21284) );
  AOI22_X1 U24227 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(keyinput193), .B1(
        BUF2_REG_14__SCAN_IN), .B2(keyinput247), .ZN(n21278) );
  OAI221_X1 U24228 ( .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput193), .C1(
        BUF2_REG_14__SCAN_IN), .C2(keyinput247), .A(n21278), .ZN(n21283) );
  AOI22_X1 U24229 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput239), 
        .B1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B2(keyinput144), .ZN(n21279) );
  OAI221_X1 U24230 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput239), 
        .C1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .C2(keyinput144), .A(n21279), 
        .ZN(n21282) );
  AOI22_X1 U24231 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput146), .B1(
        P2_LWORD_REG_8__SCAN_IN), .B2(keyinput197), .ZN(n21280) );
  OAI221_X1 U24232 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput146), .C1(
        P2_LWORD_REG_8__SCAN_IN), .C2(keyinput197), .A(n21280), .ZN(n21281) );
  NOR4_X1 U24233 ( .A1(n21284), .A2(n21283), .A3(n21282), .A4(n21281), .ZN(
        n21315) );
  AOI22_X1 U24234 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(keyinput131), .B1(
        DATAI_24_), .B2(keyinput219), .ZN(n21285) );
  OAI221_X1 U24235 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(keyinput131), .C1(
        DATAI_24_), .C2(keyinput219), .A(n21285), .ZN(n21292) );
  AOI22_X1 U24236 ( .A1(BUF1_REG_15__SCAN_IN), .A2(keyinput252), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(keyinput161), .ZN(n21286) );
  OAI221_X1 U24237 ( .B1(BUF1_REG_15__SCAN_IN), .B2(keyinput252), .C1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .C2(keyinput161), .A(n21286), .ZN(
        n21291) );
  AOI22_X1 U24238 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(keyinput173), .B1(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput205), .ZN(n21287) );
  OAI221_X1 U24239 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(keyinput173), .C1(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(keyinput205), .A(n21287), 
        .ZN(n21290) );
  AOI22_X1 U24240 ( .A1(DATAI_4_), .A2(keyinput236), .B1(
        P1_INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput213), .ZN(n21288) );
  OAI221_X1 U24241 ( .B1(DATAI_4_), .B2(keyinput236), .C1(
        P1_INSTQUEUE_REG_14__1__SCAN_IN), .C2(keyinput213), .A(n21288), .ZN(
        n21289) );
  NOR4_X1 U24242 ( .A1(n21292), .A2(n21291), .A3(n21290), .A4(n21289), .ZN(
        n21314) );
  AOI22_X1 U24243 ( .A1(BS16), .A2(keyinput172), .B1(
        P3_INSTQUEUE_REG_9__2__SCAN_IN), .B2(keyinput156), .ZN(n21293) );
  OAI221_X1 U24244 ( .B1(BS16), .B2(keyinput172), .C1(
        P3_INSTQUEUE_REG_9__2__SCAN_IN), .C2(keyinput156), .A(n21293), .ZN(
        n21300) );
  AOI22_X1 U24245 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(keyinput143), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput166), .ZN(n21294) );
  OAI221_X1 U24246 ( .B1(P1_DATAO_REG_18__SCAN_IN), .B2(keyinput143), .C1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(keyinput166), .A(n21294), .ZN(
        n21299) );
  AOI22_X1 U24247 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(keyinput227), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(keyinput153), .ZN(n21295) );
  OAI221_X1 U24248 ( .B1(P1_DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput227), .C1(
        P3_EAX_REG_4__SCAN_IN), .C2(keyinput153), .A(n21295), .ZN(n21298) );
  AOI22_X1 U24249 ( .A1(P3_ADDRESS_REG_8__SCAN_IN), .A2(keyinput234), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(keyinput206), .ZN(n21296) );
  OAI221_X1 U24250 ( .B1(P3_ADDRESS_REG_8__SCAN_IN), .B2(keyinput234), .C1(
        P1_LWORD_REG_6__SCAN_IN), .C2(keyinput206), .A(n21296), .ZN(n21297) );
  NOR4_X1 U24251 ( .A1(n21300), .A2(n21299), .A3(n21298), .A4(n21297), .ZN(
        n21313) );
  AOI22_X1 U24252 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(keyinput202), .B1(
        P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput225), .ZN(n21301) );
  OAI221_X1 U24253 ( .B1(P1_DATAO_REG_5__SCAN_IN), .B2(keyinput202), .C1(
        P2_INSTQUEUE_REG_14__1__SCAN_IN), .C2(keyinput225), .A(n21301), .ZN(
        n21311) );
  AOI22_X1 U24254 ( .A1(P3_DATAO_REG_16__SCAN_IN), .A2(keyinput249), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(keyinput244), .ZN(n21302) );
  OAI221_X1 U24255 ( .B1(P3_DATAO_REG_16__SCAN_IN), .B2(keyinput249), .C1(
        P2_EAX_REG_13__SCAN_IN), .C2(keyinput244), .A(n21302), .ZN(n21310) );
  INV_X1 U24256 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n21304) );
  AOI22_X1 U24257 ( .A1(n21305), .A2(keyinput208), .B1(keyinput180), .B2(
        n21304), .ZN(n21303) );
  OAI221_X1 U24258 ( .B1(n21305), .B2(keyinput208), .C1(n21304), .C2(
        keyinput180), .A(n21303), .ZN(n21309) );
  INV_X1 U24259 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n21307) );
  AOI22_X1 U24260 ( .A1(n21307), .A2(keyinput207), .B1(keyinput210), .B2(
        n21541), .ZN(n21306) );
  OAI221_X1 U24261 ( .B1(n21307), .B2(keyinput207), .C1(n21541), .C2(
        keyinput210), .A(n21306), .ZN(n21308) );
  NOR4_X1 U24262 ( .A1(n21311), .A2(n21310), .A3(n21309), .A4(n21308), .ZN(
        n21312) );
  NAND4_X1 U24263 ( .A1(n21315), .A2(n21314), .A3(n21313), .A4(n21312), .ZN(
        n21421) );
  AOI22_X1 U24264 ( .A1(n21318), .A2(keyinput250), .B1(n21317), .B2(
        keyinput155), .ZN(n21316) );
  OAI221_X1 U24265 ( .B1(n21318), .B2(keyinput250), .C1(n21317), .C2(
        keyinput155), .A(n21316), .ZN(n21326) );
  INV_X1 U24266 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n21320) );
  AOI22_X1 U24267 ( .A1(n21499), .A2(keyinput130), .B1(keyinput169), .B2(
        n21320), .ZN(n21319) );
  OAI221_X1 U24268 ( .B1(n21499), .B2(keyinput130), .C1(n21320), .C2(
        keyinput169), .A(n21319), .ZN(n21325) );
  AOI22_X1 U24269 ( .A1(n21522), .A2(keyinput176), .B1(n13555), .B2(
        keyinput238), .ZN(n21321) );
  OAI221_X1 U24270 ( .B1(n21522), .B2(keyinput176), .C1(n13555), .C2(
        keyinput238), .A(n21321), .ZN(n21324) );
  AOI22_X1 U24271 ( .A1(n21430), .A2(keyinput204), .B1(n21517), .B2(
        keyinput179), .ZN(n21322) );
  OAI221_X1 U24272 ( .B1(n21430), .B2(keyinput204), .C1(n21517), .C2(
        keyinput179), .A(n21322), .ZN(n21323) );
  NOR4_X1 U24273 ( .A1(n21326), .A2(n21325), .A3(n21324), .A4(n21323), .ZN(
        n21364) );
  INV_X1 U24274 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n21459) );
  INV_X1 U24275 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n21442) );
  AOI22_X1 U24276 ( .A1(n21459), .A2(keyinput203), .B1(keyinput175), .B2(
        n21442), .ZN(n21327) );
  OAI221_X1 U24277 ( .B1(n21459), .B2(keyinput203), .C1(n21442), .C2(
        keyinput175), .A(n21327), .ZN(n21335) );
  AOI22_X1 U24278 ( .A1(n21456), .A2(keyinput189), .B1(keyinput135), .B2(
        n21502), .ZN(n21328) );
  OAI221_X1 U24279 ( .B1(n21456), .B2(keyinput189), .C1(n21502), .C2(
        keyinput135), .A(n21328), .ZN(n21334) );
  INV_X1 U24280 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n21535) );
  AOI22_X1 U24281 ( .A1(n21535), .A2(keyinput138), .B1(keyinput230), .B2(
        n21330), .ZN(n21329) );
  OAI221_X1 U24282 ( .B1(n21535), .B2(keyinput138), .C1(n21330), .C2(
        keyinput230), .A(n21329), .ZN(n21333) );
  AOI22_X1 U24283 ( .A1(n12009), .A2(keyinput174), .B1(keyinput209), .B2(
        n21509), .ZN(n21331) );
  OAI221_X1 U24284 ( .B1(n12009), .B2(keyinput174), .C1(n21509), .C2(
        keyinput209), .A(n21331), .ZN(n21332) );
  NOR4_X1 U24285 ( .A1(n21335), .A2(n21334), .A3(n21333), .A4(n21332), .ZN(
        n21363) );
  INV_X1 U24286 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n21337) );
  AOI22_X1 U24287 ( .A1(n21337), .A2(keyinput129), .B1(keyinput145), .B2(
        n21437), .ZN(n21336) );
  OAI221_X1 U24288 ( .B1(n21337), .B2(keyinput129), .C1(n21437), .C2(
        keyinput145), .A(n21336), .ZN(n21347) );
  AOI22_X1 U24289 ( .A1(n21339), .A2(keyinput199), .B1(n21466), .B2(
        keyinput218), .ZN(n21338) );
  OAI221_X1 U24290 ( .B1(n21339), .B2(keyinput199), .C1(n21466), .C2(
        keyinput218), .A(n21338), .ZN(n21346) );
  AOI22_X1 U24291 ( .A1(n21341), .A2(keyinput233), .B1(n21429), .B2(
        keyinput224), .ZN(n21340) );
  OAI221_X1 U24292 ( .B1(n21341), .B2(keyinput233), .C1(n21429), .C2(
        keyinput224), .A(n21340), .ZN(n21345) );
  INV_X1 U24293 ( .A(P3_LWORD_REG_10__SCAN_IN), .ZN(n21343) );
  AOI22_X1 U24294 ( .A1(n21469), .A2(keyinput187), .B1(keyinput201), .B2(
        n21343), .ZN(n21342) );
  OAI221_X1 U24295 ( .B1(n21469), .B2(keyinput187), .C1(n21343), .C2(
        keyinput201), .A(n21342), .ZN(n21344) );
  NOR4_X1 U24296 ( .A1(n21347), .A2(n21346), .A3(n21345), .A4(n21344), .ZN(
        n21362) );
  AOI22_X1 U24297 ( .A1(n21349), .A2(keyinput186), .B1(n13315), .B2(
        keyinput248), .ZN(n21348) );
  OAI221_X1 U24298 ( .B1(n21349), .B2(keyinput186), .C1(n13315), .C2(
        keyinput248), .A(n21348), .ZN(n21360) );
  INV_X1 U24299 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n21352) );
  INV_X1 U24300 ( .A(P3_UWORD_REG_12__SCAN_IN), .ZN(n21351) );
  AOI22_X1 U24301 ( .A1(n21352), .A2(keyinput242), .B1(n21351), .B2(
        keyinput160), .ZN(n21350) );
  OAI221_X1 U24302 ( .B1(n21352), .B2(keyinput242), .C1(n21351), .C2(
        keyinput160), .A(n21350), .ZN(n21359) );
  XNOR2_X1 U24303 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput251), .ZN(
        n21355) );
  XNOR2_X1 U24304 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B(keyinput255), .ZN(
        n21354) );
  XNOR2_X1 U24305 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(keyinput240), 
        .ZN(n21353) );
  NAND3_X1 U24306 ( .A1(n21355), .A2(n21354), .A3(n21353), .ZN(n21358) );
  XNOR2_X1 U24307 ( .A(n21356), .B(keyinput226), .ZN(n21357) );
  NOR4_X1 U24308 ( .A1(n21360), .A2(n21359), .A3(n21358), .A4(n21357), .ZN(
        n21361) );
  NAND4_X1 U24309 ( .A1(n21364), .A2(n21363), .A3(n21362), .A4(n21361), .ZN(
        n21420) );
  AOI22_X1 U24310 ( .A1(n21367), .A2(keyinput188), .B1(n21366), .B2(
        keyinput132), .ZN(n21365) );
  OAI221_X1 U24311 ( .B1(n21367), .B2(keyinput188), .C1(n21366), .C2(
        keyinput132), .A(n21365), .ZN(n21376) );
  INV_X1 U24312 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n21369) );
  AOI22_X1 U24313 ( .A1(n21369), .A2(keyinput136), .B1(n21526), .B2(
        keyinput149), .ZN(n21368) );
  OAI221_X1 U24314 ( .B1(n21369), .B2(keyinput136), .C1(n21526), .C2(
        keyinput149), .A(n21368), .ZN(n21375) );
  INV_X1 U24315 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n21371) );
  INV_X1 U24316 ( .A(READY1), .ZN(n21506) );
  AOI22_X1 U24317 ( .A1(n21371), .A2(keyinput177), .B1(keyinput142), .B2(
        n21506), .ZN(n21370) );
  OAI221_X1 U24318 ( .B1(n21371), .B2(keyinput177), .C1(n21506), .C2(
        keyinput142), .A(n21370), .ZN(n21374) );
  AOI22_X1 U24319 ( .A1(n13596), .A2(keyinput168), .B1(keyinput216), .B2(
        n21444), .ZN(n21372) );
  OAI221_X1 U24320 ( .B1(n13596), .B2(keyinput168), .C1(n21444), .C2(
        keyinput216), .A(n21372), .ZN(n21373) );
  NOR4_X1 U24321 ( .A1(n21376), .A2(n21375), .A3(n21374), .A4(n21373), .ZN(
        n21418) );
  AOI22_X1 U24322 ( .A1(n21378), .A2(keyinput237), .B1(keyinput137), .B2(
        n21473), .ZN(n21377) );
  OAI221_X1 U24323 ( .B1(n21378), .B2(keyinput237), .C1(n21473), .C2(
        keyinput137), .A(n21377), .ZN(n21388) );
  INV_X1 U24324 ( .A(DATAI_31_), .ZN(n21380) );
  AOI22_X1 U24325 ( .A1(n21505), .A2(keyinput243), .B1(n21380), .B2(
        keyinput245), .ZN(n21379) );
  OAI221_X1 U24326 ( .B1(n21505), .B2(keyinput243), .C1(n21380), .C2(
        keyinput245), .A(n21379), .ZN(n21387) );
  AOI22_X1 U24327 ( .A1(n21382), .A2(keyinput162), .B1(n21537), .B2(
        keyinput212), .ZN(n21381) );
  OAI221_X1 U24328 ( .B1(n21382), .B2(keyinput162), .C1(n21537), .C2(
        keyinput212), .A(n21381), .ZN(n21386) );
  INV_X1 U24329 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n21538) );
  XOR2_X1 U24330 ( .A(n21538), .B(keyinput133), .Z(n21384) );
  XNOR2_X1 U24331 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B(keyinput163), .ZN(
        n21383) );
  NAND2_X1 U24332 ( .A1(n21384), .A2(n21383), .ZN(n21385) );
  NOR4_X1 U24333 ( .A1(n21388), .A2(n21387), .A3(n21386), .A4(n21385), .ZN(
        n21417) );
  INV_X1 U24334 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21391) );
  AOI22_X1 U24335 ( .A1(n21391), .A2(keyinput196), .B1(keyinput170), .B2(
        n21390), .ZN(n21389) );
  OAI221_X1 U24336 ( .B1(n21391), .B2(keyinput196), .C1(n21390), .C2(
        keyinput170), .A(n21389), .ZN(n21402) );
  AOI22_X1 U24337 ( .A1(n13180), .A2(keyinput254), .B1(keyinput183), .B2(
        n21393), .ZN(n21392) );
  OAI221_X1 U24338 ( .B1(n13180), .B2(keyinput254), .C1(n21393), .C2(
        keyinput183), .A(n21392), .ZN(n21401) );
  AOI22_X1 U24339 ( .A1(n21395), .A2(keyinput159), .B1(n12382), .B2(
        keyinput223), .ZN(n21394) );
  OAI221_X1 U24340 ( .B1(n21395), .B2(keyinput159), .C1(n12382), .C2(
        keyinput223), .A(n21394), .ZN(n21400) );
  AOI22_X1 U24341 ( .A1(n21398), .A2(keyinput184), .B1(n21397), .B2(
        keyinput165), .ZN(n21396) );
  OAI221_X1 U24342 ( .B1(n21398), .B2(keyinput184), .C1(n21397), .C2(
        keyinput165), .A(n21396), .ZN(n21399) );
  NOR4_X1 U24343 ( .A1(n21402), .A2(n21401), .A3(n21400), .A4(n21399), .ZN(
        n21416) );
  AOI22_X1 U24344 ( .A1(n21404), .A2(keyinput171), .B1(n11869), .B2(
        keyinput185), .ZN(n21403) );
  OAI221_X1 U24345 ( .B1(n21404), .B2(keyinput171), .C1(n11869), .C2(
        keyinput185), .A(n21403), .ZN(n21414) );
  INV_X1 U24346 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n21407) );
  INV_X1 U24347 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n21406) );
  AOI22_X1 U24348 ( .A1(n21407), .A2(keyinput220), .B1(n21406), .B2(
        keyinput229), .ZN(n21405) );
  OAI221_X1 U24349 ( .B1(n21407), .B2(keyinput220), .C1(n21406), .C2(
        keyinput229), .A(n21405), .ZN(n21413) );
  AOI22_X1 U24350 ( .A1(n21443), .A2(keyinput134), .B1(n21409), .B2(
        keyinput154), .ZN(n21408) );
  OAI221_X1 U24351 ( .B1(n21443), .B2(keyinput134), .C1(n21409), .C2(
        keyinput154), .A(n21408), .ZN(n21412) );
  AOI22_X1 U24352 ( .A1(n21488), .A2(keyinput151), .B1(keyinput194), .B2(
        n21485), .ZN(n21410) );
  OAI221_X1 U24353 ( .B1(n21488), .B2(keyinput151), .C1(n21485), .C2(
        keyinput194), .A(n21410), .ZN(n21411) );
  NOR4_X1 U24354 ( .A1(n21414), .A2(n21413), .A3(n21412), .A4(n21411), .ZN(
        n21415) );
  NAND4_X1 U24355 ( .A1(n21418), .A2(n21417), .A3(n21416), .A4(n21415), .ZN(
        n21419) );
  NOR4_X1 U24356 ( .A1(n21422), .A2(n21421), .A3(n21420), .A4(n21419), .ZN(
        n21627) );
  AOI22_X1 U24357 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(keyinput104), .B1(
        P3_EAX_REG_25__SCAN_IN), .B2(keyinput19), .ZN(n21423) );
  OAI221_X1 U24358 ( .B1(P2_UWORD_REG_3__SCAN_IN), .B2(keyinput104), .C1(
        P3_EAX_REG_25__SCAN_IN), .C2(keyinput19), .A(n21423), .ZN(n21434) );
  AOI22_X1 U24359 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(keyinput49), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(keyinput80), .ZN(n21424) );
  OAI221_X1 U24360 ( .B1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B2(keyinput49), 
        .C1(P2_EAX_REG_28__SCAN_IN), .C2(keyinput80), .A(n21424), .ZN(n21433)
         );
  AOI22_X1 U24361 ( .A1(n21427), .A2(keyinput20), .B1(keyinput39), .B2(n21426), 
        .ZN(n21425) );
  OAI221_X1 U24362 ( .B1(n21427), .B2(keyinput20), .C1(n21426), .C2(keyinput39), .A(n21425), .ZN(n21432) );
  AOI22_X1 U24363 ( .A1(n21430), .A2(keyinput76), .B1(n21429), .B2(keyinput96), 
        .ZN(n21428) );
  OAI221_X1 U24364 ( .B1(n21430), .B2(keyinput76), .C1(n21429), .C2(keyinput96), .A(n21428), .ZN(n21431) );
  NOR4_X1 U24365 ( .A1(n21434), .A2(n21433), .A3(n21432), .A4(n21431), .ZN(
        n21483) );
  AOI22_X1 U24366 ( .A1(n21437), .A2(keyinput17), .B1(n21436), .B2(keyinput12), 
        .ZN(n21435) );
  OAI221_X1 U24367 ( .B1(n21437), .B2(keyinput17), .C1(n21436), .C2(keyinput12), .A(n21435), .ZN(n21450) );
  AOI22_X1 U24368 ( .A1(n21440), .A2(keyinput93), .B1(keyinput74), .B2(n21439), 
        .ZN(n21438) );
  OAI221_X1 U24369 ( .B1(n21440), .B2(keyinput93), .C1(n21439), .C2(keyinput74), .A(n21438), .ZN(n21449) );
  AOI22_X1 U24370 ( .A1(n21443), .A2(keyinput6), .B1(n21442), .B2(keyinput47), 
        .ZN(n21441) );
  OAI221_X1 U24371 ( .B1(n21443), .B2(keyinput6), .C1(n21442), .C2(keyinput47), 
        .A(n21441), .ZN(n21448) );
  XOR2_X1 U24372 ( .A(n21444), .B(keyinput88), .Z(n21446) );
  XNOR2_X1 U24373 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B(keyinput127), .ZN(
        n21445) );
  NAND2_X1 U24374 ( .A1(n21446), .A2(n21445), .ZN(n21447) );
  NOR4_X1 U24375 ( .A1(n21450), .A2(n21449), .A3(n21448), .A4(n21447), .ZN(
        n21482) );
  INV_X1 U24376 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n21453) );
  AOI22_X1 U24377 ( .A1(n21453), .A2(keyinput78), .B1(keyinput87), .B2(n21452), 
        .ZN(n21451) );
  OAI221_X1 U24378 ( .B1(n21453), .B2(keyinput78), .C1(n21452), .C2(keyinput87), .A(n21451), .ZN(n21464) );
  AOI22_X1 U24379 ( .A1(n21456), .A2(keyinput61), .B1(keyinput107), .B2(n21455), .ZN(n21454) );
  OAI221_X1 U24380 ( .B1(n21456), .B2(keyinput61), .C1(n21455), .C2(
        keyinput107), .A(n21454), .ZN(n21463) );
  INV_X1 U24381 ( .A(DATAI_24_), .ZN(n21458) );
  AOI22_X1 U24382 ( .A1(n21459), .A2(keyinput75), .B1(keyinput91), .B2(n21458), 
        .ZN(n21457) );
  OAI221_X1 U24383 ( .B1(n21459), .B2(keyinput75), .C1(n21458), .C2(keyinput91), .A(n21457), .ZN(n21462) );
  AOI22_X1 U24384 ( .A1(n13315), .A2(keyinput120), .B1(keyinput126), .B2(
        n13180), .ZN(n21460) );
  OAI221_X1 U24385 ( .B1(n13315), .B2(keyinput120), .C1(n13180), .C2(
        keyinput126), .A(n21460), .ZN(n21461) );
  NOR4_X1 U24386 ( .A1(n21464), .A2(n21463), .A3(n21462), .A4(n21461), .ZN(
        n21481) );
  AOI22_X1 U24387 ( .A1(n21467), .A2(keyinput28), .B1(keyinput90), .B2(n21466), 
        .ZN(n21465) );
  OAI221_X1 U24388 ( .B1(n21467), .B2(keyinput28), .C1(n21466), .C2(keyinput90), .A(n21465), .ZN(n21479) );
  INV_X1 U24389 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n21470) );
  AOI22_X1 U24390 ( .A1(n21470), .A2(keyinput97), .B1(keyinput59), .B2(n21469), 
        .ZN(n21468) );
  OAI221_X1 U24391 ( .B1(n21470), .B2(keyinput97), .C1(n21469), .C2(keyinput59), .A(n21468), .ZN(n21478) );
  INV_X1 U24392 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n21472) );
  AOI22_X1 U24393 ( .A1(n21473), .A2(keyinput9), .B1(keyinput69), .B2(n21472), 
        .ZN(n21471) );
  OAI221_X1 U24394 ( .B1(n21473), .B2(keyinput9), .C1(n21472), .C2(keyinput69), 
        .A(n21471), .ZN(n21477) );
  XOR2_X1 U24395 ( .A(n12382), .B(keyinput95), .Z(n21475) );
  XNOR2_X1 U24396 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput123), .ZN(
        n21474) );
  NAND2_X1 U24397 ( .A1(n21475), .A2(n21474), .ZN(n21476) );
  NOR4_X1 U24398 ( .A1(n21479), .A2(n21478), .A3(n21477), .A4(n21476), .ZN(
        n21480) );
  NAND4_X1 U24399 ( .A1(n21483), .A2(n21482), .A3(n21481), .A4(n21480), .ZN(
        n21626) );
  AOI22_X1 U24400 ( .A1(n13596), .A2(keyinput40), .B1(keyinput66), .B2(n21485), 
        .ZN(n21484) );
  OAI221_X1 U24401 ( .B1(n13596), .B2(keyinput40), .C1(n21485), .C2(keyinput66), .A(n21484), .ZN(n21497) );
  AOI22_X1 U24402 ( .A1(n13603), .A2(keyinput100), .B1(n21487), .B2(keyinput77), .ZN(n21486) );
  OAI221_X1 U24403 ( .B1(n13603), .B2(keyinput100), .C1(n21487), .C2(
        keyinput77), .A(n21486), .ZN(n21491) );
  XNOR2_X1 U24404 ( .A(n21488), .B(keyinput23), .ZN(n21490) );
  XOR2_X1 U24405 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B(keyinput63), .Z(
        n21489) );
  OR3_X1 U24406 ( .A1(n21491), .A2(n21490), .A3(n21489), .ZN(n21496) );
  AOI22_X1 U24407 ( .A1(n21494), .A2(keyinput3), .B1(n21493), .B2(keyinput65), 
        .ZN(n21492) );
  OAI221_X1 U24408 ( .B1(n21494), .B2(keyinput3), .C1(n21493), .C2(keyinput65), 
        .A(n21492), .ZN(n21495) );
  NOR3_X1 U24409 ( .A1(n21497), .A2(n21496), .A3(n21495), .ZN(n21549) );
  AOI22_X1 U24410 ( .A1(n21500), .A2(keyinput30), .B1(keyinput2), .B2(n21499), 
        .ZN(n21498) );
  OAI221_X1 U24411 ( .B1(n21500), .B2(keyinput30), .C1(n21499), .C2(keyinput2), 
        .A(n21498), .ZN(n21513) );
  AOI22_X1 U24412 ( .A1(n21503), .A2(keyinput106), .B1(n21502), .B2(keyinput7), 
        .ZN(n21501) );
  OAI221_X1 U24413 ( .B1(n21503), .B2(keyinput106), .C1(n21502), .C2(keyinput7), .A(n21501), .ZN(n21512) );
  AOI22_X1 U24414 ( .A1(n21506), .A2(keyinput14), .B1(keyinput115), .B2(n21505), .ZN(n21504) );
  OAI221_X1 U24415 ( .B1(n21506), .B2(keyinput14), .C1(n21505), .C2(
        keyinput115), .A(n21504), .ZN(n21511) );
  INV_X1 U24416 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21508) );
  AOI22_X1 U24417 ( .A1(n21509), .A2(keyinput81), .B1(n21508), .B2(keyinput16), 
        .ZN(n21507) );
  OAI221_X1 U24418 ( .B1(n21509), .B2(keyinput81), .C1(n21508), .C2(keyinput16), .A(n21507), .ZN(n21510) );
  NOR4_X1 U24419 ( .A1(n21513), .A2(n21512), .A3(n21511), .A4(n21510), .ZN(
        n21548) );
  INV_X1 U24420 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n21515) );
  AOI22_X1 U24421 ( .A1(n21516), .A2(keyinput118), .B1(n21515), .B2(keyinput29), .ZN(n21514) );
  OAI221_X1 U24422 ( .B1(n21516), .B2(keyinput118), .C1(n21515), .C2(
        keyinput29), .A(n21514), .ZN(n21520) );
  XOR2_X1 U24423 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B(keyinput64), .Z(
        n21519) );
  XNOR2_X1 U24424 ( .A(n21517), .B(keyinput51), .ZN(n21518) );
  OR3_X1 U24425 ( .A1(n21520), .A2(n21519), .A3(n21518), .ZN(n21529) );
  AOI22_X1 U24426 ( .A1(n21523), .A2(keyinput45), .B1(n21522), .B2(keyinput48), 
        .ZN(n21521) );
  OAI221_X1 U24427 ( .B1(n21523), .B2(keyinput45), .C1(n21522), .C2(keyinput48), .A(n21521), .ZN(n21528) );
  AOI22_X1 U24428 ( .A1(n21526), .A2(keyinput21), .B1(keyinput18), .B2(n21525), 
        .ZN(n21524) );
  OAI221_X1 U24429 ( .B1(n21526), .B2(keyinput21), .C1(n21525), .C2(keyinput18), .A(n21524), .ZN(n21527) );
  NOR3_X1 U24430 ( .A1(n21529), .A2(n21528), .A3(n21527), .ZN(n21547) );
  AOI22_X1 U24431 ( .A1(n21532), .A2(keyinput13), .B1(n21531), .B2(keyinput25), 
        .ZN(n21530) );
  OAI221_X1 U24432 ( .B1(n21532), .B2(keyinput13), .C1(n21531), .C2(keyinput25), .A(n21530), .ZN(n21545) );
  AOI22_X1 U24433 ( .A1(n21535), .A2(keyinput10), .B1(n21534), .B2(keyinput116), .ZN(n21533) );
  OAI221_X1 U24434 ( .B1(n21535), .B2(keyinput10), .C1(n21534), .C2(
        keyinput116), .A(n21533), .ZN(n21544) );
  AOI22_X1 U24435 ( .A1(n21538), .A2(keyinput5), .B1(n21537), .B2(keyinput84), 
        .ZN(n21536) );
  OAI221_X1 U24436 ( .B1(n21538), .B2(keyinput5), .C1(n21537), .C2(keyinput84), 
        .A(n21536), .ZN(n21543) );
  AOI22_X1 U24437 ( .A1(n21541), .A2(keyinput82), .B1(n21540), .B2(keyinput112), .ZN(n21539) );
  OAI221_X1 U24438 ( .B1(n21541), .B2(keyinput82), .C1(n21540), .C2(
        keyinput112), .A(n21539), .ZN(n21542) );
  NOR4_X1 U24439 ( .A1(n21545), .A2(n21544), .A3(n21543), .A4(n21542), .ZN(
        n21546) );
  NAND4_X1 U24440 ( .A1(n21549), .A2(n21548), .A3(n21547), .A4(n21546), .ZN(
        n21625) );
  OAI22_X1 U24441 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(keyinput1), .B1(
        keyinput50), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21550) );
  AOI221_X1 U24442 ( .B1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput1), .C1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .C2(keyinput50), .A(n21550), .ZN(
        n21557) );
  OAI22_X1 U24443 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(keyinput42), .B1(
        BUF1_REG_15__SCAN_IN), .B2(keyinput124), .ZN(n21551) );
  AOI221_X1 U24444 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(keyinput42), .C1(
        keyinput124), .C2(BUF1_REG_15__SCAN_IN), .A(n21551), .ZN(n21556) );
  OAI22_X1 U24445 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(keyinput37), .B1(
        keyinput56), .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n21552) );
  AOI221_X1 U24446 ( .B1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput37), 
        .C1(P2_DATAO_REG_18__SCAN_IN), .C2(keyinput56), .A(n21552), .ZN(n21555) );
  OAI22_X1 U24447 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(keyinput89), .B1(
        keyinput103), .B2(P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21553) );
  AOI221_X1 U24448 ( .B1(P3_EAX_REG_27__SCAN_IN), .B2(keyinput89), .C1(
        P1_DATAWIDTH_REG_2__SCAN_IN), .C2(keyinput103), .A(n21553), .ZN(n21554) );
  NAND4_X1 U24449 ( .A1(n21557), .A2(n21556), .A3(n21555), .A4(n21554), .ZN(
        n21585) );
  OAI22_X1 U24450 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(keyinput68), .B1(
        P3_INSTQUEUE_REG_6__4__SCAN_IN), .B2(keyinput79), .ZN(n21558) );
  AOI221_X1 U24451 ( .B1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput68), 
        .C1(keyinput79), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(n21558), .ZN(
        n21565) );
  OAI22_X1 U24452 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(keyinput36), 
        .B1(keyinput99), .B2(P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n21559) );
  AOI221_X1 U24453 ( .B1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(keyinput36), 
        .C1(P1_DATAWIDTH_REG_5__SCAN_IN), .C2(keyinput99), .A(n21559), .ZN(
        n21564) );
  OAI22_X1 U24454 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(keyinput72), 
        .B1(P2_DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput83), .ZN(n21560) );
  AOI221_X1 U24455 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput72), 
        .C1(keyinput83), .C2(P2_DATAWIDTH_REG_10__SCAN_IN), .A(n21560), .ZN(
        n21563) );
  OAI22_X1 U24456 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(keyinput125), .B1(
        keyinput67), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21561) );
  AOI221_X1 U24457 ( .B1(P2_ADDRESS_REG_7__SCAN_IN), .B2(keyinput125), .C1(
        P3_INSTQUEUE_REG_14__4__SCAN_IN), .C2(keyinput67), .A(n21561), .ZN(
        n21562) );
  NAND4_X1 U24458 ( .A1(n21565), .A2(n21564), .A3(n21563), .A4(n21562), .ZN(
        n21584) );
  OAI22_X1 U24459 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput35), 
        .B1(keyinput4), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n21566) );
  AOI221_X1 U24460 ( .B1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput35), 
        .C1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .C2(keyinput4), .A(n21566), .ZN(
        n21573) );
  OAI22_X1 U24461 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(keyinput38), 
        .B1(keyinput31), .B2(BUF2_REG_30__SCAN_IN), .ZN(n21567) );
  AOI221_X1 U24462 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput38), 
        .C1(BUF2_REG_30__SCAN_IN), .C2(keyinput31), .A(n21567), .ZN(n21572) );
  OAI22_X1 U24463 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput43), .B1(
        keyinput55), .B2(P1_DATAWIDTH_REG_28__SCAN_IN), .ZN(n21568) );
  AOI221_X1 U24464 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput43), .C1(
        P1_DATAWIDTH_REG_28__SCAN_IN), .C2(keyinput55), .A(n21568), .ZN(n21571) );
  OAI22_X1 U24465 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(keyinput57), .B1(
        P3_INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput101), .ZN(n21569) );
  AOI221_X1 U24466 ( .B1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B2(keyinput57), 
        .C1(keyinput101), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(n21569), 
        .ZN(n21570) );
  NAND4_X1 U24467 ( .A1(n21573), .A2(n21572), .A3(n21571), .A4(n21570), .ZN(
        n21583) );
  OAI22_X1 U24468 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(keyinput114), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput58), .ZN(n21574) );
  AOI221_X1 U24469 ( .B1(P3_DATAO_REG_17__SCAN_IN), .B2(keyinput114), .C1(
        keyinput58), .C2(P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21574), .ZN(n21581) );
  OAI22_X1 U24470 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(keyinput86), .B1(
        P2_D_C_N_REG_SCAN_IN), .B2(keyinput105), .ZN(n21575) );
  AOI221_X1 U24471 ( .B1(P2_EBX_REG_11__SCAN_IN), .B2(keyinput86), .C1(
        keyinput105), .C2(P2_D_C_N_REG_SCAN_IN), .A(n21575), .ZN(n21580) );
  OAI22_X1 U24472 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(keyinput113), 
        .B1(P3_EBX_REG_13__SCAN_IN), .B2(keyinput22), .ZN(n21576) );
  AOI221_X1 U24473 ( .B1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput113), 
        .C1(keyinput22), .C2(P3_EBX_REG_13__SCAN_IN), .A(n21576), .ZN(n21579)
         );
  OAI22_X1 U24474 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(keyinput52), 
        .B1(keyinput122), .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n21577) );
  AOI221_X1 U24475 ( .B1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput52), 
        .C1(P1_DATAO_REG_29__SCAN_IN), .C2(keyinput122), .A(n21577), .ZN(
        n21578) );
  NAND4_X1 U24476 ( .A1(n21581), .A2(n21580), .A3(n21579), .A4(n21578), .ZN(
        n21582) );
  NOR4_X1 U24477 ( .A1(n21585), .A2(n21584), .A3(n21583), .A4(n21582), .ZN(
        n21623) );
  OAI22_X1 U24478 ( .A1(P2_ADDRESS_REG_5__SCAN_IN), .A2(keyinput53), .B1(
        keyinput121), .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n21586) );
  AOI221_X1 U24479 ( .B1(P2_ADDRESS_REG_5__SCAN_IN), .B2(keyinput53), .C1(
        P3_DATAO_REG_16__SCAN_IN), .C2(keyinput121), .A(n21586), .ZN(n21593)
         );
  OAI22_X1 U24480 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(keyinput109), .B1(
        BUF1_REG_3__SCAN_IN), .B2(keyinput34), .ZN(n21587) );
  AOI221_X1 U24481 ( .B1(P2_ADDRESS_REG_18__SCAN_IN), .B2(keyinput109), .C1(
        keyinput34), .C2(BUF1_REG_3__SCAN_IN), .A(n21587), .ZN(n21592) );
  OAI22_X1 U24482 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(keyinput46), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(keyinput32), .ZN(n21588) );
  AOI221_X1 U24483 ( .B1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B2(keyinput46), 
        .C1(keyinput32), .C2(P3_UWORD_REG_12__SCAN_IN), .A(n21588), .ZN(n21591) );
  OAI22_X1 U24484 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(keyinput33), .B1(
        keyinput108), .B2(DATAI_4_), .ZN(n21589) );
  AOI221_X1 U24485 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(keyinput33), 
        .C1(DATAI_4_), .C2(keyinput108), .A(n21589), .ZN(n21590) );
  NAND4_X1 U24486 ( .A1(n21593), .A2(n21592), .A3(n21591), .A4(n21590), .ZN(
        n21621) );
  OAI22_X1 U24487 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(keyinput41), .B1(
        keyinput70), .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n21594) );
  AOI221_X1 U24488 ( .B1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B2(keyinput41), 
        .C1(P1_UWORD_REG_4__SCAN_IN), .C2(keyinput70), .A(n21594), .ZN(n21601)
         );
  OAI22_X1 U24489 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(keyinput54), 
        .B1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput26), .ZN(n21595) );
  AOI221_X1 U24490 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput54), 
        .C1(keyinput26), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(n21595), .ZN(
        n21600) );
  OAI22_X1 U24491 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(keyinput11), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(keyinput62), .ZN(n21596) );
  AOI221_X1 U24492 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(keyinput11), .C1(
        keyinput62), .C2(P1_EAX_REG_19__SCAN_IN), .A(n21596), .ZN(n21599) );
  OAI22_X1 U24493 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(keyinput110), 
        .B1(keyinput119), .B2(BUF2_REG_14__SCAN_IN), .ZN(n21597) );
  AOI221_X1 U24494 ( .B1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B2(keyinput110), 
        .C1(BUF2_REG_14__SCAN_IN), .C2(keyinput119), .A(n21597), .ZN(n21598)
         );
  NAND4_X1 U24495 ( .A1(n21601), .A2(n21600), .A3(n21599), .A4(n21598), .ZN(
        n21620) );
  OAI22_X1 U24496 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(keyinput98), 
        .B1(P3_LWORD_REG_10__SCAN_IN), .B2(keyinput73), .ZN(n21602) );
  AOI221_X1 U24497 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput98), 
        .C1(keyinput73), .C2(P3_LWORD_REG_10__SCAN_IN), .A(n21602), .ZN(n21609) );
  OAI22_X1 U24498 ( .A1(BUF2_REG_15__SCAN_IN), .A2(keyinput8), .B1(BS16), .B2(
        keyinput44), .ZN(n21603) );
  AOI221_X1 U24499 ( .B1(BUF2_REG_15__SCAN_IN), .B2(keyinput8), .C1(keyinput44), .C2(BS16), .A(n21603), .ZN(n21608) );
  OAI22_X1 U24500 ( .A1(DATAI_31_), .A2(keyinput117), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(keyinput102), .ZN(n21604) );
  AOI221_X1 U24501 ( .B1(DATAI_31_), .B2(keyinput117), .C1(keyinput102), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n21604), .ZN(n21607) );
  OAI22_X1 U24502 ( .A1(BUF1_REG_9__SCAN_IN), .A2(keyinput0), .B1(keyinput92), 
        .B2(P2_READREQUEST_REG_SCAN_IN), .ZN(n21605) );
  AOI221_X1 U24503 ( .B1(BUF1_REG_9__SCAN_IN), .B2(keyinput0), .C1(
        P2_READREQUEST_REG_SCAN_IN), .C2(keyinput92), .A(n21605), .ZN(n21606)
         );
  NAND4_X1 U24504 ( .A1(n21609), .A2(n21608), .A3(n21607), .A4(n21606), .ZN(
        n21619) );
  OAI22_X1 U24505 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(keyinput94), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(keyinput60), .ZN(n21610) );
  AOI221_X1 U24506 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(keyinput94), .C1(
        keyinput60), .C2(P3_EBX_REG_3__SCAN_IN), .A(n21610), .ZN(n21617) );
  OAI22_X1 U24507 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(keyinput24), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(keyinput15), .ZN(n21611) );
  AOI221_X1 U24508 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput24), .C1(
        keyinput15), .C2(P1_DATAO_REG_18__SCAN_IN), .A(n21611), .ZN(n21616) );
  OAI22_X1 U24509 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(keyinput85), 
        .B1(P3_DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput71), .ZN(n21612) );
  AOI221_X1 U24510 ( .B1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput85), 
        .C1(keyinput71), .C2(P3_DATAWIDTH_REG_5__SCAN_IN), .A(n21612), .ZN(
        n21615) );
  OAI22_X1 U24511 ( .A1(P2_EAX_REG_19__SCAN_IN), .A2(keyinput27), .B1(
        keyinput111), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n21613) );
  AOI221_X1 U24512 ( .B1(P2_EAX_REG_19__SCAN_IN), .B2(keyinput27), .C1(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(keyinput111), .A(n21613), .ZN(
        n21614) );
  NAND4_X1 U24513 ( .A1(n21617), .A2(n21616), .A3(n21615), .A4(n21614), .ZN(
        n21618) );
  NOR4_X1 U24514 ( .A1(n21621), .A2(n21620), .A3(n21619), .A4(n21618), .ZN(
        n21622) );
  NAND2_X1 U24515 ( .A1(n21623), .A2(n21622), .ZN(n21624) );
  NOR4_X1 U24516 ( .A1(n21627), .A2(n21626), .A3(n21625), .A4(n21624), .ZN(
        n21628) );
  XNOR2_X1 U24517 ( .A(n21629), .B(n21628), .ZN(P3_U3018) );
  INV_X1 U13020 ( .A(n11407), .ZN(n16194) );
  INV_X2 U11359 ( .A(n16194), .ZN(n15002) );
  CLKBUF_X1 U11282 ( .A(n9852), .Z(n9853) );
  AND2_X1 U11293 ( .A1(n11832), .A2(n13805), .ZN(n11848) );
  CLKBUF_X2 U11306 ( .A(n12957), .Z(n9821) );
  CLKBUF_X1 U11316 ( .A(n10547), .Z(n20523) );
  CLKBUF_X1 U11338 ( .A(n11723), .Z(n11732) );
  NAND2_X2 U11341 ( .A1(n13974), .A2(n20501), .ZN(n21231) );
  XNOR2_X1 U11346 ( .A(n11343), .B(n20455), .ZN(n14147) );
  CLKBUF_X1 U11361 ( .A(n19485), .Z(n19466) );
  CLKBUF_X1 U11365 ( .A(n11784), .Z(n16615) );
  CLKBUF_X1 U11381 ( .A(n18945), .Z(n9866) );
  CLKBUF_X1 U11382 ( .A(n16785), .Z(n16800) );
  INV_X1 U11496 ( .A(n10150), .ZN(n9824) );
  CLKBUF_X1 U11617 ( .A(n17773), .Z(n17782) );
endmodule

